// Benchmark "systemcaes" written by ABC on Wed Apr 29 13:53:47 2015

module systemcaes ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379,
    pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389,
    pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399,
    pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409,
    pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419,
    pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429,
    pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459,
    pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469,
    pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479,
    pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489,
    pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499,
    pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509,
    pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519,
    pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549,
    pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559,
    pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569,
    pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579,
    pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589,
    pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599,
    pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609,
    pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639,
    pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649,
    pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659,
    pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669,
    pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679,
    pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689,
    pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699,
    pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729,
    pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739,
    pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749,
    pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759,
    pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769,
    pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779,
    pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789,
    pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818, pi819,
    pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828, pi829,
    pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838, pi839,
    pi840, pi841, pi842, pi843, pi844, pi845, pi846, pi847, pi848, pi849,
    pi850, pi851, pi852, pi853, pi854, pi855, pi856, pi857, pi858, pi859,
    pi860, pi861, pi862, pi863, pi864, pi865, pi866, pi867, pi868, pi869,
    pi870, pi871, pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879,
    pi880, pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908, pi909,
    pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917, pi918, pi919,
    pi920, pi921, pi922, pi923, pi924, pi925, pi926, pi927, pi928, pi929,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667, po668, po669,
    po670, po671, po672, po673, po674, po675, po676, po677, po678, po679,
    po680, po681, po682, po683, po684, po685, po686, po687, po688, po689,
    po690, po691, po692, po693, po694, po695, po696, po697, po698, po699,
    po700, po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728, po729,
    po730, po731, po732, po733, po734, po735, po736, po737, po738, po739,
    po740, po741, po742, po743, po744, po745, po746, po747, po748, po749,
    po750, po751, po752, po753, po754, po755, po756, po757, po758, po759,
    po760, po761, po762, po763, po764, po765, po766, po767, po768, po769,
    po770, po771, po772, po773, po774, po775, po776, po777, po778, po779,
    po780, po781, po782, po783, po784, po785, po786, po787, po788, po789,
    po790, po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378,
    pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388,
    pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398,
    pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408,
    pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418,
    pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428,
    pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438,
    pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468,
    pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478,
    pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488,
    pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498,
    pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508,
    pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518,
    pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528,
    pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558,
    pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568,
    pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578,
    pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588,
    pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598,
    pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608,
    pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618,
    pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648,
    pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658,
    pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668,
    pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678,
    pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688,
    pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698,
    pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708,
    pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738,
    pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748,
    pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758,
    pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768,
    pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778,
    pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788,
    pi789, pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798,
    pi799, pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828,
    pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838,
    pi839, pi840, pi841, pi842, pi843, pi844, pi845, pi846, pi847, pi848,
    pi849, pi850, pi851, pi852, pi853, pi854, pi855, pi856, pi857, pi858,
    pi859, pi860, pi861, pi862, pi863, pi864, pi865, pi866, pi867, pi868,
    pi869, pi870, pi871, pi872, pi873, pi874, pi875, pi876, pi877, pi878,
    pi879, pi880, pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888,
    pi889, pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917, pi918,
    pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926, pi927, pi928,
    pi929;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403, po404, po405, po406, po407, po408, po409,
    po410, po411, po412, po413, po414, po415, po416, po417, po418, po419,
    po420, po421, po422, po423, po424, po425, po426, po427, po428, po429,
    po430, po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458, po459,
    po460, po461, po462, po463, po464, po465, po466, po467, po468, po469,
    po470, po471, po472, po473, po474, po475, po476, po477, po478, po479,
    po480, po481, po482, po483, po484, po485, po486, po487, po488, po489,
    po490, po491, po492, po493, po494, po495, po496, po497, po498, po499,
    po500, po501, po502, po503, po504, po505, po506, po507, po508, po509,
    po510, po511, po512, po513, po514, po515, po516, po517, po518, po519,
    po520, po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548, po549,
    po550, po551, po552, po553, po554, po555, po556, po557, po558, po559,
    po560, po561, po562, po563, po564, po565, po566, po567, po568, po569,
    po570, po571, po572, po573, po574, po575, po576, po577, po578, po579,
    po580, po581, po582, po583, po584, po585, po586, po587, po588, po589,
    po590, po591, po592, po593, po594, po595, po596, po597, po598, po599,
    po600, po601, po602, po603, po604, po605, po606, po607, po608, po609,
    po610, po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638, po639,
    po640, po641, po642, po643, po644, po645, po646, po647, po648, po649,
    po650, po651, po652, po653, po654, po655, po656, po657, po658, po659,
    po660, po661, po662, po663, po664, po665, po666, po667, po668, po669,
    po670, po671, po672, po673, po674, po675, po676, po677, po678, po679,
    po680, po681, po682, po683, po684, po685, po686, po687, po688, po689,
    po690, po691, po692, po693, po694, po695, po696, po697, po698, po699,
    po700, po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728, po729,
    po730, po731, po732, po733, po734, po735, po736, po737, po738, po739,
    po740, po741, po742, po743, po744, po745, po746, po747, po748, po749,
    po750, po751, po752, po753, po754, po755, po756, po757, po758, po759,
    po760, po761, po762, po763, po764, po765, po766, po767, po768, po769,
    po770, po771, po772, po773, po774, po775, po776, po777, po778, po779,
    po780, po781, po782, po783, po784, po785, po786, po787, po788, po789,
    po790, po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818;
  wire n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
    n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
    n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2063, n2064, n2066, n2067, n2068, n2069, n2071, n2072, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2151, n2152, n2154, n2155, n2156,
    n2157, n2158, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2213, n2214, n2215, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2287, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2375, n2376,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2397, n2398,
    n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
    n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
    n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
    n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
    n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
    n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
    n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
    n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3611,
    n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
    n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3767,
    n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3782, n3783, n3784, n3785, n3786, n3787, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3843, n3844, n3845, n3846, n3847, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
    n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3900, n3901, n3902,
    n3903, n3904, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
    n4002, n4003, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4040, n4041, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4065, n4066, n4067,
    n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4180, n4181, n4182, n4183, n4184, n4186, n4187, n4189,
    n4190, n4191, n4192, n4193, n4194, n4196, n4197, n4198, n4199, n4200,
    n4202, n4203, n4204, n4205, n4206, n4207, n4209, n4210, n4211, n4212,
    n4213, n4214, n4216, n4217, n4218, n4219, n4220, n4222, n4223, n4224,
    n4225, n4226, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
    n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
    n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4337, n4338, n4339, n4340, n4341, n4342, n4344, n4345, n4346, n4347,
    n4348, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4360, n4361, n4362, n4363, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4405,
    n4406, n4407, n4408, n4409, n4410, n4411, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4692, n4693,
    n4694, n4695, n4696, n4698, n4699, n4700, n4701, n4702, n4704, n4705,
    n4706, n4707, n4708, n4710, n4711, n4712, n4713, n4714, n4716, n4717,
    n4719, n4720, n4721, n4722, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4735, n4736, n4737, n4738, n4739, n4741,
    n4742, n4743, n4744, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
    n4764, n4765, n4766, n4768, n4769, n4770, n4771, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4784, n4785, n4786,
    n4787, n4788, n4790, n4791, n4792, n4793, n4794, n4796, n4797, n4798,
    n4799, n4800, n4802, n4803, n4804, n4805, n4806, n4808, n4809, n4810,
    n4811, n4812, n4814, n4815, n4816, n4817, n4818, n4820, n4821, n4822,
    n4823, n4824, n4826, n4827, n4828, n4829, n4830, n4832, n4833, n4834,
    n4835, n4836, n4838, n4839, n4840, n4841, n4842, n4844, n4845, n4846,
    n4847, n4848, n4850, n4851, n4852, n4853, n4854, n4856, n4857, n4858,
    n4859, n4861, n4862, n4864, n4865, n4867, n4868, n4870, n4871, n4872,
    n4873, n4875, n4876, n4878, n4879, n4880, n4881, n4883, n4884, n4885,
    n4886, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4931,
    n4932, n4933, n4934, n4936, n4937, n4938, n4939, n4941, n4942, n4943,
    n4944, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
    n4955, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5012, n5013, n5014, n5015, n5017, n5018, n5019, n5020, n5022,
    n5023, n5025, n5026, n5027, n5028, n5030, n5031, n5032, n5033, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5046,
    n5047, n5048, n5049, n5051, n5052, n5053, n5054, n5055, n5057, n5058,
    n5059, n5060, n5061, n5063, n5064, n5065, n5066, n5067, n5069, n5070,
    n5071, n5072, n5073, n5075, n5076, n5078, n5079, n5080, n5081, n5082,
    n5083, n5084, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100, n5102, n5103, n5104, n5105,
    n5106, n5107, n5108, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
    n5117, n5118, n5119, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5154, n5155, n5157, n5158, n5159, n5160, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5184,
    n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5206,
    n5207, n5208, n5209, n5210, n5212, n5213, n5214, n5215, n5216, n5218,
    n5219, n5220, n5221, n5222, n5224, n5225, n5226, n5227, n5229, n5230,
    n5231, n5232, n5233, n5235, n5236, n5238, n5239, n5240, n5241, n5243,
    n5244, n5245, n5246, n5248, n5249, n5251, n5252, n5253, n5254, n5256,
    n5257, n5258, n5259, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
    n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
    n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
    n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
    n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
    n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
    n5450, n5451, n5452, n5453, n5454, n5455, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
    n5501, n5502, n5503, n5504, n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5707, n5708, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
    n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
    n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
    n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
    n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5856, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
    n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
    n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997, n5998, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6144, n6145,
    n6147, n6148, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
    n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
    n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
    n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
    n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6486, n6487, n6489, n6490, n6492, n6493, n6495, n6496, n6498,
    n6499, n6501, n6502, n6504, n6505, n6507, n6508, n6510, n6511, n6513,
    n6514, n6516, n6517, n6519, n6520, n6522, n6523, n6525, n6526, n6528,
    n6529, n6531, n6532, n6534, n6535, n6537, n6538, n6540, n6541, n6543,
    n6544, n6546, n6547, n6549, n6550, n6552, n6553, n6555, n6556, n6558,
    n6559, n6561, n6562, n6564, n6565, n6567, n6568, n6570, n6571, n6573,
    n6574, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702, n6704, n6705, n6706, n6707,
    n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
    n6738, n6739, n6740, n6741, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
    n6779, n6780, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
    n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
    n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
    n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
    n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7094, n7095, n7096, n7097,
    n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
    n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
    n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
    n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
    n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
    n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
    n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
    n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
    n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
    n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
    n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
    n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
    n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
    n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872, n7874, n7875, n7876, n7877,
    n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
    n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
    n7908, n7909, n7910, n7911, n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7952, n7953, n7955, n7956, n7958, n7959, n7961, n7962,
    n7964, n7965, n7967, n7968, n7970, n7971, n7973, n7974, n7976, n7977,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8018, n8019,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8060, n8061,
    n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
    n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
    n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
    n8092, n8093, n8094, n8095, n8096, n8097, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
    n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
    n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
    n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
    n8482, n8483, n8484, n8485, n8486, n8487, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8528, n8529, n8530, n8531, n8532, n8533,
    n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
    n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
    n8564, n8565, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
    n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
    n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682, n8684, n8685, n8686, n8687,
    n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
    n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
    n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
    n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8840, n8841,
    n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
    n8872, n8873, n8874, n8875, n8876, n8877, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
    n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
    n9108, n9109, n9110, n9111, n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9230, n9231,
    n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
    n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9308, n9309, n9311, n9312, n9314, n9315,
    n9317, n9318, n9320, n9321, n9323, n9324, n9326, n9327, n9329, n9330,
    n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
    n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
    n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9449, n9450, n9451, n9452, n9453, n9454,
    n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
    n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
    n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
    n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
    n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
    n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
    n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
    n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
    n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
    n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
    n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
    n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
    n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
    n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
    n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
    n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
    n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
    n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
    n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
    n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
    n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
    n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
    n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
    n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
    n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
    n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
    n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
    n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
    n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
    n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
    n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
    n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
    n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
    n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
    n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
    n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
    n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
    n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
    n10289, n10290, n10291, n10292, n10293, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
    n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
    n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
    n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10352, n10353,
    n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
    n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
    n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
    n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
    n10464, n10465, n10466, n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
    n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
    n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10663, n10664, n10665, n10666, n10667,
    n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
    n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
    n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
    n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
    n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
    n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
    n10852, n10853, n10854, n10855, n10856, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
    n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
    n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
    n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
    n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
    n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051, n11053, n11054, n11055,
    n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
    n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11092,
    n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
    n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
    n11166, n11167, n11168, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
    n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
    n11203, n11204, n11205, n11206, n11207, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
    n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
    n11360, n11361, n11362, n11363, n11365, n11366, n11367, n11368, n11369,
    n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
    n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
    n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
    n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
    n11480, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
    n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11521, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
    n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
    n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
    n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
    n11674, n11675, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
    n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
    n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
    n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11794,
    n11795, n11797, n11798, n11800, n11801, n11803, n11804, n11805, n11806,
    n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
    n11844, n11845, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
    n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
    n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
    n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
    n11881, n11882, n11883, n11884, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923, n11925, n11926, n11928,
    n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
    n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
    n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
    n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
    n11965, n11967, n11968, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12009, n12010, n12011, n12012,
    n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
    n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
    n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
    n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
    n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
    n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
    n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
    n12160, n12161, n12162, n12163, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
    n12197, n12198, n12199, n12200, n12201, n12202, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12243,
    n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
    n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
    n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
    n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
    n12280, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
    n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
    n12317, n12318, n12319, n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
    n12438, n12439, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
    n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
    n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
    n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
    n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
    n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
    n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
    n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
    n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
    n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
    n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
    n12565, n12566, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
    n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
    n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
    n12611, n12612, n12613, n12614, n12615, n12616, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12656, n12657,
    n12659, n12660, n12662, n12663, n12665, n12666, n12668, n12669, n12671,
    n12672, n12674, n12675, n12677, n12678, n12679, n12680, n12681, n12682,
    n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
    n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
    n12710, n12711, n12712, n12713, n12715, n12716, n12718, n12719, n12720,
    n12721, n12722, n12724, n12725, n12726, n12727, n12729, n12730, n12731,
    n12732, n12734, n12735, n12736, n12737, n12738, n12740, n12741, n12742,
    n12743, n12745, n12746, n12747, n12748, n12750, n12751, n12752, n12753,
    n12755, n12756, n12757, n12758, n12760, n12761, n12763, n12764, n12766,
    n12767, n12769, n12770, n12772, n12773, n12775, n12777, n12778, n12780,
    n12781, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833, n12835, n12836, n12837,
    n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
    n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
    n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
    n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12907, n12908, n12909, n12910, n12911, n12912,
    n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
    n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12930, n12931,
    n12932, n12933, n12935, n12936, n12937, n12938, n12940, n12941, n12942,
    n12943, n12945, n12946, n12947, n12948, n12950, n12951, n12952, n12953,
    n12955, n12956, n12957, n12958, n12960, n12961, n12962, n12963, n12964,
    n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
    n12974, n12975, n12976, n12977, n12978, n12980, n12981, n12982, n12983,
    n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
    n13003, n13004, n13005, n13006, n13008, n13009, n13010, n13011, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
    n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13065, n13066, n13067, n13068, n13069,
    n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
    n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
    n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13097,
    n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
    n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13129, n13130, n13131, n13132, n13133, n13134,
    n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
    n13182, n13183, n13184, n13185, n13186, n13187, n13189, n13190, n13191,
    n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
    n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
    n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
    n13219, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
    n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13279, n13280, n13281, n13282, n13283, n13284,
    n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
    n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
    n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13343, n13344, n13345, n13347, n13348, n13350, n13351,
    n13353, n13354, n13356, n13357, n13358, n13359, n13361, n13362, n13363,
    n13364, n13366, n13367, n13368, n13369, n13371, n13372, n13373, n13374,
    n13376, n13377, n13378, n13379, n13381, n13382, n13383, n13384, n13386,
    n13387, n13388, n13389, n13391, n13392, n13393, n13394, n13396, n13397,
    n13398, n13399, n13401, n13402, n13403, n13404, n13406, n13407, n13408,
    n13409, n13411, n13412, n13413, n13414, n13416, n13417, n13418, n13419,
    n13421, n13422, n13423, n13424, n13426, n13427, n13428, n13429, n13431,
    n13432, n13433, n13434, n13436, n13437, n13438, n13439, n13441, n13442,
    n13443, n13444, n13446, n13447, n13448, n13449, n13451, n13452, n13453,
    n13454, n13456, n13457, n13458, n13459, n13461, n13462, n13463, n13464,
    n13466, n13467, n13468, n13469, n13471, n13472, n13474, n13475, n13476,
    n13477, n13479, n13480, n13481, n13482, n13484, n13485, n13486, n13487,
    n13489, n13490, n13491, n13492, n13494, n13495, n13496, n13497, n13499,
    n13500, n13501, n13502, n13504, n13505, n13506, n13507, n13509, n13510,
    n13511, n13512, n13514, n13515, n13516, n13517, n13519, n13520, n13521,
    n13522, n13524, n13525, n13526, n13527, n13529, n13530, n13531, n13532,
    n13534, n13535, n13536, n13537, n13539, n13540, n13541, n13542, n13544,
    n13545, n13546, n13547, n13549, n13550, n13552, n13553, n13555, n13556,
    n13558, n13559, n13560, n13561, n13563, n13564, n13565, n13566, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
    n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
    n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
    n13624, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
    n13672, n13673, n13675, n13676, n13678, n13679, n13681, n13682, n13684,
    n13685, n13687, n13688, n13690, n13691, n13693, n13694, n13696, n13697,
    n13698, n13699, n13701, n13702, n13704, n13705, n13706, n13707, n13709,
    n13710, n13711, n13712, n13714, n13715, n13717, n13718, n13720, n13721,
    n13722, n13723, n13725, n13726, n13728, n13729, n13731, n13732, n13734,
    n13735, n13736, n13737, n13739, n13740, n13741, n13742, n13744, n13745,
    n13747, n13748, n13750, n13751, n13753, n13754, n13756, n13757, n13758,
    n13759, n13761, n13762, n13764, n13765, n13767, n13768, n13769, n13770,
    n13772, n13773, n13775, n13776, n13778, n13779, n13781, n13782, n13784,
    n13785, n13786, n13788, n13789, n13790, n13792, n13793, n13794, n13796,
    n13797, n13798, n13800, n13801, n13802, n13804, n13805, n13806, n13807,
    n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
    n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
    n13826, n13827, n13829, n13831, n13832, n13833, n13834, n13835, n13836,
    n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
    n13846, n13847, n13848, n13849, n13850, n13852, n13853, n13854, n13855,
    n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
    n13865, n13866, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13889, n13890, n13891, n13892, n13893,
    n13894, n13895, n13896, n13897, n13899, n13900, n13902, n13903, n13904,
    n13906, n13907, n13909, n13910, n13911, n13914, n13915, n13916, n13917,
    n13918, n13920, n13921, n13922, n13923, n13924, n13926, n13927, n13928,
    n13929, n13931, n13932, n13933, n13934, n13935, n13936, n13938, n13940,
    n13942, n13944, n13946, n13948, n13950, n13952, n13954, n13956, n13958,
    n13960, n13962, n13964, n13966, n13968, n13970, n13972, n13974, n13976,
    n13978, n13980, n13982, n13984, n13986, n13988, n13990, n13992, n13994,
    n13996, n13998, n14000, n14002, n14004, n14006, n14008, n14010, n14012,
    n14014, n14016, n14018, n14020, n14022, n14024, n14026, n14028, n14030,
    n14032, n14034, n14036, n14038, n14040, n14042, n14044, n14046, n14048,
    n14050, n14052, n14054, n14056, n14058, n14060, n14062, n14064, n14066,
    n14068, n14070, n14072, n14074, n14076, n14078, n14080, n14082, n14084,
    n14086, n14088, n14090, n14092, n14094, n14096, n14098, n14100, n14102,
    n14104, n14106, n14108, n14110, n14112, n14114, n14116, n14118, n14120,
    n14122, n14124, n14126, n14128, n14130, n14132, n14133;
  assign n1751 = ~pi555 & ~pi557;
  assign n1752 = ~pi556 & n1751;
  assign n1753 = ~pi558 & n1752;
  assign n1754 = pi559 & n1753;
  assign n1755 = ~pi551 & ~pi552;
  assign n1756 = ~pi550 & n1755;
  assign n1757 = pi000 & ~n1756;
  assign n1758 = pi813 & n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = n1754 & ~n1759;
  assign n1761 = pi559 & ~n1753;
  assign n1762 = pi813 & n1761;
  assign n1763 = pi390 & pi557;
  assign n1764 = ~pi390 & ~pi557;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = pi551 & pi558;
  assign n1767 = ~pi551 & ~pi558;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = ~n1765 & ~n1768;
  assign n1770 = pi552 & pi556;
  assign n1771 = ~pi552 & ~pi556;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = pi550 & pi555;
  assign n1774 = ~pi550 & ~pi555;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1772 & ~n1775;
  assign n1777 = n1769 & n1776;
  assign n1778 = pi665 & ~n1777;
  assign n1779 = pi000 & n1778;
  assign n1780 = ~n1759 & ~n1778;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = ~n1761 & ~n1781;
  assign n1783 = ~n1762 & ~n1782;
  assign n1784 = ~n1754 & ~n1783;
  assign n1785 = ~n1760 & ~n1784;
  assign n1786 = pi845 & n1761;
  assign n1787 = ~n1761 & n1778;
  assign n1788 = pi012 & n1787;
  assign n1789 = ~n1786 & ~n1788;
  assign n1790 = ~n1754 & ~n1789;
  assign n1791 = ~n1761 & ~n1778;
  assign n1792 = ~n1754 & ~n1791;
  assign n1793 = pi845 & n1756;
  assign n1794 = pi012 & ~n1756;
  assign n1795 = ~n1793 & ~n1794;
  assign n1796 = ~n1792 & ~n1795;
  assign n1797 = ~n1790 & ~n1796;
  assign n1798 = pi005 & pi006;
  assign n1799 = pi005 & pi008;
  assign n1800 = pi006 & n1799;
  assign n1801 = n1798 & ~n1800;
  assign n1802 = ~n1798 & n1800;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = pi005 & pi007;
  assign n1805 = ~pi006 & n1804;
  assign n1806 = pi006 & ~n1804;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = pi007 & pi008;
  assign n1809 = ~n1799 & n1808;
  assign n1810 = n1799 & ~n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n1807 & n1811;
  assign n1813 = n1807 & ~n1811;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = ~n1803 & n1814;
  assign n1816 = n1803 & ~n1814;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = ~pi178 & pi195;
  assign n1819 = pi178 & ~pi195;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = ~n1817 & ~n1820;
  assign n1822 = pi006 & pi008;
  assign n1823 = pi006 & n1808;
  assign n1824 = ~n1822 & n1823;
  assign n1825 = n1822 & ~n1823;
  assign n1826 = ~n1824 & ~n1825;
  assign n1827 = pi006 & ~n1808;
  assign n1828 = ~pi006 & n1808;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~pi007 & n1799;
  assign n1831 = pi007 & ~n1799;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = n1829 & ~n1832;
  assign n1834 = ~n1829 & n1832;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~n1826 & n1835;
  assign n1837 = n1826 & ~n1835;
  assign n1838 = ~n1836 & ~n1837;
  assign n1839 = pi164 & ~pi195;
  assign n1840 = ~pi164 & pi195;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~n1838 & ~n1841;
  assign n1843 = ~n1821 & n1842;
  assign n1844 = n1821 & ~n1842;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~pi164 & ~pi190;
  assign n1847 = pi164 & pi190;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = pi006 & pi007;
  assign n1850 = n1798 & ~n1849;
  assign n1851 = ~n1798 & n1849;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~pi005 & ~pi007;
  assign n1854 = ~n1804 & ~n1853;
  assign n1855 = n1806 & ~n1854;
  assign n1856 = ~n1806 & ~n1853;
  assign n1857 = ~n1804 & n1856;
  assign n1858 = ~n1855 & ~n1857;
  assign n1859 = n1822 & n1858;
  assign n1860 = ~n1822 & ~n1858;
  assign n1861 = ~n1859 & ~n1860;
  assign n1862 = ~n1852 & n1861;
  assign n1863 = n1852 & ~n1861;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = n1848 & ~n1864;
  assign n1866 = ~n1804 & n1808;
  assign n1867 = n1804 & ~n1808;
  assign n1868 = ~n1866 & ~n1867;
  assign n1869 = pi007 & n1799;
  assign n1870 = pi008 & n1858;
  assign n1871 = ~pi008 & ~n1858;
  assign n1872 = ~n1870 & ~n1871;
  assign n1873 = ~n1869 & n1872;
  assign n1874 = n1869 & ~n1872;
  assign n1875 = ~n1873 & ~n1874;
  assign n1876 = n1868 & n1875;
  assign n1877 = ~n1868 & ~n1875;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = pi190 & ~n1878;
  assign n1880 = pi164 & ~n1838;
  assign n1881 = pi190 & ~n1864;
  assign n1882 = ~n1880 & n1881;
  assign n1883 = n1880 & ~n1881;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = pi195 & ~n1817;
  assign n1886 = pi178 & ~n1878;
  assign n1887 = n1885 & n1886;
  assign n1888 = ~n1885 & ~n1886;
  assign n1889 = ~n1887 & ~n1888;
  assign n1890 = ~n1884 & n1889;
  assign n1891 = n1884 & ~n1889;
  assign n1892 = ~n1890 & ~n1891;
  assign n1893 = ~n1879 & n1892;
  assign n1894 = n1879 & ~n1892;
  assign n1895 = ~n1893 & ~n1894;
  assign n1896 = ~n1865 & n1895;
  assign n1897 = n1865 & ~n1895;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n1845 & n1898;
  assign n1900 = n1845 & ~n1898;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = pi190 & ~n1838;
  assign n1903 = ~n1820 & ~n1864;
  assign n1904 = ~n1902 & n1903;
  assign n1905 = n1902 & ~n1903;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = pi164 & ~n1817;
  assign n1908 = pi195 & ~n1878;
  assign n1909 = ~n1907 & n1908;
  assign n1910 = n1907 & ~n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1906 & n1911;
  assign n1913 = n1906 & ~n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = n1817 & n1838;
  assign n1916 = ~n1817 & ~n1838;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = pi192 & n1917;
  assign n1919 = n1838 & ~n1864;
  assign n1920 = ~n1838 & n1864;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = pi110 & ~n1921;
  assign n1923 = ~n1918 & n1922;
  assign n1924 = n1918 & ~n1922;
  assign n1925 = ~n1923 & ~n1924;
  assign n1926 = pi132 & ~n1817;
  assign n1927 = n1864 & n1878;
  assign n1928 = ~n1864 & ~n1878;
  assign n1929 = ~n1927 & ~n1928;
  assign n1930 = pi165 & n1929;
  assign n1931 = n1926 & n1930;
  assign n1932 = ~n1926 & ~n1930;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = n1925 & n1933;
  assign n1935 = ~n1925 & ~n1933;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = n1914 & n1936;
  assign n1938 = ~n1914 & ~n1936;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = n1901 & ~n1939;
  assign n1941 = ~n1901 & n1939;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = ~n1841 & ~n1864;
  assign n1944 = ~n1820 & ~n1838;
  assign n1945 = ~n1943 & n1944;
  assign n1946 = n1943 & ~n1944;
  assign n1947 = ~n1945 & ~n1946;
  assign n1948 = pi164 & ~n1878;
  assign n1949 = pi190 & ~n1817;
  assign n1950 = n1948 & ~n1949;
  assign n1951 = ~n1948 & n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = n1845 & n1898;
  assign n1954 = ~n1845 & ~n1898;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n1936 & n1955;
  assign n1957 = n1936 & ~n1955;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = n1952 & n1958;
  assign n1960 = ~n1952 & ~n1958;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = n1947 & n1961;
  assign n1963 = ~n1947 & ~n1961;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = ~n1942 & n1964;
  assign n1966 = n1942 & ~n1964;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = pi110 & ~n1838;
  assign n1969 = pi192 & ~n1817;
  assign n1970 = ~n1968 & n1969;
  assign n1971 = n1968 & ~n1969;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = pi165 & ~n1864;
  assign n1974 = pi132 & ~n1878;
  assign n1975 = ~n1973 & n1974;
  assign n1976 = n1973 & ~n1974;
  assign n1977 = ~n1975 & ~n1976;
  assign n1978 = ~n1892 & ~n1977;
  assign n1979 = n1892 & n1977;
  assign n1980 = ~n1978 & ~n1979;
  assign n1981 = n1972 & n1980;
  assign n1982 = ~n1972 & ~n1980;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = ~n1901 & ~n1914;
  assign n1985 = n1901 & n1914;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = n1983 & n1986;
  assign n1988 = ~n1983 & ~n1986;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = pi192 & ~n1921;
  assign n1991 = pi110 & n1929;
  assign n1992 = ~n1990 & n1991;
  assign n1993 = n1990 & ~n1991;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = pi132 & ~n1838;
  assign n1996 = pi165 & ~n1817;
  assign n1997 = ~n1995 & n1996;
  assign n1998 = n1995 & ~n1996;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = n1994 & ~n1999;
  assign n2001 = ~n1994 & n1999;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~n1901 & ~n2002;
  assign n2004 = n1901 & n2002;
  assign n2005 = ~n2003 & ~n2004;
  assign n2006 = ~n1914 & n2005;
  assign n2007 = n1914 & ~n2005;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~n1989 & n2008;
  assign n2010 = ~n1983 & n1986;
  assign n2011 = n1983 & ~n1986;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n2008 & ~n2012;
  assign n2014 = ~n2009 & ~n2013;
  assign n2015 = n1967 & ~n2014;
  assign n2016 = ~n1967 & n2014;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~pi553 & ~pi554;
  assign n2019 = ~pi668 & n2018;
  assign n2020 = ~n1754 & n1778;
  assign n2021 = ~n1754 & n1761;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = n2019 & ~n2022;
  assign n2024 = ~pi553 & ~pi668;
  assign n2025 = pi554 & ~n2024;
  assign n2026 = ~n2019 & ~n2025;
  assign n2027 = ~n2023 & ~n2026;
  assign n2028 = pi673 & n2027;
  assign n2029 = ~n2017 & ~n2028;
  assign n2030 = ~n1964 & n2028;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = pi909 & n1761;
  assign n2033 = pi909 & n1756;
  assign n2034 = ~pi133 & ~n1756;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = ~n1778 & ~n2035;
  assign n2037 = ~pi133 & n1778;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~n1761 & ~n2038;
  assign n2040 = ~n2032 & ~n2039;
  assign n2041 = ~n1754 & ~n2040;
  assign n2042 = n1754 & ~n2035;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = n2031 & ~n2043;
  assign n2045 = ~n2031 & n2043;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = pi877 & n1756;
  assign n2048 = pi045 & ~n1756;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = ~n1778 & ~n2049;
  assign n2051 = pi045 & n1778;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = ~n1761 & ~n2052;
  assign n2054 = pi877 & n1761;
  assign n2055 = ~n2053 & ~n2054;
  assign n2056 = ~n1754 & ~n2055;
  assign n2057 = n1754 & ~n2049;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = ~n2046 & n2058;
  assign n2060 = ~n2045 & ~n2058;
  assign n2061 = ~n2044 & n2060;
  assign po187 = n2059 | n2061;
  assign n2063 = ~n1797 & ~po187;
  assign n2064 = n1797 & po187;
  assign po144 = n2063 | n2064;
  assign n2066 = ~n1785 & ~po144;
  assign n2067 = n1785 & po144;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~pi553 & pi554;
  assign po814 = ~pi668 & n2069;
  assign n2071 = ~n2068 & po814;
  assign n2072 = pi000 & ~po814;
  assign po132 = n2071 | n2072;
  assign n2074 = pi001 & ~n1756;
  assign n2075 = pi814 & n1756;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = n1754 & ~n2076;
  assign n2078 = pi814 & n1761;
  assign n2079 = pi001 & n1778;
  assign n2080 = ~n1778 & ~n2076;
  assign n2081 = ~n2079 & ~n2080;
  assign n2082 = ~n1761 & ~n2081;
  assign n2083 = ~n2078 & ~n2082;
  assign n2084 = ~n1754 & ~n2083;
  assign n2085 = ~n2077 & ~n2084;
  assign n2086 = pi846 & n1761;
  assign n2087 = pi013 & n1787;
  assign n2088 = ~n2086 & ~n2087;
  assign n2089 = ~n1754 & ~n2088;
  assign n2090 = pi846 & n1756;
  assign n2091 = pi013 & ~n1756;
  assign n2092 = ~n2090 & ~n2091;
  assign n2093 = ~n1792 & ~n2092;
  assign n2094 = ~n2089 & ~n2093;
  assign n2095 = pi110 & ~n1817;
  assign n2096 = pi192 & n1929;
  assign n2097 = ~n2095 & n2096;
  assign n2098 = n2095 & ~n2096;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = pi165 & ~n1838;
  assign n2101 = pi132 & ~n1864;
  assign n2102 = n2100 & n2101;
  assign n2103 = ~n2100 & ~n2101;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = n2099 & n2104;
  assign n2106 = ~n2099 & ~n2104;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = n1942 & ~n2107;
  assign n2109 = ~n1942 & n2107;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n1989 & n2110;
  assign n2112 = ~n2012 & ~n2110;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n1967 & n2113;
  assign n2115 = n1967 & ~n2113;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = ~n2028 & ~n2116;
  assign n2118 = n2028 & ~n2110;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = pi910 & n1761;
  assign n2121 = pi910 & n1756;
  assign n2122 = ~pi134 & ~n1756;
  assign n2123 = ~n2121 & ~n2122;
  assign n2124 = ~n1778 & ~n2123;
  assign n2125 = ~pi134 & n1778;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n1761 & ~n2126;
  assign n2128 = ~n2120 & ~n2127;
  assign n2129 = ~n1754 & ~n2128;
  assign n2130 = n1754 & ~n2123;
  assign n2131 = ~n2129 & ~n2130;
  assign n2132 = n2119 & ~n2131;
  assign n2133 = ~n2119 & n2131;
  assign n2134 = ~n2132 & ~n2133;
  assign n2135 = pi878 & n1756;
  assign n2136 = pi044 & ~n1756;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n1778 & ~n2137;
  assign n2139 = pi044 & n1778;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = ~n1761 & ~n2140;
  assign n2142 = pi878 & n1761;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = ~n1754 & ~n2143;
  assign n2145 = n1754 & ~n2137;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = ~n2134 & n2146;
  assign n2148 = ~n2133 & ~n2146;
  assign n2149 = ~n2132 & n2148;
  assign po185 = n2147 | n2149;
  assign n2151 = ~n2094 & ~po185;
  assign n2152 = n2094 & po185;
  assign po147 = n2151 | n2152;
  assign n2154 = ~n2085 & ~po147;
  assign n2155 = n2085 & po147;
  assign n2156 = ~n2154 & ~n2155;
  assign n2157 = po814 & ~n2156;
  assign n2158 = pi001 & ~po814;
  assign po133 = n2157 | n2158;
  assign n2160 = pi014 & ~n1756;
  assign n2161 = pi847 & n1756;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~n1792 & ~n2162;
  assign n2164 = pi847 & n1761;
  assign n2165 = pi014 & n1787;
  assign n2166 = ~n2164 & ~n2165;
  assign n2167 = ~n1754 & ~n2166;
  assign n2168 = ~n2163 & ~n2167;
  assign n2169 = pi167 & n1778;
  assign n2170 = pi911 & n1756;
  assign n2171 = pi167 & ~n1756;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = ~n1778 & ~n2172;
  assign n2174 = ~n2169 & ~n2173;
  assign n2175 = ~n1761 & ~n2174;
  assign n2176 = pi911 & n1761;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = ~n1754 & n2177;
  assign n2179 = n1754 & n2172;
  assign n2180 = ~n2178 & ~n2179;
  assign n2181 = n1967 & n1986;
  assign n2182 = ~n1967 & ~n1986;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = ~n2005 & n2110;
  assign n2185 = n2005 & ~n2110;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2028 & n2186;
  assign n2188 = ~n2183 & n2187;
  assign n2189 = ~n2005 & n2028;
  assign n2190 = ~n2028 & ~n2186;
  assign n2191 = ~n2182 & n2190;
  assign n2192 = ~n2181 & n2191;
  assign n2193 = ~n2189 & ~n2192;
  assign n2194 = ~n2188 & n2193;
  assign n2195 = n2180 & n2194;
  assign n2196 = ~n2180 & ~n2194;
  assign po315 = n2195 | n2196;
  assign n2198 = pi879 & n1756;
  assign n2199 = pi048 & ~n1756;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = ~n1778 & ~n2200;
  assign n2202 = pi048 & n1778;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = ~n1761 & ~n2203;
  assign n2205 = pi879 & n1761;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = ~n1754 & ~n2206;
  assign n2208 = n1754 & ~n2200;
  assign n2209 = ~n2207 & ~n2208;
  assign n2210 = ~po315 & ~n2209;
  assign n2211 = po315 & n2209;
  assign po191 = n2210 | n2211;
  assign n2213 = n2168 & po191;
  assign n2214 = ~n2168 & ~n2211;
  assign n2215 = ~n2210 & n2214;
  assign po149 = n2213 | n2215;
  assign n2217 = pi815 & n1756;
  assign n2218 = pi002 & ~n1756;
  assign n2219 = ~n2217 & ~n2218;
  assign n2220 = n1754 & ~n2219;
  assign n2221 = pi815 & n1761;
  assign n2222 = ~n1778 & ~n2219;
  assign n2223 = pi002 & n1778;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~n1761 & ~n2224;
  assign n2226 = ~n2221 & ~n2225;
  assign n2227 = ~n1754 & ~n2226;
  assign n2228 = ~n2220 & ~n2227;
  assign n2229 = po149 & n2228;
  assign n2230 = ~n2213 & ~n2228;
  assign n2231 = ~n2215 & n2230;
  assign n2232 = ~n2229 & ~n2231;
  assign n2233 = po814 & ~n2232;
  assign n2234 = pi002 & ~po814;
  assign po134 = n2233 | n2234;
  assign n2236 = pi166 & n1778;
  assign n2237 = pi912 & n1756;
  assign n2238 = pi166 & ~n1756;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~n1778 & ~n2239;
  assign n2241 = ~n2236 & ~n2240;
  assign n2242 = ~n1761 & ~n2241;
  assign n2243 = pi912 & n1761;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = ~n1754 & n2244;
  assign n2246 = n1754 & n2239;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n1892 & n2107;
  assign n2249 = ~n1892 & ~n2107;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = ~n1939 & n2002;
  assign n2252 = n1939 & ~n2002;
  assign n2253 = ~n2251 & ~n2252;
  assign n2254 = ~n2250 & n2253;
  assign n2255 = n2250 & ~n2253;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = n2028 & n2256;
  assign n2258 = ~n1967 & n2256;
  assign n2259 = n1967 & ~n2256;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = n2186 & ~n2260;
  assign n2262 = ~n2028 & n2261;
  assign n2263 = n2190 & n2260;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = ~n2257 & n2264;
  assign n2266 = n2247 & n2265;
  assign n2267 = ~n2247 & ~n2265;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = pi880 & n1756;
  assign n2270 = pi049 & ~n1756;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = n1754 & ~n2271;
  assign n2273 = ~n1778 & ~n2271;
  assign n2274 = pi049 & n1778;
  assign n2275 = ~n2273 & ~n2274;
  assign n2276 = ~n1761 & ~n2275;
  assign n2277 = pi880 & n1761;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~n1754 & ~n2278;
  assign n2280 = ~n2272 & ~n2279;
  assign n2281 = n2268 & ~n2280;
  assign n2282 = ~n2257 & ~n2263;
  assign n2283 = ~n2262 & n2282;
  assign n2284 = n2247 & n2283;
  assign n2285 = ~n2247 & ~n2283;
  assign po313 = n2284 | n2285;
  assign n2287 = n2280 & po313;
  assign po193 = n2281 | n2287;
  assign n2289 = pi848 & n1761;
  assign n2290 = pi015 & n1787;
  assign n2291 = ~n2289 & ~n2290;
  assign n2292 = ~n1754 & ~n2291;
  assign n2293 = pi015 & ~n1756;
  assign n2294 = pi848 & n1756;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = ~n1792 & ~n2295;
  assign n2297 = ~n2292 & ~n2296;
  assign n2298 = ~po193 & ~n2297;
  assign n2299 = po193 & n2297;
  assign po151 = n2298 | n2299;
  assign n2301 = pi816 & n1756;
  assign n2302 = pi003 & ~n1756;
  assign n2303 = ~n2301 & ~n2302;
  assign n2304 = n1754 & ~n2303;
  assign n2305 = pi816 & n1761;
  assign n2306 = ~n1778 & ~n2303;
  assign n2307 = pi003 & n1778;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n1761 & ~n2308;
  assign n2310 = ~n2305 & ~n2309;
  assign n2311 = ~n1754 & ~n2310;
  assign n2312 = ~n2304 & ~n2311;
  assign n2313 = po151 & n2312;
  assign n2314 = ~po151 & ~n2312;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = po814 & ~n2315;
  assign n2317 = pi003 & ~po814;
  assign po135 = n2316 | n2317;
  assign n2319 = pi016 & ~n1756;
  assign n2320 = pi849 & n1756;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = ~n1792 & ~n2321;
  assign n2323 = pi849 & n1761;
  assign n2324 = pi016 & n1787;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = ~n1754 & ~n2325;
  assign n2327 = ~n2322 & ~n2326;
  assign n2328 = n2008 & ~n2256;
  assign n2329 = ~n2008 & n2256;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = ~n1964 & n2186;
  assign n2332 = n1964 & ~n2186;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = ~n2028 & n2333;
  assign n2335 = n2330 & n2334;
  assign n2336 = ~n2028 & ~n2256;
  assign n2337 = n2008 & ~n2336;
  assign n2338 = ~n2028 & n2256;
  assign n2339 = ~n2008 & ~n2338;
  assign n2340 = ~n2337 & ~n2339;
  assign n2341 = ~n2008 & n2028;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = ~n2334 & ~n2342;
  assign n2344 = ~n2335 & ~n2343;
  assign n2345 = pi913 & n1761;
  assign n2346 = pi913 & n1756;
  assign n2347 = ~pi155 & ~n1756;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n1778 & ~n2348;
  assign n2350 = ~pi155 & n1778;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n1761 & ~n2351;
  assign n2353 = ~n2345 & ~n2352;
  assign n2354 = ~n1754 & ~n2353;
  assign n2355 = n1754 & ~n2348;
  assign n2356 = ~n2354 & ~n2355;
  assign n2357 = ~n2344 & n2356;
  assign n2358 = n2344 & ~n2356;
  assign n2359 = ~n2357 & ~n2358;
  assign n2360 = pi881 & n1756;
  assign n2361 = pi057 & ~n1756;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = ~n1778 & ~n2362;
  assign n2364 = pi057 & n1778;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n1761 & ~n2365;
  assign n2367 = pi881 & n1761;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n1754 & ~n2368;
  assign n2370 = n1754 & ~n2362;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = n2359 & ~n2371;
  assign n2373 = ~n2359 & n2371;
  assign po203 = n2372 | n2373;
  assign n2375 = n2327 & po203;
  assign n2376 = ~n2327 & ~po203;
  assign po153 = n2375 | n2376;
  assign n2378 = ~pi817 & n1756;
  assign n2379 = ~pi004 & ~n1756;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = n1754 & n2380;
  assign n2382 = pi817 & n1761;
  assign n2383 = ~n1778 & n2380;
  assign n2384 = pi004 & n1778;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = ~n1761 & ~n2385;
  assign n2387 = ~n2382 & ~n2386;
  assign n2388 = ~n1754 & ~n2387;
  assign n2389 = ~n2381 & ~n2388;
  assign n2390 = po153 & ~n2389;
  assign n2391 = ~n2375 & n2389;
  assign n2392 = ~n2376 & n2391;
  assign n2393 = ~n2390 & ~n2392;
  assign n2394 = po814 & n2393;
  assign n2395 = pi004 & ~po814;
  assign po136 = n2394 | n2395;
  assign n2397 = pi668 & n2018;
  assign n2398 = ~n2312 & n2397;
  assign n2399 = pi824 & n1756;
  assign n2400 = pi221 & ~n1756;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = n1754 & n2401;
  assign n2403 = ~n1778 & ~n2401;
  assign n2404 = pi221 & n1778;
  assign n2405 = ~n2403 & ~n2404;
  assign n2406 = ~n1761 & ~n2405;
  assign n2407 = pi824 & n1761;
  assign n2408 = ~n1754 & ~n2407;
  assign n2409 = ~n2406 & n2408;
  assign n2410 = ~n2402 & ~n2409;
  assign n2411 = ~pi554 & ~pi668;
  assign n2412 = pi553 & n2411;
  assign n2413 = n2410 & n2412;
  assign n2414 = ~pi832 & n1756;
  assign n2415 = ~pi199 & ~n1756;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = n1754 & n2416;
  assign n2418 = pi832 & n1761;
  assign n2419 = ~n1778 & n2416;
  assign n2420 = pi199 & n1778;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = ~n1761 & ~n2421;
  assign n2423 = ~n2418 & ~n2422;
  assign n2424 = ~n1754 & ~n2423;
  assign n2425 = ~n2417 & ~n2424;
  assign n2426 = n2023 & ~n2425;
  assign n2427 = pi808 & n1756;
  assign n2428 = pi209 & ~n1756;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = n1754 & n2429;
  assign n2431 = ~n1778 & ~n2429;
  assign n2432 = pi209 & n1778;
  assign n2433 = ~n2431 & ~n2432;
  assign n2434 = ~n1761 & ~n2433;
  assign n2435 = pi808 & n1761;
  assign n2436 = ~n1754 & ~n2435;
  assign n2437 = ~n2434 & n2436;
  assign n2438 = ~n2430 & ~n2437;
  assign n2439 = pi553 & ~pi554;
  assign n2440 = pi668 & n2439;
  assign n2441 = n2438 & n2440;
  assign n2442 = ~n2426 & ~n2441;
  assign n2443 = ~n2413 & n2442;
  assign n2444 = ~n2398 & n2443;
  assign n2445 = ~n2027 & ~n2444;
  assign n2446 = pi555 & pi558;
  assign n2447 = ~pi556 & ~pi557;
  assign n2448 = n2446 & n2447;
  assign n2449 = pi673 & ~n2448;
  assign n2450 = pi598 & n2449;
  assign n2451 = pi370 & ~n2449;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = ~pi565 & pi566;
  assign n2454 = pi563 & ~pi567;
  assign n2455 = n2453 & n2454;
  assign n2456 = ~n2452 & n2455;
  assign n2457 = pi658 & n2449;
  assign n2458 = pi381 & ~n2449;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = pi563 & pi567;
  assign n2461 = pi565 & ~pi566;
  assign n2462 = n2460 & n2461;
  assign n2463 = ~n2459 & n2462;
  assign n2464 = ~n2456 & ~n2463;
  assign n2465 = ~pi565 & ~pi566;
  assign n2466 = n2454 & n2465;
  assign n2467 = pi391 & ~n2449;
  assign n2468 = pi629 & n2449;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = n2466 & ~n2469;
  assign n2471 = pi573 & n2449;
  assign n2472 = pi284 & ~n2449;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = ~pi563 & pi567;
  assign n2475 = n2465 & n2474;
  assign n2476 = ~n2473 & n2475;
  assign n2477 = ~n2470 & ~n2476;
  assign n2478 = pi533 & n2449;
  assign n2479 = pi360 & ~n2449;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = pi565 & pi566;
  assign n2482 = n2454 & n2481;
  assign n2483 = ~n2480 & n2482;
  assign n2484 = pi639 & n2449;
  assign n2485 = pi320 & ~n2449;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = ~pi563 & ~pi567;
  assign n2488 = n2453 & n2487;
  assign n2489 = ~n2486 & n2488;
  assign n2490 = ~n2483 & ~n2489;
  assign n2491 = pi577 & n2449;
  assign n2492 = pi361 & ~n2449;
  assign n2493 = ~n2491 & ~n2492;
  assign n2494 = pi566 & n2460;
  assign n2495 = ~pi565 & n2494;
  assign n2496 = ~n2493 & n2495;
  assign n2497 = pi640 & n2449;
  assign n2498 = pi398 & ~n2449;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = n2454 & n2461;
  assign n2501 = ~n2499 & n2500;
  assign n2502 = ~n2496 & ~n2501;
  assign n2503 = pi601 & n2449;
  assign n2504 = pi280 & ~n2449;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = n2465 & n2487;
  assign n2507 = ~n2505 & n2506;
  assign n2508 = pi593 & n2449;
  assign n2509 = pi260 & ~n2449;
  assign n2510 = ~n2508 & ~n2509;
  assign n2511 = n2453 & n2474;
  assign n2512 = ~n2510 & n2511;
  assign n2513 = ~n2507 & ~n2512;
  assign n2514 = pi538 & n2449;
  assign n2515 = pi256 & ~n2449;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = pi565 & n2494;
  assign n2518 = ~n2516 & n2517;
  assign n2519 = pi622 & n2449;
  assign n2520 = pi278 & ~n2449;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2461 & n2474;
  assign n2523 = ~n2521 & n2522;
  assign n2524 = ~n2518 & ~n2523;
  assign n2525 = n2513 & n2524;
  assign n2526 = n2502 & n2525;
  assign n2527 = n2490 & n2526;
  assign n2528 = pi539 & n2449;
  assign n2529 = pi329 & ~n2449;
  assign n2530 = ~n2528 & ~n2529;
  assign n2531 = n2474 & n2481;
  assign n2532 = ~n2530 & n2531;
  assign n2533 = pi534 & n2449;
  assign n2534 = pi311 & ~n2449;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = n2481 & n2487;
  assign n2537 = ~n2535 & n2536;
  assign n2538 = ~n2532 & ~n2537;
  assign n2539 = n2527 & n2538;
  assign n2540 = ~pi566 & n2487;
  assign n2541 = pi565 & n2540;
  assign n2542 = pi302 & ~n2449;
  assign n2543 = pi619 & n2449;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = n2541 & ~n2544;
  assign n2546 = pi570 & n2449;
  assign n2547 = pi362 & ~n2449;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = n2460 & n2465;
  assign n2550 = ~n2548 & n2549;
  assign n2551 = ~n2545 & ~n2550;
  assign n2552 = n2539 & n2551;
  assign n2553 = n2477 & n2552;
  assign n2554 = n2464 & n2553;
  assign n2555 = ~pi565 & n2540;
  assign n2556 = pi568 & n2555;
  assign n2557 = ~pi565 & ~pi568;
  assign n2558 = n2540 & n2557;
  assign n2559 = ~n2556 & ~n2558;
  assign n2560 = ~n2554 & n2559;
  assign n2561 = ~n2505 & n2558;
  assign n2562 = pi673 & n1753;
  assign n2563 = ~pi673 & n2448;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = ~pi562 & ~n2564;
  assign n2566 = pi435 & n2448;
  assign n2567 = pi673 & n2566;
  assign n2568 = ~pi666 & pi673;
  assign n2569 = ~pi435 & ~pi673;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2567 & ~n2570;
  assign n2572 = ~n2565 & ~n2571;
  assign n2573 = n2561 & n2572;
  assign n2574 = ~n2560 & ~n2573;
  assign n2575 = n2027 & ~n2574;
  assign n2576 = ~n2445 & ~n2575;
  assign n2577 = pi606 & n2449;
  assign n2578 = pi377 & ~n2449;
  assign n2579 = ~n2577 & ~n2578;
  assign n2580 = n2549 & ~n2579;
  assign n2581 = pi587 & n2449;
  assign n2582 = pi343 & ~n2449;
  assign n2583 = ~n2581 & ~n2582;
  assign n2584 = n2462 & ~n2583;
  assign n2585 = ~n2580 & ~n2584;
  assign n2586 = pi403 & ~n2449;
  assign n2587 = pi651 & n2449;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = n2466 & ~n2588;
  assign n2590 = pi571 & n2449;
  assign n2591 = pi265 & ~n2449;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = n2475 & ~n2592;
  assign n2594 = ~n2589 & ~n2593;
  assign n2595 = pi588 & n2449;
  assign n2596 = pi354 & ~n2449;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = n2495 & ~n2597;
  assign n2599 = pi596 & n2449;
  assign n2600 = pi383 & ~n2449;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = n2500 & ~n2601;
  assign n2603 = ~n2598 & ~n2602;
  assign n2604 = pi518 & n2449;
  assign n2605 = pi386 & ~n2449;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2482 & ~n2606;
  assign n2608 = pi600 & n2449;
  assign n2609 = pi392 & ~n2449;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = n2488 & ~n2610;
  assign n2612 = ~n2607 & ~n2611;
  assign n2613 = pi653 & n2449;
  assign n2614 = pi324 & ~n2449;
  assign n2615 = ~n2613 & ~n2614;
  assign n2616 = n2506 & ~n2615;
  assign n2617 = pi659 & n2449;
  assign n2618 = pi304 & ~n2449;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = n2511 & ~n2619;
  assign n2621 = ~n2616 & ~n2620;
  assign n2622 = pi520 & n2449;
  assign n2623 = pi303 & ~n2449;
  assign n2624 = ~n2622 & ~n2623;
  assign n2625 = n2517 & ~n2624;
  assign n2626 = pi652 & n2449;
  assign n2627 = pi271 & ~n2449;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = n2522 & ~n2628;
  assign n2630 = ~n2625 & ~n2629;
  assign n2631 = n2621 & n2630;
  assign n2632 = n2612 & n2631;
  assign n2633 = n2603 & n2632;
  assign n2634 = pi521 & n2449;
  assign n2635 = pi258 & ~n2449;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = n2536 & ~n2636;
  assign n2638 = pi523 & n2449;
  assign n2639 = pi323 & ~n2449;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = n2531 & ~n2640;
  assign n2642 = ~n2637 & ~n2641;
  assign n2643 = n2633 & n2642;
  assign n2644 = pi286 & ~n2449;
  assign n2645 = pi586 & n2449;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = n2541 & ~n2646;
  assign n2648 = pi635 & n2449;
  assign n2649 = pi367 & ~n2449;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2455 & ~n2650;
  assign n2652 = ~n2647 & ~n2651;
  assign n2653 = n2643 & n2652;
  assign n2654 = n2594 & n2653;
  assign n2655 = n2585 & n2654;
  assign n2656 = n2559 & ~n2655;
  assign n2657 = n2558 & ~n2615;
  assign n2658 = n2572 & n2657;
  assign n2659 = ~n2656 & ~n2658;
  assign n2660 = n2027 & ~n2659;
  assign n2661 = ~pi811 & n1756;
  assign n2662 = ~pi011 & ~n1756;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n1754 & n2663;
  assign n2665 = pi811 & n1761;
  assign n2666 = ~n1778 & n2663;
  assign n2667 = pi011 & n1778;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n1761 & ~n2668;
  assign n2670 = ~n2665 & ~n2669;
  assign n2671 = ~n1754 & ~n2670;
  assign n2672 = ~n2664 & ~n2671;
  assign n2673 = n2397 & ~n2672;
  assign n2674 = pi211 & ~n1756;
  assign n2675 = pi803 & n1756;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = n1754 & ~n2676;
  assign n2678 = pi803 & n1761;
  assign n2679 = pi211 & n1778;
  assign n2680 = ~n1778 & ~n2676;
  assign n2681 = ~n2679 & ~n2680;
  assign n2682 = ~n1761 & ~n2681;
  assign n2683 = ~n2678 & ~n2682;
  assign n2684 = ~n1754 & ~n2683;
  assign n2685 = ~n2677 & ~n2684;
  assign n2686 = n2440 & ~n2685;
  assign n2687 = pi819 & n1761;
  assign n2688 = pi216 & n1778;
  assign n2689 = pi216 & ~n1756;
  assign n2690 = pi819 & n1756;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = ~n1778 & ~n2691;
  assign n2693 = ~n2688 & ~n2692;
  assign n2694 = ~n1761 & ~n2693;
  assign n2695 = ~n2687 & ~n2694;
  assign n2696 = ~n1754 & ~n2695;
  assign n2697 = n1754 & ~n2691;
  assign n2698 = ~n2696 & ~n2697;
  assign n2699 = n2412 & ~n2698;
  assign n2700 = ~n2686 & ~n2699;
  assign n2701 = ~pi827 & n1756;
  assign n2702 = ~pi202 & ~n1756;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = n1754 & n2703;
  assign n2705 = pi827 & n1761;
  assign n2706 = ~n1778 & n2703;
  assign n2707 = pi202 & n1778;
  assign n2708 = ~n2706 & ~n2707;
  assign n2709 = ~n1761 & ~n2708;
  assign n2710 = ~n2705 & ~n2709;
  assign n2711 = ~n1754 & ~n2710;
  assign n2712 = ~n2704 & ~n2711;
  assign n2713 = n2023 & ~n2712;
  assign n2714 = n2700 & ~n2713;
  assign n2715 = ~n2673 & n2714;
  assign n2716 = ~n2027 & ~n2715;
  assign n2717 = ~n2660 & ~n2716;
  assign n2718 = pi572 & n2449;
  assign n2719 = pi276 & ~n2449;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = n2475 & ~n2720;
  assign n2722 = pi610 & n2449;
  assign n2723 = pi371 & ~n2449;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = n2455 & ~n2724;
  assign n2726 = ~n2721 & ~n2725;
  assign n2727 = pi468 & n2449;
  assign n2728 = pi309 & ~n2449;
  assign n2729 = ~n2727 & ~n2728;
  assign n2730 = n2536 & ~n2729;
  assign n2731 = pi466 & n2449;
  assign n2732 = pi327 & ~n2449;
  assign n2733 = ~n2731 & ~n2732;
  assign n2734 = n2531 & ~n2733;
  assign n2735 = ~n2730 & ~n2734;
  assign n2736 = pi630 & n2449;
  assign n2737 = pi384 & ~n2449;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = n2500 & ~n2738;
  assign n2740 = pi637 & n2449;
  assign n2741 = pi275 & ~n2449;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = n2522 & ~n2742;
  assign n2744 = ~n2739 & ~n2743;
  assign n2745 = pi467 & n2449;
  assign n2746 = pi355 & ~n2449;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n2482 & ~n2747;
  assign n2749 = pi469 & n2449;
  assign n2750 = pi326 & ~n2449;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = n2517 & ~n2751;
  assign n2753 = ~n2748 & ~n2752;
  assign n2754 = pi642 & n2449;
  assign n2755 = pi300 & ~n2449;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = n2506 & ~n2756;
  assign n2758 = pi627 & n2449;
  assign n2759 = pi401 & ~n2449;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = n2495 & ~n2760;
  assign n2762 = ~n2757 & ~n2761;
  assign n2763 = pi654 & n2449;
  assign n2764 = pi316 & ~n2449;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = n2488 & ~n2765;
  assign n2767 = pi608 & n2449;
  assign n2768 = pi257 & ~n2449;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = n2511 & ~n2769;
  assign n2771 = ~n2766 & ~n2770;
  assign n2772 = n2762 & n2771;
  assign n2773 = n2753 & n2772;
  assign n2774 = n2744 & n2773;
  assign n2775 = pi616 & n2449;
  assign n2776 = pi378 & ~n2449;
  assign n2777 = ~n2775 & ~n2776;
  assign n2778 = n2462 & ~n2777;
  assign n2779 = pi656 & n2449;
  assign n2780 = pi253 & ~n2449;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = n2541 & ~n2781;
  assign n2783 = ~n2778 & ~n2782;
  assign n2784 = n2774 & n2783;
  assign n2785 = pi365 & ~n2449;
  assign n2786 = pi597 & n2449;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = n2466 & ~n2787;
  assign n2789 = pi664 & n2449;
  assign n2790 = pi342 & ~n2449;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = n2549 & ~n2791;
  assign n2793 = ~n2788 & ~n2792;
  assign n2794 = n2784 & n2793;
  assign n2795 = n2735 & n2794;
  assign n2796 = n2726 & n2795;
  assign n2797 = n2559 & ~n2796;
  assign n2798 = n2558 & ~n2756;
  assign n2799 = n2572 & n2798;
  assign n2800 = ~n2797 & ~n2799;
  assign n2801 = n2027 & ~n2800;
  assign n2802 = ~pi806 & n1756;
  assign n2803 = ~pi207 & ~n1756;
  assign n2804 = ~n2802 & ~n2803;
  assign n2805 = n1754 & n2804;
  assign n2806 = pi806 & n1761;
  assign n2807 = ~n1778 & n2804;
  assign n2808 = pi207 & n1778;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n1761 & ~n2809;
  assign n2811 = ~n2806 & ~n2810;
  assign n2812 = ~n1754 & ~n2811;
  assign n2813 = ~n2805 & ~n2812;
  assign n2814 = n2440 & ~n2813;
  assign n2815 = pi196 & ~n1756;
  assign n2816 = pi830 & n1756;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n1778 & ~n2817;
  assign n2819 = pi196 & n1778;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = ~n1761 & ~n2820;
  assign n2822 = pi830 & n1761;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = ~n1754 & ~n2823;
  assign n2825 = n1754 & ~n2817;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = n2023 & ~n2826;
  assign n2828 = ~n2085 & n2397;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = pi822 & n1756;
  assign n2831 = pi222 & ~n1756;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n1778 & ~n2832;
  assign n2834 = pi222 & n1778;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = ~n1761 & ~n2835;
  assign n2837 = pi822 & n1761;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n1754 & ~n2838;
  assign n2840 = n1754 & ~n2832;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = n2412 & ~n2841;
  assign n2843 = n2829 & ~n2842;
  assign n2844 = ~n2814 & n2843;
  assign n2845 = ~n2027 & ~n2844;
  assign n2846 = ~n2801 & ~n2845;
  assign n2847 = n2717 & ~n2846;
  assign n2848 = ~n2717 & n2846;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = ~n2576 & ~n2849;
  assign n2851 = n2576 & ~n2848;
  assign n2852 = ~n2847 & n2851;
  assign n2853 = ~n2850 & ~n2852;
  assign n2854 = n2028 & n2853;
  assign n2855 = ~n2389 & n2397;
  assign n2856 = ~pi833 & n1756;
  assign n2857 = ~pi201 & ~n1756;
  assign n2858 = ~n2856 & ~n2857;
  assign n2859 = n1754 & n2858;
  assign n2860 = pi833 & n1761;
  assign n2861 = ~n1778 & n2858;
  assign n2862 = pi201 & n1778;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = ~n1761 & ~n2863;
  assign n2865 = ~n2860 & ~n2864;
  assign n2866 = ~n1754 & ~n2865;
  assign n2867 = ~n2859 & ~n2866;
  assign n2868 = n2023 & ~n2867;
  assign n2869 = pi825 & n1761;
  assign n2870 = pi212 & n1778;
  assign n2871 = pi212 & ~n1756;
  assign n2872 = pi825 & n1756;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = ~n1778 & ~n2873;
  assign n2875 = ~n2870 & ~n2874;
  assign n2876 = ~n1761 & ~n2875;
  assign n2877 = ~n2869 & ~n2876;
  assign n2878 = ~n1754 & ~n2877;
  assign n2879 = n1754 & ~n2873;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = n2412 & ~n2880;
  assign n2882 = ~pi809 & n1756;
  assign n2883 = ~pi213 & ~n1756;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = n1754 & n2884;
  assign n2886 = pi809 & n1761;
  assign n2887 = ~n1778 & n2884;
  assign n2888 = pi213 & n1778;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = ~n1761 & ~n2889;
  assign n2891 = ~n2886 & ~n2890;
  assign n2892 = ~n1754 & ~n2891;
  assign n2893 = ~n2885 & ~n2892;
  assign n2894 = n2440 & ~n2893;
  assign n2895 = ~n2881 & ~n2894;
  assign n2896 = ~n2868 & n2895;
  assign n2897 = ~n2855 & n2896;
  assign n2898 = ~n2027 & ~n2897;
  assign n2899 = n2027 & n2559;
  assign n2900 = pi589 & n2449;
  assign n2901 = pi399 & ~n2449;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = n2495 & ~n2902;
  assign n2904 = pi618 & n2449;
  assign n2905 = pi385 & ~n2449;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = n2500 & ~n2906;
  assign n2908 = ~n2903 & ~n2907;
  assign n2909 = pi547 & n2449;
  assign n2910 = pi363 & ~n2449;
  assign n2911 = ~n2909 & ~n2910;
  assign n2912 = n2482 & ~n2911;
  assign n2913 = pi661 & n2449;
  assign n2914 = pi321 & ~n2449;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n2488 & ~n2915;
  assign n2917 = ~n2912 & ~n2916;
  assign n2918 = pi660 & n2449;
  assign n2919 = pi281 & ~n2449;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n2506 & ~n2920;
  assign n2922 = pi662 & n2449;
  assign n2923 = pi261 & ~n2449;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = n2511 & ~n2924;
  assign n2926 = ~n2921 & ~n2925;
  assign n2927 = pi546 & n2449;
  assign n2928 = pi308 & ~n2449;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = n2517 & ~n2929;
  assign n2931 = pi605 & n2449;
  assign n2932 = pi279 & ~n2449;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = n2522 & ~n2933;
  assign n2935 = ~n2930 & ~n2934;
  assign n2936 = n2926 & n2935;
  assign n2937 = n2917 & n2936;
  assign n2938 = n2908 & n2937;
  assign n2939 = pi375 & ~n2449;
  assign n2940 = pi614 & n2449;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n2466 & ~n2941;
  assign n2943 = pi649 & n2449;
  assign n2944 = pi254 & ~n2449;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = n2475 & ~n2945;
  assign n2947 = ~n2942 & ~n2946;
  assign n2948 = pi548 & n2449;
  assign n2949 = pi313 & ~n2449;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n2536 & ~n2950;
  assign n2952 = pi549 & n2449;
  assign n2953 = pi331 & ~n2449;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = n2531 & ~n2954;
  assign n2956 = ~n2951 & ~n2955;
  assign n2957 = pi611 & n2449;
  assign n2958 = pi344 & ~n2449;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = n2549 & ~n2959;
  assign n2961 = pi632 & n2449;
  assign n2962 = pi372 & ~n2449;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n2455 & ~n2963;
  assign n2965 = ~n2960 & ~n2964;
  assign n2966 = pi255 & ~n2449;
  assign n2967 = pi646 & n2449;
  assign n2968 = ~n2966 & ~n2967;
  assign n2969 = n2541 & ~n2968;
  assign n2970 = pi617 & n2449;
  assign n2971 = pi382 & ~n2449;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = n2462 & ~n2972;
  assign n2974 = ~n2969 & ~n2973;
  assign n2975 = n2965 & n2974;
  assign n2976 = n2956 & n2975;
  assign n2977 = n2947 & n2976;
  assign n2978 = n2938 & n2977;
  assign n2979 = n2899 & ~n2978;
  assign n2980 = ~n2898 & ~n2979;
  assign n2981 = n2027 & n2572;
  assign n2982 = n2558 & n2981;
  assign n2983 = ~n2920 & n2982;
  assign n2984 = n2980 & ~n2983;
  assign n2985 = ~n2028 & ~n2984;
  assign n2986 = ~n2854 & ~n2985;
  assign n2987 = pi826 & n1756;
  assign n2988 = pi200 & ~n1756;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = ~n1778 & ~n2989;
  assign n2991 = pi200 & n1778;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = ~n1761 & ~n2992;
  assign n2994 = pi826 & n1761;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = ~n1754 & ~n2995;
  assign n2997 = n1754 & ~n2989;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = n2023 & ~n2998;
  assign n3000 = pi818 & n1756;
  assign n3001 = pi217 & ~n1756;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = n1754 & n3002;
  assign n3004 = pi818 & n1761;
  assign n3005 = ~n1754 & ~n3004;
  assign n3006 = ~n1778 & ~n3002;
  assign n3007 = pi217 & n1778;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = ~n1761 & ~n3008;
  assign n3010 = n3005 & ~n3009;
  assign n3011 = ~n3003 & ~n3010;
  assign n3012 = n2412 & n3011;
  assign n3013 = ~n2999 & ~n3012;
  assign n3014 = ~pi810 & n1756;
  assign n3015 = ~pi009 & ~n1756;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = n1754 & n3016;
  assign n3018 = ~n1778 & n3016;
  assign n3019 = pi009 & n1778;
  assign n3020 = ~n3018 & ~n3019;
  assign n3021 = ~n1761 & ~n3020;
  assign n3022 = pi810 & n1761;
  assign n3023 = ~n3021 & ~n3022;
  assign n3024 = ~n1754 & ~n3023;
  assign n3025 = ~n3017 & ~n3024;
  assign n3026 = n2397 & ~n3025;
  assign n3027 = pi802 & n1756;
  assign n3028 = pi210 & ~n1756;
  assign n3029 = ~n3027 & ~n3028;
  assign n3030 = ~n1778 & ~n3029;
  assign n3031 = pi210 & n1778;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = ~n1761 & ~n3032;
  assign n3034 = pi802 & n1761;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = ~n1754 & ~n3035;
  assign n3037 = n1754 & ~n3029;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = n2440 & ~n3038;
  assign n3040 = ~n3026 & ~n3039;
  assign n3041 = n3013 & n3040;
  assign n3042 = ~n2027 & ~n3041;
  assign n3043 = pi643 & n2449;
  assign n3044 = pi374 & ~n2449;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n2462 & ~n3045;
  assign n3047 = pi541 & n2449;
  assign n3048 = pi306 & ~n2449;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = n2536 & ~n3049;
  assign n3051 = ~n3046 & ~n3050;
  assign n3052 = pi352 & ~n2449;
  assign n3053 = pi574 & n2449;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = n2466 & ~n3054;
  assign n3056 = pi620 & n2449;
  assign n3057 = pi376 & ~n2449;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = n2549 & ~n3058;
  assign n3060 = ~n3055 & ~n3059;
  assign n3061 = pi648 & n2449;
  assign n3062 = pi299 & ~n2449;
  assign n3063 = ~n3061 & ~n3062;
  assign n3064 = n2522 & ~n3063;
  assign n3065 = pi540 & n2449;
  assign n3066 = pi266 & ~n2449;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = n2517 & ~n3067;
  assign n3069 = ~n3064 & ~n3068;
  assign n3070 = pi582 & n2449;
  assign n3071 = pi307 & ~n2449;
  assign n3072 = ~n3070 & ~n3071;
  assign n3073 = n2511 & ~n3072;
  assign n3074 = pi599 & n2449;
  assign n3075 = pi373 & ~n2449;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n2488 & ~n3076;
  assign n3078 = ~n3073 & ~n3077;
  assign n3079 = pi647 & n2449;
  assign n3080 = pi322 & ~n2449;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n2506 & ~n3081;
  assign n3083 = pi595 & n2449;
  assign n3084 = pi353 & ~n2449;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = n2495 & ~n3085;
  assign n3087 = ~n3082 & ~n3086;
  assign n3088 = pi535 & n2449;
  assign n3089 = pi400 & ~n2449;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n2482 & ~n3090;
  assign n3092 = pi583 & n2449;
  assign n3093 = pi408 & ~n2449;
  assign n3094 = ~n3092 & ~n3093;
  assign n3095 = n2500 & ~n3094;
  assign n3096 = ~n3091 & ~n3095;
  assign n3097 = n3087 & n3096;
  assign n3098 = n3078 & n3097;
  assign n3099 = n3069 & n3098;
  assign n3100 = pi623 & n2449;
  assign n3101 = pi366 & ~n2449;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = n2455 & ~n3102;
  assign n3104 = pi604 & n2449;
  assign n3105 = pi330 & ~n2449;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = n2541 & ~n3106;
  assign n3108 = ~n3103 & ~n3107;
  assign n3109 = n3099 & n3108;
  assign n3110 = pi527 & n2449;
  assign n3111 = pi264 & ~n2449;
  assign n3112 = ~n3110 & ~n3111;
  assign n3113 = n2531 & ~n3112;
  assign n3114 = pi569 & n2449;
  assign n3115 = pi310 & ~n2449;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n2475 & ~n3116;
  assign n3118 = ~n3113 & ~n3117;
  assign n3119 = n3109 & n3118;
  assign n3120 = n3060 & n3119;
  assign n3121 = n3051 & n3120;
  assign n3122 = n2559 & ~n3121;
  assign n3123 = n2558 & ~n3081;
  assign n3124 = n2572 & n3123;
  assign n3125 = ~n3122 & ~n3124;
  assign n3126 = n2027 & ~n3125;
  assign n3127 = ~n3042 & ~n3126;
  assign n3128 = pi218 & ~n1756;
  assign n3129 = pi821 & n1756;
  assign n3130 = ~n3128 & ~n3129;
  assign n3131 = n1754 & ~n3130;
  assign n3132 = pi821 & n1761;
  assign n3133 = ~n1778 & ~n3130;
  assign n3134 = pi218 & n1778;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n1761 & ~n3135;
  assign n3137 = ~n3132 & ~n3136;
  assign n3138 = ~n1754 & ~n3137;
  assign n3139 = ~n3131 & ~n3138;
  assign n3140 = n2412 & ~n3139;
  assign n3141 = ~pi829 & n1756;
  assign n3142 = ~pi197 & ~n1756;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = n1754 & n3143;
  assign n3145 = pi829 & n1761;
  assign n3146 = pi197 & n1778;
  assign n3147 = ~n1778 & n3143;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = ~n1761 & ~n3148;
  assign n3150 = ~n3145 & ~n3149;
  assign n3151 = ~n1754 & ~n3150;
  assign n3152 = ~n3144 & ~n3151;
  assign n3153 = n2023 & ~n3152;
  assign n3154 = ~n3140 & ~n3153;
  assign n3155 = pi805 & n1761;
  assign n3156 = pi206 & n1778;
  assign n3157 = pi206 & ~n1756;
  assign n3158 = pi805 & n1756;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = ~n1778 & ~n3159;
  assign n3161 = ~n3156 & ~n3160;
  assign n3162 = ~n1761 & ~n3161;
  assign n3163 = ~n3155 & ~n3162;
  assign n3164 = ~n1754 & ~n3163;
  assign n3165 = n1754 & ~n3159;
  assign n3166 = ~n3164 & ~n3165;
  assign n3167 = n2440 & ~n3166;
  assign n3168 = ~n1785 & n2397;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = n3154 & n3169;
  assign n3171 = ~n2027 & ~n3170;
  assign n3172 = pi636 & n2449;
  assign n3173 = pi268 & ~n2449;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = n2475 & ~n3174;
  assign n3176 = pi510 & n2449;
  assign n3177 = pi319 & ~n2449;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = n2531 & ~n3178;
  assign n3180 = ~n3175 & ~n3179;
  assign n3181 = pi581 & n2449;
  assign n3182 = pi379 & ~n2449;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = n2549 & ~n3183;
  assign n3185 = pi625 & n2449;
  assign n3186 = pi368 & ~n2449;
  assign n3187 = ~n3185 & ~n3186;
  assign n3188 = n2455 & ~n3187;
  assign n3189 = ~n3184 & ~n3188;
  assign n3190 = pi633 & n2449;
  assign n3191 = pi405 & ~n2449;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = n2500 & ~n3192;
  assign n3194 = pi644 & n2449;
  assign n3195 = pi341 & ~n2449;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = n2511 & ~n3196;
  assign n3198 = ~n3193 & ~n3197;
  assign n3199 = pi576 & n2449;
  assign n3200 = pi357 & ~n2449;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = n2495 & ~n3201;
  assign n3203 = pi607 & n2449;
  assign n3204 = pi274 & ~n2449;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = n2522 & ~n3205;
  assign n3207 = ~n3202 & ~n3206;
  assign n3208 = pi624 & n2449;
  assign n3209 = pi272 & ~n2449;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n2506 & ~n3210;
  assign n3212 = pi584 & n2449;
  assign n3213 = pi315 & ~n2449;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = n2488 & ~n3214;
  assign n3216 = ~n3211 & ~n3215;
  assign n3217 = pi511 & n2449;
  assign n3218 = pi404 & ~n2449;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = n2482 & ~n3219;
  assign n3221 = pi493 & n2449;
  assign n3222 = pi270 & ~n2449;
  assign n3223 = ~n3221 & ~n3222;
  assign n3224 = n2517 & ~n3223;
  assign n3225 = ~n3220 & ~n3224;
  assign n3226 = n3216 & n3225;
  assign n3227 = n3207 & n3226;
  assign n3228 = n3198 & n3227;
  assign n3229 = pi509 & n2449;
  assign n3230 = pi340 & ~n2449;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = n2536 & ~n3231;
  assign n3233 = pi621 & n2449;
  assign n3234 = pi364 & ~n2449;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = n2466 & ~n3235;
  assign n3237 = ~n3232 & ~n3236;
  assign n3238 = n3228 & n3237;
  assign n3239 = pi287 & ~n2449;
  assign n3240 = pi631 & n2449;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = n2541 & ~n3241;
  assign n3243 = pi663 & n2449;
  assign n3244 = pi346 & ~n2449;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = n2462 & ~n3245;
  assign n3247 = ~n3242 & ~n3246;
  assign n3248 = n3238 & n3247;
  assign n3249 = n3189 & n3248;
  assign n3250 = n3180 & n3249;
  assign n3251 = n2559 & ~n3250;
  assign n3252 = n2558 & ~n3210;
  assign n3253 = n2572 & n3252;
  assign n3254 = ~n3251 & ~n3253;
  assign n3255 = n2027 & ~n3254;
  assign n3256 = ~n3171 & ~n3255;
  assign n3257 = ~n2576 & n3256;
  assign n3258 = n2576 & ~n3256;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = ~n3127 & n3259;
  assign n3261 = n3127 & ~n3259;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = n2028 & ~n3262;
  assign n3264 = ~n2028 & ~n2717;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = ~n2986 & n3265;
  assign n3267 = n2986 & ~n3265;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = n2849 & ~n2984;
  assign n3270 = ~n2849 & n2984;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = n2028 & n3271;
  assign n3273 = pi650 & n2449;
  assign n3274 = pi317 & ~n2449;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = n2462 & ~n3275;
  assign n3277 = pi525 & n2449;
  assign n3278 = pi282 & ~n2449;
  assign n3279 = ~n3277 & ~n3278;
  assign n3280 = n2531 & ~n3279;
  assign n3281 = ~n3276 & ~n3280;
  assign n3282 = pi397 & ~n2449;
  assign n3283 = pi657 & n2449;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = n2466 & ~n3284;
  assign n3286 = pi591 & n2449;
  assign n3287 = pi267 & ~n2449;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = n2475 & ~n3288;
  assign n3290 = ~n3285 & ~n3289;
  assign n3291 = pi634 & n2449;
  assign n3292 = pi356 & ~n2449;
  assign n3293 = ~n3291 & ~n3292;
  assign n3294 = n2495 & ~n3293;
  assign n3295 = pi641 & n2449;
  assign n3296 = pi406 & ~n2449;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = n2500 & ~n3297;
  assign n3299 = ~n3294 & ~n3298;
  assign n3300 = pi519 & n2449;
  assign n3301 = pi407 & ~n2449;
  assign n3302 = ~n3300 & ~n3301;
  assign n3303 = n2482 & ~n3302;
  assign n3304 = pi602 & n2449;
  assign n3305 = pi314 & ~n2449;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = n2488 & ~n3306;
  assign n3308 = ~n3303 & ~n3307;
  assign n3309 = pi594 & n2449;
  assign n3310 = pi269 & ~n2449;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = n2506 & ~n3311;
  assign n3313 = pi603 & n2449;
  assign n3314 = pi305 & ~n2449;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = n2511 & ~n3315;
  assign n3317 = ~n3312 & ~n3316;
  assign n3318 = pi524 & n2449;
  assign n3319 = pi312 & ~n2449;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = n2517 & ~n3320;
  assign n3322 = pi638 & n2449;
  assign n3323 = pi273 & ~n2449;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = n2522 & ~n3324;
  assign n3326 = ~n3321 & ~n3325;
  assign n3327 = n3317 & n3326;
  assign n3328 = n3308 & n3327;
  assign n3329 = n3299 & n3328;
  assign n3330 = pi522 & n2449;
  assign n3331 = pi262 & ~n2449;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = n2536 & ~n3332;
  assign n3334 = pi626 & n2449;
  assign n3335 = pi285 & ~n2449;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = n2541 & ~n3336;
  assign n3338 = ~n3333 & ~n3337;
  assign n3339 = n3329 & n3338;
  assign n3340 = pi579 & n2449;
  assign n3341 = pi345 & ~n2449;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = n2549 & ~n3342;
  assign n3344 = pi580 & n2449;
  assign n3345 = pi395 & ~n2449;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = n2455 & ~n3346;
  assign n3348 = ~n3343 & ~n3347;
  assign n3349 = n3339 & n3348;
  assign n3350 = n3290 & n3349;
  assign n3351 = n3281 & n3350;
  assign n3352 = n2559 & ~n3351;
  assign n3353 = n2558 & ~n3311;
  assign n3354 = n2572 & n3353;
  assign n3355 = ~n3352 & ~n3354;
  assign n3356 = n2027 & ~n3355;
  assign n3357 = ~pi828 & n1756;
  assign n3358 = ~pi203 & ~n1756;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = n1754 & n3359;
  assign n3361 = pi828 & n1761;
  assign n3362 = ~n1778 & n3359;
  assign n3363 = pi203 & n1778;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n1761 & ~n3364;
  assign n3366 = ~n3361 & ~n3365;
  assign n3367 = ~n1754 & ~n3366;
  assign n3368 = ~n3360 & ~n3367;
  assign n3369 = n2023 & ~n3368;
  assign n3370 = pi820 & n1761;
  assign n3371 = pi219 & n1778;
  assign n3372 = pi219 & ~n1756;
  assign n3373 = pi820 & n1756;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = ~n1778 & ~n3374;
  assign n3376 = ~n3371 & ~n3375;
  assign n3377 = ~n1761 & ~n3376;
  assign n3378 = ~n3370 & ~n3377;
  assign n3379 = ~n1754 & ~n3378;
  assign n3380 = n1754 & ~n3374;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = n2412 & ~n3381;
  assign n3383 = pi804 & n1761;
  assign n3384 = pi205 & n1778;
  assign n3385 = pi205 & ~n1756;
  assign n3386 = pi804 & n1756;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n1778 & ~n3387;
  assign n3389 = ~n3384 & ~n3388;
  assign n3390 = ~n1761 & ~n3389;
  assign n3391 = ~n3383 & ~n3390;
  assign n3392 = ~n1754 & ~n3391;
  assign n3393 = n1754 & ~n3387;
  assign n3394 = ~n3392 & ~n3393;
  assign n3395 = n2440 & ~n3394;
  assign n3396 = pi812 & n1761;
  assign n3397 = pi010 & n1778;
  assign n3398 = pi010 & ~n1756;
  assign n3399 = pi812 & n1756;
  assign n3400 = ~n3398 & ~n3399;
  assign n3401 = ~n1778 & ~n3400;
  assign n3402 = ~n3397 & ~n3401;
  assign n3403 = ~n1761 & ~n3402;
  assign n3404 = ~n3396 & ~n3403;
  assign n3405 = ~n1754 & ~n3404;
  assign n3406 = n1754 & ~n3400;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = n2397 & ~n3407;
  assign n3409 = ~n3395 & ~n3408;
  assign n3410 = ~n3382 & n3409;
  assign n3411 = ~n3369 & n3410;
  assign n3412 = ~n2027 & ~n3411;
  assign n3413 = ~n3356 & ~n3412;
  assign n3414 = ~n2028 & ~n3413;
  assign n3415 = ~n3272 & ~n3414;
  assign n3416 = ~n3265 & ~n3415;
  assign n3417 = n3265 & n3415;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = ~n3268 & ~n3418;
  assign n3420 = n3268 & n3418;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = ~n2984 & n3413;
  assign n3423 = n2984 & ~n3413;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n2846 & n3424;
  assign n3426 = n2846 & ~n3424;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n2028 & ~n3427;
  assign n3429 = ~pi831 & n1756;
  assign n3430 = ~pi198 & ~n1756;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = n1754 & n3431;
  assign n3433 = pi831 & n1761;
  assign n3434 = ~n1778 & n3431;
  assign n3435 = pi198 & n1778;
  assign n3436 = ~n3434 & ~n3435;
  assign n3437 = ~n1761 & ~n3436;
  assign n3438 = ~n3433 & ~n3437;
  assign n3439 = ~n1754 & ~n3438;
  assign n3440 = ~n3432 & ~n3439;
  assign n3441 = n2023 & ~n3440;
  assign n3442 = ~pi807 & n1756;
  assign n3443 = ~pi208 & ~n1756;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = ~n1778 & n3444;
  assign n3446 = pi208 & n1778;
  assign n3447 = ~n3445 & ~n3446;
  assign n3448 = ~n1761 & ~n3447;
  assign n3449 = pi807 & n1761;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~n1754 & n3450;
  assign n3452 = n1754 & ~n3444;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = n2440 & n3453;
  assign n3455 = ~n3441 & ~n3454;
  assign n3456 = pi823 & n1756;
  assign n3457 = pi220 & ~n1756;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = n1754 & ~n3458;
  assign n3460 = ~n1778 & ~n3458;
  assign n3461 = pi220 & n1778;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = ~n1761 & ~n3462;
  assign n3464 = pi823 & n1761;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = ~n1754 & ~n3465;
  assign n3467 = ~n3459 & ~n3466;
  assign n3468 = n2412 & ~n3467;
  assign n3469 = n3455 & ~n3468;
  assign n3470 = ~n2228 & n2397;
  assign n3471 = n3469 & ~n3470;
  assign n3472 = ~n2027 & ~n3471;
  assign n3473 = pi609 & n2449;
  assign n3474 = pi380 & ~n2449;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = n2462 & ~n3475;
  assign n3477 = pi628 & n2449;
  assign n3478 = pi351 & ~n2449;
  assign n3479 = ~n3477 & ~n3478;
  assign n3480 = n2549 & ~n3479;
  assign n3481 = ~n3476 & ~n3480;
  assign n3482 = pi301 & ~n2449;
  assign n3483 = pi645 & n2449;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = n2541 & ~n3484;
  assign n3486 = pi543 & n2449;
  assign n3487 = pi263 & ~n2449;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = n2536 & ~n3488;
  assign n3490 = ~n3485 & ~n3489;
  assign n3491 = pi613 & n2449;
  assign n3492 = pi402 & ~n2449;
  assign n3493 = ~n3491 & ~n3492;
  assign n3494 = n2500 & ~n3493;
  assign n3495 = pi590 & n2449;
  assign n3496 = pi318 & ~n2449;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = n2488 & ~n3497;
  assign n3499 = ~n3494 & ~n3498;
  assign n3500 = pi531 & n2449;
  assign n3501 = pi358 & ~n2449;
  assign n3502 = ~n3500 & ~n3501;
  assign n3503 = n2482 & ~n3502;
  assign n3504 = pi544 & n2449;
  assign n3505 = pi297 & ~n2449;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = n2517 & ~n3506;
  assign n3508 = ~n3503 & ~n3507;
  assign n3509 = pi615 & n2449;
  assign n3510 = pi277 & ~n2449;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = n2506 & ~n3511;
  assign n3513 = pi585 & n2449;
  assign n3514 = pi359 & ~n2449;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = n2495 & ~n3515;
  assign n3517 = ~n3512 & ~n3516;
  assign n3518 = pi592 & n2449;
  assign n3519 = pi259 & ~n2449;
  assign n3520 = ~n3518 & ~n3519;
  assign n3521 = n2511 & ~n3520;
  assign n3522 = pi575 & n2449;
  assign n3523 = pi325 & ~n2449;
  assign n3524 = ~n3522 & ~n3523;
  assign n3525 = n2522 & ~n3524;
  assign n3526 = ~n3521 & ~n3525;
  assign n3527 = n3517 & n3526;
  assign n3528 = n3508 & n3527;
  assign n3529 = n3499 & n3528;
  assign n3530 = pi530 & n2449;
  assign n3531 = pi283 & ~n2449;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = n2531 & ~n3532;
  assign n3534 = pi612 & n2449;
  assign n3535 = pi328 & ~n2449;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = n2475 & ~n3536;
  assign n3538 = ~n3533 & ~n3537;
  assign n3539 = n3529 & n3538;
  assign n3540 = pi393 & ~n2449;
  assign n3541 = pi655 & n2449;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = n2466 & ~n3542;
  assign n3544 = pi578 & n2449;
  assign n3545 = pi369 & ~n2449;
  assign n3546 = ~n3544 & ~n3545;
  assign n3547 = n2455 & ~n3546;
  assign n3548 = ~n3543 & ~n3547;
  assign n3549 = n3539 & n3548;
  assign n3550 = n3490 & n3549;
  assign n3551 = n3481 & n3550;
  assign n3552 = n2559 & ~n3551;
  assign n3553 = n2558 & ~n3511;
  assign n3554 = n2572 & n3553;
  assign n3555 = ~n3552 & ~n3554;
  assign n3556 = n2027 & ~n3555;
  assign n3557 = ~n3472 & ~n3556;
  assign n3558 = ~n2028 & ~n3557;
  assign n3559 = ~n3428 & ~n3558;
  assign n3560 = ~n2986 & n3559;
  assign n3561 = n2986 & ~n3559;
  assign po344 = n3560 | n3561;
  assign n3563 = ~n3421 & po344;
  assign n3564 = ~n2028 & ~n3256;
  assign n3565 = ~n3127 & n3557;
  assign n3566 = n3127 & ~n3557;
  assign n3567 = ~n3565 & ~n3566;
  assign n3568 = n3413 & n3567;
  assign n3569 = ~n3413 & ~n3567;
  assign n3570 = ~n3568 & ~n3569;
  assign n3571 = n2028 & n3570;
  assign n3572 = ~n3564 & ~n3571;
  assign n3573 = ~n3415 & ~n3572;
  assign n3574 = n3415 & ~n3564;
  assign n3575 = ~n3571 & n3574;
  assign n3576 = ~n3573 & ~n3575;
  assign n3577 = po344 & n3576;
  assign n3578 = n3415 & n3572;
  assign n3579 = ~n3573 & ~n3578;
  assign n3580 = ~po344 & ~n3579;
  assign po311 = ~n3577 & ~n3580;
  assign n3582 = ~n2717 & n3259;
  assign n3583 = n2717 & ~n3259;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585 = n2028 & ~n3584;
  assign n3586 = ~n2028 & ~n2846;
  assign n3587 = ~n3585 & ~n3586;
  assign n3588 = ~n3415 & n3587;
  assign n3589 = n3415 & ~n3587;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = ~n3268 & n3590;
  assign n3592 = n3268 & ~n3590;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = po311 & ~n3593;
  assign n3595 = ~n3563 & n3594;
  assign n3596 = n3563 & ~n3594;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = ~n2028 & ~n2576;
  assign n3599 = n2028 & n3256;
  assign n3600 = ~n3567 & n3599;
  assign n3601 = ~n3256 & n3567;
  assign n3602 = n2028 & n3601;
  assign n3603 = ~n3600 & ~n3602;
  assign n3604 = ~n3598 & n3603;
  assign n3605 = n3587 & ~n3604;
  assign n3606 = ~n3587 & n3604;
  assign n3607 = ~n3605 & ~n3606;
  assign n3608 = ~n3559 & n3607;
  assign n3609 = n3559 & ~n3607;
  assign po327 = n3608 | n3609;
  assign n3611 = n3418 & po327;
  assign n3612 = ~n3424 & ~n3557;
  assign n3613 = n3424 & n3557;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = n2028 & n3614;
  assign n3616 = ~n2028 & n3127;
  assign n3617 = ~n3615 & ~n3616;
  assign n3618 = n3607 & n3617;
  assign n3619 = ~n3607 & ~n3617;
  assign n3620 = ~n3618 & ~n3619;
  assign n3621 = ~n3559 & n3620;
  assign n3622 = n3559 & ~n3620;
  assign n3623 = ~n3621 & ~n3622;
  assign n3624 = ~n3590 & n3623;
  assign n3625 = n3590 & ~n3623;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = n3268 & ~n3607;
  assign n3628 = ~n3268 & n3607;
  assign po339 = n3627 | n3628;
  assign n3630 = ~n3626 & po339;
  assign n3631 = ~n3611 & n3630;
  assign n3632 = n3611 & ~n3630;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = ~po311 & po327;
  assign n3635 = po311 & ~po327;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = po311 & n3636;
  assign n3638 = ~po311 & ~n3636;
  assign n3639 = ~n3637 & ~n3638;
  assign n3640 = n3268 & ~n3639;
  assign n3641 = ~po311 & n3636;
  assign n3642 = po311 & ~n3636;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = ~n3268 & ~n3643;
  assign n3645 = ~n3640 & ~n3644;
  assign n3646 = ~n3633 & n3645;
  assign n3647 = n3633 & ~n3645;
  assign n3648 = ~n3646 & ~n3647;
  assign n3649 = ~n3597 & n3648;
  assign n3650 = n3597 & ~n3648;
  assign po137 = n3649 | n3650;
  assign n3652 = ~n3268 & po339;
  assign n3653 = n3418 & po311;
  assign n3654 = n3652 & ~n3653;
  assign n3655 = ~n3652 & n3653;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~n3590 & ~po327;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = n3656 & n3657;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = po344 & ~n3626;
  assign n3662 = ~po344 & ~po339;
  assign n3663 = po344 & po339;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = po344 & ~n3664;
  assign n3666 = ~po344 & po339;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = ~n3639 & n3667;
  assign n3669 = ~n3643 & ~n3667;
  assign n3670 = ~n3668 & ~n3669;
  assign n3671 = n3661 & n3670;
  assign n3672 = ~n3661 & ~n3670;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = ~n3660 & n3673;
  assign n3675 = n3660 & ~n3673;
  assign po138 = n3674 | n3675;
  assign n3677 = ~n3268 & po327;
  assign n3678 = n3418 & po339;
  assign n3679 = ~n3677 & n3678;
  assign n3680 = n3677 & ~n3678;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = po344 & ~n3593;
  assign n3683 = po311 & ~n3626;
  assign n3684 = ~n3682 & n3683;
  assign n3685 = n3682 & ~n3683;
  assign n3686 = ~n3684 & ~n3685;
  assign n3687 = ~n3681 & n3686;
  assign n3688 = n3681 & ~n3686;
  assign n3689 = ~n3687 & ~n3688;
  assign n3690 = n3418 & n3590;
  assign n3691 = ~n3418 & ~n3590;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = ~n3639 & ~n3664;
  assign n3694 = ~n3643 & n3664;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = ~n3692 & n3695;
  assign n3697 = n3692 & ~n3695;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = ~n3689 & n3698;
  assign n3700 = n3689 & ~n3698;
  assign po139 = n3699 | n3700;
  assign n3702 = po327 & ~n3623;
  assign n3703 = ~n3590 & po339;
  assign n3704 = ~n3702 & n3703;
  assign n3705 = n3702 & ~n3703;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = n3418 & po344;
  assign n3708 = ~n3268 & po311;
  assign n3709 = ~n3707 & n3708;
  assign n3710 = n3707 & ~n3708;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = n3706 & ~n3711;
  assign n3713 = ~n3706 & n3711;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = ~n3268 & n3623;
  assign n3716 = n3268 & ~n3623;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = po311 & n3667;
  assign n3719 = ~po311 & ~n3667;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = n3717 & n3720;
  assign n3722 = ~n3717 & ~n3720;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3714 & ~n3723;
  assign n3725 = n3714 & n3723;
  assign po140 = n3724 | n3725;
  assign n3727 = pi874 & n1761;
  assign n3728 = pi056 & n1787;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~n1754 & ~n3729;
  assign n3731 = pi056 & ~n1756;
  assign n3732 = pi874 & n1756;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n1792 & ~n3733;
  assign n3735 = ~n3730 & ~n3734;
  assign n3736 = n1983 & n2028;
  assign n3737 = ~n2008 & ~n2256;
  assign n3738 = n2008 & n2256;
  assign n3739 = ~n3737 & ~n3738;
  assign n3740 = ~n2028 & n3739;
  assign n3741 = ~n1983 & n2186;
  assign n3742 = n1983 & ~n2186;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = n3740 & ~n3743;
  assign n3745 = ~n2028 & n2330;
  assign n3746 = n3743 & n3745;
  assign n3747 = ~n3744 & ~n3746;
  assign n3748 = ~n3736 & n3747;
  assign n3749 = pi906 & n1761;
  assign n3750 = pi906 & n1756;
  assign n3751 = ~pi136 & ~n1756;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n1778 & ~n3752;
  assign n3754 = ~pi136 & n1778;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n1761 & ~n3755;
  assign n3757 = ~n3749 & ~n3756;
  assign n3758 = ~n1754 & ~n3757;
  assign n3759 = n1754 & ~n3752;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = ~n3748 & n3760;
  assign n3762 = n3748 & ~n3760;
  assign n3763 = ~n3761 & ~n3762;
  assign n3764 = n3735 & n3763;
  assign n3765 = ~n3735 & ~n3763;
  assign po201 = ~n3764 & ~n3765;
  assign n3767 = pi842 & n1761;
  assign n3768 = pi842 & n1756;
  assign n3769 = pi017 & ~n1756;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = ~n1778 & ~n3770;
  assign n3772 = pi017 & n1778;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~n1761 & ~n3773;
  assign n3775 = ~n3767 & ~n3774;
  assign n3776 = ~n1754 & ~n3775;
  assign n3777 = n1754 & ~n3770;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = ~po201 & ~n3778;
  assign n3780 = po201 & n3778;
  assign po155 = n3779 | n3780;
  assign n3782 = ~n3025 & po155;
  assign n3783 = n3025 & ~n3779;
  assign n3784 = ~n3780 & n3783;
  assign n3785 = ~n3782 & ~n3784;
  assign n3786 = po814 & n3785;
  assign n3787 = pi009 & ~po814;
  assign po141 = n3786 | n3787;
  assign n3789 = pi844 & n1761;
  assign n3790 = pi042 & n1787;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~n1754 & ~n3791;
  assign n3793 = pi844 & n1756;
  assign n3794 = pi042 & ~n1756;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = ~n1792 & ~n3795;
  assign n3797 = ~n3792 & ~n3796;
  assign n3798 = pi908 & n1761;
  assign n3799 = pi908 & n1756;
  assign n3800 = ~pi188 & ~n1756;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~n1778 & ~n3801;
  assign n3803 = ~pi188 & n1778;
  assign n3804 = ~n3802 & ~n3803;
  assign n3805 = ~n1761 & ~n3804;
  assign n3806 = ~n3798 & ~n3805;
  assign n3807 = ~n1754 & ~n3806;
  assign n3808 = n1754 & ~n3801;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = n1942 & ~n1989;
  assign n3811 = ~n1942 & ~n2012;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~n3739 & n3812;
  assign n3814 = ~n2028 & ~n3813;
  assign n3815 = ~n2330 & ~n3812;
  assign n3816 = n3814 & ~n3815;
  assign n3817 = n1942 & n2028;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = n3809 & n3818;
  assign n3820 = pi876 & n1756;
  assign n3821 = ~pi046 & ~n1756;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = ~n1778 & ~n3822;
  assign n3824 = ~pi046 & n1778;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = ~n1761 & ~n3825;
  assign n3827 = pi876 & n1761;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = ~n1754 & ~n3828;
  assign n3830 = n1754 & ~n3822;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = ~n3819 & ~n3831;
  assign n3833 = ~n3809 & ~n3818;
  assign n3834 = n3832 & ~n3833;
  assign n3835 = ~n3797 & ~n3834;
  assign n3836 = ~n3819 & ~n3833;
  assign n3837 = n3831 & ~n3836;
  assign n3838 = n3835 & ~n3837;
  assign n3839 = ~n3831 & n3836;
  assign n3840 = ~n3837 & ~n3839;
  assign n3841 = n3797 & ~n3840;
  assign po181 = n3838 | n3841;
  assign n3843 = n3407 & po181;
  assign n3844 = ~n3407 & ~po181;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = po814 & ~n3845;
  assign n3847 = pi010 & ~po814;
  assign po142 = n3846 | n3847;
  assign n3849 = pi843 & n1761;
  assign n3850 = pi843 & n1756;
  assign n3851 = pi043 & ~n1756;
  assign n3852 = ~n3850 & ~n3851;
  assign n3853 = ~n1778 & ~n3852;
  assign n3854 = pi043 & n1778;
  assign n3855 = ~n3853 & ~n3854;
  assign n3856 = ~n1761 & ~n3855;
  assign n3857 = ~n3849 & ~n3856;
  assign n3858 = ~n1754 & ~n3857;
  assign n3859 = n1754 & ~n3852;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = n2005 & ~n2012;
  assign n3862 = ~n1989 & ~n2005;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n3739 & n3863;
  assign n3865 = ~n2330 & ~n3863;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = ~n2028 & ~n3866;
  assign n3868 = ~n1986 & n2028;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = pi907 & n1761;
  assign n3871 = pi907 & n1756;
  assign n3872 = ~pi176 & ~n1756;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n1778 & ~n3873;
  assign n3875 = ~pi176 & n1778;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = ~n1761 & ~n3876;
  assign n3878 = ~n3870 & ~n3877;
  assign n3879 = ~n1754 & ~n3878;
  assign n3880 = n1754 & ~n3873;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = n3869 & ~n3881;
  assign n3883 = ~n3869 & n3881;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = ~pi047 & n1787;
  assign n3886 = pi875 & n1761;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = ~n1754 & ~n3887;
  assign n3889 = pi875 & n1756;
  assign n3890 = ~pi047 & ~n1756;
  assign n3891 = ~n3889 & ~n3890;
  assign n3892 = ~n1792 & ~n3891;
  assign n3893 = ~n3888 & ~n3892;
  assign n3894 = n3884 & ~n3893;
  assign n3895 = ~n3884 & n3893;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3860 & n3896;
  assign n3898 = n3860 & ~n3896;
  assign po183 = n3897 | n3898;
  assign n3900 = n2672 & ~po183;
  assign n3901 = ~n2672 & po183;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = po814 & n3902;
  assign n3904 = pi011 & ~po814;
  assign po143 = n3903 | n3904;
  assign n3906 = pi565 & ~n2540;
  assign n3907 = ~n2555 & ~n3906;
  assign n3908 = ~pi568 & n2506;
  assign n3909 = pi563 & ~n3908;
  assign n3910 = n3907 & n3909;
  assign n3911 = pi568 & ~n2506;
  assign n3912 = ~n3908 & ~n3911;
  assign n3913 = pi566 & ~n2487;
  assign n3914 = ~n2540 & ~n3913;
  assign n3915 = n3912 & n3914;
  assign n3916 = ~n3908 & n3915;
  assign n3917 = ~n2460 & ~n2487;
  assign n3918 = n3916 & ~n3917;
  assign n3919 = n3910 & n3918;
  assign n3920 = pi018 & ~n3919;
  assign n3921 = ~n2194 & n3919;
  assign n3922 = ~n3920 & ~n3921;
  assign n3923 = n2559 & ~n3922;
  assign n3924 = pi022 & n2556;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = pi018 & n2558;
  assign po157 = ~n3925 | n3926;
  assign n3928 = pi019 & ~n3919;
  assign n3929 = ~n2265 & n3919;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n2559 & ~n3930;
  assign n3932 = pi023 & n2556;
  assign n3933 = ~n3931 & ~n3932;
  assign n3934 = pi019 & n2558;
  assign po158 = ~n3933 | n3934;
  assign n3936 = ~n3908 & ~n3914;
  assign n3937 = n3912 & n3936;
  assign n3938 = ~n3917 & n3937;
  assign n3939 = ~n3907 & n3909;
  assign n3940 = n3938 & n3939;
  assign n3941 = pi020 & ~n3940;
  assign n3942 = ~n2194 & n3940;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = n2559 & ~n3943;
  assign n3945 = pi024 & n2556;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = pi020 & n2558;
  assign po159 = ~n3946 | n3947;
  assign n3949 = pi021 & ~n3940;
  assign n3950 = ~n2265 & n3940;
  assign n3951 = ~n3949 & ~n3950;
  assign n3952 = n2559 & ~n3951;
  assign n3953 = pi025 & n2556;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = pi021 & n2558;
  assign po160 = ~n3954 | n3955;
  assign n3957 = n3918 & n3939;
  assign n3958 = pi022 & ~n3957;
  assign n3959 = ~n2194 & n3957;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = n2559 & ~n3960;
  assign n3962 = pi018 & n2556;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = pi022 & n2558;
  assign po161 = ~n3963 | n3964;
  assign n3966 = pi023 & ~n3957;
  assign n3967 = ~n2265 & n3957;
  assign n3968 = ~n3966 & ~n3967;
  assign n3969 = n2559 & ~n3968;
  assign n3970 = pi019 & n2556;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = pi023 & n2558;
  assign po162 = ~n3971 | n3972;
  assign n3974 = n3910 & n3938;
  assign n3975 = pi024 & ~n3974;
  assign n3976 = ~n2194 & n3974;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = n2559 & ~n3977;
  assign n3979 = pi020 & n2556;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = pi024 & n2558;
  assign po163 = ~n3980 | n3981;
  assign n3983 = pi025 & ~n3974;
  assign n3984 = ~n2265 & n3974;
  assign n3985 = ~n3983 & ~n3984;
  assign n3986 = n2559 & ~n3985;
  assign n3987 = pi021 & n2556;
  assign n3988 = ~n3986 & ~n3987;
  assign n3989 = pi025 & n2558;
  assign po164 = ~n3988 | n3989;
  assign n3991 = ~pi673 & ~n2265;
  assign n3992 = pi038 & pi673;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = n2556 & ~n3993;
  assign n3995 = pi026 & n2558;
  assign n3996 = ~pi563 & ~n3908;
  assign n3997 = n3907 & n3996;
  assign n3998 = n3918 & n3997;
  assign n3999 = pi026 & ~n3998;
  assign n4000 = ~n2265 & n3998;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n2559 & ~n4001;
  assign n4003 = ~n3995 & ~n4002;
  assign po165 = n3994 | ~n4003;
  assign n4005 = ~pi673 & ~n2194;
  assign n4006 = pi039 & pi673;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = n2556 & ~n4007;
  assign n4009 = pi027 & n2558;
  assign n4010 = pi027 & ~n3998;
  assign n4011 = ~n2194 & n3998;
  assign n4012 = ~n4010 & ~n4011;
  assign n4013 = n2559 & ~n4012;
  assign n4014 = ~n4009 & ~n4013;
  assign po166 = n4008 | ~n4014;
  assign n4016 = pi031 & pi673;
  assign n4017 = pi041 & ~pi673;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = n2556 & ~n4018;
  assign n4020 = pi028 & n2558;
  assign n4021 = n3916 & n3917;
  assign n4022 = n3997 & n4021;
  assign n4023 = pi028 & ~n4022;
  assign n4024 = ~n2265 & n4022;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = n2559 & ~n4025;
  assign n4027 = ~n4020 & ~n4026;
  assign po167 = n4019 | ~n4027;
  assign n4029 = pi030 & pi673;
  assign n4030 = pi040 & ~pi673;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = n2556 & ~n4031;
  assign n4033 = pi029 & n2558;
  assign n4034 = pi029 & ~n4022;
  assign n4035 = ~n2194 & n4022;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = n2559 & ~n4036;
  assign n4038 = ~n4033 & ~n4037;
  assign po168 = n4032 | ~n4038;
  assign n4040 = pi034 & pi673;
  assign n4041 = pi029 & ~pi673;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = n2556 & ~n4042;
  assign n4044 = pi030 & n2558;
  assign n4045 = ~n3907 & n3996;
  assign n4046 = n3917 & n3937;
  assign n4047 = n4045 & n4046;
  assign n4048 = pi030 & ~n4047;
  assign n4049 = ~n2194 & n4047;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = n2559 & ~n4050;
  assign n4052 = ~n4044 & ~n4051;
  assign po169 = n4043 | ~n4052;
  assign n4054 = pi035 & pi673;
  assign n4055 = pi028 & ~pi673;
  assign n4056 = ~n4054 & ~n4055;
  assign n4057 = n2556 & ~n4056;
  assign n4058 = pi031 & n2558;
  assign n4059 = pi031 & ~n4047;
  assign n4060 = ~n2265 & n4047;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = n2559 & ~n4061;
  assign n4063 = ~n4058 & ~n4062;
  assign po170 = n4057 | ~n4063;
  assign n4065 = pi039 & ~pi673;
  assign n4066 = pi673 & ~n2194;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = n2556 & ~n4067;
  assign n4069 = pi032 & n2558;
  assign n4070 = n3918 & n4045;
  assign n4071 = pi032 & ~n4070;
  assign n4072 = ~n2194 & n4070;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = n2559 & ~n4073;
  assign n4075 = ~n4069 & ~n4074;
  assign po171 = n4068 | ~n4075;
  assign n4077 = pi038 & ~pi673;
  assign n4078 = pi673 & ~n2265;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = n2556 & ~n4079;
  assign n4081 = pi033 & n2558;
  assign n4082 = pi033 & ~n4070;
  assign n4083 = ~n2265 & n4070;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = n2559 & ~n4084;
  assign n4086 = ~n4081 & ~n4085;
  assign po172 = n4080 | ~n4086;
  assign n4088 = pi030 & ~pi673;
  assign n4089 = pi040 & pi673;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = n2556 & ~n4090;
  assign n4092 = pi034 & n2558;
  assign n4093 = n4021 & n4045;
  assign n4094 = pi034 & ~n4093;
  assign n4095 = ~n2194 & n4093;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = n2559 & ~n4096;
  assign n4098 = ~n4092 & ~n4097;
  assign po173 = n4091 | ~n4098;
  assign n4100 = pi031 & ~pi673;
  assign n4101 = pi041 & pi673;
  assign n4102 = ~n4100 & ~n4101;
  assign n4103 = n2556 & ~n4102;
  assign n4104 = pi035 & n2558;
  assign n4105 = pi035 & ~n4093;
  assign n4106 = ~n2265 & n4093;
  assign n4107 = ~n4105 & ~n4106;
  assign n4108 = n2559 & ~n4107;
  assign n4109 = ~n4104 & ~n4108;
  assign po174 = n4103 | ~n4109;
  assign n4111 = pi027 & pi673;
  assign n4112 = pi032 & ~pi673;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = n2556 & ~n4113;
  assign n4115 = pi036 & n2558;
  assign n4116 = n3938 & n4045;
  assign n4117 = pi036 & ~n4116;
  assign n4118 = ~n2194 & n4116;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = n2559 & ~n4119;
  assign n4121 = ~n4115 & ~n4120;
  assign po175 = n4114 | ~n4121;
  assign n4123 = pi026 & pi673;
  assign n4124 = pi033 & ~pi673;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = n2556 & ~n4125;
  assign n4127 = pi037 & n2558;
  assign n4128 = pi037 & ~n4116;
  assign n4129 = ~n2265 & n4116;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = n2559 & ~n4130;
  assign n4132 = ~n4127 & ~n4131;
  assign po176 = n4126 | ~n4132;
  assign n4134 = pi026 & ~pi673;
  assign n4135 = pi033 & pi673;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = n2556 & ~n4136;
  assign n4138 = pi038 & n2558;
  assign n4139 = n3938 & n3997;
  assign n4140 = pi038 & ~n4139;
  assign n4141 = ~n2265 & n4139;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = n2559 & ~n4142;
  assign n4144 = ~n4138 & ~n4143;
  assign po177 = n4137 | ~n4144;
  assign n4146 = pi027 & ~pi673;
  assign n4147 = pi032 & pi673;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = n2556 & ~n4148;
  assign n4150 = pi039 & n2558;
  assign n4151 = pi039 & ~n4139;
  assign n4152 = ~n2194 & n4139;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = n2559 & ~n4153;
  assign n4155 = ~n4150 & ~n4154;
  assign po178 = n4149 | ~n4155;
  assign n4157 = pi034 & ~pi673;
  assign n4158 = pi029 & pi673;
  assign n4159 = ~n4157 & ~n4158;
  assign n4160 = n2556 & ~n4159;
  assign n4161 = pi040 & n2558;
  assign n4162 = n3997 & n4046;
  assign n4163 = pi040 & ~n4162;
  assign n4164 = ~n2194 & n4162;
  assign n4165 = ~n4163 & ~n4164;
  assign n4166 = n2559 & ~n4165;
  assign n4167 = ~n4161 & ~n4166;
  assign po179 = n4160 | ~n4167;
  assign n4169 = pi035 & ~pi673;
  assign n4170 = pi028 & pi673;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = n2556 & ~n4171;
  assign n4173 = pi041 & n2558;
  assign n4174 = pi041 & ~n4162;
  assign n4175 = ~n2265 & n4162;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n2559 & ~n4176;
  assign n4178 = ~n4173 & ~n4177;
  assign po180 = n4172 | ~n4178;
  assign n4180 = ~pi046 & ~po814;
  assign n4181 = n3831 & n3836;
  assign n4182 = ~n3831 & ~n3836;
  assign n4183 = ~n4181 & ~n4182;
  assign n4184 = po814 & n4183;
  assign po189 = n4180 | n4184;
  assign n4186 = ~pi047 & ~po814;
  assign n4187 = po814 & ~n3896;
  assign po190 = n4186 | n4187;
  assign n4189 = pi050 & ~n2559;
  assign n4190 = n3910 & n4021;
  assign n4191 = ~n2194 & n4190;
  assign n4192 = pi050 & ~n4190;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = n2559 & ~n4193;
  assign po195 = n4189 | n4194;
  assign n4196 = pi051 & ~n2559;
  assign n4197 = ~n2265 & n4190;
  assign n4198 = pi051 & ~n4190;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = n2559 & ~n4199;
  assign po196 = n4196 | n4200;
  assign n4202 = pi052 & ~n2559;
  assign n4203 = n3939 & n4046;
  assign n4204 = ~n2194 & n4203;
  assign n4205 = pi052 & ~n4203;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = n2559 & ~n4206;
  assign po197 = n4202 | n4207;
  assign n4209 = pi053 & ~n2559;
  assign n4210 = n3910 & n4046;
  assign n4211 = ~n2265 & n4210;
  assign n4212 = pi053 & ~n4210;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = n2559 & ~n4213;
  assign po198 = n4209 | n4214;
  assign n4216 = pi054 & ~n2559;
  assign n4217 = ~n2265 & n4203;
  assign n4218 = pi054 & ~n4203;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = n2559 & ~n4219;
  assign po199 = n4216 | n4220;
  assign n4222 = pi055 & ~n2559;
  assign n4223 = ~n2194 & n4210;
  assign n4224 = pi055 & ~n4210;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = n2559 & ~n4225;
  assign po200 = n4222 | n4226;
  assign n4228 = ~n3748 & n3919;
  assign n4229 = pi058 & ~n3919;
  assign n4230 = ~n4228 & ~n4229;
  assign n4231 = n2559 & ~n4230;
  assign n4232 = pi059 & n2556;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = pi058 & n2558;
  assign po205 = ~n4233 | n4234;
  assign n4236 = ~n3748 & n3957;
  assign n4237 = pi059 & ~n3957;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = n2559 & ~n4238;
  assign n4240 = pi058 & n2556;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = pi059 & n2558;
  assign po206 = ~n4241 | n4242;
  assign n4244 = ~n3748 & n3974;
  assign n4245 = pi060 & ~n3974;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = n2559 & ~n4246;
  assign n4248 = pi061 & n2556;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = pi060 & n2558;
  assign po207 = ~n4249 | n4250;
  assign n4252 = ~n3748 & n3940;
  assign n4253 = pi061 & ~n3940;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = n2559 & ~n4254;
  assign n4256 = pi060 & n2556;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = pi061 & n2558;
  assign po208 = ~n4257 | n4258;
  assign n4260 = ~pi062 & ~n4116;
  assign n4261 = ~n3748 & n4116;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = n2559 & ~n4262;
  assign n4264 = ~pi062 & n2558;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = pi092 & ~pi673;
  assign n4267 = pi067 & pi673;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n2556 & ~n4268;
  assign po209 = ~n4265 | n4269;
  assign n4271 = ~n3748 & n4022;
  assign n4272 = pi063 & ~n4022;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = n2559 & ~n4273;
  assign n4275 = pi063 & n2558;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = pi064 & pi673;
  assign n4278 = pi066 & ~pi673;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = n2556 & ~n4279;
  assign po210 = ~n4276 | n4280;
  assign n4282 = pi064 & ~n4047;
  assign n4283 = ~n3748 & n4047;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = n2559 & ~n4284;
  assign n4286 = pi064 & n2558;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = pi068 & pi673;
  assign n4289 = pi063 & ~pi673;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n2556 & ~n4290;
  assign po211 = ~n4287 | n4291;
  assign n4293 = ~n3748 & n4139;
  assign n4294 = pi065 & ~n4139;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = n2559 & ~n4295;
  assign n4297 = pi065 & n2558;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = pi092 & pi673;
  assign n4300 = pi067 & ~pi673;
  assign n4301 = ~n4299 & ~n4300;
  assign n4302 = n2556 & ~n4301;
  assign po212 = ~n4298 | n4302;
  assign n4304 = ~n3748 & n4162;
  assign n4305 = pi066 & ~n4162;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = n2559 & ~n4306;
  assign n4308 = pi066 & n2558;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = pi068 & ~pi673;
  assign n4311 = pi063 & pi673;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = n2556 & ~n4312;
  assign po213 = ~n4309 | n4313;
  assign n4315 = ~n3748 & n3998;
  assign n4316 = pi067 & ~n3998;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = n2559 & ~n4317;
  assign n4319 = pi067 & n2558;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = ~pi673 & ~n3748;
  assign n4322 = pi065 & pi673;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = n2556 & ~n4323;
  assign po214 = ~n4320 | n4324;
  assign n4326 = pi068 & ~n4093;
  assign n4327 = ~n3748 & n4093;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = n2559 & ~n4328;
  assign n4330 = pi068 & n2558;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = pi064 & ~pi673;
  assign n4333 = pi066 & pi673;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = n2556 & ~n4334;
  assign po215 = ~n4331 | n4335;
  assign n4337 = pi069 & ~n2559;
  assign n4338 = n3939 & n4021;
  assign n4339 = ~n2194 & n4338;
  assign n4340 = pi069 & ~n4338;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = n2559 & ~n4341;
  assign po216 = n4337 | n4342;
  assign n4344 = pi070 & ~n2559;
  assign n4345 = ~n2265 & n4338;
  assign n4346 = pi070 & ~n4338;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = n2559 & ~n4347;
  assign po217 = n4344 | n4348;
  assign n4350 = ~n2194 & n2440;
  assign n4351 = ~po814 & ~n2440;
  assign n4352 = ~n2397 & n4351;
  assign n4353 = ~n2412 & n4352;
  assign n4354 = ~n2412 & ~n4353;
  assign n4355 = ~pi071 & ~n4354;
  assign n4356 = ~n4350 & ~n4355;
  assign n4357 = ~po814 & ~n2397;
  assign n4358 = ~pi071 & ~n4357;
  assign po218 = ~n4356 | n4358;
  assign n4360 = ~n2265 & n2440;
  assign n4361 = ~pi072 & ~n4354;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = ~pi072 & ~n4357;
  assign po219 = ~n4362 | n4363;
  assign n4365 = ~n2031 & n3919;
  assign n4366 = pi073 & ~n3919;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = n2559 & ~n4367;
  assign n4369 = pi080 & n2556;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = pi073 & n2558;
  assign po220 = ~n4370 | n4371;
  assign n4373 = ~n2119 & n3919;
  assign n4374 = pi074 & ~n3919;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = n2559 & ~n4375;
  assign n4377 = pi079 & n2556;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = pi074 & n2558;
  assign po221 = ~n4378 | n4379;
  assign n4381 = ~n2344 & n3919;
  assign n4382 = pi075 & ~n3919;
  assign n4383 = ~n4381 & ~n4382;
  assign n4384 = n2559 & ~n4383;
  assign n4385 = pi081 & n2556;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = pi075 & n2558;
  assign po222 = ~n4386 | n4387;
  assign n4389 = ~n2031 & n3940;
  assign n4390 = pi076 & ~n3940;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = n2559 & ~n4391;
  assign n4393 = pi082 & n2556;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = pi076 & n2558;
  assign po223 = ~n4394 | n4395;
  assign n4397 = ~n2119 & n3940;
  assign n4398 = pi077 & ~n3940;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = n2559 & ~n4399;
  assign n4401 = pi083 & n2556;
  assign n4402 = ~n4400 & ~n4401;
  assign n4403 = pi077 & n2558;
  assign po224 = ~n4402 | n4403;
  assign n4405 = ~n2344 & n3940;
  assign n4406 = pi078 & ~n3940;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = n2559 & ~n4407;
  assign n4409 = pi084 & n2556;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = pi078 & n2558;
  assign po225 = ~n4410 | n4411;
  assign n4413 = ~n2119 & n3957;
  assign n4414 = pi079 & ~n3957;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = n2559 & ~n4415;
  assign n4417 = pi074 & n2556;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = pi079 & n2558;
  assign po226 = ~n4418 | n4419;
  assign n4421 = ~n2031 & n3957;
  assign n4422 = pi080 & ~n3957;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = n2559 & ~n4423;
  assign n4425 = pi073 & n2556;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = pi080 & n2558;
  assign po227 = ~n4426 | n4427;
  assign n4429 = ~n2344 & n3957;
  assign n4430 = pi081 & ~n3957;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n2559 & ~n4431;
  assign n4433 = pi075 & n2556;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = pi081 & n2558;
  assign po228 = ~n4434 | n4435;
  assign n4437 = ~n2031 & n3974;
  assign n4438 = pi082 & ~n3974;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = n2559 & ~n4439;
  assign n4441 = pi076 & n2556;
  assign n4442 = ~n4440 & ~n4441;
  assign n4443 = pi082 & n2558;
  assign po229 = ~n4442 | n4443;
  assign n4445 = ~n2119 & n3974;
  assign n4446 = pi083 & ~n3974;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n2559 & ~n4447;
  assign n4449 = pi077 & n2556;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = pi083 & n2558;
  assign po230 = ~n4450 | n4451;
  assign n4453 = ~n2344 & n3974;
  assign n4454 = pi084 & ~n3974;
  assign n4455 = ~n4453 & ~n4454;
  assign n4456 = n2559 & ~n4455;
  assign n4457 = pi078 & n2556;
  assign n4458 = ~n4456 & ~n4457;
  assign n4459 = pi084 & n2558;
  assign po231 = ~n4458 | n4459;
  assign n4461 = ~n2344 & n3998;
  assign n4462 = pi085 & ~n3998;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = n2559 & ~n4463;
  assign n4465 = pi085 & n2558;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~pi673 & ~n2344;
  assign n4468 = pi102 & pi673;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = n2556 & ~n4469;
  assign po232 = ~n4466 | n4470;
  assign n4472 = ~n2031 & n4022;
  assign n4473 = pi086 & ~n4022;
  assign n4474 = ~n4472 & ~n4473;
  assign n4475 = n2559 & ~n4474;
  assign n4476 = pi086 & n2558;
  assign n4477 = ~n4475 & ~n4476;
  assign n4478 = pi090 & pi673;
  assign n4479 = pi104 & ~pi673;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481 = n2556 & ~n4480;
  assign po233 = ~n4477 | n4481;
  assign n4483 = ~n2119 & n4022;
  assign n4484 = pi087 & ~n4022;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = n2559 & ~n4485;
  assign n4487 = pi087 & n2558;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = pi089 & pi673;
  assign n4490 = pi103 & ~pi673;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = n2556 & ~n4491;
  assign po234 = ~n4488 | n4492;
  assign n4494 = ~n2344 & n4022;
  assign n4495 = pi088 & ~n4022;
  assign n4496 = ~n4494 & ~n4495;
  assign n4497 = n2559 & ~n4496;
  assign n4498 = pi088 & n2558;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = pi091 & pi673;
  assign n4501 = pi105 & ~pi673;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = n2556 & ~n4502;
  assign po235 = ~n4499 | n4503;
  assign n4505 = pi089 & ~n4047;
  assign n4506 = ~n2119 & n4047;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = n2559 & ~n4507;
  assign n4509 = pi089 & n2558;
  assign n4510 = ~n4508 & ~n4509;
  assign n4511 = pi095 & pi673;
  assign n4512 = pi087 & ~pi673;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = n2556 & ~n4513;
  assign po236 = ~n4510 | n4514;
  assign n4516 = pi090 & ~n4047;
  assign n4517 = ~n2031 & n4047;
  assign n4518 = ~n4516 & ~n4517;
  assign n4519 = n2559 & ~n4518;
  assign n4520 = pi090 & n2558;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = pi094 & pi673;
  assign n4523 = pi086 & ~pi673;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n2556 & ~n4524;
  assign po237 = ~n4521 | n4525;
  assign n4527 = pi091 & ~n4047;
  assign n4528 = ~n2344 & n4047;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = n2559 & ~n4529;
  assign n4531 = pi091 & n2558;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = pi096 & pi673;
  assign n4534 = pi088 & ~pi673;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = n2556 & ~n4535;
  assign po238 = ~n4532 | n4536;
  assign n4538 = pi065 & ~pi673;
  assign n4539 = pi673 & ~n3748;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = n2556 & ~n4540;
  assign n4542 = pi092 & n2558;
  assign n4543 = ~n4541 & ~n4542;
  assign n4544 = pi092 & ~n4070;
  assign n4545 = ~n3748 & n4070;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = n2559 & ~n4546;
  assign po239 = ~n4543 | n4547;
  assign n4549 = pi093 & ~n4116;
  assign n4550 = ~n2119 & n4116;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = n2559 & ~n4551;
  assign n4553 = pi093 & n2558;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = pi112 & pi673;
  assign n4556 = pi097 & ~pi673;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = n2556 & ~n4557;
  assign po240 = ~n4554 | n4558;
  assign n4560 = pi094 & ~n4093;
  assign n4561 = ~n2031 & n4093;
  assign n4562 = ~n4560 & ~n4561;
  assign n4563 = n2559 & ~n4562;
  assign n4564 = pi094 & n2558;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = pi090 & ~pi673;
  assign n4567 = pi104 & pi673;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = n2556 & ~n4568;
  assign po241 = ~n4565 | n4569;
  assign n4571 = pi095 & ~n4093;
  assign n4572 = ~n2119 & n4093;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = n2559 & ~n4573;
  assign n4575 = pi095 & n2558;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = pi089 & ~pi673;
  assign n4578 = pi103 & pi673;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = n2556 & ~n4579;
  assign po242 = ~n4576 | n4580;
  assign n4582 = pi096 & ~n4093;
  assign n4583 = ~n2344 & n4093;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = n2559 & ~n4584;
  assign n4586 = pi096 & n2558;
  assign n4587 = ~n4585 & ~n4586;
  assign n4588 = pi091 & ~pi673;
  assign n4589 = pi105 & pi673;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n2556 & ~n4590;
  assign po243 = ~n4587 | n4591;
  assign n4593 = pi097 & ~n4070;
  assign n4594 = ~n2119 & n4070;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = n2559 & ~n4595;
  assign n4597 = pi097 & n2558;
  assign n4598 = ~n4596 & ~n4597;
  assign n4599 = pi673 & ~n2119;
  assign n4600 = pi098 & ~pi673;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = n2556 & ~n4601;
  assign po244 = ~n4598 | n4602;
  assign n4604 = ~n2119 & n4139;
  assign n4605 = pi098 & ~n4139;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = n2559 & ~n4606;
  assign n4608 = pi098 & n2558;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = pi112 & ~pi673;
  assign n4611 = pi097 & pi673;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = n2556 & ~n4612;
  assign po245 = ~n4609 | n4613;
  assign n4615 = ~n2031 & n4139;
  assign n4616 = pi099 & ~n4139;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = n2559 & ~n4617;
  assign n4619 = pi099 & n2558;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = pi115 & pi673;
  assign n4622 = pi118 & ~pi673;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = n2556 & ~n4623;
  assign po246 = ~n4620 | n4624;
  assign n4626 = pi100 & ~n4116;
  assign n4627 = ~n2031 & n4116;
  assign n4628 = ~n4626 & ~n4627;
  assign n4629 = n2559 & ~n4628;
  assign n4630 = pi100 & n2558;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = pi115 & ~pi673;
  assign n4633 = pi118 & pi673;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = n2556 & ~n4634;
  assign po247 = ~n4631 | n4635;
  assign n4637 = pi101 & ~n4116;
  assign n4638 = ~n2344 & n4116;
  assign n4639 = ~n4637 & ~n4638;
  assign n4640 = n2559 & ~n4639;
  assign n4641 = pi101 & n2558;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = pi116 & ~pi673;
  assign n4644 = pi085 & pi673;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = n2556 & ~n4645;
  assign po248 = ~n4642 | n4646;
  assign n4648 = ~n2344 & n4139;
  assign n4649 = pi102 & ~n4139;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = n2559 & ~n4650;
  assign n4652 = pi102 & n2558;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = pi116 & pi673;
  assign n4655 = pi085 & ~pi673;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = n2556 & ~n4656;
  assign po249 = ~n4653 | n4657;
  assign n4659 = ~n2119 & n4162;
  assign n4660 = pi103 & ~n4162;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = n2559 & ~n4661;
  assign n4663 = pi103 & n2558;
  assign n4664 = ~n4662 & ~n4663;
  assign n4665 = pi095 & ~pi673;
  assign n4666 = pi087 & pi673;
  assign n4667 = ~n4665 & ~n4666;
  assign n4668 = n2556 & ~n4667;
  assign po250 = ~n4664 | n4668;
  assign n4670 = ~n2031 & n4162;
  assign n4671 = pi104 & ~n4162;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = n2559 & ~n4672;
  assign n4674 = pi104 & n2558;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = pi094 & ~pi673;
  assign n4677 = pi086 & pi673;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = n2556 & ~n4678;
  assign po251 = ~n4675 | n4679;
  assign n4681 = ~n2344 & n4162;
  assign n4682 = pi105 & ~n4162;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = n2559 & ~n4683;
  assign n4685 = pi105 & n2558;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = pi096 & ~pi673;
  assign n4688 = pi088 & pi673;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = n2556 & ~n4689;
  assign po252 = ~n4686 | n4690;
  assign n4692 = pi106 & ~n2559;
  assign n4693 = ~n3748 & n4190;
  assign n4694 = pi106 & ~n4190;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = n2559 & ~n4695;
  assign po253 = n4692 | n4696;
  assign n4698 = pi107 & ~n2559;
  assign n4699 = ~n3748 & n4203;
  assign n4700 = pi107 & ~n4203;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = n2559 & ~n4701;
  assign po254 = n4698 | n4702;
  assign n4704 = pi108 & ~n2559;
  assign n4705 = ~n3748 & n4338;
  assign n4706 = pi108 & ~n4338;
  assign n4707 = ~n4705 & ~n4706;
  assign n4708 = n2559 & ~n4707;
  assign po255 = n4704 | n4708;
  assign n4710 = pi109 & ~n2559;
  assign n4711 = ~n3748 & n4210;
  assign n4712 = pi109 & ~n4210;
  assign n4713 = ~n4711 & ~n4712;
  assign n4714 = n2559 & ~n4713;
  assign po256 = n4710 | n4714;
  assign n4716 = ~n3268 & ~po311;
  assign n4717 = n3268 & po311;
  assign po257 = n4716 | n4717;
  assign n4719 = ~pi111 & ~n4354;
  assign n4720 = ~n2265 & n2397;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = ~pi111 & ~n4351;
  assign po258 = ~n4721 | n4722;
  assign n4724 = ~pi673 & ~n2119;
  assign n4725 = pi098 & pi673;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = n2556 & ~n4726;
  assign n4728 = pi112 & n2558;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = ~n2119 & n3998;
  assign n4731 = pi112 & ~n3998;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733 = n2559 & ~n4732;
  assign po259 = ~n4729 | n4733;
  assign n4735 = ~n2440 & ~n4353;
  assign n4736 = ~pi113 & ~n4735;
  assign n4737 = ~n2265 & n2412;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = ~pi113 & ~n4357;
  assign po260 = ~n4738 | n4739;
  assign n4741 = ~pi114 & ~n4735;
  assign n4742 = ~n2194 & n2412;
  assign n4743 = ~n4741 & ~n4742;
  assign n4744 = ~pi114 & ~n4357;
  assign po261 = ~n4743 | n4744;
  assign n4746 = pi099 & ~pi673;
  assign n4747 = pi673 & ~n2031;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = n2556 & ~n4748;
  assign n4750 = pi115 & n2558;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n2031 & n4070;
  assign n4753 = pi115 & ~n4070;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = n2559 & ~n4754;
  assign po262 = ~n4751 | n4755;
  assign n4757 = pi102 & ~pi673;
  assign n4758 = pi673 & ~n2344;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = n2556 & ~n4759;
  assign n4761 = pi116 & n2558;
  assign n4762 = ~n4760 & ~n4761;
  assign n4763 = ~n2344 & n4070;
  assign n4764 = pi116 & ~n4070;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = n2559 & ~n4765;
  assign po263 = ~n4762 | n4766;
  assign n4768 = ~pi117 & ~n4354;
  assign n4769 = ~n2194 & n2397;
  assign n4770 = ~n4768 & ~n4769;
  assign n4771 = ~pi117 & ~n4351;
  assign po264 = ~n4770 | n4771;
  assign n4773 = ~pi673 & ~n2031;
  assign n4774 = pi099 & pi673;
  assign n4775 = ~n4773 & ~n4774;
  assign n4776 = n2556 & ~n4775;
  assign n4777 = pi118 & n2558;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = ~n2031 & n3998;
  assign n4780 = pi118 & ~n3998;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = n2559 & ~n4781;
  assign po265 = ~n4778 | n4782;
  assign n4784 = pi119 & ~n2559;
  assign n4785 = ~n2031 & n4190;
  assign n4786 = pi119 & ~n4190;
  assign n4787 = ~n4785 & ~n4786;
  assign n4788 = n2559 & ~n4787;
  assign po266 = n4784 | n4788;
  assign n4790 = pi120 & ~n2559;
  assign n4791 = ~n2119 & n4190;
  assign n4792 = pi120 & ~n4190;
  assign n4793 = ~n4791 & ~n4792;
  assign n4794 = n2559 & ~n4793;
  assign po267 = n4790 | n4794;
  assign n4796 = pi121 & ~n2559;
  assign n4797 = ~n2344 & n4190;
  assign n4798 = pi121 & ~n4190;
  assign n4799 = ~n4797 & ~n4798;
  assign n4800 = n2559 & ~n4799;
  assign po268 = n4796 | n4800;
  assign n4802 = pi122 & ~n2559;
  assign n4803 = ~n2031 & n4203;
  assign n4804 = pi122 & ~n4203;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = n2559 & ~n4805;
  assign po269 = n4802 | n4806;
  assign n4808 = pi123 & ~n2559;
  assign n4809 = ~n2119 & n4203;
  assign n4810 = pi123 & ~n4203;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = n2559 & ~n4811;
  assign po270 = n4808 | n4812;
  assign n4814 = pi124 & ~n2559;
  assign n4815 = ~n2344 & n4203;
  assign n4816 = pi124 & ~n4203;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n2559 & ~n4817;
  assign po271 = n4814 | n4818;
  assign n4820 = pi125 & ~n2559;
  assign n4821 = ~n2031 & n4338;
  assign n4822 = pi125 & ~n4338;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = n2559 & ~n4823;
  assign po272 = n4820 | n4824;
  assign n4826 = pi126 & ~n2559;
  assign n4827 = ~n2119 & n4338;
  assign n4828 = pi126 & ~n4338;
  assign n4829 = ~n4827 & ~n4828;
  assign n4830 = n2559 & ~n4829;
  assign po273 = n4826 | n4830;
  assign n4832 = pi127 & ~n2559;
  assign n4833 = ~n2344 & n4338;
  assign n4834 = pi127 & ~n4338;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = n2559 & ~n4835;
  assign po274 = n4832 | n4836;
  assign n4838 = pi128 & ~n2559;
  assign n4839 = ~n2344 & n4210;
  assign n4840 = pi128 & ~n4210;
  assign n4841 = ~n4839 & ~n4840;
  assign n4842 = n2559 & ~n4841;
  assign po275 = n4838 | n4842;
  assign n4844 = pi129 & ~n2559;
  assign n4845 = ~n2031 & n4210;
  assign n4846 = pi129 & ~n4210;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = n2559 & ~n4847;
  assign po276 = n4844 | n4848;
  assign n4850 = pi130 & ~n2559;
  assign n4851 = ~n2119 & n4210;
  assign n4852 = pi130 & ~n4210;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = n2559 & ~n4853;
  assign po277 = n4850 | n4854;
  assign n4856 = n2440 & ~n3748;
  assign n4857 = ~pi131 & ~n4354;
  assign n4858 = ~n4856 & ~n4857;
  assign n4859 = ~pi131 & ~n4357;
  assign po278 = ~n4858 | n4859;
  assign n4861 = ~po327 & ~n3623;
  assign n4862 = po327 & n3623;
  assign po279 = n4861 | n4862;
  assign n4864 = ~pi133 & ~po814;
  assign n4865 = ~n2046 & po814;
  assign po280 = n4864 | n4865;
  assign n4867 = ~pi134 & ~po814;
  assign n4868 = po814 & ~n2134;
  assign po281 = n4867 | n4868;
  assign n4870 = ~n2119 & n2440;
  assign n4871 = ~pi135 & ~n4354;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = ~pi135 & ~n4357;
  assign po282 = ~n4872 | n4873;
  assign n4875 = ~pi136 & ~po814;
  assign n4876 = po814 & ~n3763;
  assign po283 = n4875 | n4876;
  assign n4878 = ~n2344 & n2440;
  assign n4879 = ~pi137 & ~n4354;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = ~pi137 & ~n4357;
  assign po284 = ~n4880 | n4881;
  assign n4883 = ~n2031 & n2440;
  assign n4884 = ~pi138 & ~n4354;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = ~pi138 & ~n4357;
  assign po285 = ~n4885 | n4886;
  assign n4888 = n3818 & n3919;
  assign n4889 = pi139 & ~n3919;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n2559 & ~n4890;
  assign n4892 = pi142 & n2556;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = pi139 & n2558;
  assign po286 = ~n4893 | n4894;
  assign n4896 = n3818 & n3940;
  assign n4897 = pi140 & ~n3940;
  assign n4898 = ~n4896 & ~n4897;
  assign n4899 = n2559 & ~n4898;
  assign n4900 = pi141 & n2556;
  assign n4901 = ~n4899 & ~n4900;
  assign n4902 = pi140 & n2558;
  assign po287 = ~n4901 | n4902;
  assign n4904 = n3818 & n3974;
  assign n4905 = pi141 & ~n3974;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = n2559 & ~n4906;
  assign n4908 = pi140 & n2556;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = pi141 & n2558;
  assign po288 = ~n4909 | n4910;
  assign n4912 = n3818 & n3957;
  assign n4913 = pi142 & ~n3957;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = n2559 & ~n4914;
  assign n4916 = pi139 & n2556;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = pi142 & n2558;
  assign po289 = ~n4917 | n4918;
  assign n4920 = n3818 & n4022;
  assign n4921 = pi143 & ~n4022;
  assign n4922 = ~n4920 & ~n4921;
  assign n4923 = n2559 & ~n4922;
  assign n4924 = pi143 & n2558;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = pi147 & pi673;
  assign n4927 = pi151 & ~pi673;
  assign n4928 = ~n4926 & ~n4927;
  assign n4929 = n2556 & ~n4928;
  assign po290 = ~n4925 | n4929;
  assign n4931 = ~pi144 & ~n4354;
  assign n4932 = n2397 & ~n3748;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = ~pi144 & ~n4351;
  assign po291 = ~n4933 | n4934;
  assign n4936 = ~pi145 & ~n4735;
  assign n4937 = ~n2031 & n2412;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = ~pi145 & ~n4357;
  assign po292 = ~n4938 | n4939;
  assign n4941 = ~pi146 & ~n4735;
  assign n4942 = ~n2119 & n2412;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = ~pi146 & ~n4357;
  assign po293 = ~n4943 | n4944;
  assign n4946 = pi147 & ~n4047;
  assign n4947 = n3818 & n4047;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = n2559 & ~n4948;
  assign n4950 = pi147 & n2558;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = pi149 & pi673;
  assign n4953 = pi143 & ~pi673;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = n2556 & ~n4954;
  assign po294 = ~n4951 | n4955;
  assign n4957 = pi148 & ~n4116;
  assign n4958 = n3818 & n4116;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = n2559 & ~n4959;
  assign n4961 = pi148 & n2558;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = pi158 & ~pi673;
  assign n4964 = pi152 & pi673;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = n2556 & ~n4965;
  assign po295 = ~n4962 | n4966;
  assign n4968 = pi149 & ~n4093;
  assign n4969 = n3818 & n4093;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = n2559 & ~n4970;
  assign n4972 = pi149 & n2558;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = pi147 & ~pi673;
  assign n4975 = pi151 & pi673;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = n2556 & ~n4976;
  assign po296 = ~n4973 | n4977;
  assign n4979 = n3818 & n4139;
  assign n4980 = pi150 & ~n4139;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n2559 & ~n4981;
  assign n4983 = pi150 & n2558;
  assign n4984 = ~n4982 & ~n4983;
  assign n4985 = pi158 & pi673;
  assign n4986 = pi152 & ~pi673;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = n2556 & ~n4987;
  assign po297 = ~n4984 | n4988;
  assign n4990 = n3818 & n4162;
  assign n4991 = pi151 & ~n4162;
  assign n4992 = ~n4990 & ~n4991;
  assign n4993 = n2559 & ~n4992;
  assign n4994 = pi151 & n2558;
  assign n4995 = ~n4993 & ~n4994;
  assign n4996 = pi149 & ~pi673;
  assign n4997 = pi143 & pi673;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n2556 & ~n4998;
  assign po298 = ~n4995 | n4999;
  assign n5001 = n3818 & n3998;
  assign n5002 = pi152 & ~n3998;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = n2559 & ~n5003;
  assign n5005 = pi152 & n2558;
  assign n5006 = ~n5004 & ~n5005;
  assign n5007 = ~pi673 & n3818;
  assign n5008 = pi150 & pi673;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = n2556 & ~n5009;
  assign po299 = ~n5006 | n5010;
  assign n5012 = ~pi153 & ~n4735;
  assign n5013 = n2412 & ~n3748;
  assign n5014 = ~n5012 & ~n5013;
  assign n5015 = ~pi153 & ~n4357;
  assign po300 = ~n5014 | n5015;
  assign n5017 = ~pi154 & ~n4354;
  assign n5018 = ~n2119 & n2397;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = ~pi154 & ~n4351;
  assign po301 = ~n5019 | n5020;
  assign n5022 = ~pi155 & ~po814;
  assign n5023 = po814 & ~n2359;
  assign po302 = n5022 | n5023;
  assign n5025 = ~pi156 & ~n4354;
  assign n5026 = ~n2031 & n2397;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~pi156 & ~n4351;
  assign po303 = ~n5027 | n5028;
  assign n5030 = ~pi157 & ~n4354;
  assign n5031 = ~n2344 & n2397;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = ~pi157 & ~n4351;
  assign po304 = ~n5032 | n5033;
  assign n5035 = pi150 & ~pi673;
  assign n5036 = pi673 & n3818;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = n2556 & ~n5037;
  assign n5039 = pi158 & n2558;
  assign n5040 = ~n5038 & ~n5039;
  assign n5041 = n3818 & n4070;
  assign n5042 = pi158 & ~n4070;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = n2559 & ~n5043;
  assign po305 = ~n5040 | n5044;
  assign n5046 = ~pi159 & ~n4735;
  assign n5047 = ~n2344 & n2412;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = ~pi159 & ~n4357;
  assign po306 = ~n5048 | n5049;
  assign n5051 = pi160 & ~n2559;
  assign n5052 = n3818 & n4190;
  assign n5053 = pi160 & ~n4190;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = n2559 & ~n5054;
  assign po307 = n5051 | n5055;
  assign n5057 = pi161 & ~n2559;
  assign n5058 = n3818 & n4203;
  assign n5059 = pi161 & ~n4203;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = n2559 & ~n5060;
  assign po308 = n5057 | n5061;
  assign n5063 = pi162 & ~n2559;
  assign n5064 = n3818 & n4338;
  assign n5065 = pi162 & ~n4338;
  assign n5066 = ~n5064 & ~n5065;
  assign n5067 = n2559 & ~n5066;
  assign po309 = n5063 | n5067;
  assign n5069 = pi163 & ~n2559;
  assign n5070 = n3818 & n4210;
  assign n5071 = pi163 & ~n4210;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = n2559 & ~n5072;
  assign po310 = n5069 | n5073;
  assign n5075 = n3418 & ~po339;
  assign n5076 = ~n3418 & po339;
  assign po312 = n5075 | n5076;
  assign n5078 = ~n3869 & n3919;
  assign n5079 = pi168 & ~n3919;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = n2559 & ~n5080;
  assign n5082 = pi169 & n2556;
  assign n5083 = ~n5081 & ~n5082;
  assign n5084 = pi168 & n2558;
  assign po317 = ~n5083 | n5084;
  assign n5086 = ~n3869 & n3957;
  assign n5087 = pi169 & ~n3957;
  assign n5088 = ~n5086 & ~n5087;
  assign n5089 = n2559 & ~n5088;
  assign n5090 = pi168 & n2556;
  assign n5091 = ~n5089 & ~n5090;
  assign n5092 = pi169 & n2558;
  assign po318 = ~n5091 | n5092;
  assign n5094 = ~n3869 & n3974;
  assign n5095 = pi170 & ~n3974;
  assign n5096 = ~n5094 & ~n5095;
  assign n5097 = n2559 & ~n5096;
  assign n5098 = pi171 & n2556;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = pi170 & n2558;
  assign po319 = ~n5099 | n5100;
  assign n5102 = ~n3869 & n3940;
  assign n5103 = pi171 & ~n3940;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = n2559 & ~n5104;
  assign n5106 = pi170 & n2556;
  assign n5107 = ~n5105 & ~n5106;
  assign n5108 = pi171 & n2558;
  assign po320 = ~n5107 | n5108;
  assign n5110 = pi172 & ~n4047;
  assign n5111 = ~n3869 & n4047;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n2559 & ~n5112;
  assign n5114 = pi172 & n2558;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = pi180 & pi673;
  assign n5117 = pi181 & ~pi673;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = n2556 & ~n5118;
  assign po321 = ~n5115 | n5119;
  assign n5121 = ~pi173 & ~n4116;
  assign n5122 = ~n3869 & n4116;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = n2559 & ~n5123;
  assign n5125 = ~pi173 & n2558;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = pi182 & ~pi673;
  assign n5128 = pi175 & pi673;
  assign n5129 = ~n5127 & ~n5128;
  assign n5130 = n2556 & ~n5129;
  assign po322 = ~n5126 | n5130;
  assign n5132 = ~n3869 & n4139;
  assign n5133 = pi174 & ~n4139;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = n2559 & ~n5134;
  assign n5136 = pi174 & n2558;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = pi182 & pi673;
  assign n5139 = pi175 & ~pi673;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = n2556 & ~n5140;
  assign po323 = ~n5137 | n5141;
  assign n5143 = ~n3869 & n3998;
  assign n5144 = pi175 & ~n3998;
  assign n5145 = ~n5143 & ~n5144;
  assign n5146 = n2559 & ~n5145;
  assign n5147 = pi175 & n2558;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = ~pi673 & ~n3869;
  assign n5150 = pi174 & pi673;
  assign n5151 = ~n5149 & ~n5150;
  assign n5152 = n2556 & ~n5151;
  assign po324 = ~n5148 | n5152;
  assign n5154 = ~pi176 & ~po814;
  assign n5155 = po814 & ~n3884;
  assign po325 = n5154 | n5155;
  assign n5157 = n2440 & n3818;
  assign n5158 = ~pi177 & ~n4354;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = ~pi177 & ~n4357;
  assign po326 = ~n5159 | n5160;
  assign n5162 = ~n3869 & n4162;
  assign n5163 = pi179 & ~n4162;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = n2559 & ~n5164;
  assign n5166 = pi179 & n2558;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = pi180 & ~pi673;
  assign n5169 = pi181 & pi673;
  assign n5170 = ~n5168 & ~n5169;
  assign n5171 = n2556 & ~n5170;
  assign po328 = ~n5167 | n5171;
  assign n5173 = pi180 & ~n4093;
  assign n5174 = ~n3869 & n4093;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = n2559 & ~n5175;
  assign n5177 = pi180 & n2558;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = pi172 & ~pi673;
  assign n5180 = pi179 & pi673;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = n2556 & ~n5181;
  assign po329 = ~n5178 | n5182;
  assign n5184 = ~n3869 & n4022;
  assign n5185 = pi181 & ~n4022;
  assign n5186 = ~n5184 & ~n5185;
  assign n5187 = n2559 & ~n5186;
  assign n5188 = pi181 & n2558;
  assign n5189 = ~n5187 & ~n5188;
  assign n5190 = pi172 & pi673;
  assign n5191 = pi179 & ~pi673;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = n2556 & ~n5192;
  assign po330 = ~n5189 | n5193;
  assign n5195 = pi174 & ~pi673;
  assign n5196 = pi673 & ~n3869;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = n2556 & ~n5197;
  assign n5199 = pi182 & n2558;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = ~n3869 & n4070;
  assign n5202 = pi182 & ~n4070;
  assign n5203 = ~n5201 & ~n5202;
  assign n5204 = n2559 & ~n5203;
  assign po331 = ~n5200 | n5204;
  assign n5206 = ~pi183 & ~n2559;
  assign n5207 = ~n3869 & n4338;
  assign n5208 = ~pi183 & ~n4338;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n2559 & ~n5209;
  assign po332 = n5206 | n5210;
  assign n5212 = ~pi184 & ~n2559;
  assign n5213 = ~n3869 & n4210;
  assign n5214 = ~pi184 & ~n4210;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = n2559 & ~n5215;
  assign po333 = n5212 | n5216;
  assign n5218 = ~pi185 & ~n2559;
  assign n5219 = ~n3869 & n4203;
  assign n5220 = ~pi185 & ~n4203;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = n2559 & ~n5221;
  assign po334 = n5218 | n5222;
  assign n5224 = ~pi186 & ~n4354;
  assign n5225 = n2397 & n3818;
  assign n5226 = ~n5224 & ~n5225;
  assign n5227 = ~pi186 & ~n4351;
  assign po335 = ~n5226 | n5227;
  assign n5229 = ~pi187 & ~n2559;
  assign n5230 = ~n3869 & n4190;
  assign n5231 = ~pi187 & ~n4190;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = n2559 & ~n5232;
  assign po336 = n5229 | n5233;
  assign n5235 = ~pi188 & ~po814;
  assign n5236 = po814 & ~n3836;
  assign po337 = n5235 | n5236;
  assign n5238 = ~pi189 & ~n4735;
  assign n5239 = n2412 & n3818;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = ~pi189 & ~n4357;
  assign po338 = ~n5240 | n5241;
  assign n5243 = n2440 & ~n3869;
  assign n5244 = ~pi191 & ~n4354;
  assign n5245 = ~n5243 & ~n5244;
  assign n5246 = ~pi191 & ~n4357;
  assign po340 = ~n5245 | n5246;
  assign n5248 = ~po344 & ~n3590;
  assign n5249 = po344 & n3590;
  assign po341 = n5248 | n5249;
  assign n5251 = ~pi193 & ~n4354;
  assign n5252 = n2397 & ~n3869;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~pi193 & ~n4351;
  assign po342 = ~n5253 | n5254;
  assign n5256 = ~pi194 & ~n4735;
  assign n5257 = n2412 & ~n3869;
  assign n5258 = ~n5256 & ~n5257;
  assign n5259 = ~pi194 & ~n4357;
  assign po343 = ~n5258 | n5259;
  assign n5261 = pi196 & ~po814;
  assign n5262 = pi862 & n1761;
  assign n5263 = ~pi204 & n1787;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = ~n1754 & ~n5264;
  assign n5266 = pi862 & n1756;
  assign n5267 = ~pi204 & ~n1756;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n1792 & ~n5268;
  assign n5270 = ~n5265 & ~n5269;
  assign n5271 = pi894 & n1756;
  assign n5272 = ~pi228 & ~n1756;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = ~n1778 & ~n5273;
  assign n5275 = ~pi228 & n1778;
  assign n5276 = ~n5274 & ~n5275;
  assign n5277 = ~n1761 & ~n5276;
  assign n5278 = pi894 & n1761;
  assign n5279 = ~n5277 & ~n5278;
  assign n5280 = ~n1754 & ~n5279;
  assign n5281 = n1754 & ~n5273;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~pi390 & n1778;
  assign n5284 = pi390 & ~n1778;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n1761 & n5285;
  assign n5287 = ~n1754 & ~n5286;
  assign n5288 = pi390 & n1754;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n1754 & ~n1761;
  assign n5291 = pi390 & pi550;
  assign n5292 = ~pi390 & ~pi550;
  assign n5293 = n1778 & ~n5292;
  assign n5294 = ~n5291 & n5293;
  assign n5295 = pi550 & ~n1778;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = n5290 & ~n5296;
  assign n5298 = pi550 & n1754;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = pi552 & n5291;
  assign n5301 = pi551 & n5300;
  assign n5302 = ~pi551 & ~n5300;
  assign n5303 = ~n5301 & ~n5302;
  assign n5304 = n1778 & n5303;
  assign n5305 = pi551 & ~n1778;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = n5290 & ~n5306;
  assign n5308 = pi551 & n1754;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = pi552 & n1754;
  assign n5311 = ~pi552 & ~n5291;
  assign n5312 = n1778 & ~n5311;
  assign n5313 = ~n5300 & n5312;
  assign n5314 = pi552 & ~n1778;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = n5290 & ~n5315;
  assign n5317 = ~n5310 & ~n5316;
  assign n5318 = ~n5309 & n5317;
  assign n5319 = n5299 & n5318;
  assign n5320 = ~n5289 & n5319;
  assign n5321 = n5309 & ~n5317;
  assign n5322 = ~n5289 & n5321;
  assign n5323 = n5299 & n5322;
  assign n5324 = ~n5320 & ~n5323;
  assign n5325 = n5289 & n5318;
  assign n5326 = ~n5299 & n5325;
  assign n5327 = n5324 & ~n5326;
  assign n5328 = pi926 & n1756;
  assign n5329 = pi288 & ~n1756;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = n1754 & ~n5330;
  assign n5332 = pi288 & n1787;
  assign n5333 = n1791 & ~n5330;
  assign n5334 = pi926 & n1761;
  assign n5335 = ~n5333 & ~n5334;
  assign n5336 = ~n5332 & n5335;
  assign n5337 = ~n1754 & ~n5336;
  assign n5338 = ~n5331 & ~n5337;
  assign n5339 = ~pi154 & ~n5338;
  assign n5340 = pi154 & n5338;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = n5327 & n5341;
  assign n5343 = ~n5327 & ~n5341;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = ~n5282 & n5344;
  assign n5346 = n5282 & ~n5344;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = n5270 & n5347;
  assign n5349 = ~n5270 & ~n5347;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = n2826 & n5350;
  assign n5352 = ~n2826 & ~n5350;
  assign n5353 = ~n5351 & ~n5352;
  assign n5354 = po814 & ~n5353;
  assign po345 = n5261 | n5354;
  assign n5356 = pi197 & ~po814;
  assign n5357 = pi861 & n1761;
  assign n5358 = ~pi215 & n1787;
  assign n5359 = ~n5357 & ~n5358;
  assign n5360 = ~n1754 & ~n5359;
  assign n5361 = pi861 & n1756;
  assign n5362 = ~pi215 & ~n1756;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = ~n1792 & ~n5363;
  assign n5365 = ~n5360 & ~n5364;
  assign n5366 = pi238 & n1778;
  assign n5367 = pi893 & n1756;
  assign n5368 = pi238 & ~n1756;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = ~n1778 & ~n5369;
  assign n5371 = ~n5366 & ~n5370;
  assign n5372 = ~n1761 & ~n5371;
  assign n5373 = pi893 & n1761;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n1754 & ~n5374;
  assign n5376 = n1754 & ~n5369;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = n5289 & n5321;
  assign n5379 = n5299 & n5378;
  assign n5380 = ~n5320 & ~n5379;
  assign n5381 = pi925 & n1761;
  assign n5382 = pi333 & n1787;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = ~n1754 & ~n5383;
  assign n5385 = pi925 & n1756;
  assign n5386 = pi333 & ~n1756;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = ~n1792 & ~n5387;
  assign n5389 = ~n5384 & ~n5388;
  assign n5390 = ~pi156 & ~n5389;
  assign n5391 = pi156 & n5389;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = n5380 & n5392;
  assign n5394 = ~n5380 & ~n5392;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~n5377 & n5395;
  assign n5397 = n5377 & ~n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = ~n5365 & n5398;
  assign n5400 = n5365 & ~n5398;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = ~n3152 & n5401;
  assign n5403 = n3152 & ~n5401;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = po814 & ~n5404;
  assign po346 = n5356 | n5405;
  assign n5407 = pi198 & ~po814;
  assign n5408 = pi863 & n1761;
  assign n5409 = ~pi214 & n1787;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n1754 & ~n5410;
  assign n5412 = pi863 & n1756;
  assign n5413 = ~pi214 & ~n1756;
  assign n5414 = ~n5412 & ~n5413;
  assign n5415 = ~n1792 & ~n5414;
  assign n5416 = ~n5411 & ~n5415;
  assign n5417 = pi895 & n1761;
  assign n5418 = pi895 & n1756;
  assign n5419 = ~pi239 & ~n1756;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = ~n1778 & ~n5420;
  assign n5422 = ~pi239 & n1778;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = ~n1761 & ~n5423;
  assign n5425 = ~n5417 & ~n5424;
  assign n5426 = ~n1754 & ~n5425;
  assign n5427 = n1754 & ~n5420;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~n5299 & n5378;
  assign n5430 = ~n5326 & ~n5429;
  assign n5431 = pi927 & n1761;
  assign n5432 = pi332 & n1787;
  assign n5433 = ~n5431 & ~n5432;
  assign n5434 = ~n1754 & ~n5433;
  assign n5435 = pi927 & n1756;
  assign n5436 = pi332 & ~n1756;
  assign n5437 = ~n5435 & ~n5436;
  assign n5438 = ~n1792 & ~n5437;
  assign n5439 = ~n5434 & ~n5438;
  assign n5440 = ~pi117 & ~n5439;
  assign n5441 = pi117 & n5439;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = n5430 & n5442;
  assign n5444 = ~n5430 & ~n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n5428 & n5445;
  assign n5447 = ~n5428 & ~n5445;
  assign n5448 = ~n5446 & ~n5447;
  assign n5449 = n5416 & n5448;
  assign n5450 = ~n5416 & ~n5448;
  assign n5451 = ~n5449 & ~n5450;
  assign n5452 = ~n3440 & n5451;
  assign n5453 = n3440 & ~n5451;
  assign n5454 = ~n5452 & ~n5453;
  assign n5455 = po814 & ~n5454;
  assign po347 = n5407 | n5455;
  assign n5457 = pi199 & ~po814;
  assign n5458 = pi864 & n1761;
  assign n5459 = ~pi226 & n1787;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = ~n1754 & ~n5460;
  assign n5462 = pi864 & n1756;
  assign n5463 = ~pi226 & ~n1756;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = ~n1792 & ~n5464;
  assign n5466 = ~n5461 & ~n5465;
  assign n5467 = pi249 & n1778;
  assign n5468 = pi896 & n1756;
  assign n5469 = pi249 & ~n1756;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = ~n1778 & ~n5470;
  assign n5472 = ~n5467 & ~n5471;
  assign n5473 = ~n1761 & ~n5472;
  assign n5474 = pi896 & n1761;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = ~n1754 & ~n5475;
  assign n5477 = n1754 & ~n5470;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = ~n5299 & n5322;
  assign n5480 = pi928 & n1761;
  assign n5481 = pi394 & n1787;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = ~n1754 & ~n5482;
  assign n5484 = pi928 & n1756;
  assign n5485 = pi394 & ~n1756;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n1792 & ~n5486;
  assign n5488 = ~n5483 & ~n5487;
  assign n5489 = ~pi111 & ~n5488;
  assign n5490 = pi111 & n5488;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = ~n5479 & n5491;
  assign n5493 = n5479 & ~n5491;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = ~n5478 & n5494;
  assign n5496 = n5478 & ~n5494;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = ~n5466 & n5497;
  assign n5499 = n5466 & ~n5497;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = ~n2425 & n5500;
  assign n5502 = n2425 & ~n5500;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = po814 & ~n5503;
  assign po348 = n5457 | n5504;
  assign n5506 = pi200 & ~po814;
  assign n5507 = pi858 & n1761;
  assign n5508 = ~pi227 & n1787;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n1754 & ~n5509;
  assign n5511 = pi858 & n1756;
  assign n5512 = ~pi227 & ~n1756;
  assign n5513 = ~n5511 & ~n5512;
  assign n5514 = ~n1792 & ~n5513;
  assign n5515 = ~n5510 & ~n5514;
  assign n5516 = pi248 & n1778;
  assign n5517 = pi890 & n1756;
  assign n5518 = pi248 & ~n1756;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = ~n1778 & ~n5519;
  assign n5521 = ~n5516 & ~n5520;
  assign n5522 = ~n1761 & ~n5521;
  assign n5523 = pi890 & n1761;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n1754 & ~n5524;
  assign n5526 = n1754 & ~n5519;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = ~n5289 & n5317;
  assign n5529 = n5299 & n5528;
  assign n5530 = pi922 & n1761;
  assign n5531 = pi387 & n1787;
  assign n5532 = ~n5530 & ~n5531;
  assign n5533 = ~n1754 & ~n5532;
  assign n5534 = pi922 & n1756;
  assign n5535 = pi387 & ~n1756;
  assign n5536 = ~n5534 & ~n5535;
  assign n5537 = ~n1792 & ~n5536;
  assign n5538 = ~n5533 & ~n5537;
  assign n5539 = ~pi144 & ~n5538;
  assign n5540 = pi144 & n5538;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = ~n5529 & n5541;
  assign n5543 = n5529 & ~n5541;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = ~n5527 & n5544;
  assign n5546 = n5527 & ~n5544;
  assign n5547 = ~n5545 & ~n5546;
  assign n5548 = ~n5515 & n5547;
  assign n5549 = n5515 & ~n5547;
  assign n5550 = ~n5548 & ~n5549;
  assign n5551 = ~n2998 & n5550;
  assign n5552 = n2998 & ~n5550;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = po814 & ~n5553;
  assign po349 = n5506 | n5554;
  assign n5556 = pi201 & ~po814;
  assign n5557 = pi865 & n1761;
  assign n5558 = ~pi225 & n1787;
  assign n5559 = ~n5557 & ~n5558;
  assign n5560 = ~n1754 & ~n5559;
  assign n5561 = pi865 & n1756;
  assign n5562 = ~pi225 & ~n1756;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = ~n1792 & ~n5563;
  assign n5565 = ~n5560 & ~n5564;
  assign n5566 = pi250 & n1778;
  assign n5567 = pi897 & n1756;
  assign n5568 = pi250 & ~n1756;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = ~n1778 & ~n5569;
  assign n5571 = ~n5566 & ~n5570;
  assign n5572 = ~n1761 & ~n5571;
  assign n5573 = pi897 & n1761;
  assign n5574 = ~n5572 & ~n5573;
  assign n5575 = ~n1754 & ~n5574;
  assign n5576 = n1754 & ~n5569;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = n5299 & n5325;
  assign n5579 = pi929 & n1761;
  assign n5580 = pi389 & n1787;
  assign n5581 = ~n5579 & ~n5580;
  assign n5582 = ~n1754 & ~n5581;
  assign n5583 = pi929 & n1756;
  assign n5584 = pi389 & ~n1756;
  assign n5585 = ~n5583 & ~n5584;
  assign n5586 = ~n1792 & ~n5585;
  assign n5587 = ~n5582 & ~n5586;
  assign n5588 = ~pi157 & ~n5587;
  assign n5589 = pi157 & n5587;
  assign n5590 = ~n5588 & ~n5589;
  assign n5591 = ~n5578 & n5590;
  assign n5592 = n5578 & ~n5590;
  assign n5593 = ~n5591 & ~n5592;
  assign n5594 = ~n5577 & n5593;
  assign n5595 = n5577 & ~n5593;
  assign n5596 = ~n5594 & ~n5595;
  assign n5597 = ~n5565 & n5596;
  assign n5598 = n5565 & ~n5596;
  assign n5599 = ~n5597 & ~n5598;
  assign n5600 = ~n2867 & n5599;
  assign n5601 = n2867 & ~n5599;
  assign n5602 = ~n5600 & ~n5601;
  assign n5603 = po814 & ~n5602;
  assign po350 = n5556 | n5603;
  assign n5605 = pi202 & ~po814;
  assign n5606 = pi859 & n1761;
  assign n5607 = ~pi223 & n1787;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n1754 & ~n5608;
  assign n5610 = pi859 & n1756;
  assign n5611 = ~pi223 & ~n1756;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = ~n1792 & ~n5612;
  assign n5614 = ~n5609 & ~n5613;
  assign n5615 = pi251 & n1778;
  assign n5616 = pi891 & n1756;
  assign n5617 = pi251 & ~n1756;
  assign n5618 = ~n5616 & ~n5617;
  assign n5619 = ~n1778 & ~n5618;
  assign n5620 = ~n5615 & ~n5619;
  assign n5621 = ~n1761 & ~n5620;
  assign n5622 = pi891 & n1761;
  assign n5623 = ~n5621 & ~n5622;
  assign n5624 = ~n1754 & ~n5623;
  assign n5625 = n1754 & ~n5618;
  assign n5626 = ~n5624 & ~n5625;
  assign n5627 = ~n5299 & n5317;
  assign n5628 = n5289 & n5627;
  assign n5629 = ~n5320 & ~n5628;
  assign n5630 = pi923 & n1761;
  assign n5631 = pi388 & n1787;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = ~n1754 & ~n5632;
  assign n5634 = pi923 & n1756;
  assign n5635 = pi388 & ~n1756;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n1792 & ~n5636;
  assign n5638 = ~n5633 & ~n5637;
  assign n5639 = ~pi193 & ~n5638;
  assign n5640 = pi193 & n5638;
  assign n5641 = ~n5639 & ~n5640;
  assign n5642 = n5629 & n5641;
  assign n5643 = ~n5629 & ~n5641;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = ~n5626 & n5644;
  assign n5646 = n5626 & ~n5644;
  assign n5647 = ~n5645 & ~n5646;
  assign n5648 = ~n5614 & n5647;
  assign n5649 = n5614 & ~n5647;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = ~n2712 & n5650;
  assign n5652 = n2712 & ~n5650;
  assign n5653 = ~n5651 & ~n5652;
  assign n5654 = po814 & ~n5653;
  assign po351 = n5605 | n5654;
  assign n5656 = pi203 & ~po814;
  assign n5657 = pi860 & n1761;
  assign n5658 = ~pi224 & n1787;
  assign n5659 = ~n5657 & ~n5658;
  assign n5660 = ~n1754 & ~n5659;
  assign n5661 = pi860 & n1756;
  assign n5662 = ~pi224 & ~n1756;
  assign n5663 = ~n5661 & ~n5662;
  assign n5664 = ~n1792 & ~n5663;
  assign n5665 = ~n5660 & ~n5664;
  assign n5666 = pi892 & n1761;
  assign n5667 = pi892 & n1756;
  assign n5668 = ~pi247 & ~n1756;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = ~n1778 & ~n5669;
  assign n5671 = ~pi247 & n1778;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = ~n1761 & ~n5672;
  assign n5674 = ~n5666 & ~n5673;
  assign n5675 = ~n1754 & ~n5674;
  assign n5676 = n1754 & ~n5669;
  assign n5677 = ~n5675 & ~n5676;
  assign n5678 = ~n5289 & n5309;
  assign n5679 = n5627 & n5678;
  assign n5680 = ~n5326 & ~n5679;
  assign n5681 = pi924 & n1761;
  assign n5682 = pi396 & n1787;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = ~n1754 & ~n5683;
  assign n5685 = pi924 & n1756;
  assign n5686 = pi396 & ~n1756;
  assign n5687 = ~n5685 & ~n5686;
  assign n5688 = ~n1792 & ~n5687;
  assign n5689 = ~n5684 & ~n5688;
  assign n5690 = ~pi186 & ~n5689;
  assign n5691 = pi186 & n5689;
  assign n5692 = ~n5690 & ~n5691;
  assign n5693 = n5680 & n5692;
  assign n5694 = ~n5680 & ~n5692;
  assign n5695 = ~n5693 & ~n5694;
  assign n5696 = n5677 & n5695;
  assign n5697 = ~n5677 & ~n5695;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = n5665 & n5698;
  assign n5700 = ~n5665 & ~n5698;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = ~n3368 & n5701;
  assign n5703 = n3368 & ~n5701;
  assign n5704 = ~n5702 & ~n5703;
  assign n5705 = po814 & ~n5704;
  assign po352 = n5656 | n5705;
  assign n5707 = po814 & n5350;
  assign n5708 = ~pi204 & ~po814;
  assign po353 = n5707 | n5708;
  assign n5710 = pi205 & ~po814;
  assign n5711 = pi292 & n1778;
  assign n5712 = pi868 & n1756;
  assign n5713 = pi292 & ~n1756;
  assign n5714 = ~n5712 & ~n5713;
  assign n5715 = ~n1778 & ~n5714;
  assign n5716 = ~n5711 & ~n5715;
  assign n5717 = ~n1761 & ~n5716;
  assign n5718 = pi868 & n1761;
  assign n5719 = ~n5717 & ~n5718;
  assign n5720 = ~n1754 & ~n5719;
  assign n5721 = n1754 & ~n5714;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = pi900 & n1761;
  assign n5724 = pi414 & ~n1756;
  assign n5725 = pi900 & n1756;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n1778 & ~n5726;
  assign n5728 = pi414 & n1778;
  assign n5729 = ~n5727 & ~n5728;
  assign n5730 = ~n1761 & ~n5729;
  assign n5731 = ~n5723 & ~n5730;
  assign n5732 = ~n1754 & ~n5731;
  assign n5733 = n1754 & ~n5726;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = pi189 & ~n5734;
  assign n5736 = ~pi189 & n5734;
  assign n5737 = ~n5735 & ~n5736;
  assign n5738 = ~n5722 & n5737;
  assign n5739 = n5722 & ~n5737;
  assign n5740 = ~n5738 & ~n5739;
  assign n5741 = pi836 & n1761;
  assign n5742 = ~pi231 & n1787;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = ~n1754 & ~n5743;
  assign n5745 = pi836 & n1756;
  assign n5746 = ~pi231 & ~n1756;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~n1792 & ~n5747;
  assign n5749 = ~n5744 & ~n5748;
  assign n5750 = ~n5740 & ~n5749;
  assign n5751 = n5740 & n5749;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = n3394 & n5752;
  assign n5754 = ~n3394 & ~n5752;
  assign n5755 = ~n5753 & ~n5754;
  assign n5756 = po814 & ~n5755;
  assign po354 = n5710 | n5756;
  assign n5758 = pi206 & ~po814;
  assign n5759 = pi837 & n1761;
  assign n5760 = pi837 & n1756;
  assign n5761 = ~pi232 & ~n1756;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = ~n1778 & ~n5762;
  assign n5764 = ~pi232 & n1778;
  assign n5765 = ~n5763 & ~n5764;
  assign n5766 = ~n1761 & ~n5765;
  assign n5767 = ~n5759 & ~n5766;
  assign n5768 = ~n1754 & ~n5767;
  assign n5769 = n1754 & ~n5762;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = pi869 & n1756;
  assign n5772 = pi291 & ~n1756;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = n1754 & ~n5773;
  assign n5775 = pi291 & n1787;
  assign n5776 = n1791 & ~n5773;
  assign n5777 = pi869 & n1761;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = ~n5775 & n5778;
  assign n5780 = ~n1754 & ~n5779;
  assign n5781 = ~n5774 & ~n5780;
  assign n5782 = pi901 & n1761;
  assign n5783 = pi901 & n1756;
  assign n5784 = pi437 & ~n1756;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~n1778 & ~n5785;
  assign n5787 = pi437 & n1778;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = ~n1761 & ~n5788;
  assign n5790 = ~n5782 & ~n5789;
  assign n5791 = ~n1754 & ~n5790;
  assign n5792 = n1754 & ~n5785;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = pi145 & ~n5793;
  assign n5795 = ~pi145 & n5793;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = n5781 & ~n5796;
  assign n5798 = ~n5781 & n5796;
  assign n5799 = ~n5797 & ~n5798;
  assign n5800 = n5770 & n5799;
  assign n5801 = ~n5770 & ~n5799;
  assign n5802 = ~n5800 & ~n5801;
  assign n5803 = n3166 & n5802;
  assign n5804 = ~n3166 & ~n5802;
  assign n5805 = ~n5803 & ~n5804;
  assign n5806 = po814 & ~n5805;
  assign po355 = n5758 | n5806;
  assign n5808 = pi207 & ~po814;
  assign n5809 = pi838 & n1761;
  assign n5810 = pi838 & n1756;
  assign n5811 = ~pi233 & ~n1756;
  assign n5812 = ~n5810 & ~n5811;
  assign n5813 = ~n1778 & ~n5812;
  assign n5814 = ~pi233 & n1778;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n1761 & ~n5815;
  assign n5817 = ~n5809 & ~n5816;
  assign n5818 = ~n1754 & ~n5817;
  assign n5819 = n1754 & ~n5812;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = pi902 & n1761;
  assign n5822 = pi902 & n1756;
  assign n5823 = pi415 & ~n1756;
  assign n5824 = ~n5822 & ~n5823;
  assign n5825 = ~n1778 & ~n5824;
  assign n5826 = pi415 & n1778;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = ~n1761 & ~n5827;
  assign n5829 = ~n5821 & ~n5828;
  assign n5830 = ~n1754 & ~n5829;
  assign n5831 = n1754 & ~n5824;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = pi146 & ~n5832;
  assign n5834 = ~pi146 & n5832;
  assign n5835 = ~n5833 & ~n5834;
  assign n5836 = pi870 & n1761;
  assign n5837 = pi293 & n1787;
  assign n5838 = ~n5836 & ~n5837;
  assign n5839 = ~n1754 & ~n5838;
  assign n5840 = pi870 & n1756;
  assign n5841 = pi293 & ~n1756;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n1792 & ~n5842;
  assign n5844 = ~n5839 & ~n5843;
  assign n5845 = ~n5835 & n5844;
  assign n5846 = n5835 & ~n5844;
  assign n5847 = ~n5845 & ~n5846;
  assign n5848 = n5820 & n5847;
  assign n5849 = ~n5820 & ~n5847;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = n2813 & n5850;
  assign n5852 = ~n2813 & ~n5850;
  assign n5853 = ~n5851 & ~n5852;
  assign n5854 = po814 & ~n5853;
  assign po356 = n5808 | n5854;
  assign n5856 = pi208 & ~po814;
  assign n5857 = pi839 & n1761;
  assign n5858 = pi839 & n1756;
  assign n5859 = ~pi237 & ~n1756;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~n1778 & ~n5860;
  assign n5862 = ~pi237 & n1778;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = ~n1761 & ~n5863;
  assign n5865 = ~n5857 & ~n5864;
  assign n5866 = ~n1754 & ~n5865;
  assign n5867 = n1754 & ~n5860;
  assign n5868 = ~n5866 & ~n5867;
  assign n5869 = pi903 & n1761;
  assign n5870 = pi903 & n1756;
  assign n5871 = pi416 & ~n1756;
  assign n5872 = ~n5870 & ~n5871;
  assign n5873 = ~n1778 & ~n5872;
  assign n5874 = pi416 & n1778;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n1761 & ~n5875;
  assign n5877 = ~n5869 & ~n5876;
  assign n5878 = ~n1754 & ~n5877;
  assign n5879 = n1754 & ~n5872;
  assign n5880 = ~n5878 & ~n5879;
  assign n5881 = pi114 & ~n5880;
  assign n5882 = ~pi114 & n5880;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = pi871 & n1761;
  assign n5885 = pi252 & n1787;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = ~n1754 & ~n5886;
  assign n5888 = pi871 & n1756;
  assign n5889 = pi252 & ~n1756;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = ~n1792 & ~n5890;
  assign n5892 = ~n5887 & ~n5891;
  assign n5893 = ~n5883 & n5892;
  assign n5894 = n5883 & ~n5892;
  assign n5895 = ~n5893 & ~n5894;
  assign n5896 = n5868 & n5895;
  assign n5897 = ~n5868 & ~n5895;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = ~n3453 & n5898;
  assign n5900 = n3453 & ~n5898;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = po814 & ~n5901;
  assign po357 = n5856 | n5902;
  assign n5904 = pi209 & ~po814;
  assign n5905 = pi840 & n1761;
  assign n5906 = pi840 & n1756;
  assign n5907 = ~pi234 & ~n1756;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = ~n1778 & ~n5908;
  assign n5910 = ~pi234 & n1778;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = ~n1761 & ~n5911;
  assign n5913 = ~n5905 & ~n5912;
  assign n5914 = ~n1754 & ~n5913;
  assign n5915 = n1754 & ~n5908;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = pi904 & n1761;
  assign n5918 = pi904 & n1756;
  assign n5919 = pi417 & ~n1756;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n1778 & ~n5920;
  assign n5922 = pi417 & n1778;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~n1761 & ~n5923;
  assign n5925 = ~n5917 & ~n5924;
  assign n5926 = ~n1754 & ~n5925;
  assign n5927 = n1754 & ~n5920;
  assign n5928 = ~n5926 & ~n5927;
  assign n5929 = pi113 & ~n5928;
  assign n5930 = ~pi113 & n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = pi872 & n1761;
  assign n5933 = pi294 & n1787;
  assign n5934 = ~n5932 & ~n5933;
  assign n5935 = ~n1754 & ~n5934;
  assign n5936 = pi872 & n1756;
  assign n5937 = pi294 & ~n1756;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = ~n1792 & ~n5938;
  assign n5940 = ~n5935 & ~n5939;
  assign n5941 = ~n5931 & n5940;
  assign n5942 = n5931 & ~n5940;
  assign n5943 = ~n5941 & ~n5942;
  assign n5944 = n5916 & n5943;
  assign n5945 = ~n5916 & ~n5943;
  assign n5946 = ~n5944 & ~n5945;
  assign n5947 = ~n2438 & n5946;
  assign n5948 = n2438 & ~n5946;
  assign n5949 = ~n5947 & ~n5948;
  assign n5950 = po814 & ~n5949;
  assign po358 = n5904 | n5950;
  assign n5952 = pi210 & ~po814;
  assign n5953 = pi289 & n1778;
  assign n5954 = pi866 & n1756;
  assign n5955 = pi289 & ~n1756;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~n1778 & ~n5956;
  assign n5958 = ~n5953 & ~n5957;
  assign n5959 = ~n1761 & ~n5958;
  assign n5960 = pi866 & n1761;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~n1754 & ~n5961;
  assign n5963 = n1754 & ~n5956;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = pi898 & n1761;
  assign n5966 = pi898 & n1756;
  assign n5967 = pi413 & ~n1756;
  assign n5968 = ~n5966 & ~n5967;
  assign n5969 = ~n1778 & ~n5968;
  assign n5970 = pi413 & n1778;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = ~n1761 & ~n5971;
  assign n5973 = ~n5965 & ~n5972;
  assign n5974 = ~n1754 & ~n5973;
  assign n5975 = n1754 & ~n5968;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = pi153 & ~n5976;
  assign n5978 = ~pi153 & n5976;
  assign n5979 = ~n5977 & ~n5978;
  assign n5980 = ~n5964 & n5979;
  assign n5981 = n5964 & ~n5979;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = pi834 & n1761;
  assign n5984 = ~pi229 & n1787;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = ~n1754 & ~n5985;
  assign n5987 = pi834 & n1756;
  assign n5988 = ~pi229 & ~n1756;
  assign n5989 = ~n5987 & ~n5988;
  assign n5990 = ~n1792 & ~n5989;
  assign n5991 = ~n5986 & ~n5990;
  assign n5992 = ~n5982 & ~n5991;
  assign n5993 = n5982 & n5991;
  assign n5994 = ~n5992 & ~n5993;
  assign n5995 = n3038 & n5994;
  assign n5996 = ~n3038 & ~n5994;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = po814 & ~n5997;
  assign po359 = n5952 | n5998;
  assign n6000 = pi211 & ~po814;
  assign n6001 = pi290 & n1778;
  assign n6002 = pi867 & n1756;
  assign n6003 = pi290 & ~n1756;
  assign n6004 = ~n6002 & ~n6003;
  assign n6005 = ~n1778 & ~n6004;
  assign n6006 = ~n6001 & ~n6005;
  assign n6007 = ~n1761 & ~n6006;
  assign n6008 = pi867 & n1761;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = ~n1754 & ~n6009;
  assign n6011 = n1754 & ~n6004;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = pi899 & n1761;
  assign n6014 = pi899 & n1756;
  assign n6015 = pi409 & ~n1756;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = ~n1778 & ~n6016;
  assign n6018 = pi409 & n1778;
  assign n6019 = ~n6017 & ~n6018;
  assign n6020 = ~n1761 & ~n6019;
  assign n6021 = ~n6013 & ~n6020;
  assign n6022 = ~n1754 & ~n6021;
  assign n6023 = n1754 & ~n6016;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = pi194 & ~n6024;
  assign n6026 = ~pi194 & n6024;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = ~n6012 & n6027;
  assign n6029 = n6012 & ~n6027;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = pi835 & n1761;
  assign n6032 = ~pi230 & n1787;
  assign n6033 = ~n6031 & ~n6032;
  assign n6034 = ~n1754 & ~n6033;
  assign n6035 = pi835 & n1756;
  assign n6036 = ~pi230 & ~n1756;
  assign n6037 = ~n6035 & ~n6036;
  assign n6038 = ~n1792 & ~n6037;
  assign n6039 = ~n6034 & ~n6038;
  assign n6040 = ~n6030 & ~n6039;
  assign n6041 = n6030 & n6039;
  assign n6042 = ~n6040 & ~n6041;
  assign n6043 = n2685 & n6042;
  assign n6044 = ~n2685 & ~n6042;
  assign n6045 = ~n6043 & ~n6044;
  assign n6046 = po814 & ~n6045;
  assign po360 = n6000 | n6046;
  assign n6048 = pi212 & ~po814;
  assign n6049 = pi296 & n1778;
  assign n6050 = pi889 & n1756;
  assign n6051 = pi296 & ~n1756;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = ~n1778 & ~n6052;
  assign n6054 = ~n6049 & ~n6053;
  assign n6055 = ~n1761 & ~n6054;
  assign n6056 = pi889 & n1761;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n1754 & ~n6057;
  assign n6059 = n1754 & ~n6052;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = pi921 & n1761;
  assign n6062 = pi921 & n1756;
  assign n6063 = pi419 & ~n1756;
  assign n6064 = ~n6062 & ~n6063;
  assign n6065 = ~n1778 & ~n6064;
  assign n6066 = pi419 & n1778;
  assign n6067 = ~n6065 & ~n6066;
  assign n6068 = ~n1761 & ~n6067;
  assign n6069 = ~n6061 & ~n6068;
  assign n6070 = ~n1754 & ~n6069;
  assign n6071 = n1754 & ~n6064;
  assign n6072 = ~n6070 & ~n6071;
  assign n6073 = pi137 & ~n6072;
  assign n6074 = ~pi137 & n6072;
  assign n6075 = ~n6073 & ~n6074;
  assign n6076 = ~n6060 & n6075;
  assign n6077 = n6060 & ~n6075;
  assign n6078 = ~n6076 & ~n6077;
  assign n6079 = pi857 & n1761;
  assign n6080 = ~pi236 & n1787;
  assign n6081 = ~n6079 & ~n6080;
  assign n6082 = ~n1754 & ~n6081;
  assign n6083 = pi857 & n1756;
  assign n6084 = ~pi236 & ~n1756;
  assign n6085 = ~n6083 & ~n6084;
  assign n6086 = ~n1792 & ~n6085;
  assign n6087 = ~n6082 & ~n6086;
  assign n6088 = ~n6078 & ~n6087;
  assign n6089 = n6078 & n6087;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = n2880 & n6090;
  assign n6092 = ~n2880 & ~n6090;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = po814 & ~n6093;
  assign po361 = n6048 | n6094;
  assign n6096 = pi213 & ~po814;
  assign n6097 = pi841 & n1761;
  assign n6098 = pi841 & n1756;
  assign n6099 = ~pi235 & ~n1756;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n1778 & ~n6100;
  assign n6102 = ~pi235 & n1778;
  assign n6103 = ~n6101 & ~n6102;
  assign n6104 = ~n1761 & ~n6103;
  assign n6105 = ~n6097 & ~n6104;
  assign n6106 = ~n1754 & ~n6105;
  assign n6107 = n1754 & ~n6100;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = pi905 & n1761;
  assign n6110 = pi905 & n1756;
  assign n6111 = pi418 & ~n1756;
  assign n6112 = ~n6110 & ~n6111;
  assign n6113 = ~n1778 & ~n6112;
  assign n6114 = pi418 & n1778;
  assign n6115 = ~n6113 & ~n6114;
  assign n6116 = ~n1761 & ~n6115;
  assign n6117 = ~n6109 & ~n6116;
  assign n6118 = ~n1754 & ~n6117;
  assign n6119 = n1754 & ~n6112;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121 = pi159 & ~n6120;
  assign n6122 = ~pi159 & n6120;
  assign n6123 = ~n6121 & ~n6122;
  assign n6124 = pi873 & n1761;
  assign n6125 = pi295 & n1787;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = ~n1754 & ~n6126;
  assign n6128 = pi873 & n1756;
  assign n6129 = pi295 & ~n1756;
  assign n6130 = ~n6128 & ~n6129;
  assign n6131 = ~n1792 & ~n6130;
  assign n6132 = ~n6127 & ~n6131;
  assign n6133 = ~n6123 & n6132;
  assign n6134 = n6123 & ~n6132;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = n6108 & n6135;
  assign n6137 = ~n6108 & ~n6135;
  assign n6138 = ~n6136 & ~n6137;
  assign n6139 = n2893 & n6138;
  assign n6140 = ~n2893 & ~n6138;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = po814 & ~n6141;
  assign po362 = n6096 | n6142;
  assign n6144 = ~pi214 & ~po814;
  assign n6145 = po814 & ~n5451;
  assign po363 = n6144 | n6145;
  assign n6147 = ~pi215 & ~po814;
  assign n6148 = po814 & ~n5401;
  assign po364 = n6147 | n6148;
  assign n6150 = pi216 & ~po814;
  assign n6151 = pi298 & n1778;
  assign n6152 = pi883 & n1756;
  assign n6153 = pi298 & ~n1756;
  assign n6154 = ~n6152 & ~n6153;
  assign n6155 = ~n1778 & ~n6154;
  assign n6156 = ~n6151 & ~n6155;
  assign n6157 = ~n1761 & ~n6156;
  assign n6158 = pi883 & n1761;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = ~n1754 & ~n6159;
  assign n6161 = n1754 & ~n6154;
  assign n6162 = ~n6160 & ~n6161;
  assign n6163 = pi915 & n1761;
  assign n6164 = pi915 & n1756;
  assign n6165 = pi421 & ~n1756;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = ~n1778 & ~n6166;
  assign n6168 = pi421 & n1778;
  assign n6169 = ~n6167 & ~n6168;
  assign n6170 = ~n1761 & ~n6169;
  assign n6171 = ~n6163 & ~n6170;
  assign n6172 = ~n1754 & ~n6171;
  assign n6173 = n1754 & ~n6166;
  assign n6174 = ~n6172 & ~n6173;
  assign n6175 = pi191 & ~n6174;
  assign n6176 = ~pi191 & n6174;
  assign n6177 = ~n6175 & ~n6176;
  assign n6178 = ~n6162 & n6177;
  assign n6179 = n6162 & ~n6177;
  assign n6180 = ~n6178 & ~n6179;
  assign n6181 = pi851 & n1761;
  assign n6182 = ~pi240 & n1787;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = ~n1754 & ~n6183;
  assign n6185 = pi851 & n1756;
  assign n6186 = ~pi240 & ~n1756;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = ~n1792 & ~n6187;
  assign n6189 = ~n6184 & ~n6188;
  assign n6190 = ~n6180 & ~n6189;
  assign n6191 = n6180 & n6189;
  assign n6192 = ~n6190 & ~n6191;
  assign n6193 = n2698 & n6192;
  assign n6194 = ~n2698 & ~n6192;
  assign n6195 = ~n6193 & ~n6194;
  assign n6196 = po814 & ~n6195;
  assign po365 = n6150 | n6196;
  assign n6198 = pi217 & ~po814;
  assign n6199 = pi334 & n1778;
  assign n6200 = pi882 & n1756;
  assign n6201 = pi334 & ~n1756;
  assign n6202 = ~n6200 & ~n6201;
  assign n6203 = ~n1778 & ~n6202;
  assign n6204 = ~n6199 & ~n6203;
  assign n6205 = ~n1761 & ~n6204;
  assign n6206 = pi882 & n1761;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = ~n1754 & ~n6207;
  assign n6209 = n1754 & ~n6202;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = pi914 & n1761;
  assign n6212 = pi914 & n1756;
  assign n6213 = pi430 & ~n1756;
  assign n6214 = ~n6212 & ~n6213;
  assign n6215 = ~n1778 & ~n6214;
  assign n6216 = pi430 & n1778;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = ~n1761 & ~n6217;
  assign n6219 = ~n6211 & ~n6218;
  assign n6220 = ~n1754 & ~n6219;
  assign n6221 = n1754 & ~n6214;
  assign n6222 = ~n6220 & ~n6221;
  assign n6223 = pi131 & ~n6222;
  assign n6224 = ~pi131 & n6222;
  assign n6225 = ~n6223 & ~n6224;
  assign n6226 = ~n6210 & n6225;
  assign n6227 = n6210 & ~n6225;
  assign n6228 = ~n6226 & ~n6227;
  assign n6229 = pi850 & n1761;
  assign n6230 = ~pi245 & n1787;
  assign n6231 = ~n6229 & ~n6230;
  assign n6232 = ~n1754 & ~n6231;
  assign n6233 = pi850 & n1756;
  assign n6234 = ~pi245 & ~n1756;
  assign n6235 = ~n6233 & ~n6234;
  assign n6236 = ~n1792 & ~n6235;
  assign n6237 = ~n6232 & ~n6236;
  assign n6238 = ~n6228 & ~n6237;
  assign n6239 = n6228 & n6237;
  assign n6240 = ~n6238 & ~n6239;
  assign n6241 = ~n3011 & n6240;
  assign n6242 = n3011 & ~n6240;
  assign n6243 = ~n6241 & ~n6242;
  assign n6244 = po814 & ~n6243;
  assign po366 = n6198 | n6244;
  assign n6246 = pi218 & ~po814;
  assign n6247 = pi335 & n1778;
  assign n6248 = pi885 & n1756;
  assign n6249 = pi335 & ~n1756;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n1778 & ~n6250;
  assign n6252 = ~n6247 & ~n6251;
  assign n6253 = ~n1761 & ~n6252;
  assign n6254 = pi885 & n1761;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n1754 & ~n6255;
  assign n6257 = n1754 & ~n6250;
  assign n6258 = ~n6256 & ~n6257;
  assign n6259 = pi917 & n1761;
  assign n6260 = pi917 & n1756;
  assign n6261 = pi431 & ~n1756;
  assign n6262 = ~n6260 & ~n6261;
  assign n6263 = ~n1778 & ~n6262;
  assign n6264 = pi431 & n1778;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = ~n1761 & ~n6265;
  assign n6267 = ~n6259 & ~n6266;
  assign n6268 = ~n1754 & ~n6267;
  assign n6269 = n1754 & ~n6262;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = pi138 & ~n6270;
  assign n6272 = ~pi138 & n6270;
  assign n6273 = ~n6271 & ~n6272;
  assign n6274 = ~n6258 & n6273;
  assign n6275 = n6258 & ~n6273;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = pi853 & n1761;
  assign n6278 = ~pi242 & n1787;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~n1754 & ~n6279;
  assign n6281 = pi853 & n1756;
  assign n6282 = ~pi242 & ~n1756;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~n1792 & ~n6283;
  assign n6285 = ~n6280 & ~n6284;
  assign n6286 = ~n6276 & ~n6285;
  assign n6287 = n6276 & n6285;
  assign n6288 = ~n6286 & ~n6287;
  assign n6289 = n3139 & n6288;
  assign n6290 = ~n3139 & ~n6288;
  assign n6291 = ~n6289 & ~n6290;
  assign n6292 = po814 & ~n6291;
  assign po367 = n6246 | n6292;
  assign n6294 = pi219 & ~po814;
  assign n6295 = pi338 & n1778;
  assign n6296 = pi884 & n1756;
  assign n6297 = pi338 & ~n1756;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = ~n1778 & ~n6298;
  assign n6300 = ~n6295 & ~n6299;
  assign n6301 = ~n1761 & ~n6300;
  assign n6302 = pi884 & n1761;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = ~n1754 & ~n6303;
  assign n6305 = n1754 & ~n6298;
  assign n6306 = ~n6304 & ~n6305;
  assign n6307 = pi916 & n1761;
  assign n6308 = pi916 & n1756;
  assign n6309 = pi433 & ~n1756;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~n1778 & ~n6310;
  assign n6312 = pi433 & n1778;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~n1761 & ~n6313;
  assign n6315 = ~n6307 & ~n6314;
  assign n6316 = ~n1754 & ~n6315;
  assign n6317 = n1754 & ~n6310;
  assign n6318 = ~n6316 & ~n6317;
  assign n6319 = pi177 & ~n6318;
  assign n6320 = ~pi177 & n6318;
  assign n6321 = ~n6319 & ~n6320;
  assign n6322 = ~n6306 & n6321;
  assign n6323 = n6306 & ~n6321;
  assign n6324 = ~n6322 & ~n6323;
  assign n6325 = pi852 & n1761;
  assign n6326 = ~pi241 & n1787;
  assign n6327 = ~n6325 & ~n6326;
  assign n6328 = ~n1754 & ~n6327;
  assign n6329 = pi852 & n1756;
  assign n6330 = ~pi241 & ~n1756;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = ~n1792 & ~n6331;
  assign n6333 = ~n6328 & ~n6332;
  assign n6334 = ~n6324 & ~n6333;
  assign n6335 = n6324 & n6333;
  assign n6336 = ~n6334 & ~n6335;
  assign n6337 = n3381 & n6336;
  assign n6338 = ~n3381 & ~n6336;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = po814 & ~n6339;
  assign po368 = n6294 | n6340;
  assign n6342 = pi220 & ~po814;
  assign n6343 = pi337 & n1778;
  assign n6344 = pi887 & n1756;
  assign n6345 = pi337 & ~n1756;
  assign n6346 = ~n6344 & ~n6345;
  assign n6347 = ~n1778 & ~n6346;
  assign n6348 = ~n6343 & ~n6347;
  assign n6349 = ~n1761 & ~n6348;
  assign n6350 = pi887 & n1761;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = ~n1754 & ~n6351;
  assign n6353 = n1754 & ~n6346;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = pi919 & n1761;
  assign n6356 = pi919 & n1756;
  assign n6357 = pi436 & ~n1756;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = ~n1778 & ~n6358;
  assign n6360 = pi436 & n1778;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n1761 & ~n6361;
  assign n6363 = ~n6355 & ~n6362;
  assign n6364 = ~n1754 & ~n6363;
  assign n6365 = n1754 & ~n6358;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = pi071 & ~n6366;
  assign n6368 = ~pi071 & n6366;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = ~n6354 & n6369;
  assign n6371 = n6354 & ~n6369;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = pi855 & n1761;
  assign n6374 = ~pi246 & n1787;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = ~n1754 & ~n6375;
  assign n6377 = pi855 & n1756;
  assign n6378 = ~pi246 & ~n1756;
  assign n6379 = ~n6377 & ~n6378;
  assign n6380 = ~n1792 & ~n6379;
  assign n6381 = ~n6376 & ~n6380;
  assign n6382 = ~n6372 & ~n6381;
  assign n6383 = n6372 & n6381;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = n3467 & n6384;
  assign n6386 = ~n3467 & ~n6384;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = po814 & ~n6387;
  assign po369 = n6342 | n6388;
  assign n6390 = pi221 & ~po814;
  assign n6391 = pi339 & n1778;
  assign n6392 = pi888 & n1756;
  assign n6393 = pi339 & ~n1756;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = ~n1778 & ~n6394;
  assign n6396 = ~n6391 & ~n6395;
  assign n6397 = ~n1761 & ~n6396;
  assign n6398 = pi888 & n1761;
  assign n6399 = ~n6397 & ~n6398;
  assign n6400 = ~n1754 & ~n6399;
  assign n6401 = n1754 & ~n6394;
  assign n6402 = ~n6400 & ~n6401;
  assign n6403 = pi920 & n1761;
  assign n6404 = pi920 & n1756;
  assign n6405 = pi434 & ~n1756;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = ~n1778 & ~n6406;
  assign n6408 = pi434 & n1778;
  assign n6409 = ~n6407 & ~n6408;
  assign n6410 = ~n1761 & ~n6409;
  assign n6411 = ~n6403 & ~n6410;
  assign n6412 = ~n1754 & ~n6411;
  assign n6413 = n1754 & ~n6406;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = pi072 & ~n6414;
  assign n6416 = ~pi072 & n6414;
  assign n6417 = ~n6415 & ~n6416;
  assign n6418 = ~n6402 & n6417;
  assign n6419 = n6402 & ~n6417;
  assign n6420 = ~n6418 & ~n6419;
  assign n6421 = pi856 & n1761;
  assign n6422 = ~pi244 & n1787;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = ~n1754 & ~n6423;
  assign n6425 = pi856 & n1756;
  assign n6426 = ~pi244 & ~n1756;
  assign n6427 = ~n6425 & ~n6426;
  assign n6428 = ~n1792 & ~n6427;
  assign n6429 = ~n6424 & ~n6428;
  assign n6430 = ~n6420 & ~n6429;
  assign n6431 = n6420 & n6429;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n2410 & n6432;
  assign n6434 = n2410 & ~n6432;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = po814 & ~n6435;
  assign po370 = n6390 | n6436;
  assign n6438 = pi222 & ~po814;
  assign n6439 = pi336 & n1778;
  assign n6440 = pi886 & n1756;
  assign n6441 = pi336 & ~n1756;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n1778 & ~n6442;
  assign n6444 = ~n6439 & ~n6443;
  assign n6445 = ~n1761 & ~n6444;
  assign n6446 = pi886 & n1761;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = ~n1754 & ~n6447;
  assign n6449 = n1754 & ~n6442;
  assign n6450 = ~n6448 & ~n6449;
  assign n6451 = pi918 & n1761;
  assign n6452 = pi918 & n1756;
  assign n6453 = pi432 & ~n1756;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n1778 & ~n6454;
  assign n6456 = pi432 & n1778;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 = ~n1761 & ~n6457;
  assign n6459 = ~n6451 & ~n6458;
  assign n6460 = ~n1754 & ~n6459;
  assign n6461 = n1754 & ~n6454;
  assign n6462 = ~n6460 & ~n6461;
  assign n6463 = pi135 & ~n6462;
  assign n6464 = ~pi135 & n6462;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n6450 & n6465;
  assign n6467 = n6450 & ~n6465;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = pi854 & n1761;
  assign n6470 = ~pi243 & n1787;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n1754 & ~n6471;
  assign n6473 = pi854 & n1756;
  assign n6474 = ~pi243 & ~n1756;
  assign n6475 = ~n6473 & ~n6474;
  assign n6476 = ~n1792 & ~n6475;
  assign n6477 = ~n6472 & ~n6476;
  assign n6478 = ~n6468 & ~n6477;
  assign n6479 = n6468 & n6477;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = n2841 & n6480;
  assign n6482 = ~n2841 & ~n6480;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = po814 & ~n6483;
  assign po371 = n6438 | n6484;
  assign n6486 = ~pi223 & ~po814;
  assign n6487 = po814 & ~n5650;
  assign po372 = n6486 | n6487;
  assign n6489 = ~pi224 & ~po814;
  assign n6490 = po814 & ~n5701;
  assign po373 = n6489 | n6490;
  assign n6492 = ~pi225 & ~po814;
  assign n6493 = po814 & ~n5599;
  assign po374 = n6492 | n6493;
  assign n6495 = ~pi226 & ~po814;
  assign n6496 = po814 & ~n5500;
  assign po375 = n6495 | n6496;
  assign n6498 = ~pi227 & ~po814;
  assign n6499 = po814 & ~n5550;
  assign po376 = n6498 | n6499;
  assign n6501 = ~pi228 & ~po814;
  assign n6502 = po814 & ~n5347;
  assign po377 = n6501 | n6502;
  assign n6504 = po814 & n5994;
  assign n6505 = ~pi229 & ~po814;
  assign po378 = n6504 | n6505;
  assign n6507 = po814 & n6042;
  assign n6508 = ~pi230 & ~po814;
  assign po379 = n6507 | n6508;
  assign n6510 = po814 & n5752;
  assign n6511 = ~pi231 & ~po814;
  assign po380 = n6510 | n6511;
  assign n6513 = po814 & n5802;
  assign n6514 = ~pi232 & ~po814;
  assign po381 = n6513 | n6514;
  assign n6516 = po814 & n5850;
  assign n6517 = ~pi233 & ~po814;
  assign po382 = n6516 | n6517;
  assign n6519 = po814 & n5946;
  assign n6520 = ~pi234 & ~po814;
  assign po383 = n6519 | n6520;
  assign n6522 = po814 & n6138;
  assign n6523 = ~pi235 & ~po814;
  assign po384 = n6522 | n6523;
  assign n6525 = po814 & n6090;
  assign n6526 = ~pi236 & ~po814;
  assign po385 = n6525 | n6526;
  assign n6528 = po814 & n5898;
  assign n6529 = ~pi237 & ~po814;
  assign po386 = n6528 | n6529;
  assign n6531 = pi238 & ~po814;
  assign n6532 = po814 & ~n5398;
  assign po387 = n6531 | n6532;
  assign n6534 = po814 & n5448;
  assign n6535 = ~pi239 & ~po814;
  assign po388 = n6534 | n6535;
  assign n6537 = po814 & n6192;
  assign n6538 = ~pi240 & ~po814;
  assign po389 = n6537 | n6538;
  assign n6540 = po814 & n6336;
  assign n6541 = ~pi241 & ~po814;
  assign po390 = n6540 | n6541;
  assign n6543 = po814 & n6288;
  assign n6544 = ~pi242 & ~po814;
  assign po391 = n6543 | n6544;
  assign n6546 = po814 & n6480;
  assign n6547 = ~pi243 & ~po814;
  assign po392 = n6546 | n6547;
  assign n6549 = po814 & n6432;
  assign n6550 = ~pi244 & ~po814;
  assign po393 = n6549 | n6550;
  assign n6552 = po814 & n6240;
  assign n6553 = ~pi245 & ~po814;
  assign po394 = n6552 | n6553;
  assign n6555 = po814 & n6384;
  assign n6556 = ~pi246 & ~po814;
  assign po395 = n6555 | n6556;
  assign n6558 = po814 & n5698;
  assign n6559 = ~pi247 & ~po814;
  assign po396 = n6558 | n6559;
  assign n6561 = pi248 & ~po814;
  assign n6562 = po814 & ~n5547;
  assign po397 = n6561 | n6562;
  assign n6564 = pi249 & ~po814;
  assign n6565 = po814 & ~n5497;
  assign po398 = n6564 | n6565;
  assign n6567 = pi250 & ~po814;
  assign n6568 = po814 & ~n5596;
  assign po399 = n6567 | n6568;
  assign n6570 = pi251 & ~po814;
  assign n6571 = po814 & ~n5647;
  assign po400 = n6570 | n6571;
  assign n6573 = pi252 & ~po814;
  assign n6574 = po814 & ~n5895;
  assign po401 = n6573 | n6574;
  assign n6576 = pi253 & n1761;
  assign n6577 = pi665 & n1777;
  assign n6578 = ~n1778 & n6577;
  assign n6579 = ~pi673 & ~n1753;
  assign n6580 = pi734 & ~n6579;
  assign n6581 = pi656 & n6579;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n2449 & ~n6582;
  assign n6584 = pi126 & n2449;
  assign n6585 = ~n6583 & ~n6584;
  assign n6586 = pi562 & n6585;
  assign n6587 = ~pi556 & pi557;
  assign n6588 = pi558 & ~pi673;
  assign n6589 = ~pi555 & n6588;
  assign n6590 = n6587 & n6589;
  assign n6591 = ~n2562 & ~n6590;
  assign n6592 = pi666 & ~pi673;
  assign n6593 = pi656 & n6592;
  assign n6594 = ~pi669 & pi673;
  assign n6595 = pi126 & n6594;
  assign n6596 = ~n6585 & ~n6594;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~n6592 & ~n6597;
  assign n6599 = ~n6593 & ~n6598;
  assign n6600 = n6591 & ~n6599;
  assign n6601 = pi126 & ~pi669;
  assign n6602 = ~n6591 & n6601;
  assign n6603 = pi669 & ~n6591;
  assign n6604 = ~n6599 & n6603;
  assign n6605 = ~n6602 & ~n6604;
  assign n6606 = ~n6600 & n6605;
  assign n6607 = n2564 & ~n6606;
  assign n6608 = pi126 & ~n2564;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = ~pi562 & n6609;
  assign n6611 = ~n6586 & ~n6610;
  assign n6612 = ~pi204 & n6611;
  assign n6613 = pi204 & ~n6611;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = n6578 & n6614;
  assign n6616 = pi253 & ~n6578;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n1761 & ~n6617;
  assign n6619 = ~n6576 & ~n6618;
  assign n6620 = ~n1754 & ~n6619;
  assign n6621 = pi862 & n6611;
  assign n6622 = ~pi862 & ~n6611;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = n1754 & n6623;
  assign po402 = n6620 | n6624;
  assign n6626 = pi254 & n1761;
  assign n6627 = pi785 & ~n6579;
  assign n6628 = pi649 & n6579;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = ~n2449 & ~n6629;
  assign n6631 = pi075 & n2449;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = pi562 & n6632;
  assign n6634 = pi649 & n6592;
  assign n6635 = pi075 & n6594;
  assign n6636 = ~n6594 & ~n6632;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = ~n6592 & ~n6637;
  assign n6639 = ~n6634 & ~n6638;
  assign n6640 = n6591 & ~n6639;
  assign n6641 = pi075 & ~pi669;
  assign n6642 = ~n6591 & n6641;
  assign n6643 = n6603 & ~n6639;
  assign n6644 = ~n6642 & ~n6643;
  assign n6645 = ~n6640 & n6644;
  assign n6646 = n2564 & ~n6645;
  assign n6647 = pi075 & ~n2564;
  assign n6648 = ~n6646 & ~n6647;
  assign n6649 = ~pi562 & n6648;
  assign n6650 = ~n6633 & ~n6649;
  assign n6651 = ~pi155 & n6650;
  assign n6652 = pi155 & ~n6650;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = n6578 & n6653;
  assign n6655 = pi254 & ~n6578;
  assign n6656 = ~n6654 & ~n6655;
  assign n6657 = ~n1761 & ~n6656;
  assign n6658 = ~n6626 & ~n6657;
  assign n6659 = ~n1754 & ~n6658;
  assign n6660 = pi913 & n6650;
  assign n6661 = ~pi913 & ~n6650;
  assign n6662 = ~n6660 & ~n6661;
  assign n6663 = n1754 & n6662;
  assign po403 = n6659 | n6663;
  assign n6665 = pi255 & n1761;
  assign n6666 = pi737 & ~n6579;
  assign n6667 = pi646 & n6579;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = ~n2449 & ~n6668;
  assign n6670 = pi127 & n2449;
  assign n6671 = ~n6669 & ~n6670;
  assign n6672 = pi562 & n6671;
  assign n6673 = pi646 & n6592;
  assign n6674 = pi127 & n6594;
  assign n6675 = ~n6594 & ~n6671;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = ~n6592 & ~n6676;
  assign n6678 = ~n6673 & ~n6677;
  assign n6679 = n6591 & ~n6678;
  assign n6680 = pi127 & ~pi669;
  assign n6681 = ~n6591 & n6680;
  assign n6682 = n6603 & ~n6678;
  assign n6683 = ~n6681 & ~n6682;
  assign n6684 = ~n6679 & n6683;
  assign n6685 = n2564 & ~n6684;
  assign n6686 = pi127 & ~n2564;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~pi562 & n6687;
  assign n6689 = ~n6672 & ~n6688;
  assign n6690 = ~pi225 & n6689;
  assign n6691 = pi225 & ~n6689;
  assign n6692 = ~n6690 & ~n6691;
  assign n6693 = n6578 & n6692;
  assign n6694 = pi255 & ~n6578;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n1761 & ~n6695;
  assign n6697 = ~n6665 & ~n6696;
  assign n6698 = ~n1754 & ~n6697;
  assign n6699 = pi865 & n6689;
  assign n6700 = ~pi865 & ~n6689;
  assign n6701 = ~n6699 & ~n6700;
  assign n6702 = n1754 & n6701;
  assign po404 = n6698 | n6702;
  assign n6704 = pi256 & n1761;
  assign n6705 = pi680 & ~n6579;
  assign n6706 = pi538 & n6579;
  assign n6707 = ~n6705 & ~n6706;
  assign n6708 = ~n2449 & ~n6707;
  assign n6709 = pi037 & n2449;
  assign n6710 = ~n6708 & ~n6709;
  assign n6711 = pi562 & n6710;
  assign n6712 = pi538 & n6592;
  assign n6713 = pi037 & n6594;
  assign n6714 = ~n6594 & ~n6710;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = ~n6592 & ~n6715;
  assign n6717 = ~n6712 & ~n6716;
  assign n6718 = n6591 & ~n6717;
  assign n6719 = pi037 & ~pi669;
  assign n6720 = ~n6591 & n6719;
  assign n6721 = n6603 & ~n6717;
  assign n6722 = ~n6720 & ~n6721;
  assign n6723 = ~n6718 & n6722;
  assign n6724 = n2564 & ~n6723;
  assign n6725 = pi037 & ~n2564;
  assign n6726 = ~n6724 & ~n6725;
  assign n6727 = ~pi562 & n6726;
  assign n6728 = ~n6711 & ~n6727;
  assign n6729 = pi209 & n6728;
  assign n6730 = ~pi209 & ~n6728;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = n6578 & n6731;
  assign n6733 = pi256 & ~n6578;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = ~n1761 & ~n6734;
  assign n6736 = ~n6704 & ~n6735;
  assign n6737 = ~n1754 & ~n6736;
  assign n6738 = pi808 & n6728;
  assign n6739 = ~pi808 & ~n6728;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = n1754 & n6740;
  assign po405 = n6737 | n6741;
  assign n6743 = pi257 & n1761;
  assign n6744 = pi750 & ~n6579;
  assign n6745 = pi608 & n6579;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = ~n2449 & ~n6746;
  assign n6748 = pi083 & n2449;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = pi562 & n6749;
  assign n6751 = pi608 & n6592;
  assign n6752 = pi083 & n6594;
  assign n6753 = ~n6594 & ~n6749;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = ~n6592 & ~n6754;
  assign n6756 = ~n6751 & ~n6755;
  assign n6757 = n6591 & ~n6756;
  assign n6758 = pi083 & ~pi669;
  assign n6759 = ~n6591 & n6758;
  assign n6760 = n6603 & ~n6756;
  assign n6761 = ~n6759 & ~n6760;
  assign n6762 = ~n6757 & n6761;
  assign n6763 = n2564 & ~n6762;
  assign n6764 = pi083 & ~n2564;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = ~pi562 & n6765;
  assign n6767 = ~n6750 & ~n6766;
  assign n6768 = pi044 & n6767;
  assign n6769 = ~pi044 & ~n6767;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = n6578 & n6770;
  assign n6772 = pi257 & ~n6578;
  assign n6773 = ~n6771 & ~n6772;
  assign n6774 = ~n1761 & ~n6773;
  assign n6775 = ~n6743 & ~n6774;
  assign n6776 = ~n1754 & ~n6775;
  assign n6777 = pi878 & n6767;
  assign n6778 = ~pi878 & ~n6767;
  assign n6779 = ~n6777 & ~n6778;
  assign n6780 = n1754 & n6779;
  assign po406 = n6776 | n6780;
  assign n6782 = pi258 & n1761;
  assign n6783 = pi699 & ~n6579;
  assign n6784 = pi521 & n6579;
  assign n6785 = ~n6783 & ~n6784;
  assign n6786 = ~n2449 & ~n6785;
  assign n6787 = ~pi185 & n2449;
  assign n6788 = ~n6786 & ~n6787;
  assign n6789 = pi562 & n6788;
  assign n6790 = pi521 & n6592;
  assign n6791 = ~pi185 & n6594;
  assign n6792 = ~n6594 & ~n6788;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~n6592 & ~n6793;
  assign n6795 = ~n6790 & ~n6794;
  assign n6796 = n6591 & ~n6795;
  assign n6797 = ~pi185 & ~pi669;
  assign n6798 = ~n6591 & n6797;
  assign n6799 = n6603 & ~n6795;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = ~n6796 & n6800;
  assign n6802 = n2564 & ~n6801;
  assign n6803 = ~pi185 & ~n2564;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = ~pi562 & n6804;
  assign n6806 = ~n6789 & ~n6805;
  assign n6807 = pi202 & n6806;
  assign n6808 = ~pi202 & ~n6806;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = n6578 & n6809;
  assign n6811 = pi258 & ~n6578;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n1761 & ~n6812;
  assign n6814 = ~n6782 & ~n6813;
  assign n6815 = ~n1754 & ~n6814;
  assign n6816 = pi827 & n6806;
  assign n6817 = ~pi827 & ~n6806;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = n1754 & n6818;
  assign po407 = n6815 | n6819;
  assign n6821 = pi259 & n1761;
  assign n6822 = pi751 & ~n6579;
  assign n6823 = pi592 & n6579;
  assign n6824 = ~n6822 & ~n6823;
  assign n6825 = ~n2449 & ~n6824;
  assign n6826 = pi024 & n2449;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828 = pi562 & n6827;
  assign n6829 = pi592 & n6592;
  assign n6830 = pi024 & n6594;
  assign n6831 = ~n6594 & ~n6827;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = ~n6592 & ~n6832;
  assign n6834 = ~n6829 & ~n6833;
  assign n6835 = n6591 & ~n6834;
  assign n6836 = pi024 & ~pi669;
  assign n6837 = ~n6591 & n6836;
  assign n6838 = n6603 & ~n6834;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = ~n6835 & n6839;
  assign n6841 = n2564 & ~n6840;
  assign n6842 = pi024 & ~n2564;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = ~pi562 & n6843;
  assign n6845 = ~n6828 & ~n6844;
  assign n6846 = pi048 & n6845;
  assign n6847 = ~pi048 & ~n6845;
  assign n6848 = ~n6846 & ~n6847;
  assign n6849 = n6578 & n6848;
  assign n6850 = pi259 & ~n6578;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = ~n1761 & ~n6851;
  assign n6853 = ~n6821 & ~n6852;
  assign n6854 = ~n1754 & ~n6853;
  assign n6855 = pi879 & n6845;
  assign n6856 = ~pi879 & ~n6845;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = n1754 & n6857;
  assign po408 = n6854 | n6858;
  assign n6860 = pi260 & n1761;
  assign n6861 = pi752 & ~n6579;
  assign n6862 = pi593 & n6579;
  assign n6863 = ~n6861 & ~n6862;
  assign n6864 = ~n2449 & ~n6863;
  assign n6865 = pi025 & n2449;
  assign n6866 = ~n6864 & ~n6865;
  assign n6867 = pi562 & n6866;
  assign n6868 = pi593 & n6592;
  assign n6869 = pi025 & n6594;
  assign n6870 = ~n6594 & ~n6866;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = ~n6592 & ~n6871;
  assign n6873 = ~n6868 & ~n6872;
  assign n6874 = n6591 & ~n6873;
  assign n6875 = pi025 & ~pi669;
  assign n6876 = ~n6591 & n6875;
  assign n6877 = n6603 & ~n6873;
  assign n6878 = ~n6876 & ~n6877;
  assign n6879 = ~n6874 & n6878;
  assign n6880 = n2564 & ~n6879;
  assign n6881 = pi025 & ~n2564;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ~pi562 & n6882;
  assign n6884 = ~n6867 & ~n6883;
  assign n6885 = pi049 & n6884;
  assign n6886 = ~pi049 & ~n6884;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888 = n6578 & n6887;
  assign n6889 = pi260 & ~n6578;
  assign n6890 = ~n6888 & ~n6889;
  assign n6891 = ~n1761 & ~n6890;
  assign n6892 = ~n6860 & ~n6891;
  assign n6893 = ~n1754 & ~n6892;
  assign n6894 = pi880 & n6884;
  assign n6895 = ~pi880 & ~n6884;
  assign n6896 = ~n6894 & ~n6895;
  assign n6897 = n1754 & n6896;
  assign po409 = n6893 | n6897;
  assign n6899 = pi261 & n1761;
  assign n6900 = pi753 & ~n6579;
  assign n6901 = pi662 & n6579;
  assign n6902 = ~n6900 & ~n6901;
  assign n6903 = ~n2449 & ~n6902;
  assign n6904 = pi084 & n2449;
  assign n6905 = ~n6903 & ~n6904;
  assign n6906 = pi562 & n6905;
  assign n6907 = pi662 & n6592;
  assign n6908 = pi084 & n6594;
  assign n6909 = ~n6594 & ~n6905;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6592 & ~n6910;
  assign n6912 = ~n6907 & ~n6911;
  assign n6913 = n6591 & ~n6912;
  assign n6914 = pi084 & ~pi669;
  assign n6915 = ~n6591 & n6914;
  assign n6916 = n6603 & ~n6912;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = ~n6913 & n6917;
  assign n6919 = n2564 & ~n6918;
  assign n6920 = pi084 & ~n2564;
  assign n6921 = ~n6919 & ~n6920;
  assign n6922 = ~pi562 & n6921;
  assign n6923 = ~n6906 & ~n6922;
  assign n6924 = pi057 & n6923;
  assign n6925 = ~pi057 & ~n6923;
  assign n6926 = ~n6924 & ~n6925;
  assign n6927 = n6578 & n6926;
  assign n6928 = pi261 & ~n6578;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = ~n1761 & ~n6929;
  assign n6931 = ~n6899 & ~n6930;
  assign n6932 = ~n1754 & ~n6931;
  assign n6933 = pi881 & n6923;
  assign n6934 = ~pi881 & ~n6923;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = n1754 & n6935;
  assign po410 = n6932 | n6936;
  assign n6938 = pi262 & n1761;
  assign n6939 = pi700 & ~n6579;
  assign n6940 = pi522 & n6579;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = ~n2449 & ~n6941;
  assign n6943 = pi161 & n2449;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = pi562 & n6944;
  assign n6946 = pi522 & n6592;
  assign n6947 = pi161 & n6594;
  assign n6948 = ~n6594 & ~n6944;
  assign n6949 = ~n6947 & ~n6948;
  assign n6950 = ~n6592 & ~n6949;
  assign n6951 = ~n6946 & ~n6950;
  assign n6952 = n6591 & ~n6951;
  assign n6953 = pi161 & ~pi669;
  assign n6954 = ~n6591 & n6953;
  assign n6955 = n6603 & ~n6951;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6952 & n6956;
  assign n6958 = n2564 & ~n6957;
  assign n6959 = pi161 & ~n2564;
  assign n6960 = ~n6958 & ~n6959;
  assign n6961 = ~pi562 & n6960;
  assign n6962 = ~n6945 & ~n6961;
  assign n6963 = pi203 & n6962;
  assign n6964 = ~pi203 & ~n6962;
  assign n6965 = ~n6963 & ~n6964;
  assign n6966 = n6578 & n6965;
  assign n6967 = pi262 & ~n6578;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = ~n1761 & ~n6968;
  assign n6970 = ~n6938 & ~n6969;
  assign n6971 = ~n1754 & ~n6970;
  assign n6972 = pi828 & n6962;
  assign n6973 = ~pi828 & ~n6962;
  assign n6974 = ~n6972 & ~n6973;
  assign n6975 = n1754 & n6974;
  assign po411 = n6971 | n6975;
  assign n6977 = pi263 & n1761;
  assign n6978 = pi703 & ~n6579;
  assign n6979 = pi543 & n6579;
  assign n6980 = ~n6978 & ~n6979;
  assign n6981 = ~n2449 & ~n6980;
  assign n6982 = pi052 & n2449;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = pi562 & n6983;
  assign n6985 = pi543 & n6592;
  assign n6986 = pi052 & n6594;
  assign n6987 = ~n6594 & ~n6983;
  assign n6988 = ~n6986 & ~n6987;
  assign n6989 = ~n6592 & ~n6988;
  assign n6990 = ~n6985 & ~n6989;
  assign n6991 = n6591 & ~n6990;
  assign n6992 = pi052 & ~pi669;
  assign n6993 = ~n6591 & n6992;
  assign n6994 = n6603 & ~n6990;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = ~n6991 & n6995;
  assign n6997 = n2564 & ~n6996;
  assign n6998 = pi052 & ~n2564;
  assign n6999 = ~n6997 & ~n6998;
  assign n7000 = ~pi562 & n6999;
  assign n7001 = ~n6984 & ~n7000;
  assign n7002 = pi198 & n7001;
  assign n7003 = ~pi198 & ~n7001;
  assign n7004 = ~n7002 & ~n7003;
  assign n7005 = n6578 & n7004;
  assign n7006 = pi263 & ~n6578;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 = ~n1761 & ~n7007;
  assign n7009 = ~n6977 & ~n7008;
  assign n7010 = ~n1754 & ~n7009;
  assign n7011 = pi831 & n7001;
  assign n7012 = ~pi831 & ~n7001;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = n1754 & n7013;
  assign po412 = n7010 | n7014;
  assign n7016 = pi264 & n1761;
  assign n7017 = pi682 & ~n6579;
  assign n7018 = pi527 & n6579;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = ~n2449 & ~n7019;
  assign n7021 = pi061 & n2449;
  assign n7022 = ~n7020 & ~n7021;
  assign n7023 = pi562 & n7022;
  assign n7024 = pi527 & n6592;
  assign n7025 = pi061 & n6594;
  assign n7026 = ~n6594 & ~n7022;
  assign n7027 = ~n7025 & ~n7026;
  assign n7028 = ~n6592 & ~n7027;
  assign n7029 = ~n7024 & ~n7028;
  assign n7030 = n6591 & ~n7029;
  assign n7031 = pi061 & ~pi669;
  assign n7032 = ~n6591 & n7031;
  assign n7033 = n6603 & ~n7029;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = ~n7030 & n7034;
  assign n7036 = n2564 & ~n7035;
  assign n7037 = pi061 & ~n2564;
  assign n7038 = ~n7036 & ~n7037;
  assign n7039 = ~pi562 & n7038;
  assign n7040 = ~n7023 & ~n7039;
  assign n7041 = pi009 & n7040;
  assign n7042 = ~pi009 & ~n7040;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = n6578 & n7043;
  assign n7045 = pi264 & ~n6578;
  assign n7046 = ~n7044 & ~n7045;
  assign n7047 = ~n1761 & ~n7046;
  assign n7048 = ~n7016 & ~n7047;
  assign n7049 = ~n1754 & ~n7048;
  assign n7050 = pi810 & n7040;
  assign n7051 = ~pi810 & ~n7040;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = n1754 & n7052;
  assign po413 = n7049 | n7053;
  assign n7055 = pi265 & n1761;
  assign n7056 = pi779 & ~n6579;
  assign n7057 = pi571 & n6579;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = ~n2449 & ~n7058;
  assign n7060 = pi168 & n2449;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = pi562 & n7061;
  assign n7063 = pi571 & n6592;
  assign n7064 = pi168 & n6594;
  assign n7065 = ~n6594 & ~n7061;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = ~n6592 & ~n7066;
  assign n7068 = ~n7063 & ~n7067;
  assign n7069 = n6591 & ~n7068;
  assign n7070 = pi168 & ~pi669;
  assign n7071 = ~n6591 & n7070;
  assign n7072 = n6603 & ~n7068;
  assign n7073 = ~n7071 & ~n7072;
  assign n7074 = ~n7069 & n7073;
  assign n7075 = n2564 & ~n7074;
  assign n7076 = pi168 & ~n2564;
  assign n7077 = ~n7075 & ~n7076;
  assign n7078 = ~pi562 & n7077;
  assign n7079 = ~n7062 & ~n7078;
  assign n7080 = ~pi176 & n7079;
  assign n7081 = pi176 & ~n7079;
  assign n7082 = ~n7080 & ~n7081;
  assign n7083 = n6578 & n7082;
  assign n7084 = pi265 & ~n6578;
  assign n7085 = ~n7083 & ~n7084;
  assign n7086 = ~n1761 & ~n7085;
  assign n7087 = ~n7055 & ~n7086;
  assign n7088 = ~n1754 & ~n7087;
  assign n7089 = pi907 & n7079;
  assign n7090 = ~pi907 & ~n7079;
  assign n7091 = ~n7089 & ~n7090;
  assign n7092 = n1754 & n7091;
  assign po414 = n7088 | n7092;
  assign n7094 = pi266 & n1761;
  assign n7095 = pi674 & ~n6579;
  assign n7096 = pi540 & n6579;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~n2449 & ~n7097;
  assign n7099 = ~pi062 & n2449;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = pi562 & n7100;
  assign n7102 = pi540 & n6592;
  assign n7103 = ~pi062 & n6594;
  assign n7104 = ~n6594 & ~n7100;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = ~n6592 & ~n7105;
  assign n7107 = ~n7102 & ~n7106;
  assign n7108 = n6591 & ~n7107;
  assign n7109 = ~pi062 & ~pi669;
  assign n7110 = ~n6591 & n7109;
  assign n7111 = n6603 & ~n7107;
  assign n7112 = ~n7110 & ~n7111;
  assign n7113 = ~n7108 & n7112;
  assign n7114 = n2564 & ~n7113;
  assign n7115 = ~pi062 & ~n2564;
  assign n7116 = ~n7114 & ~n7115;
  assign n7117 = ~pi562 & n7116;
  assign n7118 = ~n7101 & ~n7117;
  assign n7119 = pi210 & n7118;
  assign n7120 = ~pi210 & ~n7118;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = n6578 & n7121;
  assign n7123 = pi266 & ~n6578;
  assign n7124 = ~n7122 & ~n7123;
  assign n7125 = ~n1761 & ~n7124;
  assign n7126 = ~n7094 & ~n7125;
  assign n7127 = ~n1754 & ~n7126;
  assign n7128 = pi802 & n7118;
  assign n7129 = ~pi802 & ~n7118;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = n1754 & n7130;
  assign po415 = n7127 | n7131;
  assign n7133 = pi267 & n1761;
  assign n7134 = pi780 & ~n6579;
  assign n7135 = pi591 & n6579;
  assign n7136 = ~n7134 & ~n7135;
  assign n7137 = ~n2449 & ~n7136;
  assign n7138 = pi139 & n2449;
  assign n7139 = ~n7137 & ~n7138;
  assign n7140 = pi562 & n7139;
  assign n7141 = pi591 & n6592;
  assign n7142 = pi139 & n6594;
  assign n7143 = ~n6594 & ~n7139;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = ~n6592 & ~n7144;
  assign n7146 = ~n7141 & ~n7145;
  assign n7147 = n6591 & ~n7146;
  assign n7148 = pi139 & ~pi669;
  assign n7149 = ~n6591 & n7148;
  assign n7150 = n6603 & ~n7146;
  assign n7151 = ~n7149 & ~n7150;
  assign n7152 = ~n7147 & n7151;
  assign n7153 = n2564 & ~n7152;
  assign n7154 = pi139 & ~n2564;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = ~pi562 & n7155;
  assign n7157 = ~n7140 & ~n7156;
  assign n7158 = ~pi188 & n7157;
  assign n7159 = pi188 & ~n7157;
  assign n7160 = ~n7158 & ~n7159;
  assign n7161 = n6578 & n7160;
  assign n7162 = pi267 & ~n6578;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = ~n1761 & ~n7163;
  assign n7165 = ~n7133 & ~n7164;
  assign n7166 = ~n1754 & ~n7165;
  assign n7167 = pi908 & n7157;
  assign n7168 = ~pi908 & ~n7157;
  assign n7169 = ~n7167 & ~n7168;
  assign n7170 = n1754 & n7169;
  assign po416 = n7166 | n7170;
  assign n7172 = pi268 & n1761;
  assign n7173 = pi781 & ~n6579;
  assign n7174 = pi636 & n6579;
  assign n7175 = ~n7173 & ~n7174;
  assign n7176 = ~n2449 & ~n7175;
  assign n7177 = pi073 & n2449;
  assign n7178 = ~n7176 & ~n7177;
  assign n7179 = pi562 & n7178;
  assign n7180 = pi636 & n6592;
  assign n7181 = pi073 & n6594;
  assign n7182 = ~n6594 & ~n7178;
  assign n7183 = ~n7181 & ~n7182;
  assign n7184 = ~n6592 & ~n7183;
  assign n7185 = ~n7180 & ~n7184;
  assign n7186 = n6591 & ~n7185;
  assign n7187 = pi073 & ~pi669;
  assign n7188 = ~n6591 & n7187;
  assign n7189 = n6603 & ~n7185;
  assign n7190 = ~n7188 & ~n7189;
  assign n7191 = ~n7186 & n7190;
  assign n7192 = n2564 & ~n7191;
  assign n7193 = pi073 & ~n2564;
  assign n7194 = ~n7192 & ~n7193;
  assign n7195 = ~pi562 & n7194;
  assign n7196 = ~n7179 & ~n7195;
  assign n7197 = ~pi133 & n7196;
  assign n7198 = pi133 & ~n7196;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = n6578 & n7199;
  assign n7201 = pi268 & ~n6578;
  assign n7202 = ~n7200 & ~n7201;
  assign n7203 = ~n1761 & ~n7202;
  assign n7204 = ~n7172 & ~n7203;
  assign n7205 = ~n1754 & ~n7204;
  assign n7206 = pi909 & n7196;
  assign n7207 = ~pi909 & ~n7196;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = n1754 & n7208;
  assign po417 = n7205 | n7209;
  assign n7211 = pi269 & n1761;
  assign n7212 = pi796 & ~n6579;
  assign n7213 = pi594 & n6579;
  assign n7214 = ~n7212 & ~n7213;
  assign n7215 = ~n2449 & ~n7214;
  assign n7216 = pi160 & n2449;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = pi562 & n7217;
  assign n7219 = pi594 & n6592;
  assign n7220 = pi160 & n6594;
  assign n7221 = ~n6594 & ~n7217;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = ~n6592 & ~n7222;
  assign n7224 = ~n7219 & ~n7223;
  assign n7225 = n6591 & ~n7224;
  assign n7226 = pi160 & ~pi669;
  assign n7227 = ~n6591 & n7226;
  assign n7228 = n6603 & ~n7224;
  assign n7229 = ~n7227 & ~n7228;
  assign n7230 = ~n7225 & n7229;
  assign n7231 = n2564 & ~n7230;
  assign n7232 = pi160 & ~n2564;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = ~pi562 & n7233;
  assign n7235 = ~n7218 & ~n7234;
  assign n7236 = pi396 & n7235;
  assign n7237 = ~pi396 & ~n7235;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = n6578 & n7238;
  assign n7240 = pi269 & ~n6578;
  assign n7241 = ~n7239 & ~n7240;
  assign n7242 = ~n1761 & ~n7241;
  assign n7243 = ~n7211 & ~n7242;
  assign n7244 = ~n1754 & ~n7243;
  assign n7245 = pi924 & n7235;
  assign n7246 = ~pi924 & ~n7235;
  assign n7247 = ~n7245 & ~n7246;
  assign n7248 = n1754 & n7247;
  assign po418 = n7244 | n7248;
  assign n7250 = pi270 & n1761;
  assign n7251 = pi677 & ~n6579;
  assign n7252 = pi493 & n6579;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n2449 & ~n7253;
  assign n7255 = pi100 & n2449;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = pi562 & n7256;
  assign n7258 = pi493 & n6592;
  assign n7259 = pi100 & n6594;
  assign n7260 = ~n6594 & ~n7256;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = ~n6592 & ~n7261;
  assign n7263 = ~n7258 & ~n7262;
  assign n7264 = n6591 & ~n7263;
  assign n7265 = pi100 & ~pi669;
  assign n7266 = ~n6591 & n7265;
  assign n7267 = n6603 & ~n7263;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = ~n7264 & n7268;
  assign n7270 = n2564 & ~n7269;
  assign n7271 = pi100 & ~n2564;
  assign n7272 = ~n7270 & ~n7271;
  assign n7273 = ~pi562 & n7272;
  assign n7274 = ~n7257 & ~n7273;
  assign n7275 = pi206 & n7274;
  assign n7276 = ~pi206 & ~n7274;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = n6578 & n7277;
  assign n7279 = pi270 & ~n6578;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = ~n1761 & ~n7280;
  assign n7282 = ~n7250 & ~n7281;
  assign n7283 = ~n1754 & ~n7282;
  assign n7284 = pi805 & n7274;
  assign n7285 = ~pi805 & ~n7274;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = n1754 & n7286;
  assign po419 = n7283 | n7287;
  assign n7289 = pi271 & n1761;
  assign n7290 = pi715 & ~n6579;
  assign n7291 = pi652 & n6579;
  assign n7292 = ~n7290 & ~n7291;
  assign n7293 = ~n2449 & ~n7292;
  assign n7294 = pi169 & n2449;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = pi562 & n7295;
  assign n7297 = pi652 & n6592;
  assign n7298 = pi169 & n6594;
  assign n7299 = ~n6594 & ~n7295;
  assign n7300 = ~n7298 & ~n7299;
  assign n7301 = ~n6592 & ~n7300;
  assign n7302 = ~n7297 & ~n7301;
  assign n7303 = n6591 & ~n7302;
  assign n7304 = pi169 & ~pi669;
  assign n7305 = ~n6591 & n7304;
  assign n7306 = n6603 & ~n7302;
  assign n7307 = ~n7305 & ~n7306;
  assign n7308 = ~n7303 & n7307;
  assign n7309 = n2564 & ~n7308;
  assign n7310 = pi169 & ~n2564;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~pi562 & n7311;
  assign n7313 = ~n7296 & ~n7312;
  assign n7314 = pi043 & n7313;
  assign n7315 = ~pi043 & ~n7313;
  assign n7316 = ~n7314 & ~n7315;
  assign n7317 = n6578 & n7316;
  assign n7318 = pi271 & ~n6578;
  assign n7319 = ~n7317 & ~n7318;
  assign n7320 = ~n1761 & ~n7319;
  assign n7321 = ~n7289 & ~n7320;
  assign n7322 = ~n1754 & ~n7321;
  assign n7323 = pi843 & n7313;
  assign n7324 = ~pi843 & ~n7313;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = n1754 & n7325;
  assign po420 = n7322 | n7326;
  assign n7328 = pi272 & n1761;
  assign n7329 = pi797 & ~n6579;
  assign n7330 = pi624 & n6579;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = ~n2449 & ~n7331;
  assign n7333 = pi119 & n2449;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = pi562 & n7334;
  assign n7336 = pi624 & n6592;
  assign n7337 = pi119 & n6594;
  assign n7338 = ~n6594 & ~n7334;
  assign n7339 = ~n7337 & ~n7338;
  assign n7340 = ~n6592 & ~n7339;
  assign n7341 = ~n7336 & ~n7340;
  assign n7342 = n6591 & ~n7341;
  assign n7343 = pi119 & ~pi669;
  assign n7344 = ~n6591 & n7343;
  assign n7345 = n6603 & ~n7341;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = ~n7342 & n7346;
  assign n7348 = n2564 & ~n7347;
  assign n7349 = pi119 & ~n2564;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = ~pi562 & n7350;
  assign n7352 = ~n7335 & ~n7351;
  assign n7353 = pi333 & n7352;
  assign n7354 = ~pi333 & ~n7352;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = n6578 & n7355;
  assign n7357 = pi272 & ~n6578;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = ~n1761 & ~n7358;
  assign n7360 = ~n7328 & ~n7359;
  assign n7361 = ~n1754 & ~n7360;
  assign n7362 = pi925 & n7352;
  assign n7363 = ~pi925 & ~n7352;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = n1754 & n7364;
  assign po421 = n7361 | n7365;
  assign n7367 = pi273 & n1761;
  assign n7368 = pi716 & ~n6579;
  assign n7369 = pi638 & n6579;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n2449 & ~n7370;
  assign n7372 = pi142 & n2449;
  assign n7373 = ~n7371 & ~n7372;
  assign n7374 = pi562 & n7373;
  assign n7375 = pi638 & n6592;
  assign n7376 = pi142 & n6594;
  assign n7377 = ~n6594 & ~n7373;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = ~n6592 & ~n7378;
  assign n7380 = ~n7375 & ~n7379;
  assign n7381 = n6591 & ~n7380;
  assign n7382 = pi142 & ~pi669;
  assign n7383 = ~n6591 & n7382;
  assign n7384 = n6603 & ~n7380;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~n7381 & n7385;
  assign n7387 = n2564 & ~n7386;
  assign n7388 = pi142 & ~n2564;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = ~pi562 & n7389;
  assign n7391 = ~n7374 & ~n7390;
  assign n7392 = pi042 & n7391;
  assign n7393 = ~pi042 & ~n7391;
  assign n7394 = ~n7392 & ~n7393;
  assign n7395 = n6578 & n7394;
  assign n7396 = pi273 & ~n6578;
  assign n7397 = ~n7395 & ~n7396;
  assign n7398 = ~n1761 & ~n7397;
  assign n7399 = ~n7367 & ~n7398;
  assign n7400 = ~n1754 & ~n7399;
  assign n7401 = pi844 & n7391;
  assign n7402 = ~pi844 & ~n7391;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = n1754 & n7403;
  assign po422 = n7400 | n7404;
  assign n7406 = pi274 & n1761;
  assign n7407 = pi717 & ~n6579;
  assign n7408 = pi607 & n6579;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = ~n2449 & ~n7409;
  assign n7411 = pi080 & n2449;
  assign n7412 = ~n7410 & ~n7411;
  assign n7413 = pi562 & n7412;
  assign n7414 = pi607 & n6592;
  assign n7415 = pi080 & n6594;
  assign n7416 = ~n6594 & ~n7412;
  assign n7417 = ~n7415 & ~n7416;
  assign n7418 = ~n6592 & ~n7417;
  assign n7419 = ~n7414 & ~n7418;
  assign n7420 = n6591 & ~n7419;
  assign n7421 = pi080 & ~pi669;
  assign n7422 = ~n6591 & n7421;
  assign n7423 = n6603 & ~n7419;
  assign n7424 = ~n7422 & ~n7423;
  assign n7425 = ~n7420 & n7424;
  assign n7426 = n2564 & ~n7425;
  assign n7427 = pi080 & ~n2564;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = ~pi562 & n7428;
  assign n7430 = ~n7413 & ~n7429;
  assign n7431 = pi012 & n7430;
  assign n7432 = ~pi012 & ~n7430;
  assign n7433 = ~n7431 & ~n7432;
  assign n7434 = n6578 & n7433;
  assign n7435 = pi274 & ~n6578;
  assign n7436 = ~n7434 & ~n7435;
  assign n7437 = ~n1761 & ~n7436;
  assign n7438 = ~n7406 & ~n7437;
  assign n7439 = ~n1754 & ~n7438;
  assign n7440 = pi845 & n7430;
  assign n7441 = ~pi845 & ~n7430;
  assign n7442 = ~n7440 & ~n7441;
  assign n7443 = n1754 & n7442;
  assign po423 = n7439 | n7443;
  assign n7445 = pi275 & n1761;
  assign n7446 = pi718 & ~n6579;
  assign n7447 = pi637 & n6579;
  assign n7448 = ~n7446 & ~n7447;
  assign n7449 = ~n2449 & ~n7448;
  assign n7450 = pi079 & n2449;
  assign n7451 = ~n7449 & ~n7450;
  assign n7452 = pi562 & n7451;
  assign n7453 = pi637 & n6592;
  assign n7454 = pi079 & n6594;
  assign n7455 = ~n6594 & ~n7451;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~n6592 & ~n7456;
  assign n7458 = ~n7453 & ~n7457;
  assign n7459 = n6591 & ~n7458;
  assign n7460 = pi079 & ~pi669;
  assign n7461 = ~n6591 & n7460;
  assign n7462 = n6603 & ~n7458;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = ~n7459 & n7463;
  assign n7465 = n2564 & ~n7464;
  assign n7466 = pi079 & ~n2564;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~pi562 & n7467;
  assign n7469 = ~n7452 & ~n7468;
  assign n7470 = pi013 & n7469;
  assign n7471 = ~pi013 & ~n7469;
  assign n7472 = ~n7470 & ~n7471;
  assign n7473 = n6578 & n7472;
  assign n7474 = pi275 & ~n6578;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = ~n1761 & ~n7475;
  assign n7477 = ~n7445 & ~n7476;
  assign n7478 = ~n1754 & ~n7477;
  assign n7479 = pi846 & n7469;
  assign n7480 = ~pi846 & ~n7469;
  assign n7481 = ~n7479 & ~n7480;
  assign n7482 = n1754 & n7481;
  assign po424 = n7478 | n7482;
  assign n7484 = pi276 & n1761;
  assign n7485 = pi782 & ~n6579;
  assign n7486 = pi572 & n6579;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = ~n2449 & ~n7487;
  assign n7489 = pi074 & n2449;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = pi562 & n7490;
  assign n7492 = pi572 & n6592;
  assign n7493 = pi074 & n6594;
  assign n7494 = ~n6594 & ~n7490;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = ~n6592 & ~n7495;
  assign n7497 = ~n7492 & ~n7496;
  assign n7498 = n6591 & ~n7497;
  assign n7499 = pi074 & ~pi669;
  assign n7500 = ~n6591 & n7499;
  assign n7501 = n6603 & ~n7497;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = ~n7498 & n7502;
  assign n7504 = n2564 & ~n7503;
  assign n7505 = pi074 & ~n2564;
  assign n7506 = ~n7504 & ~n7505;
  assign n7507 = ~pi562 & n7506;
  assign n7508 = ~n7491 & ~n7507;
  assign n7509 = ~pi134 & n7508;
  assign n7510 = pi134 & ~n7508;
  assign n7511 = ~n7509 & ~n7510;
  assign n7512 = n6578 & n7511;
  assign n7513 = pi276 & ~n6578;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 = ~n1761 & ~n7514;
  assign n7516 = ~n7484 & ~n7515;
  assign n7517 = ~n1754 & ~n7516;
  assign n7518 = pi910 & n7508;
  assign n7519 = ~pi910 & ~n7508;
  assign n7520 = ~n7518 & ~n7519;
  assign n7521 = n1754 & n7520;
  assign po425 = n7517 | n7521;
  assign n7523 = pi277 & n1761;
  assign n7524 = pi799 & ~n6579;
  assign n7525 = pi615 & n6579;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = ~n2449 & ~n7526;
  assign n7528 = pi050 & n2449;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = pi562 & n7529;
  assign n7531 = pi615 & n6592;
  assign n7532 = pi050 & n6594;
  assign n7533 = ~n6594 & ~n7529;
  assign n7534 = ~n7532 & ~n7533;
  assign n7535 = ~n6592 & ~n7534;
  assign n7536 = ~n7531 & ~n7535;
  assign n7537 = n6591 & ~n7536;
  assign n7538 = pi050 & ~pi669;
  assign n7539 = ~n6591 & n7538;
  assign n7540 = n6603 & ~n7536;
  assign n7541 = ~n7539 & ~n7540;
  assign n7542 = ~n7537 & n7541;
  assign n7543 = n2564 & ~n7542;
  assign n7544 = pi050 & ~n2564;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~pi562 & n7545;
  assign n7547 = ~n7530 & ~n7546;
  assign n7548 = pi332 & n7547;
  assign n7549 = ~pi332 & ~n7547;
  assign n7550 = ~n7548 & ~n7549;
  assign n7551 = n6578 & n7550;
  assign n7552 = pi277 & ~n6578;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n1761 & ~n7553;
  assign n7555 = ~n7523 & ~n7554;
  assign n7556 = ~n1754 & ~n7555;
  assign n7557 = pi927 & n7547;
  assign n7558 = ~pi927 & ~n7547;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = n1754 & n7559;
  assign po426 = n7556 | n7560;
  assign n7562 = pi278 & n1761;
  assign n7563 = pi720 & ~n6579;
  assign n7564 = pi622 & n6579;
  assign n7565 = ~n7563 & ~n7564;
  assign n7566 = ~n2449 & ~n7565;
  assign n7567 = pi023 & n2449;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = pi562 & n7568;
  assign n7570 = pi622 & n6592;
  assign n7571 = pi023 & n6594;
  assign n7572 = ~n6594 & ~n7568;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = ~n6592 & ~n7573;
  assign n7575 = ~n7570 & ~n7574;
  assign n7576 = n6591 & ~n7575;
  assign n7577 = pi023 & ~pi669;
  assign n7578 = ~n6591 & n7577;
  assign n7579 = n6603 & ~n7575;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n7576 & n7580;
  assign n7582 = n2564 & ~n7581;
  assign n7583 = pi023 & ~n2564;
  assign n7584 = ~n7582 & ~n7583;
  assign n7585 = ~pi562 & n7584;
  assign n7586 = ~n7569 & ~n7585;
  assign n7587 = pi015 & n7586;
  assign n7588 = ~pi015 & ~n7586;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = n6578 & n7589;
  assign n7591 = pi278 & ~n6578;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = ~n1761 & ~n7592;
  assign n7594 = ~n7562 & ~n7593;
  assign n7595 = ~n1754 & ~n7594;
  assign n7596 = pi848 & n7586;
  assign n7597 = ~pi848 & ~n7586;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = n1754 & n7598;
  assign po427 = n7595 | n7599;
  assign n7601 = pi279 & n1761;
  assign n7602 = pi721 & ~n6579;
  assign n7603 = pi605 & n6579;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = ~n2449 & ~n7604;
  assign n7606 = pi081 & n2449;
  assign n7607 = ~n7605 & ~n7606;
  assign n7608 = pi562 & n7607;
  assign n7609 = pi605 & n6592;
  assign n7610 = pi081 & n6594;
  assign n7611 = ~n6594 & ~n7607;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n6592 & ~n7612;
  assign n7614 = ~n7609 & ~n7613;
  assign n7615 = n6591 & ~n7614;
  assign n7616 = pi081 & ~pi669;
  assign n7617 = ~n6591 & n7616;
  assign n7618 = n6603 & ~n7614;
  assign n7619 = ~n7617 & ~n7618;
  assign n7620 = ~n7615 & n7619;
  assign n7621 = n2564 & ~n7620;
  assign n7622 = pi081 & ~n2564;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = ~pi562 & n7623;
  assign n7625 = ~n7608 & ~n7624;
  assign n7626 = pi016 & n7625;
  assign n7627 = ~pi016 & ~n7625;
  assign n7628 = ~n7626 & ~n7627;
  assign n7629 = n6578 & n7628;
  assign n7630 = pi279 & ~n6578;
  assign n7631 = ~n7629 & ~n7630;
  assign n7632 = ~n1761 & ~n7631;
  assign n7633 = ~n7601 & ~n7632;
  assign n7634 = ~n1754 & ~n7633;
  assign n7635 = pi849 & n7625;
  assign n7636 = ~pi849 & ~n7625;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = n1754 & n7637;
  assign po428 = n7634 | n7638;
  assign n7640 = pi280 & n1761;
  assign n7641 = pi800 & ~n6579;
  assign n7642 = pi601 & n6579;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n2449 & ~n7643;
  assign n7645 = pi051 & n2449;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = pi562 & n7646;
  assign n7648 = pi601 & n6592;
  assign n7649 = pi051 & n6594;
  assign n7650 = ~n6594 & ~n7646;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = ~n6592 & ~n7651;
  assign n7653 = ~n7648 & ~n7652;
  assign n7654 = n6591 & ~n7653;
  assign n7655 = pi051 & ~pi669;
  assign n7656 = ~n6591 & n7655;
  assign n7657 = n6603 & ~n7653;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = ~n7654 & n7658;
  assign n7660 = n2564 & ~n7659;
  assign n7661 = pi051 & ~n2564;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = ~pi562 & n7662;
  assign n7664 = ~n7647 & ~n7663;
  assign n7665 = pi394 & n7664;
  assign n7666 = ~pi394 & ~n7664;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = n6578 & n7667;
  assign n7669 = pi280 & ~n6578;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n1761 & ~n7670;
  assign n7672 = ~n7640 & ~n7671;
  assign n7673 = ~n1754 & ~n7672;
  assign n7674 = pi928 & n7664;
  assign n7675 = ~pi928 & ~n7664;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = n1754 & n7676;
  assign po429 = n7673 | n7677;
  assign n7679 = pi281 & n1761;
  assign n7680 = pi801 & ~n6579;
  assign n7681 = pi660 & n6579;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = ~n2449 & ~n7682;
  assign n7684 = pi121 & n2449;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = pi562 & n7685;
  assign n7687 = pi660 & n6592;
  assign n7688 = pi121 & n6594;
  assign n7689 = ~n6594 & ~n7685;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 = ~n6592 & ~n7690;
  assign n7692 = ~n7687 & ~n7691;
  assign n7693 = n6591 & ~n7692;
  assign n7694 = pi121 & ~pi669;
  assign n7695 = ~n6591 & n7694;
  assign n7696 = n6603 & ~n7692;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = ~n7693 & n7697;
  assign n7699 = n2564 & ~n7698;
  assign n7700 = pi121 & ~n2564;
  assign n7701 = ~n7699 & ~n7700;
  assign n7702 = ~pi562 & n7701;
  assign n7703 = ~n7686 & ~n7702;
  assign n7704 = pi389 & n7703;
  assign n7705 = ~pi389 & ~n7703;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = n6578 & n7706;
  assign n7708 = pi281 & ~n6578;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = ~n1761 & ~n7709;
  assign n7711 = ~n7679 & ~n7710;
  assign n7712 = ~n1754 & ~n7711;
  assign n7713 = pi929 & n7703;
  assign n7714 = ~pi929 & ~n7703;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = n1754 & n7715;
  assign po430 = n7712 | n7716;
  assign n7718 = pi282 & n1761;
  assign n7719 = pi684 & ~n6579;
  assign n7720 = pi525 & n6579;
  assign n7721 = ~n7719 & ~n7720;
  assign n7722 = ~n2449 & ~n7721;
  assign n7723 = pi140 & n2449;
  assign n7724 = ~n7722 & ~n7723;
  assign n7725 = pi562 & n7724;
  assign n7726 = pi525 & n6592;
  assign n7727 = pi140 & n6594;
  assign n7728 = ~n6594 & ~n7724;
  assign n7729 = ~n7727 & ~n7728;
  assign n7730 = ~n6592 & ~n7729;
  assign n7731 = ~n7726 & ~n7730;
  assign n7732 = n6591 & ~n7731;
  assign n7733 = pi140 & ~pi669;
  assign n7734 = ~n6591 & n7733;
  assign n7735 = n6603 & ~n7731;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = ~n7732 & n7736;
  assign n7738 = n2564 & ~n7737;
  assign n7739 = pi140 & ~n2564;
  assign n7740 = ~n7738 & ~n7739;
  assign n7741 = ~pi562 & n7740;
  assign n7742 = ~n7725 & ~n7741;
  assign n7743 = pi010 & n7742;
  assign n7744 = ~pi010 & ~n7742;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = n6578 & n7745;
  assign n7747 = pi282 & ~n6578;
  assign n7748 = ~n7746 & ~n7747;
  assign n7749 = ~n1761 & ~n7748;
  assign n7750 = ~n7718 & ~n7749;
  assign n7751 = ~n1754 & ~n7750;
  assign n7752 = pi812 & n7742;
  assign n7753 = ~pi812 & ~n7742;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = n1754 & n7754;
  assign po431 = n7751 | n7755;
  assign n7757 = pi283 & n1761;
  assign n7758 = pi687 & ~n6579;
  assign n7759 = pi530 & n6579;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~n2449 & ~n7760;
  assign n7762 = pi020 & n2449;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = pi562 & n7763;
  assign n7765 = pi530 & n6592;
  assign n7766 = pi020 & n6594;
  assign n7767 = ~n6594 & ~n7763;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = ~n6592 & ~n7768;
  assign n7770 = ~n7765 & ~n7769;
  assign n7771 = n6591 & ~n7770;
  assign n7772 = pi020 & ~pi669;
  assign n7773 = ~n6591 & n7772;
  assign n7774 = n6603 & ~n7770;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = ~n7771 & n7775;
  assign n7777 = n2564 & ~n7776;
  assign n7778 = pi020 & ~n2564;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~pi562 & n7779;
  assign n7781 = ~n7764 & ~n7780;
  assign n7782 = pi002 & n7781;
  assign n7783 = ~pi002 & ~n7781;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = n6578 & n7784;
  assign n7786 = pi283 & ~n6578;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = ~n1761 & ~n7787;
  assign n7789 = ~n7757 & ~n7788;
  assign n7790 = ~n1754 & ~n7789;
  assign n7791 = pi815 & n7781;
  assign n7792 = ~pi815 & ~n7781;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = n1754 & n7793;
  assign po432 = n7790 | n7794;
  assign n7796 = pi284 & n1761;
  assign n7797 = pi784 & ~n6579;
  assign n7798 = pi573 & n6579;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = ~n2449 & ~n7799;
  assign n7801 = pi019 & n2449;
  assign n7802 = ~n7800 & ~n7801;
  assign n7803 = pi562 & n7802;
  assign n7804 = pi573 & n6592;
  assign n7805 = pi019 & n6594;
  assign n7806 = ~n6594 & ~n7802;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = ~n6592 & ~n7807;
  assign n7809 = ~n7804 & ~n7808;
  assign n7810 = n6591 & ~n7809;
  assign n7811 = pi019 & ~pi669;
  assign n7812 = ~n6591 & n7811;
  assign n7813 = n6603 & ~n7809;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n7810 & n7814;
  assign n7816 = n2564 & ~n7815;
  assign n7817 = pi019 & ~n2564;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~pi562 & n7818;
  assign n7820 = ~n7803 & ~n7819;
  assign n7821 = pi166 & n7820;
  assign n7822 = ~pi166 & ~n7820;
  assign n7823 = ~n7821 & ~n7822;
  assign n7824 = n6578 & n7823;
  assign n7825 = pi284 & ~n6578;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = ~n1761 & ~n7826;
  assign n7828 = ~n7796 & ~n7827;
  assign n7829 = ~n1754 & ~n7828;
  assign n7830 = pi912 & n7820;
  assign n7831 = ~pi912 & ~n7820;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = n1754 & n7832;
  assign po433 = n7829 | n7833;
  assign n7835 = pi285 & n1761;
  assign n7836 = pi732 & ~n6579;
  assign n7837 = pi626 & n6579;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = ~n2449 & ~n7838;
  assign n7840 = pi162 & n2449;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = pi562 & n7841;
  assign n7843 = pi626 & n6592;
  assign n7844 = pi162 & n6594;
  assign n7845 = ~n6594 & ~n7841;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = ~n6592 & ~n7846;
  assign n7848 = ~n7843 & ~n7847;
  assign n7849 = n6591 & ~n7848;
  assign n7850 = pi162 & ~pi669;
  assign n7851 = ~n6591 & n7850;
  assign n7852 = n6603 & ~n7848;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = ~n7849 & n7853;
  assign n7855 = n2564 & ~n7854;
  assign n7856 = pi162 & ~n2564;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~pi562 & n7857;
  assign n7859 = ~n7842 & ~n7858;
  assign n7860 = ~pi224 & n7859;
  assign n7861 = pi224 & ~n7859;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = n6578 & n7862;
  assign n7864 = pi285 & ~n6578;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = ~n1761 & ~n7865;
  assign n7867 = ~n7835 & ~n7866;
  assign n7868 = ~n1754 & ~n7867;
  assign n7869 = pi860 & n7859;
  assign n7870 = ~pi860 & ~n7859;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = n1754 & n7871;
  assign po434 = n7868 | n7872;
  assign n7874 = pi286 & n1761;
  assign n7875 = pi731 & ~n6579;
  assign n7876 = pi586 & n6579;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = ~n2449 & ~n7877;
  assign n7879 = ~pi183 & n2449;
  assign n7880 = ~n7878 & ~n7879;
  assign n7881 = pi562 & n7880;
  assign n7882 = pi586 & n6592;
  assign n7883 = ~pi183 & n6594;
  assign n7884 = ~n6594 & ~n7880;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n6592 & ~n7885;
  assign n7887 = ~n7882 & ~n7886;
  assign n7888 = n6591 & ~n7887;
  assign n7889 = ~pi183 & ~pi669;
  assign n7890 = ~n6591 & n7889;
  assign n7891 = n6603 & ~n7887;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = ~n7888 & n7892;
  assign n7894 = n2564 & ~n7893;
  assign n7895 = ~pi183 & ~n2564;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = ~pi562 & n7896;
  assign n7898 = ~n7881 & ~n7897;
  assign n7899 = ~pi223 & n7898;
  assign n7900 = pi223 & ~n7898;
  assign n7901 = ~n7899 & ~n7900;
  assign n7902 = n6578 & n7901;
  assign n7903 = pi286 & ~n6578;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n1761 & ~n7904;
  assign n7906 = ~n7874 & ~n7905;
  assign n7907 = ~n1754 & ~n7906;
  assign n7908 = pi859 & n7898;
  assign n7909 = ~pi859 & ~n7898;
  assign n7910 = ~n7908 & ~n7909;
  assign n7911 = n1754 & n7910;
  assign po435 = n7907 | n7911;
  assign n7913 = pi287 & n1761;
  assign n7914 = pi733 & ~n6579;
  assign n7915 = pi631 & n6579;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n2449 & ~n7916;
  assign n7918 = pi125 & n2449;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = pi562 & n7919;
  assign n7921 = pi631 & n6592;
  assign n7922 = pi125 & n6594;
  assign n7923 = ~n6594 & ~n7919;
  assign n7924 = ~n7922 & ~n7923;
  assign n7925 = ~n6592 & ~n7924;
  assign n7926 = ~n7921 & ~n7925;
  assign n7927 = n6591 & ~n7926;
  assign n7928 = pi125 & ~pi669;
  assign n7929 = ~n6591 & n7928;
  assign n7930 = n6603 & ~n7926;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = ~n7927 & n7931;
  assign n7933 = n2564 & ~n7932;
  assign n7934 = pi125 & ~n2564;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~pi562 & n7935;
  assign n7937 = ~n7920 & ~n7936;
  assign n7938 = ~pi215 & n7937;
  assign n7939 = pi215 & ~n7937;
  assign n7940 = ~n7938 & ~n7939;
  assign n7941 = n6578 & n7940;
  assign n7942 = pi287 & ~n6578;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = ~n1761 & ~n7943;
  assign n7945 = ~n7913 & ~n7944;
  assign n7946 = ~n1754 & ~n7945;
  assign n7947 = pi861 & n7937;
  assign n7948 = ~pi861 & ~n7937;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = n1754 & n7949;
  assign po436 = n7946 | n7950;
  assign n7952 = pi288 & ~po814;
  assign n7953 = po814 & ~n5344;
  assign po437 = n7952 | n7953;
  assign n7955 = pi289 & ~po814;
  assign n7956 = po814 & ~n5982;
  assign po438 = n7955 | n7956;
  assign n7958 = pi290 & ~po814;
  assign n7959 = po814 & ~n6030;
  assign po439 = n7958 | n7959;
  assign n7961 = pi291 & ~po814;
  assign n7962 = po814 & ~n5799;
  assign po440 = n7961 | n7962;
  assign n7964 = pi292 & ~po814;
  assign n7965 = po814 & ~n5740;
  assign po441 = n7964 | n7965;
  assign n7967 = pi293 & ~po814;
  assign n7968 = po814 & ~n5847;
  assign po442 = n7967 | n7968;
  assign n7970 = pi294 & ~po814;
  assign n7971 = po814 & ~n5943;
  assign po443 = n7970 | n7971;
  assign n7973 = pi295 & ~po814;
  assign n7974 = po814 & ~n6135;
  assign po444 = n7973 | n7974;
  assign n7976 = pi296 & ~po814;
  assign n7977 = po814 & ~n6078;
  assign po445 = n7976 | n7977;
  assign n7979 = pi297 & n1761;
  assign n7980 = pi679 & ~n6579;
  assign n7981 = pi544 & n6579;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = ~n2449 & ~n7982;
  assign n7984 = pi036 & n2449;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = pi562 & n7985;
  assign n7987 = pi544 & n6592;
  assign n7988 = pi036 & n6594;
  assign n7989 = ~n6594 & ~n7985;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = ~n6592 & ~n7990;
  assign n7992 = ~n7987 & ~n7991;
  assign n7993 = n6591 & ~n7992;
  assign n7994 = pi036 & ~pi669;
  assign n7995 = ~n6591 & n7994;
  assign n7996 = n6603 & ~n7992;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = ~n7993 & n7997;
  assign n7999 = n2564 & ~n7998;
  assign n8000 = pi036 & ~n2564;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = ~pi562 & n8001;
  assign n8003 = ~n7986 & ~n8002;
  assign n8004 = pi208 & n8003;
  assign n8005 = ~pi208 & ~n8003;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = n6578 & n8006;
  assign n8008 = pi297 & ~n6578;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~n1761 & ~n8009;
  assign n8011 = ~n7979 & ~n8010;
  assign n8012 = ~n1754 & ~n8011;
  assign n8013 = pi807 & n8003;
  assign n8014 = ~pi807 & ~n8003;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = n1754 & n8015;
  assign po446 = n8012 | n8016;
  assign n8018 = pi298 & ~po814;
  assign n8019 = po814 & ~n6180;
  assign po447 = n8018 | n8019;
  assign n8021 = pi299 & n1761;
  assign n8022 = pi714 & ~n6579;
  assign n8023 = pi648 & n6579;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = ~n2449 & ~n8024;
  assign n8026 = pi059 & n2449;
  assign n8027 = ~n8025 & ~n8026;
  assign n8028 = pi562 & n8027;
  assign n8029 = pi648 & n6592;
  assign n8030 = pi059 & n6594;
  assign n8031 = ~n6594 & ~n8027;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = ~n6592 & ~n8032;
  assign n8034 = ~n8029 & ~n8033;
  assign n8035 = n6591 & ~n8034;
  assign n8036 = pi059 & ~pi669;
  assign n8037 = ~n6591 & n8036;
  assign n8038 = n6603 & ~n8034;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = ~n8035 & n8039;
  assign n8041 = n2564 & ~n8040;
  assign n8042 = pi059 & ~n2564;
  assign n8043 = ~n8041 & ~n8042;
  assign n8044 = ~pi562 & n8043;
  assign n8045 = ~n8028 & ~n8044;
  assign n8046 = pi017 & n8045;
  assign n8047 = ~pi017 & ~n8045;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = n6578 & n8048;
  assign n8050 = pi299 & ~n6578;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = ~n1761 & ~n8051;
  assign n8053 = ~n8021 & ~n8052;
  assign n8054 = ~n1754 & ~n8053;
  assign n8055 = pi842 & n8045;
  assign n8056 = ~pi842 & ~n8045;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = n1754 & n8057;
  assign po448 = n8054 | n8058;
  assign n8060 = pi300 & n1761;
  assign n8061 = pi798 & ~n6579;
  assign n8062 = pi642 & n6579;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n2449 & ~n8063;
  assign n8065 = pi120 & n2449;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = pi562 & n8066;
  assign n8068 = pi642 & n6592;
  assign n8069 = pi120 & n6594;
  assign n8070 = ~n6594 & ~n8066;
  assign n8071 = ~n8069 & ~n8070;
  assign n8072 = ~n6592 & ~n8071;
  assign n8073 = ~n8068 & ~n8072;
  assign n8074 = n6591 & ~n8073;
  assign n8075 = pi120 & ~pi669;
  assign n8076 = ~n6591 & n8075;
  assign n8077 = n6603 & ~n8073;
  assign n8078 = ~n8076 & ~n8077;
  assign n8079 = ~n8074 & n8078;
  assign n8080 = n2564 & ~n8079;
  assign n8081 = pi120 & ~n2564;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = ~pi562 & n8082;
  assign n8084 = ~n8067 & ~n8083;
  assign n8085 = pi288 & n8084;
  assign n8086 = ~pi288 & ~n8084;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = n6578 & n8087;
  assign n8089 = pi300 & ~n6578;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = ~n1761 & ~n8090;
  assign n8092 = ~n8060 & ~n8091;
  assign n8093 = ~n1754 & ~n8092;
  assign n8094 = pi926 & n8084;
  assign n8095 = ~pi926 & ~n8084;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = n1754 & n8096;
  assign po449 = n8093 | n8097;
  assign n8099 = pi301 & n1761;
  assign n8100 = pi735 & ~n6579;
  assign n8101 = pi645 & n6579;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n2449 & ~n8102;
  assign n8104 = pi069 & n2449;
  assign n8105 = ~n8103 & ~n8104;
  assign n8106 = pi562 & n8105;
  assign n8107 = pi645 & n6592;
  assign n8108 = pi069 & n6594;
  assign n8109 = ~n6594 & ~n8105;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = ~n6592 & ~n8110;
  assign n8112 = ~n8107 & ~n8111;
  assign n8113 = n6591 & ~n8112;
  assign n8114 = pi069 & ~pi669;
  assign n8115 = ~n6591 & n8114;
  assign n8116 = n6603 & ~n8112;
  assign n8117 = ~n8115 & ~n8116;
  assign n8118 = ~n8113 & n8117;
  assign n8119 = n2564 & ~n8118;
  assign n8120 = pi069 & ~n2564;
  assign n8121 = ~n8119 & ~n8120;
  assign n8122 = ~pi562 & n8121;
  assign n8123 = ~n8106 & ~n8122;
  assign n8124 = ~pi214 & n8123;
  assign n8125 = pi214 & ~n8123;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = n6578 & n8126;
  assign n8128 = pi301 & ~n6578;
  assign n8129 = ~n8127 & ~n8128;
  assign n8130 = ~n1761 & ~n8129;
  assign n8131 = ~n8099 & ~n8130;
  assign n8132 = ~n1754 & ~n8131;
  assign n8133 = pi863 & n8123;
  assign n8134 = ~pi863 & ~n8123;
  assign n8135 = ~n8133 & ~n8134;
  assign n8136 = n1754 & n8135;
  assign po450 = n8132 | n8136;
  assign n8138 = pi302 & n1761;
  assign n8139 = pi736 & ~n6579;
  assign n8140 = pi619 & n6579;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = ~n2449 & ~n8141;
  assign n8143 = pi070 & n2449;
  assign n8144 = ~n8142 & ~n8143;
  assign n8145 = pi562 & n8144;
  assign n8146 = pi619 & n6592;
  assign n8147 = pi070 & n6594;
  assign n8148 = ~n6594 & ~n8144;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = ~n6592 & ~n8149;
  assign n8151 = ~n8146 & ~n8150;
  assign n8152 = n6591 & ~n8151;
  assign n8153 = pi070 & ~pi669;
  assign n8154 = ~n6591 & n8153;
  assign n8155 = n6603 & ~n8151;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n8152 & n8156;
  assign n8158 = n2564 & ~n8157;
  assign n8159 = pi070 & ~n2564;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~pi562 & n8160;
  assign n8162 = ~n8145 & ~n8161;
  assign n8163 = ~pi226 & n8162;
  assign n8164 = pi226 & ~n8162;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = n6578 & n8165;
  assign n8167 = pi302 & ~n6578;
  assign n8168 = ~n8166 & ~n8167;
  assign n8169 = ~n1761 & ~n8168;
  assign n8170 = ~n8138 & ~n8169;
  assign n8171 = ~n1754 & ~n8170;
  assign n8172 = pi864 & n8162;
  assign n8173 = ~pi864 & ~n8162;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = n1754 & n8174;
  assign po451 = n8171 | n8175;
  assign n8177 = pi303 & n1761;
  assign n8178 = pi675 & ~n6579;
  assign n8179 = pi520 & n6579;
  assign n8180 = ~n8178 & ~n8179;
  assign n8181 = ~n2449 & ~n8180;
  assign n8182 = ~pi173 & n2449;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = pi562 & n8183;
  assign n8185 = pi520 & n6592;
  assign n8186 = ~pi173 & n6594;
  assign n8187 = ~n6594 & ~n8183;
  assign n8188 = ~n8186 & ~n8187;
  assign n8189 = ~n6592 & ~n8188;
  assign n8190 = ~n8185 & ~n8189;
  assign n8191 = n6591 & ~n8190;
  assign n8192 = ~pi173 & ~pi669;
  assign n8193 = ~n6591 & n8192;
  assign n8194 = n6603 & ~n8190;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n8191 & n8195;
  assign n8197 = n2564 & ~n8196;
  assign n8198 = ~pi173 & ~n2564;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = ~pi562 & n8199;
  assign n8201 = ~n8184 & ~n8200;
  assign n8202 = pi211 & n8201;
  assign n8203 = ~pi211 & ~n8201;
  assign n8204 = ~n8202 & ~n8203;
  assign n8205 = n6578 & n8204;
  assign n8206 = pi303 & ~n6578;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n1761 & ~n8207;
  assign n8209 = ~n8177 & ~n8208;
  assign n8210 = ~n1754 & ~n8209;
  assign n8211 = pi803 & n8201;
  assign n8212 = ~pi803 & ~n8201;
  assign n8213 = ~n8211 & ~n8212;
  assign n8214 = n1754 & n8213;
  assign po452 = n8210 | n8214;
  assign n8216 = pi304 & n1761;
  assign n8217 = pi747 & ~n6579;
  assign n8218 = pi659 & n6579;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = ~n2449 & ~n8219;
  assign n8221 = pi170 & n2449;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = pi562 & n8222;
  assign n8224 = pi659 & n6592;
  assign n8225 = pi170 & n6594;
  assign n8226 = ~n6594 & ~n8222;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~n6592 & ~n8227;
  assign n8229 = ~n8224 & ~n8228;
  assign n8230 = n6591 & ~n8229;
  assign n8231 = pi170 & ~pi669;
  assign n8232 = ~n6591 & n8231;
  assign n8233 = n6603 & ~n8229;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8230 & n8234;
  assign n8236 = n2564 & ~n8235;
  assign n8237 = pi170 & ~n2564;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~pi562 & n8238;
  assign n8240 = ~n8223 & ~n8239;
  assign n8241 = ~pi047 & n8240;
  assign n8242 = pi047 & ~n8240;
  assign n8243 = ~n8241 & ~n8242;
  assign n8244 = n6578 & n8243;
  assign n8245 = pi304 & ~n6578;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~n1761 & ~n8246;
  assign n8248 = ~n8216 & ~n8247;
  assign n8249 = ~n1754 & ~n8248;
  assign n8250 = pi875 & n8240;
  assign n8251 = ~pi875 & ~n8240;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = n1754 & n8252;
  assign po453 = n8249 | n8253;
  assign n8255 = pi305 & n1761;
  assign n8256 = pi748 & ~n6579;
  assign n8257 = pi603 & n6579;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = ~n2449 & ~n8258;
  assign n8260 = pi141 & n2449;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = pi562 & n8261;
  assign n8263 = pi603 & n6592;
  assign n8264 = pi141 & n6594;
  assign n8265 = ~n6594 & ~n8261;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = ~n6592 & ~n8266;
  assign n8268 = ~n8263 & ~n8267;
  assign n8269 = n6591 & ~n8268;
  assign n8270 = pi141 & ~pi669;
  assign n8271 = ~n6591 & n8270;
  assign n8272 = n6603 & ~n8268;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = ~n8269 & n8273;
  assign n8275 = n2564 & ~n8274;
  assign n8276 = pi141 & ~n2564;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = ~pi562 & n8277;
  assign n8279 = ~n8262 & ~n8278;
  assign n8280 = ~pi046 & n8279;
  assign n8281 = pi046 & ~n8279;
  assign n8282 = ~n8280 & ~n8281;
  assign n8283 = n6578 & n8282;
  assign n8284 = pi305 & ~n6578;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = ~n1761 & ~n8285;
  assign n8287 = ~n8255 & ~n8286;
  assign n8288 = ~n1754 & ~n8287;
  assign n8289 = pi876 & n8279;
  assign n8290 = ~pi876 & ~n8279;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = n1754 & n8291;
  assign po454 = n8288 | n8292;
  assign n8294 = pi306 & n1761;
  assign n8295 = pi698 & ~n6579;
  assign n8296 = pi541 & n6579;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = ~n2449 & ~n8297;
  assign n8299 = pi107 & n2449;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = pi562 & n8300;
  assign n8302 = pi541 & n6592;
  assign n8303 = pi107 & n6594;
  assign n8304 = ~n6594 & ~n8300;
  assign n8305 = ~n8303 & ~n8304;
  assign n8306 = ~n6592 & ~n8305;
  assign n8307 = ~n8302 & ~n8306;
  assign n8308 = n6591 & ~n8307;
  assign n8309 = pi107 & ~pi669;
  assign n8310 = ~n6591 & n8309;
  assign n8311 = n6603 & ~n8307;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = ~n8308 & n8312;
  assign n8314 = n2564 & ~n8313;
  assign n8315 = pi107 & ~n2564;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = ~pi562 & n8316;
  assign n8318 = ~n8301 & ~n8317;
  assign n8319 = pi200 & n8318;
  assign n8320 = ~pi200 & ~n8318;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = n6578 & n8321;
  assign n8323 = pi306 & ~n6578;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = ~n1761 & ~n8324;
  assign n8326 = ~n8294 & ~n8325;
  assign n8327 = ~n1754 & ~n8326;
  assign n8328 = pi826 & n8318;
  assign n8329 = ~pi826 & ~n8318;
  assign n8330 = ~n8328 & ~n8329;
  assign n8331 = n1754 & n8330;
  assign po455 = n8327 | n8331;
  assign n8333 = pi307 & n1761;
  assign n8334 = pi746 & ~n6579;
  assign n8335 = pi582 & n6579;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n2449 & ~n8336;
  assign n8338 = pi060 & n2449;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = pi562 & n8339;
  assign n8341 = pi582 & n6592;
  assign n8342 = pi060 & n6594;
  assign n8343 = ~n6594 & ~n8339;
  assign n8344 = ~n8342 & ~n8343;
  assign n8345 = ~n6592 & ~n8344;
  assign n8346 = ~n8341 & ~n8345;
  assign n8347 = n6591 & ~n8346;
  assign n8348 = pi060 & ~pi669;
  assign n8349 = ~n6591 & n8348;
  assign n8350 = n6603 & ~n8346;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~n8347 & n8351;
  assign n8353 = n2564 & ~n8352;
  assign n8354 = pi060 & ~n2564;
  assign n8355 = ~n8353 & ~n8354;
  assign n8356 = ~pi562 & n8355;
  assign n8357 = ~n8340 & ~n8356;
  assign n8358 = pi056 & n8357;
  assign n8359 = ~pi056 & ~n8357;
  assign n8360 = ~n8358 & ~n8359;
  assign n8361 = n6578 & n8360;
  assign n8362 = pi307 & ~n6578;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n1761 & ~n8363;
  assign n8365 = ~n8333 & ~n8364;
  assign n8366 = ~n1754 & ~n8365;
  assign n8367 = pi874 & n8357;
  assign n8368 = ~pi874 & ~n8357;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n1754 & n8369;
  assign po456 = n8366 | n8370;
  assign n8372 = pi308 & n1761;
  assign n8373 = pi681 & ~n6579;
  assign n8374 = pi546 & n6579;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = ~n2449 & ~n8375;
  assign n8377 = pi101 & n2449;
  assign n8378 = ~n8376 & ~n8377;
  assign n8379 = pi562 & n8378;
  assign n8380 = pi546 & n6592;
  assign n8381 = pi101 & n6594;
  assign n8382 = ~n6594 & ~n8378;
  assign n8383 = ~n8381 & ~n8382;
  assign n8384 = ~n6592 & ~n8383;
  assign n8385 = ~n8380 & ~n8384;
  assign n8386 = n6591 & ~n8385;
  assign n8387 = pi101 & ~pi669;
  assign n8388 = ~n6591 & n8387;
  assign n8389 = n6603 & ~n8385;
  assign n8390 = ~n8388 & ~n8389;
  assign n8391 = ~n8386 & n8390;
  assign n8392 = n2564 & ~n8391;
  assign n8393 = pi101 & ~n2564;
  assign n8394 = ~n8392 & ~n8393;
  assign n8395 = ~pi562 & n8394;
  assign n8396 = ~n8379 & ~n8395;
  assign n8397 = pi213 & n8396;
  assign n8398 = ~pi213 & ~n8396;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = n6578 & n8399;
  assign n8401 = pi308 & ~n6578;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = ~n1761 & ~n8402;
  assign n8404 = ~n8372 & ~n8403;
  assign n8405 = ~n1754 & ~n8404;
  assign n8406 = pi809 & n8396;
  assign n8407 = ~pi809 & ~n8396;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = n1754 & n8408;
  assign po457 = n8405 | n8409;
  assign n8411 = pi309 & n1761;
  assign n8412 = pi702 & ~n6579;
  assign n8413 = pi468 & n6579;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = ~n2449 & ~n8414;
  assign n8416 = pi123 & n2449;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = pi562 & n8417;
  assign n8419 = pi468 & n6592;
  assign n8420 = pi123 & n6594;
  assign n8421 = ~n6594 & ~n8417;
  assign n8422 = ~n8420 & ~n8421;
  assign n8423 = ~n6592 & ~n8422;
  assign n8424 = ~n8419 & ~n8423;
  assign n8425 = n6591 & ~n8424;
  assign n8426 = pi123 & ~pi669;
  assign n8427 = ~n6591 & n8426;
  assign n8428 = n6603 & ~n8424;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~n8425 & n8429;
  assign n8431 = n2564 & ~n8430;
  assign n8432 = pi123 & ~n2564;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = ~pi562 & n8433;
  assign n8435 = ~n8418 & ~n8434;
  assign n8436 = pi196 & n8435;
  assign n8437 = ~pi196 & ~n8435;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = n6578 & n8438;
  assign n8440 = pi309 & ~n6578;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = ~n1761 & ~n8441;
  assign n8443 = ~n8411 & ~n8442;
  assign n8444 = ~n1754 & ~n8443;
  assign n8445 = pi830 & n8435;
  assign n8446 = ~pi830 & ~n8435;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = n1754 & n8447;
  assign po458 = n8444 | n8448;
  assign n8450 = pi310 & n1761;
  assign n8451 = pi778 & ~n6579;
  assign n8452 = pi569 & n6579;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = ~n2449 & ~n8453;
  assign n8455 = pi058 & n2449;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = pi562 & n8456;
  assign n8458 = pi569 & n6592;
  assign n8459 = pi058 & n6594;
  assign n8460 = ~n6594 & ~n8456;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = ~n6592 & ~n8461;
  assign n8463 = ~n8458 & ~n8462;
  assign n8464 = n6591 & ~n8463;
  assign n8465 = pi058 & ~pi669;
  assign n8466 = ~n6591 & n8465;
  assign n8467 = n6603 & ~n8463;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = ~n8464 & n8468;
  assign n8470 = n2564 & ~n8469;
  assign n8471 = pi058 & ~n2564;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = ~pi562 & n8472;
  assign n8474 = ~n8457 & ~n8473;
  assign n8475 = ~pi136 & n8474;
  assign n8476 = pi136 & ~n8474;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = n6578 & n8477;
  assign n8479 = pi310 & ~n6578;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = ~n1761 & ~n8480;
  assign n8482 = ~n8450 & ~n8481;
  assign n8483 = ~n1754 & ~n8482;
  assign n8484 = pi906 & n8474;
  assign n8485 = ~pi906 & ~n8474;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = n1754 & n8486;
  assign po459 = n8483 | n8487;
  assign n8489 = pi311 & n1761;
  assign n8490 = pi704 & ~n6579;
  assign n8491 = pi534 & n6579;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = ~n2449 & ~n8492;
  assign n8494 = pi054 & n2449;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = pi562 & n8495;
  assign n8497 = pi534 & n6592;
  assign n8498 = pi054 & n6594;
  assign n8499 = ~n6594 & ~n8495;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = ~n6592 & ~n8500;
  assign n8502 = ~n8497 & ~n8501;
  assign n8503 = n6591 & ~n8502;
  assign n8504 = pi054 & ~pi669;
  assign n8505 = ~n6591 & n8504;
  assign n8506 = n6603 & ~n8502;
  assign n8507 = ~n8505 & ~n8506;
  assign n8508 = ~n8503 & n8507;
  assign n8509 = n2564 & ~n8508;
  assign n8510 = pi054 & ~n2564;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = ~pi562 & n8511;
  assign n8513 = ~n8496 & ~n8512;
  assign n8514 = pi199 & n8513;
  assign n8515 = ~pi199 & ~n8513;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = n6578 & n8516;
  assign n8518 = pi311 & ~n6578;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = ~n1761 & ~n8519;
  assign n8521 = ~n8489 & ~n8520;
  assign n8522 = ~n1754 & ~n8521;
  assign n8523 = pi832 & n8513;
  assign n8524 = ~pi832 & ~n8513;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = n1754 & n8525;
  assign po460 = n8522 | n8526;
  assign n8528 = pi312 & n1761;
  assign n8529 = pi676 & ~n6579;
  assign n8530 = pi524 & n6579;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = ~n2449 & ~n8531;
  assign n8533 = pi148 & n2449;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = pi562 & n8534;
  assign n8536 = pi524 & n6592;
  assign n8537 = pi148 & n6594;
  assign n8538 = ~n6594 & ~n8534;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = ~n6592 & ~n8539;
  assign n8541 = ~n8536 & ~n8540;
  assign n8542 = n6591 & ~n8541;
  assign n8543 = pi148 & ~pi669;
  assign n8544 = ~n6591 & n8543;
  assign n8545 = n6603 & ~n8541;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = ~n8542 & n8546;
  assign n8548 = n2564 & ~n8547;
  assign n8549 = pi148 & ~n2564;
  assign n8550 = ~n8548 & ~n8549;
  assign n8551 = ~pi562 & n8550;
  assign n8552 = ~n8535 & ~n8551;
  assign n8553 = pi205 & n8552;
  assign n8554 = ~pi205 & ~n8552;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = n6578 & n8555;
  assign n8557 = pi312 & ~n6578;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = ~n1761 & ~n8558;
  assign n8560 = ~n8528 & ~n8559;
  assign n8561 = ~n1754 & ~n8560;
  assign n8562 = pi804 & n8552;
  assign n8563 = ~pi804 & ~n8552;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = n1754 & n8564;
  assign po461 = n8561 | n8565;
  assign n8567 = pi313 & n1761;
  assign n8568 = pi705 & ~n6579;
  assign n8569 = pi548 & n6579;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = ~n2449 & ~n8570;
  assign n8572 = pi124 & n2449;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = pi562 & n8573;
  assign n8575 = pi548 & n6592;
  assign n8576 = pi124 & n6594;
  assign n8577 = ~n6594 & ~n8573;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n6592 & ~n8578;
  assign n8580 = ~n8575 & ~n8579;
  assign n8581 = n6591 & ~n8580;
  assign n8582 = pi124 & ~pi669;
  assign n8583 = ~n6591 & n8582;
  assign n8584 = n6603 & ~n8580;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = ~n8581 & n8585;
  assign n8587 = n2564 & ~n8586;
  assign n8588 = pi124 & ~n2564;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = ~pi562 & n8589;
  assign n8591 = ~n8574 & ~n8590;
  assign n8592 = pi201 & n8591;
  assign n8593 = ~pi201 & ~n8591;
  assign n8594 = ~n8592 & ~n8593;
  assign n8595 = n6578 & n8594;
  assign n8596 = pi313 & ~n6578;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = ~n1761 & ~n8597;
  assign n8599 = ~n8567 & ~n8598;
  assign n8600 = ~n1754 & ~n8599;
  assign n8601 = pi833 & n8591;
  assign n8602 = ~pi833 & ~n8591;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = n1754 & n8603;
  assign po462 = n8600 | n8604;
  assign n8606 = pi314 & n1761;
  assign n8607 = pi764 & ~n6579;
  assign n8608 = pi602 & n6579;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = ~n2449 & ~n8609;
  assign n8611 = pi163 & n2449;
  assign n8612 = ~n8610 & ~n8611;
  assign n8613 = pi562 & n8612;
  assign n8614 = pi602 & n6592;
  assign n8615 = pi163 & n6594;
  assign n8616 = ~n6594 & ~n8612;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = ~n6592 & ~n8617;
  assign n8619 = ~n8614 & ~n8618;
  assign n8620 = n6591 & ~n8619;
  assign n8621 = pi163 & ~pi669;
  assign n8622 = ~n6591 & n8621;
  assign n8623 = n6603 & ~n8619;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~n8620 & n8624;
  assign n8626 = n2564 & ~n8625;
  assign n8627 = pi163 & ~n2564;
  assign n8628 = ~n8626 & ~n8627;
  assign n8629 = ~pi562 & n8628;
  assign n8630 = ~n8613 & ~n8629;
  assign n8631 = ~pi247 & n8630;
  assign n8632 = pi247 & ~n8630;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = n6578 & n8633;
  assign n8635 = pi314 & ~n6578;
  assign n8636 = ~n8634 & ~n8635;
  assign n8637 = ~n1761 & ~n8636;
  assign n8638 = ~n8606 & ~n8637;
  assign n8639 = ~n1754 & ~n8638;
  assign n8640 = pi892 & n8630;
  assign n8641 = ~pi892 & ~n8630;
  assign n8642 = ~n8640 & ~n8641;
  assign n8643 = n1754 & n8642;
  assign po463 = n8639 | n8643;
  assign n8645 = pi315 & n1761;
  assign n8646 = pi765 & ~n6579;
  assign n8647 = pi584 & n6579;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n2449 & ~n8648;
  assign n8650 = pi129 & n2449;
  assign n8651 = ~n8649 & ~n8650;
  assign n8652 = pi562 & n8651;
  assign n8653 = pi584 & n6592;
  assign n8654 = pi129 & n6594;
  assign n8655 = ~n6594 & ~n8651;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = ~n6592 & ~n8656;
  assign n8658 = ~n8653 & ~n8657;
  assign n8659 = n6591 & ~n8658;
  assign n8660 = pi129 & ~pi669;
  assign n8661 = ~n6591 & n8660;
  assign n8662 = n6603 & ~n8658;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = ~n8659 & n8663;
  assign n8665 = n2564 & ~n8664;
  assign n8666 = pi129 & ~n2564;
  assign n8667 = ~n8665 & ~n8666;
  assign n8668 = ~pi562 & n8667;
  assign n8669 = ~n8652 & ~n8668;
  assign n8670 = pi238 & n8669;
  assign n8671 = ~pi238 & ~n8669;
  assign n8672 = ~n8670 & ~n8671;
  assign n8673 = n6578 & n8672;
  assign n8674 = pi315 & ~n6578;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n1761 & ~n8675;
  assign n8677 = ~n8645 & ~n8676;
  assign n8678 = ~n1754 & ~n8677;
  assign n8679 = pi893 & n8669;
  assign n8680 = ~pi893 & ~n8669;
  assign n8681 = ~n8679 & ~n8680;
  assign n8682 = n1754 & n8681;
  assign po464 = n8678 | n8682;
  assign n8684 = pi316 & n1761;
  assign n8685 = pi766 & ~n6579;
  assign n8686 = pi654 & n6579;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = ~n2449 & ~n8687;
  assign n8689 = pi130 & n2449;
  assign n8690 = ~n8688 & ~n8689;
  assign n8691 = pi562 & n8690;
  assign n8692 = pi654 & n6592;
  assign n8693 = pi130 & n6594;
  assign n8694 = ~n6594 & ~n8690;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = ~n6592 & ~n8695;
  assign n8697 = ~n8692 & ~n8696;
  assign n8698 = n6591 & ~n8697;
  assign n8699 = pi130 & ~pi669;
  assign n8700 = ~n6591 & n8699;
  assign n8701 = n6603 & ~n8697;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = ~n8698 & n8702;
  assign n8704 = n2564 & ~n8703;
  assign n8705 = pi130 & ~n2564;
  assign n8706 = ~n8704 & ~n8705;
  assign n8707 = ~pi562 & n8706;
  assign n8708 = ~n8691 & ~n8707;
  assign n8709 = ~pi228 & n8708;
  assign n8710 = pi228 & ~n8708;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = n6578 & n8711;
  assign n8713 = pi316 & ~n6578;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = ~n1761 & ~n8714;
  assign n8716 = ~n8684 & ~n8715;
  assign n8717 = ~n1754 & ~n8716;
  assign n8718 = pi894 & n8708;
  assign n8719 = ~pi894 & ~n8708;
  assign n8720 = ~n8718 & ~n8719;
  assign n8721 = n1754 & n8720;
  assign po465 = n8717 | n8721;
  assign n8723 = pi317 & n1761;
  assign n8724 = pi708 & ~n6579;
  assign n8725 = pi650 & n6579;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = ~n2449 & ~n8726;
  assign n8728 = pi158 & n2449;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = pi562 & n8729;
  assign n8731 = pi650 & n6592;
  assign n8732 = pi158 & n6594;
  assign n8733 = ~n6594 & ~n8729;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = ~n6592 & ~n8734;
  assign n8736 = ~n8731 & ~n8735;
  assign n8737 = n6591 & ~n8736;
  assign n8738 = pi158 & ~pi669;
  assign n8739 = ~n6591 & n8738;
  assign n8740 = n6603 & ~n8736;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = ~n8737 & n8741;
  assign n8743 = n2564 & ~n8742;
  assign n8744 = pi158 & ~n2564;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~pi562 & n8745;
  assign n8747 = ~n8730 & ~n8746;
  assign n8748 = ~pi231 & n8747;
  assign n8749 = pi231 & ~n8747;
  assign n8750 = ~n8748 & ~n8749;
  assign n8751 = n6578 & n8750;
  assign n8752 = pi317 & ~n6578;
  assign n8753 = ~n8751 & ~n8752;
  assign n8754 = ~n1761 & ~n8753;
  assign n8755 = ~n8723 & ~n8754;
  assign n8756 = ~n1754 & ~n8755;
  assign n8757 = pi836 & n8747;
  assign n8758 = ~pi836 & ~n8747;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = n1754 & n8759;
  assign po466 = n8756 | n8760;
  assign n8762 = pi318 & n1761;
  assign n8763 = pi767 & ~n6579;
  assign n8764 = pi590 & n6579;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = ~n2449 & ~n8765;
  assign n8767 = pi055 & n2449;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = pi562 & n8768;
  assign n8770 = pi590 & n6592;
  assign n8771 = pi055 & n6594;
  assign n8772 = ~n6594 & ~n8768;
  assign n8773 = ~n8771 & ~n8772;
  assign n8774 = ~n6592 & ~n8773;
  assign n8775 = ~n8770 & ~n8774;
  assign n8776 = n6591 & ~n8775;
  assign n8777 = pi055 & ~pi669;
  assign n8778 = ~n6591 & n8777;
  assign n8779 = n6603 & ~n8775;
  assign n8780 = ~n8778 & ~n8779;
  assign n8781 = ~n8776 & n8780;
  assign n8782 = n2564 & ~n8781;
  assign n8783 = pi055 & ~n2564;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~pi562 & n8784;
  assign n8786 = ~n8769 & ~n8785;
  assign n8787 = ~pi239 & n8786;
  assign n8788 = pi239 & ~n8786;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = n6578 & n8789;
  assign n8791 = pi318 & ~n6578;
  assign n8792 = ~n8790 & ~n8791;
  assign n8793 = ~n1761 & ~n8792;
  assign n8794 = ~n8762 & ~n8793;
  assign n8795 = ~n1754 & ~n8794;
  assign n8796 = pi895 & n8786;
  assign n8797 = ~pi895 & ~n8786;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = n1754 & n8798;
  assign po467 = n8795 | n8799;
  assign n8801 = pi319 & n1761;
  assign n8802 = pi685 & ~n6579;
  assign n8803 = pi510 & n6579;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = ~n2449 & ~n8804;
  assign n8806 = pi076 & n2449;
  assign n8807 = ~n8805 & ~n8806;
  assign n8808 = pi562 & n8807;
  assign n8809 = pi510 & n6592;
  assign n8810 = pi076 & n6594;
  assign n8811 = ~n6594 & ~n8807;
  assign n8812 = ~n8810 & ~n8811;
  assign n8813 = ~n6592 & ~n8812;
  assign n8814 = ~n8809 & ~n8813;
  assign n8815 = n6591 & ~n8814;
  assign n8816 = pi076 & ~pi669;
  assign n8817 = ~n6591 & n8816;
  assign n8818 = n6603 & ~n8814;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~n8815 & n8819;
  assign n8821 = n2564 & ~n8820;
  assign n8822 = pi076 & ~n2564;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = ~pi562 & n8823;
  assign n8825 = ~n8808 & ~n8824;
  assign n8826 = pi000 & n8825;
  assign n8827 = ~pi000 & ~n8825;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = n6578 & n8828;
  assign n8830 = pi319 & ~n6578;
  assign n8831 = ~n8829 & ~n8830;
  assign n8832 = ~n1761 & ~n8831;
  assign n8833 = ~n8801 & ~n8832;
  assign n8834 = ~n1754 & ~n8833;
  assign n8835 = pi813 & n8825;
  assign n8836 = ~pi813 & ~n8825;
  assign n8837 = ~n8835 & ~n8836;
  assign n8838 = n1754 & n8837;
  assign po468 = n8834 | n8838;
  assign n8840 = pi320 & n1761;
  assign n8841 = pi768 & ~n6579;
  assign n8842 = pi639 & n6579;
  assign n8843 = ~n8841 & ~n8842;
  assign n8844 = ~n2449 & ~n8843;
  assign n8845 = pi053 & n2449;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = pi562 & n8846;
  assign n8848 = pi639 & n6592;
  assign n8849 = pi053 & n6594;
  assign n8850 = ~n6594 & ~n8846;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = ~n6592 & ~n8851;
  assign n8853 = ~n8848 & ~n8852;
  assign n8854 = n6591 & ~n8853;
  assign n8855 = pi053 & ~pi669;
  assign n8856 = ~n6591 & n8855;
  assign n8857 = n6603 & ~n8853;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8854 & n8858;
  assign n8860 = n2564 & ~n8859;
  assign n8861 = pi053 & ~n2564;
  assign n8862 = ~n8860 & ~n8861;
  assign n8863 = ~pi562 & n8862;
  assign n8864 = ~n8847 & ~n8863;
  assign n8865 = pi249 & n8864;
  assign n8866 = ~pi249 & ~n8864;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = n6578 & n8867;
  assign n8869 = pi320 & ~n6578;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = ~n1761 & ~n8870;
  assign n8872 = ~n8840 & ~n8871;
  assign n8873 = ~n1754 & ~n8872;
  assign n8874 = pi896 & n8864;
  assign n8875 = ~pi896 & ~n8864;
  assign n8876 = ~n8874 & ~n8875;
  assign n8877 = n1754 & n8876;
  assign po469 = n8873 | n8877;
  assign n8879 = pi321 & n1761;
  assign n8880 = pi769 & ~n6579;
  assign n8881 = pi661 & n6579;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = ~n2449 & ~n8882;
  assign n8884 = pi128 & n2449;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = pi562 & n8885;
  assign n8887 = pi661 & n6592;
  assign n8888 = pi128 & n6594;
  assign n8889 = ~n6594 & ~n8885;
  assign n8890 = ~n8888 & ~n8889;
  assign n8891 = ~n6592 & ~n8890;
  assign n8892 = ~n8887 & ~n8891;
  assign n8893 = n6591 & ~n8892;
  assign n8894 = pi128 & ~pi669;
  assign n8895 = ~n6591 & n8894;
  assign n8896 = n6603 & ~n8892;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = ~n8893 & n8897;
  assign n8899 = n2564 & ~n8898;
  assign n8900 = pi128 & ~n2564;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = ~pi562 & n8901;
  assign n8903 = ~n8886 & ~n8902;
  assign n8904 = pi250 & n8903;
  assign n8905 = ~pi250 & ~n8903;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = n6578 & n8906;
  assign n8908 = pi321 & ~n6578;
  assign n8909 = ~n8907 & ~n8908;
  assign n8910 = ~n1761 & ~n8909;
  assign n8911 = ~n8879 & ~n8910;
  assign n8912 = ~n1754 & ~n8911;
  assign n8913 = pi897 & n8903;
  assign n8914 = ~pi897 & ~n8903;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = n1754 & n8915;
  assign po470 = n8912 | n8916;
  assign n8918 = pi322 & n1761;
  assign n8919 = pi794 & ~n6579;
  assign n8920 = pi647 & n6579;
  assign n8921 = ~n8919 & ~n8920;
  assign n8922 = ~n2449 & ~n8921;
  assign n8923 = pi106 & n2449;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = pi562 & n8924;
  assign n8926 = pi647 & n6592;
  assign n8927 = pi106 & n6594;
  assign n8928 = ~n6594 & ~n8924;
  assign n8929 = ~n8927 & ~n8928;
  assign n8930 = ~n6592 & ~n8929;
  assign n8931 = ~n8926 & ~n8930;
  assign n8932 = n6591 & ~n8931;
  assign n8933 = pi106 & ~pi669;
  assign n8934 = ~n6591 & n8933;
  assign n8935 = n6603 & ~n8931;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8932 & n8936;
  assign n8938 = n2564 & ~n8937;
  assign n8939 = pi106 & ~n2564;
  assign n8940 = ~n8938 & ~n8939;
  assign n8941 = ~pi562 & n8940;
  assign n8942 = ~n8925 & ~n8941;
  assign n8943 = pi387 & n8942;
  assign n8944 = ~pi387 & ~n8942;
  assign n8945 = ~n8943 & ~n8944;
  assign n8946 = n6578 & n8945;
  assign n8947 = pi322 & ~n6578;
  assign n8948 = ~n8946 & ~n8947;
  assign n8949 = ~n1761 & ~n8948;
  assign n8950 = ~n8918 & ~n8949;
  assign n8951 = ~n1754 & ~n8950;
  assign n8952 = pi922 & n8942;
  assign n8953 = ~pi922 & ~n8942;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = n1754 & n8954;
  assign po471 = n8951 | n8955;
  assign n8957 = pi323 & n1761;
  assign n8958 = pi683 & ~n6579;
  assign n8959 = pi523 & n6579;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = ~n2449 & ~n8960;
  assign n8962 = pi171 & n2449;
  assign n8963 = ~n8961 & ~n8962;
  assign n8964 = pi562 & n8963;
  assign n8965 = pi523 & n6592;
  assign n8966 = pi171 & n6594;
  assign n8967 = ~n6594 & ~n8963;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = ~n6592 & ~n8968;
  assign n8970 = ~n8965 & ~n8969;
  assign n8971 = n6591 & ~n8970;
  assign n8972 = pi171 & ~pi669;
  assign n8973 = ~n6591 & n8972;
  assign n8974 = n6603 & ~n8970;
  assign n8975 = ~n8973 & ~n8974;
  assign n8976 = ~n8971 & n8975;
  assign n8977 = n2564 & ~n8976;
  assign n8978 = pi171 & ~n2564;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = ~pi562 & n8979;
  assign n8981 = ~n8964 & ~n8980;
  assign n8982 = pi011 & n8981;
  assign n8983 = ~pi011 & ~n8981;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = n6578 & n8984;
  assign n8986 = pi323 & ~n6578;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = ~n1761 & ~n8987;
  assign n8989 = ~n8957 & ~n8988;
  assign n8990 = ~n1754 & ~n8989;
  assign n8991 = pi811 & n8981;
  assign n8992 = ~pi811 & ~n8981;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = n1754 & n8993;
  assign po472 = n8990 | n8994;
  assign n8996 = pi324 & n1761;
  assign n8997 = pi795 & ~n6579;
  assign n8998 = pi653 & n6579;
  assign n8999 = ~n8997 & ~n8998;
  assign n9000 = ~n2449 & ~n8999;
  assign n9001 = ~pi187 & n2449;
  assign n9002 = ~n9000 & ~n9001;
  assign n9003 = pi562 & n9002;
  assign n9004 = pi653 & n6592;
  assign n9005 = ~pi187 & n6594;
  assign n9006 = ~n6594 & ~n9002;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = ~n6592 & ~n9007;
  assign n9009 = ~n9004 & ~n9008;
  assign n9010 = n6591 & ~n9009;
  assign n9011 = ~pi187 & ~pi669;
  assign n9012 = ~n6591 & n9011;
  assign n9013 = n6603 & ~n9009;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~n9010 & n9014;
  assign n9016 = n2564 & ~n9015;
  assign n9017 = ~pi187 & ~n2564;
  assign n9018 = ~n9016 & ~n9017;
  assign n9019 = ~pi562 & n9018;
  assign n9020 = ~n9003 & ~n9019;
  assign n9021 = pi388 & n9020;
  assign n9022 = ~pi388 & ~n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = n6578 & n9023;
  assign n9025 = pi324 & ~n6578;
  assign n9026 = ~n9024 & ~n9025;
  assign n9027 = ~n1761 & ~n9026;
  assign n9028 = ~n8996 & ~n9027;
  assign n9029 = ~n1754 & ~n9028;
  assign n9030 = pi923 & n9020;
  assign n9031 = ~pi923 & ~n9020;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = n1754 & n9032;
  assign po473 = n9029 | n9033;
  assign n9035 = pi325 & n1761;
  assign n9036 = pi719 & ~n6579;
  assign n9037 = pi575 & n6579;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~n2449 & ~n9038;
  assign n9040 = pi022 & n2449;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = pi562 & n9041;
  assign n9043 = pi575 & n6592;
  assign n9044 = pi022 & n6594;
  assign n9045 = ~n6594 & ~n9041;
  assign n9046 = ~n9044 & ~n9045;
  assign n9047 = ~n6592 & ~n9046;
  assign n9048 = ~n9043 & ~n9047;
  assign n9049 = n6591 & ~n9048;
  assign n9050 = pi022 & ~pi669;
  assign n9051 = ~n6591 & n9050;
  assign n9052 = n6603 & ~n9048;
  assign n9053 = ~n9051 & ~n9052;
  assign n9054 = ~n9049 & n9053;
  assign n9055 = n2564 & ~n9054;
  assign n9056 = pi022 & ~n2564;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~pi562 & n9057;
  assign n9059 = ~n9042 & ~n9058;
  assign n9060 = pi014 & n9059;
  assign n9061 = ~pi014 & ~n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = n6578 & n9062;
  assign n9064 = pi325 & ~n6578;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = ~n1761 & ~n9065;
  assign n9067 = ~n9035 & ~n9066;
  assign n9068 = ~n1754 & ~n9067;
  assign n9069 = pi847 & n9059;
  assign n9070 = ~pi847 & ~n9059;
  assign n9071 = ~n9069 & ~n9070;
  assign n9072 = n1754 & n9071;
  assign po474 = n9068 | n9072;
  assign n9074 = pi326 & n1761;
  assign n9075 = pi678 & ~n6579;
  assign n9076 = pi469 & n6579;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = ~n2449 & ~n9077;
  assign n9079 = pi093 & n2449;
  assign n9080 = ~n9078 & ~n9079;
  assign n9081 = pi562 & n9080;
  assign n9082 = pi469 & n6592;
  assign n9083 = pi093 & n6594;
  assign n9084 = ~n6594 & ~n9080;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n6592 & ~n9085;
  assign n9087 = ~n9082 & ~n9086;
  assign n9088 = n6591 & ~n9087;
  assign n9089 = pi093 & ~pi669;
  assign n9090 = ~n6591 & n9089;
  assign n9091 = n6603 & ~n9087;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = ~n9088 & n9092;
  assign n9094 = n2564 & ~n9093;
  assign n9095 = pi093 & ~n2564;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = ~pi562 & n9096;
  assign n9098 = ~n9081 & ~n9097;
  assign n9099 = pi207 & n9098;
  assign n9100 = ~pi207 & ~n9098;
  assign n9101 = ~n9099 & ~n9100;
  assign n9102 = n6578 & n9101;
  assign n9103 = pi326 & ~n6578;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = ~n1761 & ~n9104;
  assign n9106 = ~n9074 & ~n9105;
  assign n9107 = ~n1754 & ~n9106;
  assign n9108 = pi806 & n9098;
  assign n9109 = ~pi806 & ~n9098;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = n1754 & n9110;
  assign po475 = n9107 | n9111;
  assign n9113 = pi327 & n1761;
  assign n9114 = pi686 & ~n6579;
  assign n9115 = pi466 & n6579;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = ~n2449 & ~n9116;
  assign n9118 = pi077 & n2449;
  assign n9119 = ~n9117 & ~n9118;
  assign n9120 = pi562 & n9119;
  assign n9121 = pi466 & n6592;
  assign n9122 = pi077 & n6594;
  assign n9123 = ~n6594 & ~n9119;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = ~n6592 & ~n9124;
  assign n9126 = ~n9121 & ~n9125;
  assign n9127 = n6591 & ~n9126;
  assign n9128 = pi077 & ~pi669;
  assign n9129 = ~n6591 & n9128;
  assign n9130 = n6603 & ~n9126;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = ~n9127 & n9131;
  assign n9133 = n2564 & ~n9132;
  assign n9134 = pi077 & ~n2564;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = ~pi562 & n9135;
  assign n9137 = ~n9120 & ~n9136;
  assign n9138 = pi001 & n9137;
  assign n9139 = ~pi001 & ~n9137;
  assign n9140 = ~n9138 & ~n9139;
  assign n9141 = n6578 & n9140;
  assign n9142 = pi327 & ~n6578;
  assign n9143 = ~n9141 & ~n9142;
  assign n9144 = ~n1761 & ~n9143;
  assign n9145 = ~n9113 & ~n9144;
  assign n9146 = ~n1754 & ~n9145;
  assign n9147 = pi814 & n9137;
  assign n9148 = ~pi814 & ~n9137;
  assign n9149 = ~n9147 & ~n9148;
  assign n9150 = n1754 & n9149;
  assign po476 = n9146 | n9150;
  assign n9152 = pi328 & n1761;
  assign n9153 = pi783 & ~n6579;
  assign n9154 = pi612 & n6579;
  assign n9155 = ~n9153 & ~n9154;
  assign n9156 = ~n2449 & ~n9155;
  assign n9157 = pi018 & n2449;
  assign n9158 = ~n9156 & ~n9157;
  assign n9159 = pi562 & n9158;
  assign n9160 = pi612 & n6592;
  assign n9161 = pi018 & n6594;
  assign n9162 = ~n6594 & ~n9158;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = ~n6592 & ~n9163;
  assign n9165 = ~n9160 & ~n9164;
  assign n9166 = n6591 & ~n9165;
  assign n9167 = pi018 & ~pi669;
  assign n9168 = ~n6591 & n9167;
  assign n9169 = n6603 & ~n9165;
  assign n9170 = ~n9168 & ~n9169;
  assign n9171 = ~n9166 & n9170;
  assign n9172 = n2564 & ~n9171;
  assign n9173 = pi018 & ~n2564;
  assign n9174 = ~n9172 & ~n9173;
  assign n9175 = ~pi562 & n9174;
  assign n9176 = ~n9159 & ~n9175;
  assign n9177 = pi167 & n9176;
  assign n9178 = ~pi167 & ~n9176;
  assign n9179 = ~n9177 & ~n9178;
  assign n9180 = n6578 & n9179;
  assign n9181 = pi328 & ~n6578;
  assign n9182 = ~n9180 & ~n9181;
  assign n9183 = ~n1761 & ~n9182;
  assign n9184 = ~n9152 & ~n9183;
  assign n9185 = ~n1754 & ~n9184;
  assign n9186 = pi911 & n9176;
  assign n9187 = ~pi911 & ~n9176;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = n1754 & n9188;
  assign po477 = n9185 | n9189;
  assign n9191 = pi329 & n1761;
  assign n9192 = pi688 & ~n6579;
  assign n9193 = pi539 & n6579;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = ~n2449 & ~n9194;
  assign n9196 = pi021 & n2449;
  assign n9197 = ~n9195 & ~n9196;
  assign n9198 = pi562 & n9197;
  assign n9199 = pi539 & n6592;
  assign n9200 = pi021 & n6594;
  assign n9201 = ~n6594 & ~n9197;
  assign n9202 = ~n9200 & ~n9201;
  assign n9203 = ~n6592 & ~n9202;
  assign n9204 = ~n9199 & ~n9203;
  assign n9205 = n6591 & ~n9204;
  assign n9206 = pi021 & ~pi669;
  assign n9207 = ~n6591 & n9206;
  assign n9208 = n6603 & ~n9204;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = ~n9205 & n9209;
  assign n9211 = n2564 & ~n9210;
  assign n9212 = pi021 & ~n2564;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~pi562 & n9213;
  assign n9215 = ~n9198 & ~n9214;
  assign n9216 = pi003 & n9215;
  assign n9217 = ~pi003 & ~n9215;
  assign n9218 = ~n9216 & ~n9217;
  assign n9219 = n6578 & n9218;
  assign n9220 = pi329 & ~n6578;
  assign n9221 = ~n9219 & ~n9220;
  assign n9222 = ~n1761 & ~n9221;
  assign n9223 = ~n9191 & ~n9222;
  assign n9224 = ~n1754 & ~n9223;
  assign n9225 = pi816 & n9215;
  assign n9226 = ~pi816 & ~n9215;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = n1754 & n9227;
  assign po478 = n9224 | n9228;
  assign n9230 = pi330 & n1761;
  assign n9231 = pi730 & ~n6579;
  assign n9232 = pi604 & n6579;
  assign n9233 = ~n9231 & ~n9232;
  assign n9234 = ~n2449 & ~n9233;
  assign n9235 = pi108 & n2449;
  assign n9236 = ~n9234 & ~n9235;
  assign n9237 = pi562 & n9236;
  assign n9238 = pi604 & n6592;
  assign n9239 = pi108 & n6594;
  assign n9240 = ~n6594 & ~n9236;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = ~n6592 & ~n9241;
  assign n9243 = ~n9238 & ~n9242;
  assign n9244 = n6591 & ~n9243;
  assign n9245 = pi108 & ~pi669;
  assign n9246 = ~n6591 & n9245;
  assign n9247 = n6603 & ~n9243;
  assign n9248 = ~n9246 & ~n9247;
  assign n9249 = ~n9244 & n9248;
  assign n9250 = n2564 & ~n9249;
  assign n9251 = pi108 & ~n2564;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = ~pi562 & n9252;
  assign n9254 = ~n9237 & ~n9253;
  assign n9255 = ~pi227 & n9254;
  assign n9256 = pi227 & ~n9254;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = n6578 & n9257;
  assign n9259 = pi330 & ~n6578;
  assign n9260 = ~n9258 & ~n9259;
  assign n9261 = ~n1761 & ~n9260;
  assign n9262 = ~n9230 & ~n9261;
  assign n9263 = ~n1754 & ~n9262;
  assign n9264 = pi858 & n9254;
  assign n9265 = ~pi858 & ~n9254;
  assign n9266 = ~n9264 & ~n9265;
  assign n9267 = n1754 & n9266;
  assign po479 = n9263 | n9267;
  assign n9269 = pi331 & n1761;
  assign n9270 = pi689 & ~n6579;
  assign n9271 = pi549 & n6579;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = ~n2449 & ~n9272;
  assign n9274 = pi078 & n2449;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = pi562 & n9275;
  assign n9277 = pi549 & n6592;
  assign n9278 = pi078 & n6594;
  assign n9279 = ~n6594 & ~n9275;
  assign n9280 = ~n9278 & ~n9279;
  assign n9281 = ~n6592 & ~n9280;
  assign n9282 = ~n9277 & ~n9281;
  assign n9283 = n6591 & ~n9282;
  assign n9284 = pi078 & ~pi669;
  assign n9285 = ~n6591 & n9284;
  assign n9286 = n6603 & ~n9282;
  assign n9287 = ~n9285 & ~n9286;
  assign n9288 = ~n9283 & n9287;
  assign n9289 = n2564 & ~n9288;
  assign n9290 = pi078 & ~n2564;
  assign n9291 = ~n9289 & ~n9290;
  assign n9292 = ~pi562 & n9291;
  assign n9293 = ~n9276 & ~n9292;
  assign n9294 = pi004 & n9293;
  assign n9295 = ~pi004 & ~n9293;
  assign n9296 = ~n9294 & ~n9295;
  assign n9297 = n6578 & n9296;
  assign n9298 = pi331 & ~n6578;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = ~n1761 & ~n9299;
  assign n9301 = ~n9269 & ~n9300;
  assign n9302 = ~n1754 & ~n9301;
  assign n9303 = pi817 & n9293;
  assign n9304 = ~pi817 & ~n9293;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = n1754 & n9305;
  assign po480 = n9302 | n9306;
  assign n9308 = pi332 & ~po814;
  assign n9309 = po814 & ~n5445;
  assign po481 = n9308 | n9309;
  assign n9311 = pi333 & ~po814;
  assign n9312 = po814 & ~n5395;
  assign po482 = n9311 | n9312;
  assign n9314 = pi334 & ~po814;
  assign n9315 = po814 & ~n6228;
  assign po483 = n9314 | n9315;
  assign n9317 = pi335 & ~po814;
  assign n9318 = po814 & ~n6276;
  assign po484 = n9317 | n9318;
  assign n9320 = pi336 & ~po814;
  assign n9321 = po814 & ~n6468;
  assign po485 = n9320 | n9321;
  assign n9323 = pi337 & ~po814;
  assign n9324 = po814 & ~n6372;
  assign po486 = n9323 | n9324;
  assign n9326 = pi338 & ~po814;
  assign n9327 = po814 & ~n6324;
  assign po487 = n9326 | n9327;
  assign n9329 = pi339 & ~po814;
  assign n9330 = po814 & ~n6420;
  assign po488 = n9329 | n9330;
  assign n9332 = pi340 & n1761;
  assign n9333 = pi701 & ~n6579;
  assign n9334 = pi509 & n6579;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = ~n2449 & ~n9335;
  assign n9337 = pi122 & n2449;
  assign n9338 = ~n9336 & ~n9337;
  assign n9339 = pi562 & n9338;
  assign n9340 = pi509 & n6592;
  assign n9341 = pi122 & n6594;
  assign n9342 = ~n6594 & ~n9338;
  assign n9343 = ~n9341 & ~n9342;
  assign n9344 = ~n6592 & ~n9343;
  assign n9345 = ~n9340 & ~n9344;
  assign n9346 = n6591 & ~n9345;
  assign n9347 = pi122 & ~pi669;
  assign n9348 = ~n6591 & n9347;
  assign n9349 = n6603 & ~n9345;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n9346 & n9350;
  assign n9352 = n2564 & ~n9351;
  assign n9353 = pi122 & ~n2564;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = ~pi562 & n9354;
  assign n9356 = ~n9339 & ~n9355;
  assign n9357 = pi197 & n9356;
  assign n9358 = ~pi197 & ~n9356;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = n6578 & n9359;
  assign n9361 = pi340 & ~n6578;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = ~n1761 & ~n9362;
  assign n9364 = ~n9332 & ~n9363;
  assign n9365 = ~n1754 & ~n9364;
  assign n9366 = pi829 & n9356;
  assign n9367 = ~pi829 & ~n9356;
  assign n9368 = ~n9366 & ~n9367;
  assign n9369 = n1754 & n9368;
  assign po489 = n9365 | n9369;
  assign n9371 = pi341 & n1761;
  assign n9372 = pi749 & ~n6579;
  assign n9373 = pi644 & n6579;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = ~n2449 & ~n9374;
  assign n9376 = pi082 & n2449;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = pi562 & n9377;
  assign n9379 = pi644 & n6592;
  assign n9380 = pi082 & n6594;
  assign n9381 = ~n6594 & ~n9377;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = ~n6592 & ~n9382;
  assign n9384 = ~n9379 & ~n9383;
  assign n9385 = n6591 & ~n9384;
  assign n9386 = pi082 & ~pi669;
  assign n9387 = ~n6591 & n9386;
  assign n9388 = n6603 & ~n9384;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n9385 & n9389;
  assign n9391 = n2564 & ~n9390;
  assign n9392 = pi082 & ~n2564;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = ~pi562 & n9393;
  assign n9395 = ~n9378 & ~n9394;
  assign n9396 = pi045 & n9395;
  assign n9397 = ~pi045 & ~n9395;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = n6578 & n9398;
  assign n9400 = pi341 & ~n6578;
  assign n9401 = ~n9399 & ~n9400;
  assign n9402 = ~n1761 & ~n9401;
  assign n9403 = ~n9371 & ~n9402;
  assign n9404 = ~n1754 & ~n9403;
  assign n9405 = pi877 & n9395;
  assign n9406 = ~pi877 & ~n9395;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = n1754 & n9407;
  assign po490 = n9404 | n9408;
  assign n9410 = pi342 & n1761;
  assign n9411 = pi774 & ~n6579;
  assign n9412 = pi664 & n6579;
  assign n9413 = ~n9411 & ~n9412;
  assign n9414 = ~n2449 & ~n9413;
  assign n9415 = pi112 & n2449;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = pi562 & n9416;
  assign n9418 = pi664 & n6592;
  assign n9419 = pi112 & n6594;
  assign n9420 = ~n6594 & ~n9416;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n6592 & ~n9421;
  assign n9423 = ~n9418 & ~n9422;
  assign n9424 = n6591 & ~n9423;
  assign n9425 = pi112 & ~pi669;
  assign n9426 = ~n6591 & n9425;
  assign n9427 = n6603 & ~n9423;
  assign n9428 = ~n9426 & ~n9427;
  assign n9429 = ~n9424 & n9428;
  assign n9430 = n2564 & ~n9429;
  assign n9431 = pi112 & ~n2564;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = ~pi562 & n9432;
  assign n9434 = ~n9417 & ~n9433;
  assign n9435 = pi415 & n9434;
  assign n9436 = ~pi415 & ~n9434;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = n6578 & n9437;
  assign n9439 = pi342 & ~n6578;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = ~n1761 & ~n9440;
  assign n9442 = ~n9410 & ~n9441;
  assign n9443 = ~n1754 & ~n9442;
  assign n9444 = pi902 & n9434;
  assign n9445 = ~pi902 & ~n9434;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = n1754 & n9446;
  assign po491 = n9443 | n9447;
  assign n9449 = pi343 & n1761;
  assign n9450 = pi707 & ~n6579;
  assign n9451 = pi587 & n6579;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = ~n2449 & ~n9452;
  assign n9454 = pi182 & n2449;
  assign n9455 = ~n9453 & ~n9454;
  assign n9456 = pi562 & n9455;
  assign n9457 = pi587 & n6592;
  assign n9458 = pi182 & n6594;
  assign n9459 = ~n6594 & ~n9455;
  assign n9460 = ~n9458 & ~n9459;
  assign n9461 = ~n6592 & ~n9460;
  assign n9462 = ~n9457 & ~n9461;
  assign n9463 = n6591 & ~n9462;
  assign n9464 = pi182 & ~pi669;
  assign n9465 = ~n6591 & n9464;
  assign n9466 = n6603 & ~n9462;
  assign n9467 = ~n9465 & ~n9466;
  assign n9468 = ~n9463 & n9467;
  assign n9469 = n2564 & ~n9468;
  assign n9470 = pi182 & ~n2564;
  assign n9471 = ~n9469 & ~n9470;
  assign n9472 = ~pi562 & n9471;
  assign n9473 = ~n9456 & ~n9472;
  assign n9474 = ~pi230 & n9473;
  assign n9475 = pi230 & ~n9473;
  assign n9476 = ~n9474 & ~n9475;
  assign n9477 = n6578 & n9476;
  assign n9478 = pi343 & ~n6578;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = ~n1761 & ~n9479;
  assign n9481 = ~n9449 & ~n9480;
  assign n9482 = ~n1754 & ~n9481;
  assign n9483 = pi835 & n9473;
  assign n9484 = ~pi835 & ~n9473;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = n1754 & n9485;
  assign po492 = n9482 | n9486;
  assign n9488 = pi344 & n1761;
  assign n9489 = pi777 & ~n6579;
  assign n9490 = pi611 & n6579;
  assign n9491 = ~n9489 & ~n9490;
  assign n9492 = ~n2449 & ~n9491;
  assign n9493 = pi085 & n2449;
  assign n9494 = ~n9492 & ~n9493;
  assign n9495 = pi562 & n9494;
  assign n9496 = pi611 & n6592;
  assign n9497 = pi085 & n6594;
  assign n9498 = ~n6594 & ~n9494;
  assign n9499 = ~n9497 & ~n9498;
  assign n9500 = ~n6592 & ~n9499;
  assign n9501 = ~n9496 & ~n9500;
  assign n9502 = n6591 & ~n9501;
  assign n9503 = pi085 & ~pi669;
  assign n9504 = ~n6591 & n9503;
  assign n9505 = n6603 & ~n9501;
  assign n9506 = ~n9504 & ~n9505;
  assign n9507 = ~n9502 & n9506;
  assign n9508 = n2564 & ~n9507;
  assign n9509 = pi085 & ~n2564;
  assign n9510 = ~n9508 & ~n9509;
  assign n9511 = ~pi562 & n9510;
  assign n9512 = ~n9495 & ~n9511;
  assign n9513 = pi418 & n9512;
  assign n9514 = ~pi418 & ~n9512;
  assign n9515 = ~n9513 & ~n9514;
  assign n9516 = n6578 & n9515;
  assign n9517 = pi344 & ~n6578;
  assign n9518 = ~n9516 & ~n9517;
  assign n9519 = ~n1761 & ~n9518;
  assign n9520 = ~n9488 & ~n9519;
  assign n9521 = ~n1754 & ~n9520;
  assign n9522 = pi905 & n9512;
  assign n9523 = ~pi905 & ~n9512;
  assign n9524 = ~n9522 & ~n9523;
  assign n9525 = n1754 & n9524;
  assign po493 = n9521 | n9525;
  assign n9527 = pi345 & n1761;
  assign n9528 = pi772 & ~n6579;
  assign n9529 = pi579 & n6579;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = ~n2449 & ~n9530;
  assign n9532 = pi152 & n2449;
  assign n9533 = ~n9531 & ~n9532;
  assign n9534 = pi562 & n9533;
  assign n9535 = pi579 & n6592;
  assign n9536 = pi152 & n6594;
  assign n9537 = ~n6594 & ~n9533;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = ~n6592 & ~n9538;
  assign n9540 = ~n9535 & ~n9539;
  assign n9541 = n6591 & ~n9540;
  assign n9542 = pi152 & ~pi669;
  assign n9543 = ~n6591 & n9542;
  assign n9544 = n6603 & ~n9540;
  assign n9545 = ~n9543 & ~n9544;
  assign n9546 = ~n9541 & n9545;
  assign n9547 = n2564 & ~n9546;
  assign n9548 = pi152 & ~n2564;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~pi562 & n9549;
  assign n9551 = ~n9534 & ~n9550;
  assign n9552 = pi414 & n9551;
  assign n9553 = ~pi414 & ~n9551;
  assign n9554 = ~n9552 & ~n9553;
  assign n9555 = n6578 & n9554;
  assign n9556 = pi345 & ~n6578;
  assign n9557 = ~n9555 & ~n9556;
  assign n9558 = ~n1761 & ~n9557;
  assign n9559 = ~n9527 & ~n9558;
  assign n9560 = ~n1754 & ~n9559;
  assign n9561 = pi900 & n9551;
  assign n9562 = ~pi900 & ~n9551;
  assign n9563 = ~n9561 & ~n9562;
  assign n9564 = n1754 & n9563;
  assign po494 = n9560 | n9564;
  assign n9566 = pi346 & n1761;
  assign n9567 = pi709 & ~n6579;
  assign n9568 = pi663 & n6579;
  assign n9569 = ~n9567 & ~n9568;
  assign n9570 = ~n2449 & ~n9569;
  assign n9571 = pi115 & n2449;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = pi562 & n9572;
  assign n9574 = pi663 & n6592;
  assign n9575 = pi115 & n6594;
  assign n9576 = ~n6594 & ~n9572;
  assign n9577 = ~n9575 & ~n9576;
  assign n9578 = ~n6592 & ~n9577;
  assign n9579 = ~n9574 & ~n9578;
  assign n9580 = n6591 & ~n9579;
  assign n9581 = pi115 & ~pi669;
  assign n9582 = ~n6591 & n9581;
  assign n9583 = n6603 & ~n9579;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = ~n9580 & n9584;
  assign n9586 = n2564 & ~n9585;
  assign n9587 = pi115 & ~n2564;
  assign n9588 = ~n9586 & ~n9587;
  assign n9589 = ~pi562 & n9588;
  assign n9590 = ~n9573 & ~n9589;
  assign n9591 = ~pi232 & n9590;
  assign n9592 = pi232 & ~n9590;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = n6578 & n9593;
  assign n9595 = pi346 & ~n6578;
  assign n9596 = ~n9594 & ~n9595;
  assign n9597 = ~n1761 & ~n9596;
  assign n9598 = ~n9566 & ~n9597;
  assign n9599 = ~n1754 & ~n9598;
  assign n9600 = pi837 & n9590;
  assign n9601 = ~pi837 & ~n9590;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = n1754 & n9602;
  assign po495 = n9599 | n9603;
  assign n9605 = ~pi560 & ~pi561;
  assign n9606 = ~pi669 & ~pi673;
  assign n9607 = pi435 & n2449;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~pi562 & ~n6591;
  assign n9610 = ~n9608 & ~n9609;
  assign n9611 = n9605 & n9610;
  assign n9612 = pi300 & n2449;
  assign n9613 = pi120 & ~n2449;
  assign n9614 = ~n9612 & ~n9613;
  assign n9615 = n9611 & ~n9614;
  assign n9616 = pi316 & n2449;
  assign n9617 = pi130 & ~n2449;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = pi560 & ~pi561;
  assign n9620 = ~n9618 & n9619;
  assign n9621 = ~n9615 & ~n9620;
  assign n9622 = ~pi560 & pi561;
  assign n9623 = pi126 & ~n2449;
  assign n9624 = pi253 & n2449;
  assign n9625 = ~n9623 & ~n9624;
  assign n9626 = n9622 & ~n9625;
  assign po815 = pi560 & pi561;
  assign n9628 = pi123 & ~n2449;
  assign n9629 = pi309 & n2449;
  assign n9630 = ~n9628 & ~n9629;
  assign n9631 = po815 & ~n9630;
  assign n9632 = ~n9626 & ~n9631;
  assign n9633 = n9621 & n9632;
  assign n9634 = pi384 & n2449;
  assign n9635 = pi095 & ~n2449;
  assign n9636 = ~n9634 & ~n9635;
  assign n9637 = n9622 & ~n9636;
  assign n9638 = pi365 & n2449;
  assign n9639 = pi087 & ~n2449;
  assign n9640 = ~n9638 & ~n9639;
  assign n9641 = n9611 & ~n9640;
  assign n9642 = pi355 & n2449;
  assign n9643 = pi089 & ~n2449;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = po815 & ~n9644;
  assign n9646 = ~n9641 & ~n9645;
  assign n9647 = pi371 & n2449;
  assign n9648 = pi103 & ~n2449;
  assign n9649 = ~n9647 & ~n9648;
  assign n9650 = n9619 & ~n9649;
  assign n9651 = n9646 & ~n9650;
  assign n9652 = ~n9637 & n9651;
  assign n9653 = pi079 & ~n2449;
  assign n9654 = pi275 & n2449;
  assign n9655 = ~n9653 & ~n9654;
  assign n9656 = n9622 & ~n9655;
  assign n9657 = pi276 & n2449;
  assign n9658 = pi074 & ~n2449;
  assign n9659 = ~n9657 & ~n9658;
  assign n9660 = n9611 & ~n9659;
  assign n9661 = ~n9656 & ~n9660;
  assign n9662 = pi257 & n2449;
  assign n9663 = pi083 & ~n2449;
  assign n9664 = ~n9662 & ~n9663;
  assign n9665 = n9619 & ~n9664;
  assign n9666 = pi327 & n2449;
  assign n9667 = pi077 & ~n2449;
  assign n9668 = ~n9666 & ~n9667;
  assign n9669 = po815 & ~n9668;
  assign n9670 = ~n9665 & ~n9669;
  assign n9671 = n9661 & n9670;
  assign n9672 = n9652 & n9671;
  assign n9673 = ~n9652 & ~n9671;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = ~n9633 & ~n9674;
  assign n9676 = n9633 & n9674;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = pi346 & n2449;
  assign n9679 = pi115 & ~n2449;
  assign n9680 = ~n9678 & ~n9679;
  assign n9681 = n9622 & ~n9680;
  assign n9682 = pi099 & ~n2449;
  assign n9683 = pi357 & n2449;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = n9619 & ~n9684;
  assign n9686 = ~n9681 & ~n9685;
  assign n9687 = pi270 & n2449;
  assign n9688 = pi100 & ~n2449;
  assign n9689 = ~n9687 & ~n9688;
  assign n9690 = po815 & ~n9689;
  assign n9691 = pi379 & n2449;
  assign n9692 = pi118 & ~n2449;
  assign n9693 = ~n9691 & ~n9692;
  assign n9694 = n9611 & ~n9693;
  assign n9695 = ~n9690 & ~n9694;
  assign n9696 = n9686 & n9695;
  assign n9697 = pi125 & ~n2449;
  assign n9698 = pi287 & n2449;
  assign n9699 = ~n9697 & ~n9698;
  assign n9700 = n9622 & ~n9699;
  assign n9701 = pi315 & n2449;
  assign n9702 = pi129 & ~n2449;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = n9619 & ~n9703;
  assign n9705 = ~n9700 & ~n9704;
  assign n9706 = pi340 & n2449;
  assign n9707 = pi122 & ~n2449;
  assign n9708 = ~n9706 & ~n9707;
  assign n9709 = po815 & ~n9708;
  assign n9710 = pi272 & n2449;
  assign n9711 = pi119 & ~n2449;
  assign n9712 = ~n9710 & ~n9711;
  assign n9713 = n9611 & ~n9712;
  assign n9714 = ~n9709 & ~n9713;
  assign n9715 = n9705 & n9714;
  assign n9716 = ~n9696 & n9715;
  assign n9717 = n9696 & ~n9715;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = pi127 & ~n2449;
  assign n9720 = pi255 & n2449;
  assign n9721 = ~n9719 & ~n9720;
  assign n9722 = n9622 & ~n9721;
  assign n9723 = pi121 & ~n2449;
  assign n9724 = pi281 & n2449;
  assign n9725 = ~n9723 & ~n9724;
  assign n9726 = n9611 & ~n9725;
  assign n9727 = ~n9722 & ~n9726;
  assign n9728 = pi313 & n2449;
  assign n9729 = pi124 & ~n2449;
  assign n9730 = ~n9728 & ~n9729;
  assign n9731 = po815 & ~n9730;
  assign n9732 = pi321 & n2449;
  assign n9733 = pi128 & ~n2449;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = n9619 & ~n9734;
  assign n9736 = ~n9731 & ~n9735;
  assign n9737 = n9727 & n9736;
  assign n9738 = pi308 & n2449;
  assign n9739 = pi101 & ~n2449;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = po815 & ~n9740;
  assign n9742 = pi085 & ~n2449;
  assign n9743 = pi344 & n2449;
  assign n9744 = ~n9742 & ~n9743;
  assign n9745 = n9611 & ~n9744;
  assign n9746 = ~n9741 & ~n9745;
  assign n9747 = pi399 & n2449;
  assign n9748 = pi102 & ~n2449;
  assign n9749 = ~n9747 & ~n9748;
  assign n9750 = n9619 & ~n9749;
  assign n9751 = pi116 & ~n2449;
  assign n9752 = pi382 & n2449;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = n9622 & ~n9753;
  assign n9755 = ~n9750 & ~n9754;
  assign n9756 = n9746 & n9755;
  assign n9757 = ~n9737 & n9756;
  assign n9758 = n9737 & ~n9756;
  assign n9759 = ~n9757 & ~n9758;
  assign n9760 = ~n9718 & n9759;
  assign n9761 = n9718 & ~n9759;
  assign n9762 = ~n9760 & ~n9761;
  assign n9763 = ~n9677 & n9762;
  assign n9764 = n9677 & ~n9762;
  assign n9765 = ~n9763 & ~n9764;
  assign n9766 = ~pi673 & ~n9765;
  assign n9767 = pi354 & n2449;
  assign n9768 = pi174 & ~n2449;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = n9619 & ~n9769;
  assign n9771 = pi377 & n2449;
  assign n9772 = pi175 & ~n2449;
  assign n9773 = ~n9771 & ~n9772;
  assign n9774 = n9611 & ~n9773;
  assign n9775 = pi182 & ~n2449;
  assign n9776 = pi343 & n2449;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = n9622 & ~n9777;
  assign n9779 = ~pi173 & ~n2449;
  assign n9780 = pi303 & n2449;
  assign n9781 = ~n9779 & ~n9780;
  assign n9782 = po815 & ~n9781;
  assign n9783 = ~n9778 & ~n9782;
  assign n9784 = ~n9774 & n9783;
  assign n9785 = ~n9770 & n9784;
  assign n9786 = ~pi185 & ~n2449;
  assign n9787 = pi258 & n2449;
  assign n9788 = ~n9786 & ~n9787;
  assign n9789 = po815 & ~n9788;
  assign n9790 = ~pi183 & ~n2449;
  assign n9791 = pi286 & n2449;
  assign n9792 = ~n9790 & ~n9791;
  assign n9793 = n9622 & ~n9792;
  assign n9794 = ~n9789 & ~n9793;
  assign n9795 = pi392 & n2449;
  assign n9796 = ~pi184 & ~n2449;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = n9619 & ~n9797;
  assign n9799 = n9794 & ~n9798;
  assign n9800 = pi324 & n2449;
  assign n9801 = ~pi187 & ~n2449;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = n9611 & ~n9802;
  assign n9804 = n9799 & ~n9803;
  assign n9805 = ~n9785 & n9804;
  assign n9806 = n9785 & ~n9804;
  assign n9807 = ~n9805 & ~n9806;
  assign n9808 = pi169 & ~n2449;
  assign n9809 = pi271 & n2449;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = n9622 & ~n9810;
  assign n9812 = pi265 & n2449;
  assign n9813 = pi168 & ~n2449;
  assign n9814 = ~n9812 & ~n9813;
  assign n9815 = n9611 & ~n9814;
  assign n9816 = ~n9811 & ~n9815;
  assign n9817 = pi304 & n2449;
  assign n9818 = pi170 & ~n2449;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = n9619 & ~n9819;
  assign n9821 = pi323 & n2449;
  assign n9822 = pi171 & ~n2449;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = po815 & ~n9823;
  assign n9825 = ~n9820 & ~n9824;
  assign n9826 = n9816 & n9825;
  assign n9827 = pi180 & ~n2449;
  assign n9828 = pi383 & n2449;
  assign n9829 = ~n9827 & ~n9828;
  assign n9830 = n9622 & ~n9829;
  assign n9831 = pi403 & n2449;
  assign n9832 = pi181 & ~n2449;
  assign n9833 = ~n9831 & ~n9832;
  assign n9834 = n9611 & ~n9833;
  assign n9835 = ~n9830 & ~n9834;
  assign n9836 = pi179 & ~n2449;
  assign n9837 = pi367 & n2449;
  assign n9838 = ~n9836 & ~n9837;
  assign n9839 = n9619 & ~n9838;
  assign n9840 = pi386 & n2449;
  assign n9841 = pi172 & ~n2449;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = po815 & ~n9842;
  assign n9844 = ~n9839 & ~n9843;
  assign n9845 = n9835 & n9844;
  assign n9846 = n9826 & n9845;
  assign n9847 = ~n9826 & ~n9845;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = n9765 & n9848;
  assign n9850 = ~n9765 & ~n9848;
  assign n9851 = ~n9849 & ~n9850;
  assign n9852 = ~n9807 & n9851;
  assign n9853 = n9807 & ~n9851;
  assign n9854 = ~n9852 & ~n9853;
  assign n9855 = pi356 & n2449;
  assign n9856 = pi150 & ~n2449;
  assign n9857 = ~n9855 & ~n9856;
  assign n9858 = n9619 & ~n9857;
  assign n9859 = pi312 & n2449;
  assign n9860 = pi148 & ~n2449;
  assign n9861 = ~n9859 & ~n9860;
  assign n9862 = po815 & ~n9861;
  assign n9863 = ~n9858 & ~n9862;
  assign n9864 = pi158 & ~n2449;
  assign n9865 = pi317 & n2449;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n9622 & ~n9866;
  assign n9868 = pi345 & n2449;
  assign n9869 = pi152 & ~n2449;
  assign n9870 = ~n9868 & ~n9869;
  assign n9871 = n9611 & ~n9870;
  assign n9872 = ~n9867 & ~n9871;
  assign n9873 = n9863 & n9872;
  assign n9874 = pi147 & ~n2449;
  assign n9875 = pi407 & n2449;
  assign n9876 = ~n9874 & ~n9875;
  assign n9877 = po815 & ~n9876;
  assign n9878 = pi397 & n2449;
  assign n9879 = pi143 & ~n2449;
  assign n9880 = ~n9878 & ~n9879;
  assign n9881 = n9611 & ~n9880;
  assign n9882 = ~n9877 & ~n9881;
  assign n9883 = pi149 & ~n2449;
  assign n9884 = pi406 & n2449;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = n9622 & ~n9885;
  assign n9887 = pi395 & n2449;
  assign n9888 = pi151 & ~n2449;
  assign n9889 = ~n9887 & ~n9888;
  assign n9890 = n9619 & ~n9889;
  assign n9891 = ~n9886 & ~n9890;
  assign n9892 = n9882 & n9891;
  assign n9893 = ~n9873 & n9892;
  assign n9894 = n9873 & ~n9892;
  assign n9895 = ~n9893 & ~n9894;
  assign n9896 = pi088 & ~n2449;
  assign n9897 = pi375 & n2449;
  assign n9898 = ~n9896 & ~n9897;
  assign n9899 = n9611 & ~n9898;
  assign n9900 = pi363 & n2449;
  assign n9901 = pi091 & ~n2449;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = po815 & ~n9902;
  assign n9904 = pi096 & ~n2449;
  assign n9905 = pi385 & n2449;
  assign n9906 = ~n9904 & ~n9905;
  assign n9907 = n9622 & ~n9906;
  assign n9908 = ~n9903 & ~n9907;
  assign n9909 = pi372 & n2449;
  assign n9910 = pi105 & ~n2449;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = n9619 & ~n9911;
  assign n9913 = n9908 & ~n9912;
  assign n9914 = ~n9899 & n9913;
  assign n9915 = ~n9756 & n9914;
  assign n9916 = n9756 & ~n9914;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = pi033 & ~n2449;
  assign n9919 = pi381 & n2449;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = n9622 & ~n9920;
  assign n9922 = pi256 & n2449;
  assign n9923 = pi037 & ~n2449;
  assign n9924 = ~n9922 & ~n9923;
  assign n9925 = po815 & ~n9924;
  assign n9926 = ~n9921 & ~n9925;
  assign n9927 = pi361 & n2449;
  assign n9928 = pi038 & ~n2449;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = n9619 & ~n9929;
  assign n9931 = pi026 & ~n2449;
  assign n9932 = pi362 & n2449;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = n9611 & ~n9933;
  assign n9935 = ~n9930 & ~n9934;
  assign n9936 = n9926 & n9935;
  assign n9937 = pi070 & ~n2449;
  assign n9938 = pi302 & n2449;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = n9622 & ~n9939;
  assign n9941 = pi320 & n2449;
  assign n9942 = pi053 & ~n2449;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = n9619 & ~n9943;
  assign n9945 = ~n9940 & ~n9944;
  assign n9946 = pi311 & n2449;
  assign n9947 = pi054 & ~n2449;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = po815 & ~n9948;
  assign n9950 = pi280 & n2449;
  assign n9951 = pi051 & ~n2449;
  assign n9952 = ~n9950 & ~n9951;
  assign n9953 = n9611 & ~n9952;
  assign n9954 = ~n9949 & ~n9953;
  assign n9955 = n9945 & n9954;
  assign n9956 = ~n9936 & n9955;
  assign n9957 = n9936 & ~n9955;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = pi035 & ~n2449;
  assign n9960 = pi398 & n2449;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = n9622 & ~n9961;
  assign n9963 = pi370 & n2449;
  assign n9964 = pi041 & ~n2449;
  assign n9965 = ~n9963 & ~n9964;
  assign n9966 = n9619 & ~n9965;
  assign n9967 = ~n9962 & ~n9966;
  assign n9968 = pi360 & n2449;
  assign n9969 = pi031 & ~n2449;
  assign n9970 = ~n9968 & ~n9969;
  assign n9971 = po815 & ~n9970;
  assign n9972 = pi028 & ~n2449;
  assign n9973 = pi391 & n2449;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = n9611 & ~n9974;
  assign n9976 = ~n9971 & ~n9975;
  assign n9977 = n9967 & n9976;
  assign n9978 = pi023 & ~n2449;
  assign n9979 = pi278 & n2449;
  assign n9980 = ~n9978 & ~n9979;
  assign n9981 = n9622 & ~n9980;
  assign n9982 = pi329 & n2449;
  assign n9983 = pi021 & ~n2449;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = po815 & ~n9984;
  assign n9986 = ~n9981 & ~n9985;
  assign n9987 = pi260 & n2449;
  assign n9988 = pi025 & ~n2449;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = n9619 & ~n9989;
  assign n9991 = pi284 & n2449;
  assign n9992 = pi019 & ~n2449;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = n9611 & ~n9993;
  assign n9995 = ~n9990 & ~n9994;
  assign n9996 = n9986 & n9995;
  assign n9997 = ~n9977 & n9996;
  assign n9998 = n9977 & ~n9996;
  assign n9999 = ~n9997 & ~n9998;
  assign n10000 = ~n9958 & n9999;
  assign n10001 = n9958 & ~n9999;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = ~n9917 & n10002;
  assign n10004 = n9917 & ~n10002;
  assign n10005 = ~n10003 & ~n10004;
  assign n10006 = ~n9936 & n9977;
  assign n10007 = n9936 & ~n9977;
  assign n10008 = ~n10006 & ~n10007;
  assign n10009 = pi358 & n2449;
  assign n10010 = pi030 & ~n2449;
  assign n10011 = ~n10009 & ~n10010;
  assign n10012 = po815 & ~n10011;
  assign n10013 = pi369 & n2449;
  assign n10014 = pi040 & ~n2449;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = n9619 & ~n10015;
  assign n10017 = ~n10012 & ~n10016;
  assign n10018 = pi034 & ~n2449;
  assign n10019 = pi402 & n2449;
  assign n10020 = ~n10018 & ~n10019;
  assign n10021 = n9622 & ~n10020;
  assign n10022 = pi393 & n2449;
  assign n10023 = pi029 & ~n2449;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n9611 & ~n10024;
  assign n10026 = ~n10021 & ~n10025;
  assign n10027 = n10017 & n10026;
  assign n10028 = pi022 & ~n2449;
  assign n10029 = pi325 & n2449;
  assign n10030 = ~n10028 & ~n10029;
  assign n10031 = n9622 & ~n10030;
  assign n10032 = pi283 & n2449;
  assign n10033 = pi020 & ~n2449;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = po815 & ~n10034;
  assign n10036 = ~n10031 & ~n10035;
  assign n10037 = pi024 & ~n2449;
  assign n10038 = pi259 & n2449;
  assign n10039 = ~n10037 & ~n10038;
  assign n10040 = n9619 & ~n10039;
  assign n10041 = pi328 & n2449;
  assign n10042 = pi018 & ~n2449;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = n9611 & ~n10043;
  assign n10045 = ~n10040 & ~n10044;
  assign n10046 = n10036 & n10045;
  assign n10047 = ~n10027 & n10046;
  assign n10048 = n10027 & ~n10046;
  assign n10049 = ~n10047 & ~n10048;
  assign n10050 = pi297 & n2449;
  assign n10051 = pi036 & ~n2449;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = po815 & ~n10052;
  assign n10054 = pi351 & n2449;
  assign n10055 = pi027 & ~n2449;
  assign n10056 = ~n10054 & ~n10055;
  assign n10057 = n9611 & ~n10056;
  assign n10058 = pi032 & ~n2449;
  assign n10059 = pi380 & n2449;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = n9622 & ~n10060;
  assign n10062 = pi039 & ~n2449;
  assign n10063 = pi359 & n2449;
  assign n10064 = ~n10062 & ~n10063;
  assign n10065 = n9619 & ~n10064;
  assign n10066 = ~n10061 & ~n10065;
  assign n10067 = ~n10057 & n10066;
  assign n10068 = ~n10053 & n10067;
  assign n10069 = pi052 & ~n2449;
  assign n10070 = pi263 & n2449;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = po815 & ~n10071;
  assign n10073 = pi069 & ~n2449;
  assign n10074 = pi301 & n2449;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076 = n9622 & ~n10075;
  assign n10077 = ~n10072 & ~n10076;
  assign n10078 = pi318 & n2449;
  assign n10079 = pi055 & ~n2449;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = n9619 & ~n10080;
  assign n10082 = pi277 & n2449;
  assign n10083 = pi050 & ~n2449;
  assign n10084 = ~n10082 & ~n10083;
  assign n10085 = n9611 & ~n10084;
  assign n10086 = ~n10081 & ~n10085;
  assign n10087 = n10077 & n10086;
  assign n10088 = ~n10068 & n10087;
  assign n10089 = n10068 & ~n10087;
  assign n10090 = ~n10088 & ~n10089;
  assign n10091 = ~n10049 & n10090;
  assign n10092 = n10049 & ~n10090;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = ~n10008 & n10093;
  assign n10095 = n10008 & ~n10093;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = ~n10005 & n10096;
  assign n10098 = n10005 & ~n10096;
  assign n10099 = ~n10097 & ~n10098;
  assign n10100 = ~n9895 & n10099;
  assign n10101 = n9895 & ~n10099;
  assign n10102 = ~n10100 & ~n10101;
  assign n10103 = ~n9854 & n10102;
  assign n10104 = n9854 & ~n10102;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = pi673 & ~n10105;
  assign n10107 = ~n9766 & ~n10106;
  assign n10108 = n9610 & ~n10107;
  assign n10109 = ~pi347 & ~n9610;
  assign n10110 = ~n10108 & ~n10109;
  assign n10111 = n9605 & ~n10110;
  assign n10112 = ~n9619 & ~n9622;
  assign n10113 = ~pi347 & ~n10112;
  assign n10114 = ~n10111 & ~n10113;
  assign n10115 = ~pi347 & po815;
  assign po496 = ~n10114 | n10115;
  assign n10117 = ~pi348 & ~n10112;
  assign n10118 = pi097 & ~n2449;
  assign n10119 = pi378 & n2449;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = n9622 & ~n10120;
  assign n10122 = pi326 & n2449;
  assign n10123 = pi093 & ~n2449;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = po815 & ~n10124;
  assign n10126 = ~n10121 & ~n10125;
  assign n10127 = pi098 & ~n2449;
  assign n10128 = pi401 & n2449;
  assign n10129 = ~n10127 & ~n10128;
  assign n10130 = n9619 & ~n10129;
  assign n10131 = pi342 & n2449;
  assign n10132 = pi112 & ~n2449;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = n9611 & ~n10133;
  assign n10135 = ~n10130 & ~n10134;
  assign n10136 = n10126 & n10135;
  assign n10137 = ~n9633 & n9652;
  assign n10138 = n9633 & ~n9652;
  assign n10139 = ~n10137 & ~n10138;
  assign n10140 = ~n10136 & n10139;
  assign n10141 = n10136 & ~n10139;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = pi341 & n2449;
  assign n10144 = pi082 & ~n2449;
  assign n10145 = ~n10143 & ~n10144;
  assign n10146 = n9619 & ~n10145;
  assign n10147 = pi080 & ~n2449;
  assign n10148 = pi274 & n2449;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = n9622 & ~n10149;
  assign n10151 = pi319 & n2449;
  assign n10152 = pi076 & ~n2449;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = po815 & ~n10153;
  assign n10155 = ~n10150 & ~n10154;
  assign n10156 = pi268 & n2449;
  assign n10157 = pi073 & ~n2449;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = n9611 & ~n10158;
  assign n10160 = n10155 & ~n10159;
  assign n10161 = ~n10146 & n10160;
  assign n10162 = n9696 & ~n10161;
  assign n10163 = ~n9696 & n10161;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = pi279 & n2449;
  assign n10166 = pi081 & ~n2449;
  assign n10167 = ~n10165 & ~n10166;
  assign n10168 = n9622 & ~n10167;
  assign n10169 = pi261 & n2449;
  assign n10170 = pi084 & ~n2449;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = n9619 & ~n10171;
  assign n10173 = ~n10168 & ~n10172;
  assign n10174 = pi331 & n2449;
  assign n10175 = pi078 & ~n2449;
  assign n10176 = ~n10174 & ~n10175;
  assign n10177 = po815 & ~n10176;
  assign n10178 = pi075 & ~n2449;
  assign n10179 = pi254 & n2449;
  assign n10180 = ~n10178 & ~n10179;
  assign n10181 = n9611 & ~n10180;
  assign n10182 = ~n10177 & ~n10181;
  assign n10183 = n10173 & n10182;
  assign n10184 = n9756 & ~n10183;
  assign n10185 = ~n9756 & n10183;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = ~n10164 & n10186;
  assign n10188 = n10164 & ~n10186;
  assign n10189 = ~n10187 & ~n10188;
  assign n10190 = ~n10142 & n10189;
  assign n10191 = n10142 & ~n10189;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = ~pi673 & ~n10192;
  assign n10194 = n9785 & n9826;
  assign n10195 = ~n9785 & ~n9826;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = n9804 & ~n9845;
  assign n10198 = ~n9804 & n9845;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = n10192 & ~n10199;
  assign n10201 = ~n10192 & n10199;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = n10196 & n10202;
  assign n10204 = ~n10196 & ~n10202;
  assign n10205 = ~n10203 & ~n10204;
  assign n10206 = pi162 & ~n2449;
  assign n10207 = pi285 & n2449;
  assign n10208 = ~n10206 & ~n10207;
  assign n10209 = n9622 & ~n10208;
  assign n10210 = pi314 & n2449;
  assign n10211 = pi163 & ~n2449;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = n9619 & ~n10212;
  assign n10214 = ~n10209 & ~n10213;
  assign n10215 = pi161 & ~n2449;
  assign n10216 = pi262 & n2449;
  assign n10217 = ~n10215 & ~n10216;
  assign n10218 = po815 & ~n10217;
  assign n10219 = pi269 & n2449;
  assign n10220 = pi160 & ~n2449;
  assign n10221 = ~n10219 & ~n10220;
  assign n10222 = n9611 & ~n10221;
  assign n10223 = ~n10218 & ~n10222;
  assign n10224 = n10214 & n10223;
  assign n10225 = pi141 & ~n2449;
  assign n10226 = pi305 & n2449;
  assign n10227 = ~n10225 & ~n10226;
  assign n10228 = n9619 & ~n10227;
  assign n10229 = pi267 & n2449;
  assign n10230 = pi139 & ~n2449;
  assign n10231 = ~n10229 & ~n10230;
  assign n10232 = n9611 & ~n10231;
  assign n10233 = ~n10228 & ~n10232;
  assign n10234 = pi142 & ~n2449;
  assign n10235 = pi273 & n2449;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = n9622 & ~n10236;
  assign n10238 = pi282 & n2449;
  assign n10239 = pi140 & ~n2449;
  assign n10240 = ~n10238 & ~n10239;
  assign n10241 = po815 & ~n10240;
  assign n10242 = ~n10237 & ~n10241;
  assign n10243 = n10233 & n10242;
  assign n10244 = ~n10224 & n10243;
  assign n10245 = n10224 & ~n10243;
  assign n10246 = ~n10244 & ~n10245;
  assign n10247 = n9737 & ~n10183;
  assign n10248 = ~n9737 & n10183;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = n9936 & ~n9996;
  assign n10251 = ~n9936 & n9996;
  assign n10252 = ~n10250 & ~n10251;
  assign n10253 = n9955 & ~n9977;
  assign n10254 = ~n9955 & n9977;
  assign n10255 = ~n10253 & ~n10254;
  assign n10256 = ~n10252 & n10255;
  assign n10257 = n10252 & ~n10255;
  assign n10258 = ~n10256 & ~n10257;
  assign n10259 = ~n10249 & n10258;
  assign n10260 = n10249 & ~n10258;
  assign n10261 = ~n10259 & ~n10260;
  assign n10262 = n9955 & ~n9996;
  assign n10263 = ~n9955 & n9996;
  assign n10264 = ~n10262 & ~n10263;
  assign n10265 = n10046 & ~n10068;
  assign n10266 = ~n10046 & n10068;
  assign n10267 = ~n10265 & ~n10266;
  assign n10268 = n10027 & ~n10087;
  assign n10269 = ~n10027 & n10087;
  assign n10270 = ~n10268 & ~n10269;
  assign n10271 = ~n10267 & n10270;
  assign n10272 = n10267 & ~n10270;
  assign n10273 = ~n10271 & ~n10272;
  assign n10274 = ~n10264 & n10273;
  assign n10275 = n10264 & ~n10273;
  assign n10276 = ~n10274 & ~n10275;
  assign n10277 = n10261 & n10276;
  assign n10278 = ~n10261 & ~n10276;
  assign n10279 = ~n10277 & ~n10278;
  assign n10280 = ~n10246 & ~n10279;
  assign n10281 = n10246 & n10279;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = ~n10205 & n10282;
  assign n10284 = n10205 & ~n10282;
  assign n10285 = ~n10283 & ~n10284;
  assign n10286 = pi673 & ~n10285;
  assign n10287 = ~n10193 & ~n10286;
  assign n10288 = n9610 & ~n10287;
  assign n10289 = ~pi348 & ~n9610;
  assign n10290 = ~n10288 & ~n10289;
  assign n10291 = n9605 & ~n10290;
  assign n10292 = ~n10117 & ~n10291;
  assign n10293 = ~pi348 & po815;
  assign po497 = ~n10292 | n10293;
  assign n10295 = ~pi349 & ~n10112;
  assign n10296 = n9633 & n10136;
  assign n10297 = ~n9633 & ~n10136;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n9671 & ~n10298;
  assign n10300 = n9671 & n10298;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = pi094 & ~n2449;
  assign n10303 = pi405 & n2449;
  assign n10304 = ~n10302 & ~n10303;
  assign n10305 = n9622 & ~n10304;
  assign n10306 = pi404 & n2449;
  assign n10307 = pi090 & ~n2449;
  assign n10308 = ~n10306 & ~n10307;
  assign n10309 = po815 & ~n10308;
  assign n10310 = ~n10305 & ~n10309;
  assign n10311 = pi104 & ~n2449;
  assign n10312 = pi368 & n2449;
  assign n10313 = ~n10311 & ~n10312;
  assign n10314 = n9619 & ~n10313;
  assign n10315 = pi364 & n2449;
  assign n10316 = pi086 & ~n2449;
  assign n10317 = ~n10315 & ~n10316;
  assign n10318 = n9611 & ~n10317;
  assign n10319 = ~n10314 & ~n10318;
  assign n10320 = n10310 & n10319;
  assign n10321 = n10161 & n10320;
  assign n10322 = ~n10161 & ~n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = n9914 & ~n10183;
  assign n10325 = ~n9914 & n10183;
  assign n10326 = ~n10324 & ~n10325;
  assign n10327 = n10323 & n10326;
  assign n10328 = ~n10323 & ~n10326;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~n10301 & n10329;
  assign n10331 = n10301 & ~n10329;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~pi673 & ~n10332;
  assign n10334 = ~n9807 & n10332;
  assign n10335 = n9807 & ~n10332;
  assign n10336 = ~n10334 & ~n10335;
  assign n10337 = n9848 & n10336;
  assign n10338 = ~n9848 & ~n10336;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = n10102 & ~n10339;
  assign n10341 = ~n10102 & n10339;
  assign n10342 = ~n10340 & ~n10341;
  assign n10343 = pi673 & ~n10342;
  assign n10344 = ~n10333 & ~n10343;
  assign n10345 = n9610 & ~n10344;
  assign n10346 = ~pi349 & ~n9610;
  assign n10347 = ~n10345 & ~n10346;
  assign n10348 = n9605 & ~n10347;
  assign n10349 = ~n10295 & ~n10348;
  assign n10350 = ~pi349 & po815;
  assign po498 = ~n10349 | n10350;
  assign n10352 = ~pi350 & ~n10112;
  assign n10353 = ~n9671 & n10136;
  assign n10354 = n9671 & ~n10136;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = ~n9652 & n10355;
  assign n10357 = n9652 & ~n10355;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n9715 & n10320;
  assign n10360 = n9715 & ~n10320;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = n9737 & n9914;
  assign n10363 = ~n9737 & ~n9914;
  assign n10364 = ~n10362 & ~n10363;
  assign n10365 = ~n10361 & ~n10364;
  assign n10366 = n10361 & n10364;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = ~n10358 & n10367;
  assign n10369 = n10358 & ~n10367;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = ~pi673 & ~n10370;
  assign n10372 = n10196 & n10370;
  assign n10373 = ~n10196 & ~n10370;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = ~n10199 & n10374;
  assign n10376 = n10199 & ~n10374;
  assign n10377 = ~n10375 & ~n10376;
  assign n10378 = n10282 & ~n10377;
  assign n10379 = ~n10282 & n10377;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = pi673 & ~n10380;
  assign n10382 = ~n10371 & ~n10381;
  assign n10383 = n9610 & ~n10382;
  assign n10384 = ~pi350 & ~n9610;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = n9605 & ~n10385;
  assign n10387 = ~n10352 & ~n10386;
  assign n10388 = ~pi350 & po815;
  assign po499 = ~n10387 | n10388;
  assign n10390 = pi351 & n1761;
  assign n10391 = pi775 & ~n6579;
  assign n10392 = pi628 & n6579;
  assign n10393 = ~n10391 & ~n10392;
  assign n10394 = ~n2449 & ~n10393;
  assign n10395 = pi027 & n2449;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = pi562 & n10396;
  assign n10398 = pi628 & n6592;
  assign n10399 = pi027 & n6594;
  assign n10400 = ~n6594 & ~n10396;
  assign n10401 = ~n10399 & ~n10400;
  assign n10402 = ~n6592 & ~n10401;
  assign n10403 = ~n10398 & ~n10402;
  assign n10404 = n6591 & ~n10403;
  assign n10405 = pi027 & ~pi669;
  assign n10406 = ~n6591 & n10405;
  assign n10407 = n6603 & ~n10403;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = ~n10404 & n10408;
  assign n10410 = n2564 & ~n10409;
  assign n10411 = pi027 & ~n2564;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = ~pi562 & n10412;
  assign n10414 = ~n10397 & ~n10413;
  assign n10415 = pi416 & n10414;
  assign n10416 = ~pi416 & ~n10414;
  assign n10417 = ~n10415 & ~n10416;
  assign n10418 = n6578 & n10417;
  assign n10419 = pi351 & ~n6578;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = ~n1761 & ~n10420;
  assign n10422 = ~n10390 & ~n10421;
  assign n10423 = ~n1754 & ~n10422;
  assign n10424 = pi903 & n10414;
  assign n10425 = ~pi903 & ~n10414;
  assign n10426 = ~n10424 & ~n10425;
  assign n10427 = n1754 & n10426;
  assign po500 = n10423 | n10427;
  assign n10429 = pi352 & n1761;
  assign n10430 = pi786 & ~n6579;
  assign n10431 = pi574 & n6579;
  assign n10432 = ~n10430 & ~n10431;
  assign n10433 = ~n2449 & ~n10432;
  assign n10434 = pi063 & n2449;
  assign n10435 = ~n10433 & ~n10434;
  assign n10436 = pi562 & n10435;
  assign n10437 = pi574 & n6592;
  assign n10438 = pi063 & n6594;
  assign n10439 = ~n6594 & ~n10435;
  assign n10440 = ~n10438 & ~n10439;
  assign n10441 = ~n6592 & ~n10440;
  assign n10442 = ~n10437 & ~n10441;
  assign n10443 = n6591 & ~n10442;
  assign n10444 = pi063 & ~pi669;
  assign n10445 = ~n6591 & n10444;
  assign n10446 = n6603 & ~n10442;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = ~n10443 & n10447;
  assign n10449 = n2564 & ~n10448;
  assign n10450 = pi063 & ~n2564;
  assign n10451 = ~n10449 & ~n10450;
  assign n10452 = ~pi562 & n10451;
  assign n10453 = ~n10436 & ~n10452;
  assign n10454 = pi430 & n10453;
  assign n10455 = ~pi430 & ~n10453;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = n6578 & n10456;
  assign n10458 = pi352 & ~n6578;
  assign n10459 = ~n10457 & ~n10458;
  assign n10460 = ~n1761 & ~n10459;
  assign n10461 = ~n10429 & ~n10460;
  assign n10462 = ~n1754 & ~n10461;
  assign n10463 = pi914 & n10453;
  assign n10464 = ~pi914 & ~n10453;
  assign n10465 = ~n10463 & ~n10464;
  assign n10466 = n1754 & n10465;
  assign po501 = n10462 | n10466;
  assign n10468 = pi353 & n1761;
  assign n10469 = pi738 & ~n6579;
  assign n10470 = pi595 & n6579;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = ~n2449 & ~n10471;
  assign n10473 = pi065 & n2449;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = pi562 & n10474;
  assign n10476 = pi595 & n6592;
  assign n10477 = pi065 & n6594;
  assign n10478 = ~n6594 & ~n10474;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = ~n6592 & ~n10479;
  assign n10481 = ~n10476 & ~n10480;
  assign n10482 = n6591 & ~n10481;
  assign n10483 = pi065 & ~pi669;
  assign n10484 = ~n6591 & n10483;
  assign n10485 = n6603 & ~n10481;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = ~n10482 & n10486;
  assign n10488 = n2564 & ~n10487;
  assign n10489 = pi065 & ~n2564;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = ~pi562 & n10490;
  assign n10492 = ~n10475 & ~n10491;
  assign n10493 = pi289 & n10492;
  assign n10494 = ~pi289 & ~n10492;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = n6578 & n10495;
  assign n10497 = pi353 & ~n6578;
  assign n10498 = ~n10496 & ~n10497;
  assign n10499 = ~n1761 & ~n10498;
  assign n10500 = ~n10468 & ~n10499;
  assign n10501 = ~n1754 & ~n10500;
  assign n10502 = pi866 & n10492;
  assign n10503 = ~pi866 & ~n10492;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = n1754 & n10504;
  assign po502 = n10501 | n10505;
  assign n10507 = pi354 & n1761;
  assign n10508 = pi739 & ~n6579;
  assign n10509 = pi588 & n6579;
  assign n10510 = ~n10508 & ~n10509;
  assign n10511 = ~n2449 & ~n10510;
  assign n10512 = pi174 & n2449;
  assign n10513 = ~n10511 & ~n10512;
  assign n10514 = pi562 & n10513;
  assign n10515 = pi588 & n6592;
  assign n10516 = pi174 & n6594;
  assign n10517 = ~n6594 & ~n10513;
  assign n10518 = ~n10516 & ~n10517;
  assign n10519 = ~n6592 & ~n10518;
  assign n10520 = ~n10515 & ~n10519;
  assign n10521 = n6591 & ~n10520;
  assign n10522 = pi174 & ~pi669;
  assign n10523 = ~n6591 & n10522;
  assign n10524 = n6603 & ~n10520;
  assign n10525 = ~n10523 & ~n10524;
  assign n10526 = ~n10521 & n10525;
  assign n10527 = n2564 & ~n10526;
  assign n10528 = pi174 & ~n2564;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = ~pi562 & n10529;
  assign n10531 = ~n10514 & ~n10530;
  assign n10532 = pi290 & n10531;
  assign n10533 = ~pi290 & ~n10531;
  assign n10534 = ~n10532 & ~n10533;
  assign n10535 = n6578 & n10534;
  assign n10536 = pi354 & ~n6578;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = ~n1761 & ~n10537;
  assign n10539 = ~n10507 & ~n10538;
  assign n10540 = ~n1754 & ~n10539;
  assign n10541 = pi867 & n10531;
  assign n10542 = ~pi867 & ~n10531;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = n1754 & n10543;
  assign po503 = n10540 | n10544;
  assign n10546 = pi355 & n1761;
  assign n10547 = pi694 & ~n6579;
  assign n10548 = pi467 & n6579;
  assign n10549 = ~n10547 & ~n10548;
  assign n10550 = ~n2449 & ~n10549;
  assign n10551 = pi089 & n2449;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = pi562 & n10552;
  assign n10554 = pi467 & n6592;
  assign n10555 = pi089 & n6594;
  assign n10556 = ~n6594 & ~n10552;
  assign n10557 = ~n10555 & ~n10556;
  assign n10558 = ~n6592 & ~n10557;
  assign n10559 = ~n10554 & ~n10558;
  assign n10560 = n6591 & ~n10559;
  assign n10561 = pi089 & ~pi669;
  assign n10562 = ~n6591 & n10561;
  assign n10563 = n6603 & ~n10559;
  assign n10564 = ~n10562 & ~n10563;
  assign n10565 = ~n10560 & n10564;
  assign n10566 = n2564 & ~n10565;
  assign n10567 = pi089 & ~n2564;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = ~pi562 & n10568;
  assign n10570 = ~n10553 & ~n10569;
  assign n10571 = pi222 & n10570;
  assign n10572 = ~pi222 & ~n10570;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = n6578 & n10573;
  assign n10575 = pi355 & ~n6578;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = ~n1761 & ~n10576;
  assign n10578 = ~n10546 & ~n10577;
  assign n10579 = ~n1754 & ~n10578;
  assign n10580 = pi822 & n10570;
  assign n10581 = ~pi822 & ~n10570;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = n1754 & n10582;
  assign po504 = n10579 | n10583;
  assign n10585 = pi356 & n1761;
  assign n10586 = pi740 & ~n6579;
  assign n10587 = pi634 & n6579;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = ~n2449 & ~n10588;
  assign n10590 = pi150 & n2449;
  assign n10591 = ~n10589 & ~n10590;
  assign n10592 = pi562 & n10591;
  assign n10593 = pi634 & n6592;
  assign n10594 = pi150 & n6594;
  assign n10595 = ~n6594 & ~n10591;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n6592 & ~n10596;
  assign n10598 = ~n10593 & ~n10597;
  assign n10599 = n6591 & ~n10598;
  assign n10600 = pi150 & ~pi669;
  assign n10601 = ~n6591 & n10600;
  assign n10602 = n6603 & ~n10598;
  assign n10603 = ~n10601 & ~n10602;
  assign n10604 = ~n10599 & n10603;
  assign n10605 = n2564 & ~n10604;
  assign n10606 = pi150 & ~n2564;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = ~pi562 & n10607;
  assign n10609 = ~n10592 & ~n10608;
  assign n10610 = pi292 & n10609;
  assign n10611 = ~pi292 & ~n10609;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = n6578 & n10612;
  assign n10614 = pi356 & ~n6578;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = ~n1761 & ~n10615;
  assign n10617 = ~n10585 & ~n10616;
  assign n10618 = ~n1754 & ~n10617;
  assign n10619 = pi868 & n10609;
  assign n10620 = ~pi868 & ~n10609;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = n1754 & n10621;
  assign po505 = n10618 | n10622;
  assign n10624 = pi357 & n1761;
  assign n10625 = pi741 & ~n6579;
  assign n10626 = pi576 & n6579;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = ~n2449 & ~n10627;
  assign n10629 = pi099 & n2449;
  assign n10630 = ~n10628 & ~n10629;
  assign n10631 = pi562 & n10630;
  assign n10632 = pi576 & n6592;
  assign n10633 = pi099 & n6594;
  assign n10634 = ~n6594 & ~n10630;
  assign n10635 = ~n10633 & ~n10634;
  assign n10636 = ~n6592 & ~n10635;
  assign n10637 = ~n10632 & ~n10636;
  assign n10638 = n6591 & ~n10637;
  assign n10639 = pi099 & ~pi669;
  assign n10640 = ~n6591 & n10639;
  assign n10641 = n6603 & ~n10637;
  assign n10642 = ~n10640 & ~n10641;
  assign n10643 = ~n10638 & n10642;
  assign n10644 = n2564 & ~n10643;
  assign n10645 = pi099 & ~n2564;
  assign n10646 = ~n10644 & ~n10645;
  assign n10647 = ~pi562 & n10646;
  assign n10648 = ~n10631 & ~n10647;
  assign n10649 = pi291 & n10648;
  assign n10650 = ~pi291 & ~n10648;
  assign n10651 = ~n10649 & ~n10650;
  assign n10652 = n6578 & n10651;
  assign n10653 = pi357 & ~n6578;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = ~n1761 & ~n10654;
  assign n10656 = ~n10624 & ~n10655;
  assign n10657 = ~n1754 & ~n10656;
  assign n10658 = pi869 & n10648;
  assign n10659 = ~pi869 & ~n10648;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = n1754 & n10660;
  assign po506 = n10657 | n10661;
  assign n10663 = pi358 & n1761;
  assign n10664 = pi695 & ~n6579;
  assign n10665 = pi531 & n6579;
  assign n10666 = ~n10664 & ~n10665;
  assign n10667 = ~n2449 & ~n10666;
  assign n10668 = pi030 & n2449;
  assign n10669 = ~n10667 & ~n10668;
  assign n10670 = pi562 & n10669;
  assign n10671 = pi531 & n6592;
  assign n10672 = pi030 & n6594;
  assign n10673 = ~n6594 & ~n10669;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = ~n6592 & ~n10674;
  assign n10676 = ~n10671 & ~n10675;
  assign n10677 = n6591 & ~n10676;
  assign n10678 = pi030 & ~pi669;
  assign n10679 = ~n6591 & n10678;
  assign n10680 = n6603 & ~n10676;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = ~n10677 & n10681;
  assign n10683 = n2564 & ~n10682;
  assign n10684 = pi030 & ~n2564;
  assign n10685 = ~n10683 & ~n10684;
  assign n10686 = ~pi562 & n10685;
  assign n10687 = ~n10670 & ~n10686;
  assign n10688 = pi220 & n10687;
  assign n10689 = ~pi220 & ~n10687;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = n6578 & n10690;
  assign n10692 = pi358 & ~n6578;
  assign n10693 = ~n10691 & ~n10692;
  assign n10694 = ~n1761 & ~n10693;
  assign n10695 = ~n10663 & ~n10694;
  assign n10696 = ~n1754 & ~n10695;
  assign n10697 = pi823 & n10687;
  assign n10698 = ~pi823 & ~n10687;
  assign n10699 = ~n10697 & ~n10698;
  assign n10700 = n1754 & n10699;
  assign po507 = n10696 | n10700;
  assign n10702 = pi359 & n1761;
  assign n10703 = pi743 & ~n6579;
  assign n10704 = pi585 & n6579;
  assign n10705 = ~n10703 & ~n10704;
  assign n10706 = ~n2449 & ~n10705;
  assign n10707 = pi039 & n2449;
  assign n10708 = ~n10706 & ~n10707;
  assign n10709 = pi562 & n10708;
  assign n10710 = pi585 & n6592;
  assign n10711 = pi039 & n6594;
  assign n10712 = ~n6594 & ~n10708;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~n6592 & ~n10713;
  assign n10715 = ~n10710 & ~n10714;
  assign n10716 = n6591 & ~n10715;
  assign n10717 = pi039 & ~pi669;
  assign n10718 = ~n6591 & n10717;
  assign n10719 = n6603 & ~n10715;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = ~n10716 & n10720;
  assign n10722 = n2564 & ~n10721;
  assign n10723 = pi039 & ~n2564;
  assign n10724 = ~n10722 & ~n10723;
  assign n10725 = ~pi562 & n10724;
  assign n10726 = ~n10709 & ~n10725;
  assign n10727 = pi252 & n10726;
  assign n10728 = ~pi252 & ~n10726;
  assign n10729 = ~n10727 & ~n10728;
  assign n10730 = n6578 & n10729;
  assign n10731 = pi359 & ~n6578;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 = ~n1761 & ~n10732;
  assign n10734 = ~n10702 & ~n10733;
  assign n10735 = ~n1754 & ~n10734;
  assign n10736 = pi871 & n10726;
  assign n10737 = ~pi871 & ~n10726;
  assign n10738 = ~n10736 & ~n10737;
  assign n10739 = n1754 & n10738;
  assign po508 = n10735 | n10739;
  assign n10741 = pi360 & n1761;
  assign n10742 = pi696 & ~n6579;
  assign n10743 = pi533 & n6579;
  assign n10744 = ~n10742 & ~n10743;
  assign n10745 = ~n2449 & ~n10744;
  assign n10746 = pi031 & n2449;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = pi562 & n10747;
  assign n10749 = pi533 & n6592;
  assign n10750 = pi031 & n6594;
  assign n10751 = ~n6594 & ~n10747;
  assign n10752 = ~n10750 & ~n10751;
  assign n10753 = ~n6592 & ~n10752;
  assign n10754 = ~n10749 & ~n10753;
  assign n10755 = n6591 & ~n10754;
  assign n10756 = pi031 & ~pi669;
  assign n10757 = ~n6591 & n10756;
  assign n10758 = n6603 & ~n10754;
  assign n10759 = ~n10757 & ~n10758;
  assign n10760 = ~n10755 & n10759;
  assign n10761 = n2564 & ~n10760;
  assign n10762 = pi031 & ~n2564;
  assign n10763 = ~n10761 & ~n10762;
  assign n10764 = ~pi562 & n10763;
  assign n10765 = ~n10748 & ~n10764;
  assign n10766 = pi221 & n10765;
  assign n10767 = ~pi221 & ~n10765;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = n6578 & n10768;
  assign n10770 = pi360 & ~n6578;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n1761 & ~n10771;
  assign n10773 = ~n10741 & ~n10772;
  assign n10774 = ~n1754 & ~n10773;
  assign n10775 = pi824 & n10765;
  assign n10776 = ~pi824 & ~n10765;
  assign n10777 = ~n10775 & ~n10776;
  assign n10778 = n1754 & n10777;
  assign po509 = n10774 | n10778;
  assign n10780 = pi361 & n1761;
  assign n10781 = pi744 & ~n6579;
  assign n10782 = pi577 & n6579;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = ~n2449 & ~n10783;
  assign n10785 = pi038 & n2449;
  assign n10786 = ~n10784 & ~n10785;
  assign n10787 = pi562 & n10786;
  assign n10788 = pi577 & n6592;
  assign n10789 = pi038 & n6594;
  assign n10790 = ~n6594 & ~n10786;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = ~n6592 & ~n10791;
  assign n10793 = ~n10788 & ~n10792;
  assign n10794 = n6591 & ~n10793;
  assign n10795 = pi038 & ~pi669;
  assign n10796 = ~n6591 & n10795;
  assign n10797 = n6603 & ~n10793;
  assign n10798 = ~n10796 & ~n10797;
  assign n10799 = ~n10794 & n10798;
  assign n10800 = n2564 & ~n10799;
  assign n10801 = pi038 & ~n2564;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~pi562 & n10802;
  assign n10804 = ~n10787 & ~n10803;
  assign n10805 = pi294 & n10804;
  assign n10806 = ~pi294 & ~n10804;
  assign n10807 = ~n10805 & ~n10806;
  assign n10808 = n6578 & n10807;
  assign n10809 = pi361 & ~n6578;
  assign n10810 = ~n10808 & ~n10809;
  assign n10811 = ~n1761 & ~n10810;
  assign n10812 = ~n10780 & ~n10811;
  assign n10813 = ~n1754 & ~n10812;
  assign n10814 = pi872 & n10804;
  assign n10815 = ~pi872 & ~n10804;
  assign n10816 = ~n10814 & ~n10815;
  assign n10817 = n1754 & n10816;
  assign po510 = n10813 | n10817;
  assign n10819 = pi362 & n1761;
  assign n10820 = pi776 & ~n6579;
  assign n10821 = pi570 & n6579;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = ~n2449 & ~n10822;
  assign n10824 = pi026 & n2449;
  assign n10825 = ~n10823 & ~n10824;
  assign n10826 = pi562 & n10825;
  assign n10827 = pi570 & n6592;
  assign n10828 = pi026 & n6594;
  assign n10829 = ~n6594 & ~n10825;
  assign n10830 = ~n10828 & ~n10829;
  assign n10831 = ~n6592 & ~n10830;
  assign n10832 = ~n10827 & ~n10831;
  assign n10833 = n6591 & ~n10832;
  assign n10834 = pi026 & ~pi669;
  assign n10835 = ~n6591 & n10834;
  assign n10836 = n6603 & ~n10832;
  assign n10837 = ~n10835 & ~n10836;
  assign n10838 = ~n10833 & n10837;
  assign n10839 = n2564 & ~n10838;
  assign n10840 = pi026 & ~n2564;
  assign n10841 = ~n10839 & ~n10840;
  assign n10842 = ~pi562 & n10841;
  assign n10843 = ~n10826 & ~n10842;
  assign n10844 = pi417 & n10843;
  assign n10845 = ~pi417 & ~n10843;
  assign n10846 = ~n10844 & ~n10845;
  assign n10847 = n6578 & n10846;
  assign n10848 = pi362 & ~n6578;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = ~n1761 & ~n10849;
  assign n10851 = ~n10819 & ~n10850;
  assign n10852 = ~n1754 & ~n10851;
  assign n10853 = pi904 & n10843;
  assign n10854 = ~pi904 & ~n10843;
  assign n10855 = ~n10853 & ~n10854;
  assign n10856 = n1754 & n10855;
  assign po511 = n10852 | n10856;
  assign n10858 = pi363 & n1761;
  assign n10859 = pi697 & ~n6579;
  assign n10860 = pi547 & n6579;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = ~n2449 & ~n10861;
  assign n10863 = pi091 & n2449;
  assign n10864 = ~n10862 & ~n10863;
  assign n10865 = pi562 & n10864;
  assign n10866 = pi547 & n6592;
  assign n10867 = pi091 & n6594;
  assign n10868 = ~n6594 & ~n10864;
  assign n10869 = ~n10867 & ~n10868;
  assign n10870 = ~n6592 & ~n10869;
  assign n10871 = ~n10866 & ~n10870;
  assign n10872 = n6591 & ~n10871;
  assign n10873 = pi091 & ~pi669;
  assign n10874 = ~n6591 & n10873;
  assign n10875 = n6603 & ~n10871;
  assign n10876 = ~n10874 & ~n10875;
  assign n10877 = ~n10872 & n10876;
  assign n10878 = n2564 & ~n10877;
  assign n10879 = pi091 & ~n2564;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = ~pi562 & n10880;
  assign n10882 = ~n10865 & ~n10881;
  assign n10883 = pi212 & n10882;
  assign n10884 = ~pi212 & ~n10882;
  assign n10885 = ~n10883 & ~n10884;
  assign n10886 = n6578 & n10885;
  assign n10887 = pi363 & ~n6578;
  assign n10888 = ~n10886 & ~n10887;
  assign n10889 = ~n1761 & ~n10888;
  assign n10890 = ~n10858 & ~n10889;
  assign n10891 = ~n1754 & ~n10890;
  assign n10892 = pi825 & n10882;
  assign n10893 = ~pi825 & ~n10882;
  assign n10894 = ~n10892 & ~n10893;
  assign n10895 = n1754 & n10894;
  assign po512 = n10891 | n10895;
  assign n10897 = pi364 & n1761;
  assign n10898 = pi789 & ~n6579;
  assign n10899 = pi621 & n6579;
  assign n10900 = ~n10898 & ~n10899;
  assign n10901 = ~n2449 & ~n10900;
  assign n10902 = pi086 & n2449;
  assign n10903 = ~n10901 & ~n10902;
  assign n10904 = pi562 & n10903;
  assign n10905 = pi621 & n6592;
  assign n10906 = pi086 & n6594;
  assign n10907 = ~n6594 & ~n10903;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = ~n6592 & ~n10908;
  assign n10910 = ~n10905 & ~n10909;
  assign n10911 = n6591 & ~n10910;
  assign n10912 = pi086 & ~pi669;
  assign n10913 = ~n6591 & n10912;
  assign n10914 = n6603 & ~n10910;
  assign n10915 = ~n10913 & ~n10914;
  assign n10916 = ~n10911 & n10915;
  assign n10917 = n2564 & ~n10916;
  assign n10918 = pi086 & ~n2564;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~pi562 & n10919;
  assign n10921 = ~n10904 & ~n10920;
  assign n10922 = pi431 & n10921;
  assign n10923 = ~pi431 & ~n10921;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = n6578 & n10924;
  assign n10926 = pi364 & ~n6578;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = ~n1761 & ~n10927;
  assign n10929 = ~n10897 & ~n10928;
  assign n10930 = ~n1754 & ~n10929;
  assign n10931 = pi917 & n10921;
  assign n10932 = ~pi917 & ~n10921;
  assign n10933 = ~n10931 & ~n10932;
  assign n10934 = n1754 & n10933;
  assign po513 = n10930 | n10934;
  assign n10936 = pi365 & n1761;
  assign n10937 = pi790 & ~n6579;
  assign n10938 = pi597 & n6579;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = ~n2449 & ~n10939;
  assign n10941 = pi087 & n2449;
  assign n10942 = ~n10940 & ~n10941;
  assign n10943 = pi562 & n10942;
  assign n10944 = pi597 & n6592;
  assign n10945 = pi087 & n6594;
  assign n10946 = ~n6594 & ~n10942;
  assign n10947 = ~n10945 & ~n10946;
  assign n10948 = ~n6592 & ~n10947;
  assign n10949 = ~n10944 & ~n10948;
  assign n10950 = n6591 & ~n10949;
  assign n10951 = pi087 & ~pi669;
  assign n10952 = ~n6591 & n10951;
  assign n10953 = n6603 & ~n10949;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = ~n10950 & n10954;
  assign n10956 = n2564 & ~n10955;
  assign n10957 = pi087 & ~n2564;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = ~pi562 & n10958;
  assign n10960 = ~n10943 & ~n10959;
  assign n10961 = pi432 & n10960;
  assign n10962 = ~pi432 & ~n10960;
  assign n10963 = ~n10961 & ~n10962;
  assign n10964 = n6578 & n10963;
  assign n10965 = pi365 & ~n6578;
  assign n10966 = ~n10964 & ~n10965;
  assign n10967 = ~n1761 & ~n10966;
  assign n10968 = ~n10936 & ~n10967;
  assign n10969 = ~n1754 & ~n10968;
  assign n10970 = pi918 & n10960;
  assign n10971 = ~pi918 & ~n10960;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = n1754 & n10972;
  assign po514 = n10969 | n10973;
  assign n10975 = pi366 & n1761;
  assign n10976 = pi754 & ~n6579;
  assign n10977 = pi623 & n6579;
  assign n10978 = ~n10976 & ~n10977;
  assign n10979 = ~n2449 & ~n10978;
  assign n10980 = pi066 & n2449;
  assign n10981 = ~n10979 & ~n10980;
  assign n10982 = pi562 & n10981;
  assign n10983 = pi623 & n6592;
  assign n10984 = pi066 & n6594;
  assign n10985 = ~n6594 & ~n10981;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = ~n6592 & ~n10986;
  assign n10988 = ~n10983 & ~n10987;
  assign n10989 = n6591 & ~n10988;
  assign n10990 = pi066 & ~pi669;
  assign n10991 = ~n6591 & n10990;
  assign n10992 = n6603 & ~n10988;
  assign n10993 = ~n10991 & ~n10992;
  assign n10994 = ~n10989 & n10993;
  assign n10995 = n2564 & ~n10994;
  assign n10996 = pi066 & ~n2564;
  assign n10997 = ~n10995 & ~n10996;
  assign n10998 = ~pi562 & n10997;
  assign n10999 = ~n10982 & ~n10998;
  assign n11000 = pi334 & n10999;
  assign n11001 = ~pi334 & ~n10999;
  assign n11002 = ~n11000 & ~n11001;
  assign n11003 = n6578 & n11002;
  assign n11004 = pi366 & ~n6578;
  assign n11005 = ~n11003 & ~n11004;
  assign n11006 = ~n1761 & ~n11005;
  assign n11007 = ~n10975 & ~n11006;
  assign n11008 = ~n1754 & ~n11007;
  assign n11009 = pi882 & n10999;
  assign n11010 = ~pi882 & ~n10999;
  assign n11011 = ~n11009 & ~n11010;
  assign n11012 = n1754 & n11011;
  assign po515 = n11008 | n11012;
  assign n11014 = pi367 & n1761;
  assign n11015 = pi755 & ~n6579;
  assign n11016 = pi635 & n6579;
  assign n11017 = ~n11015 & ~n11016;
  assign n11018 = ~n2449 & ~n11017;
  assign n11019 = pi179 & n2449;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = pi562 & n11020;
  assign n11022 = pi635 & n6592;
  assign n11023 = pi179 & n6594;
  assign n11024 = ~n6594 & ~n11020;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = ~n6592 & ~n11025;
  assign n11027 = ~n11022 & ~n11026;
  assign n11028 = n6591 & ~n11027;
  assign n11029 = pi179 & ~pi669;
  assign n11030 = ~n6591 & n11029;
  assign n11031 = n6603 & ~n11027;
  assign n11032 = ~n11030 & ~n11031;
  assign n11033 = ~n11028 & n11032;
  assign n11034 = n2564 & ~n11033;
  assign n11035 = pi179 & ~n2564;
  assign n11036 = ~n11034 & ~n11035;
  assign n11037 = ~pi562 & n11036;
  assign n11038 = ~n11021 & ~n11037;
  assign n11039 = pi298 & n11038;
  assign n11040 = ~pi298 & ~n11038;
  assign n11041 = ~n11039 & ~n11040;
  assign n11042 = n6578 & n11041;
  assign n11043 = pi367 & ~n6578;
  assign n11044 = ~n11042 & ~n11043;
  assign n11045 = ~n1761 & ~n11044;
  assign n11046 = ~n11014 & ~n11045;
  assign n11047 = ~n1754 & ~n11046;
  assign n11048 = pi883 & n11038;
  assign n11049 = ~pi883 & ~n11038;
  assign n11050 = ~n11048 & ~n11049;
  assign n11051 = n1754 & n11050;
  assign po516 = n11047 | n11051;
  assign n11053 = pi368 & n1761;
  assign n11054 = pi757 & ~n6579;
  assign n11055 = pi625 & n6579;
  assign n11056 = ~n11054 & ~n11055;
  assign n11057 = ~n2449 & ~n11056;
  assign n11058 = pi104 & n2449;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = pi562 & n11059;
  assign n11061 = pi625 & n6592;
  assign n11062 = pi104 & n6594;
  assign n11063 = ~n6594 & ~n11059;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n6592 & ~n11064;
  assign n11066 = ~n11061 & ~n11065;
  assign n11067 = n6591 & ~n11066;
  assign n11068 = pi104 & ~pi669;
  assign n11069 = ~n6591 & n11068;
  assign n11070 = n6603 & ~n11066;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = ~n11067 & n11071;
  assign n11073 = n2564 & ~n11072;
  assign n11074 = pi104 & ~n2564;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = ~pi562 & n11075;
  assign n11077 = ~n11060 & ~n11076;
  assign n11078 = pi335 & n11077;
  assign n11079 = ~pi335 & ~n11077;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = n6578 & n11080;
  assign n11082 = pi368 & ~n6578;
  assign n11083 = ~n11081 & ~n11082;
  assign n11084 = ~n1761 & ~n11083;
  assign n11085 = ~n11053 & ~n11084;
  assign n11086 = ~n1754 & ~n11085;
  assign n11087 = pi885 & n11077;
  assign n11088 = ~pi885 & ~n11077;
  assign n11089 = ~n11087 & ~n11088;
  assign n11090 = n1754 & n11089;
  assign po517 = n11086 | n11090;
  assign n11092 = pi369 & n1761;
  assign n11093 = pi759 & ~n6579;
  assign n11094 = pi578 & n6579;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = ~n2449 & ~n11095;
  assign n11097 = pi040 & n2449;
  assign n11098 = ~n11096 & ~n11097;
  assign n11099 = pi562 & n11098;
  assign n11100 = pi578 & n6592;
  assign n11101 = pi040 & n6594;
  assign n11102 = ~n6594 & ~n11098;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = ~n6592 & ~n11103;
  assign n11105 = ~n11100 & ~n11104;
  assign n11106 = n6591 & ~n11105;
  assign n11107 = pi040 & ~pi669;
  assign n11108 = ~n6591 & n11107;
  assign n11109 = n6603 & ~n11105;
  assign n11110 = ~n11108 & ~n11109;
  assign n11111 = ~n11106 & n11110;
  assign n11112 = n2564 & ~n11111;
  assign n11113 = pi040 & ~n2564;
  assign n11114 = ~n11112 & ~n11113;
  assign n11115 = ~pi562 & n11114;
  assign n11116 = ~n11099 & ~n11115;
  assign n11117 = pi337 & n11116;
  assign n11118 = ~pi337 & ~n11116;
  assign n11119 = ~n11117 & ~n11118;
  assign n11120 = n6578 & n11119;
  assign n11121 = pi369 & ~n6578;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = ~n1761 & ~n11122;
  assign n11124 = ~n11092 & ~n11123;
  assign n11125 = ~n1754 & ~n11124;
  assign n11126 = pi887 & n11116;
  assign n11127 = ~pi887 & ~n11116;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = n1754 & n11128;
  assign po518 = n11125 | n11129;
  assign n11131 = pi370 & n1761;
  assign n11132 = pi760 & ~n6579;
  assign n11133 = pi598 & n6579;
  assign n11134 = ~n11132 & ~n11133;
  assign n11135 = ~n2449 & ~n11134;
  assign n11136 = pi041 & n2449;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = pi562 & n11137;
  assign n11139 = pi598 & n6592;
  assign n11140 = pi041 & n6594;
  assign n11141 = ~n6594 & ~n11137;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = ~n6592 & ~n11142;
  assign n11144 = ~n11139 & ~n11143;
  assign n11145 = n6591 & ~n11144;
  assign n11146 = pi041 & ~pi669;
  assign n11147 = ~n6591 & n11146;
  assign n11148 = n6603 & ~n11144;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~n11145 & n11149;
  assign n11151 = n2564 & ~n11150;
  assign n11152 = pi041 & ~n2564;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = ~pi562 & n11153;
  assign n11155 = ~n11138 & ~n11154;
  assign n11156 = pi339 & n11155;
  assign n11157 = ~pi339 & ~n11155;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = n6578 & n11158;
  assign n11160 = pi370 & ~n6578;
  assign n11161 = ~n11159 & ~n11160;
  assign n11162 = ~n1761 & ~n11161;
  assign n11163 = ~n11131 & ~n11162;
  assign n11164 = ~n1754 & ~n11163;
  assign n11165 = pi888 & n11155;
  assign n11166 = ~pi888 & ~n11155;
  assign n11167 = ~n11165 & ~n11166;
  assign n11168 = n1754 & n11167;
  assign po519 = n11164 | n11168;
  assign n11170 = pi371 & n1761;
  assign n11171 = pi758 & ~n6579;
  assign n11172 = pi610 & n6579;
  assign n11173 = ~n11171 & ~n11172;
  assign n11174 = ~n2449 & ~n11173;
  assign n11175 = pi103 & n2449;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = pi562 & n11176;
  assign n11178 = pi610 & n6592;
  assign n11179 = pi103 & n6594;
  assign n11180 = ~n6594 & ~n11176;
  assign n11181 = ~n11179 & ~n11180;
  assign n11182 = ~n6592 & ~n11181;
  assign n11183 = ~n11178 & ~n11182;
  assign n11184 = n6591 & ~n11183;
  assign n11185 = pi103 & ~pi669;
  assign n11186 = ~n6591 & n11185;
  assign n11187 = n6603 & ~n11183;
  assign n11188 = ~n11186 & ~n11187;
  assign n11189 = ~n11184 & n11188;
  assign n11190 = n2564 & ~n11189;
  assign n11191 = pi103 & ~n2564;
  assign n11192 = ~n11190 & ~n11191;
  assign n11193 = ~pi562 & n11192;
  assign n11194 = ~n11177 & ~n11193;
  assign n11195 = pi336 & n11194;
  assign n11196 = ~pi336 & ~n11194;
  assign n11197 = ~n11195 & ~n11196;
  assign n11198 = n6578 & n11197;
  assign n11199 = pi371 & ~n6578;
  assign n11200 = ~n11198 & ~n11199;
  assign n11201 = ~n1761 & ~n11200;
  assign n11202 = ~n11170 & ~n11201;
  assign n11203 = ~n1754 & ~n11202;
  assign n11204 = pi886 & n11194;
  assign n11205 = ~pi886 & ~n11194;
  assign n11206 = ~n11204 & ~n11205;
  assign n11207 = n1754 & n11206;
  assign po520 = n11203 | n11207;
  assign n11209 = pi372 & n1761;
  assign n11210 = pi761 & ~n6579;
  assign n11211 = pi632 & n6579;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n2449 & ~n11212;
  assign n11214 = pi105 & n2449;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = pi562 & n11215;
  assign n11217 = pi632 & n6592;
  assign n11218 = pi105 & n6594;
  assign n11219 = ~n6594 & ~n11215;
  assign n11220 = ~n11218 & ~n11219;
  assign n11221 = ~n6592 & ~n11220;
  assign n11222 = ~n11217 & ~n11221;
  assign n11223 = n6591 & ~n11222;
  assign n11224 = pi105 & ~pi669;
  assign n11225 = ~n6591 & n11224;
  assign n11226 = n6603 & ~n11222;
  assign n11227 = ~n11225 & ~n11226;
  assign n11228 = ~n11223 & n11227;
  assign n11229 = n2564 & ~n11228;
  assign n11230 = pi105 & ~n2564;
  assign n11231 = ~n11229 & ~n11230;
  assign n11232 = ~pi562 & n11231;
  assign n11233 = ~n11216 & ~n11232;
  assign n11234 = pi296 & n11233;
  assign n11235 = ~pi296 & ~n11233;
  assign n11236 = ~n11234 & ~n11235;
  assign n11237 = n6578 & n11236;
  assign n11238 = pi372 & ~n6578;
  assign n11239 = ~n11237 & ~n11238;
  assign n11240 = ~n1761 & ~n11239;
  assign n11241 = ~n11209 & ~n11240;
  assign n11242 = ~n1754 & ~n11241;
  assign n11243 = pi889 & n11233;
  assign n11244 = ~pi889 & ~n11233;
  assign n11245 = ~n11243 & ~n11244;
  assign n11246 = n1754 & n11245;
  assign po521 = n11242 | n11246;
  assign n11248 = pi373 & n1761;
  assign n11249 = pi762 & ~n6579;
  assign n11250 = pi599 & n6579;
  assign n11251 = ~n11249 & ~n11250;
  assign n11252 = ~n2449 & ~n11251;
  assign n11253 = pi109 & n2449;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = pi562 & n11254;
  assign n11256 = pi599 & n6592;
  assign n11257 = pi109 & n6594;
  assign n11258 = ~n6594 & ~n11254;
  assign n11259 = ~n11257 & ~n11258;
  assign n11260 = ~n6592 & ~n11259;
  assign n11261 = ~n11256 & ~n11260;
  assign n11262 = n6591 & ~n11261;
  assign n11263 = pi109 & ~pi669;
  assign n11264 = ~n6591 & n11263;
  assign n11265 = n6603 & ~n11261;
  assign n11266 = ~n11264 & ~n11265;
  assign n11267 = ~n11262 & n11266;
  assign n11268 = n2564 & ~n11267;
  assign n11269 = pi109 & ~n2564;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 = ~pi562 & n11270;
  assign n11272 = ~n11255 & ~n11271;
  assign n11273 = pi248 & n11272;
  assign n11274 = ~pi248 & ~n11272;
  assign n11275 = ~n11273 & ~n11274;
  assign n11276 = n6578 & n11275;
  assign n11277 = pi373 & ~n6578;
  assign n11278 = ~n11276 & ~n11277;
  assign n11279 = ~n1761 & ~n11278;
  assign n11280 = ~n11248 & ~n11279;
  assign n11281 = ~n1754 & ~n11280;
  assign n11282 = pi890 & n11272;
  assign n11283 = ~pi890 & ~n11272;
  assign n11284 = ~n11282 & ~n11283;
  assign n11285 = n1754 & n11284;
  assign po522 = n11281 | n11285;
  assign n11287 = pi374 & n1761;
  assign n11288 = pi706 & ~n6579;
  assign n11289 = pi643 & n6579;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = ~n2449 & ~n11290;
  assign n11292 = pi092 & n2449;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = pi562 & n11293;
  assign n11295 = pi643 & n6592;
  assign n11296 = pi092 & n6594;
  assign n11297 = ~n6594 & ~n11293;
  assign n11298 = ~n11296 & ~n11297;
  assign n11299 = ~n6592 & ~n11298;
  assign n11300 = ~n11295 & ~n11299;
  assign n11301 = n6591 & ~n11300;
  assign n11302 = pi092 & ~pi669;
  assign n11303 = ~n6591 & n11302;
  assign n11304 = n6603 & ~n11300;
  assign n11305 = ~n11303 & ~n11304;
  assign n11306 = ~n11301 & n11305;
  assign n11307 = n2564 & ~n11306;
  assign n11308 = pi092 & ~n2564;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = ~pi562 & n11309;
  assign n11311 = ~n11294 & ~n11310;
  assign n11312 = ~pi229 & n11311;
  assign n11313 = pi229 & ~n11311;
  assign n11314 = ~n11312 & ~n11313;
  assign n11315 = n6578 & n11314;
  assign n11316 = pi374 & ~n6578;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = ~n1761 & ~n11317;
  assign n11319 = ~n11287 & ~n11318;
  assign n11320 = ~n1754 & ~n11319;
  assign n11321 = pi834 & n11311;
  assign n11322 = ~pi834 & ~n11311;
  assign n11323 = ~n11321 & ~n11322;
  assign n11324 = n1754 & n11323;
  assign po523 = n11320 | n11324;
  assign n11326 = pi375 & n1761;
  assign n11327 = pi793 & ~n6579;
  assign n11328 = pi614 & n6579;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~n2449 & ~n11329;
  assign n11331 = pi088 & n2449;
  assign n11332 = ~n11330 & ~n11331;
  assign n11333 = pi562 & n11332;
  assign n11334 = pi614 & n6592;
  assign n11335 = pi088 & n6594;
  assign n11336 = ~n6594 & ~n11332;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = ~n6592 & ~n11337;
  assign n11339 = ~n11334 & ~n11338;
  assign n11340 = n6591 & ~n11339;
  assign n11341 = pi088 & ~pi669;
  assign n11342 = ~n6591 & n11341;
  assign n11343 = n6603 & ~n11339;
  assign n11344 = ~n11342 & ~n11343;
  assign n11345 = ~n11340 & n11344;
  assign n11346 = n2564 & ~n11345;
  assign n11347 = pi088 & ~n2564;
  assign n11348 = ~n11346 & ~n11347;
  assign n11349 = ~pi562 & n11348;
  assign n11350 = ~n11333 & ~n11349;
  assign n11351 = pi419 & n11350;
  assign n11352 = ~pi419 & ~n11350;
  assign n11353 = ~n11351 & ~n11352;
  assign n11354 = n6578 & n11353;
  assign n11355 = pi375 & ~n6578;
  assign n11356 = ~n11354 & ~n11355;
  assign n11357 = ~n1761 & ~n11356;
  assign n11358 = ~n11326 & ~n11357;
  assign n11359 = ~n1754 & ~n11358;
  assign n11360 = pi921 & n11350;
  assign n11361 = ~pi921 & ~n11350;
  assign n11362 = ~n11360 & ~n11361;
  assign n11363 = n1754 & n11362;
  assign po524 = n11359 | n11363;
  assign n11365 = pi376 & n1761;
  assign n11366 = pi770 & ~n6579;
  assign n11367 = pi620 & n6579;
  assign n11368 = ~n11366 & ~n11367;
  assign n11369 = ~n2449 & ~n11368;
  assign n11370 = pi067 & n2449;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = pi562 & n11371;
  assign n11373 = pi620 & n6592;
  assign n11374 = pi067 & n6594;
  assign n11375 = ~n6594 & ~n11371;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = ~n6592 & ~n11376;
  assign n11378 = ~n11373 & ~n11377;
  assign n11379 = n6591 & ~n11378;
  assign n11380 = pi067 & ~pi669;
  assign n11381 = ~n6591 & n11380;
  assign n11382 = n6603 & ~n11378;
  assign n11383 = ~n11381 & ~n11382;
  assign n11384 = ~n11379 & n11383;
  assign n11385 = n2564 & ~n11384;
  assign n11386 = pi067 & ~n2564;
  assign n11387 = ~n11385 & ~n11386;
  assign n11388 = ~pi562 & n11387;
  assign n11389 = ~n11372 & ~n11388;
  assign n11390 = pi413 & n11389;
  assign n11391 = ~pi413 & ~n11389;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = n6578 & n11392;
  assign n11394 = pi376 & ~n6578;
  assign n11395 = ~n11393 & ~n11394;
  assign n11396 = ~n1761 & ~n11395;
  assign n11397 = ~n11365 & ~n11396;
  assign n11398 = ~n1754 & ~n11397;
  assign n11399 = pi898 & n11389;
  assign n11400 = ~pi898 & ~n11389;
  assign n11401 = ~n11399 & ~n11400;
  assign n11402 = n1754 & n11401;
  assign po525 = n11398 | n11402;
  assign n11404 = pi377 & n1761;
  assign n11405 = pi771 & ~n6579;
  assign n11406 = pi606 & n6579;
  assign n11407 = ~n11405 & ~n11406;
  assign n11408 = ~n2449 & ~n11407;
  assign n11409 = pi175 & n2449;
  assign n11410 = ~n11408 & ~n11409;
  assign n11411 = pi562 & n11410;
  assign n11412 = pi606 & n6592;
  assign n11413 = pi175 & n6594;
  assign n11414 = ~n6594 & ~n11410;
  assign n11415 = ~n11413 & ~n11414;
  assign n11416 = ~n6592 & ~n11415;
  assign n11417 = ~n11412 & ~n11416;
  assign n11418 = n6591 & ~n11417;
  assign n11419 = pi175 & ~pi669;
  assign n11420 = ~n6591 & n11419;
  assign n11421 = n6603 & ~n11417;
  assign n11422 = ~n11420 & ~n11421;
  assign n11423 = ~n11418 & n11422;
  assign n11424 = n2564 & ~n11423;
  assign n11425 = pi175 & ~n2564;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = ~pi562 & n11426;
  assign n11428 = ~n11411 & ~n11427;
  assign n11429 = pi409 & n11428;
  assign n11430 = ~pi409 & ~n11428;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = n6578 & n11431;
  assign n11433 = pi377 & ~n6578;
  assign n11434 = ~n11432 & ~n11433;
  assign n11435 = ~n1761 & ~n11434;
  assign n11436 = ~n11404 & ~n11435;
  assign n11437 = ~n1754 & ~n11436;
  assign n11438 = pi899 & n11428;
  assign n11439 = ~pi899 & ~n11428;
  assign n11440 = ~n11438 & ~n11439;
  assign n11441 = n1754 & n11440;
  assign po526 = n11437 | n11441;
  assign n11443 = pi378 & n1761;
  assign n11444 = pi710 & ~n6579;
  assign n11445 = pi616 & n6579;
  assign n11446 = ~n11444 & ~n11445;
  assign n11447 = ~n2449 & ~n11446;
  assign n11448 = pi097 & n2449;
  assign n11449 = ~n11447 & ~n11448;
  assign n11450 = pi562 & n11449;
  assign n11451 = pi616 & n6592;
  assign n11452 = pi097 & n6594;
  assign n11453 = ~n6594 & ~n11449;
  assign n11454 = ~n11452 & ~n11453;
  assign n11455 = ~n6592 & ~n11454;
  assign n11456 = ~n11451 & ~n11455;
  assign n11457 = n6591 & ~n11456;
  assign n11458 = pi097 & ~pi669;
  assign n11459 = ~n6591 & n11458;
  assign n11460 = n6603 & ~n11456;
  assign n11461 = ~n11459 & ~n11460;
  assign n11462 = ~n11457 & n11461;
  assign n11463 = n2564 & ~n11462;
  assign n11464 = pi097 & ~n2564;
  assign n11465 = ~n11463 & ~n11464;
  assign n11466 = ~pi562 & n11465;
  assign n11467 = ~n11450 & ~n11466;
  assign n11468 = ~pi233 & n11467;
  assign n11469 = pi233 & ~n11467;
  assign n11470 = ~n11468 & ~n11469;
  assign n11471 = n6578 & n11470;
  assign n11472 = pi378 & ~n6578;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~n1761 & ~n11473;
  assign n11475 = ~n11443 & ~n11474;
  assign n11476 = ~n1754 & ~n11475;
  assign n11477 = pi838 & n11467;
  assign n11478 = ~pi838 & ~n11467;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 = n1754 & n11479;
  assign po527 = n11476 | n11480;
  assign n11482 = pi379 & n1761;
  assign n11483 = pi773 & ~n6579;
  assign n11484 = pi581 & n6579;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = ~n2449 & ~n11485;
  assign n11487 = pi118 & n2449;
  assign n11488 = ~n11486 & ~n11487;
  assign n11489 = pi562 & n11488;
  assign n11490 = pi581 & n6592;
  assign n11491 = pi118 & n6594;
  assign n11492 = ~n6594 & ~n11488;
  assign n11493 = ~n11491 & ~n11492;
  assign n11494 = ~n6592 & ~n11493;
  assign n11495 = ~n11490 & ~n11494;
  assign n11496 = n6591 & ~n11495;
  assign n11497 = pi118 & ~pi669;
  assign n11498 = ~n6591 & n11497;
  assign n11499 = n6603 & ~n11495;
  assign n11500 = ~n11498 & ~n11499;
  assign n11501 = ~n11496 & n11500;
  assign n11502 = n2564 & ~n11501;
  assign n11503 = pi118 & ~n2564;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = ~pi562 & n11504;
  assign n11506 = ~n11489 & ~n11505;
  assign n11507 = pi437 & n11506;
  assign n11508 = ~pi437 & ~n11506;
  assign n11509 = ~n11507 & ~n11508;
  assign n11510 = n6578 & n11509;
  assign n11511 = pi379 & ~n6578;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = ~n1761 & ~n11512;
  assign n11514 = ~n11482 & ~n11513;
  assign n11515 = ~n1754 & ~n11514;
  assign n11516 = pi901 & n11506;
  assign n11517 = ~pi901 & ~n11506;
  assign n11518 = ~n11516 & ~n11517;
  assign n11519 = n1754 & n11518;
  assign po528 = n11515 | n11519;
  assign n11521 = pi380 & n1761;
  assign n11522 = pi711 & ~n6579;
  assign n11523 = pi609 & n6579;
  assign n11524 = ~n11522 & ~n11523;
  assign n11525 = ~n2449 & ~n11524;
  assign n11526 = pi032 & n2449;
  assign n11527 = ~n11525 & ~n11526;
  assign n11528 = pi562 & n11527;
  assign n11529 = pi609 & n6592;
  assign n11530 = pi032 & n6594;
  assign n11531 = ~n6594 & ~n11527;
  assign n11532 = ~n11530 & ~n11531;
  assign n11533 = ~n6592 & ~n11532;
  assign n11534 = ~n11529 & ~n11533;
  assign n11535 = n6591 & ~n11534;
  assign n11536 = pi032 & ~pi669;
  assign n11537 = ~n6591 & n11536;
  assign n11538 = n6603 & ~n11534;
  assign n11539 = ~n11537 & ~n11538;
  assign n11540 = ~n11535 & n11539;
  assign n11541 = n2564 & ~n11540;
  assign n11542 = pi032 & ~n2564;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = ~pi562 & n11543;
  assign n11545 = ~n11528 & ~n11544;
  assign n11546 = ~pi237 & n11545;
  assign n11547 = pi237 & ~n11545;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = n6578 & n11548;
  assign n11550 = pi380 & ~n6578;
  assign n11551 = ~n11549 & ~n11550;
  assign n11552 = ~n1761 & ~n11551;
  assign n11553 = ~n11521 & ~n11552;
  assign n11554 = ~n1754 & ~n11553;
  assign n11555 = pi839 & n11545;
  assign n11556 = ~pi839 & ~n11545;
  assign n11557 = ~n11555 & ~n11556;
  assign n11558 = n1754 & n11557;
  assign po529 = n11554 | n11558;
  assign n11560 = pi381 & n1761;
  assign n11561 = pi712 & ~n6579;
  assign n11562 = pi658 & n6579;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = ~n2449 & ~n11563;
  assign n11565 = pi033 & n2449;
  assign n11566 = ~n11564 & ~n11565;
  assign n11567 = pi562 & n11566;
  assign n11568 = pi658 & n6592;
  assign n11569 = pi033 & n6594;
  assign n11570 = ~n6594 & ~n11566;
  assign n11571 = ~n11569 & ~n11570;
  assign n11572 = ~n6592 & ~n11571;
  assign n11573 = ~n11568 & ~n11572;
  assign n11574 = n6591 & ~n11573;
  assign n11575 = pi033 & ~pi669;
  assign n11576 = ~n6591 & n11575;
  assign n11577 = n6603 & ~n11573;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = ~n11574 & n11578;
  assign n11580 = n2564 & ~n11579;
  assign n11581 = pi033 & ~n2564;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = ~pi562 & n11582;
  assign n11584 = ~n11567 & ~n11583;
  assign n11585 = ~pi234 & n11584;
  assign n11586 = pi234 & ~n11584;
  assign n11587 = ~n11585 & ~n11586;
  assign n11588 = n6578 & n11587;
  assign n11589 = pi381 & ~n6578;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = ~n1761 & ~n11590;
  assign n11592 = ~n11560 & ~n11591;
  assign n11593 = ~n1754 & ~n11592;
  assign n11594 = pi840 & n11584;
  assign n11595 = ~pi840 & ~n11584;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = n1754 & n11596;
  assign po530 = n11593 | n11597;
  assign n11599 = pi382 & n1761;
  assign n11600 = pi713 & ~n6579;
  assign n11601 = pi617 & n6579;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = ~n2449 & ~n11602;
  assign n11604 = pi116 & n2449;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = pi562 & n11605;
  assign n11607 = pi617 & n6592;
  assign n11608 = pi116 & n6594;
  assign n11609 = ~n6594 & ~n11605;
  assign n11610 = ~n11608 & ~n11609;
  assign n11611 = ~n6592 & ~n11610;
  assign n11612 = ~n11607 & ~n11611;
  assign n11613 = n6591 & ~n11612;
  assign n11614 = pi116 & ~pi669;
  assign n11615 = ~n6591 & n11614;
  assign n11616 = n6603 & ~n11612;
  assign n11617 = ~n11615 & ~n11616;
  assign n11618 = ~n11613 & n11617;
  assign n11619 = n2564 & ~n11618;
  assign n11620 = pi116 & ~n2564;
  assign n11621 = ~n11619 & ~n11620;
  assign n11622 = ~pi562 & n11621;
  assign n11623 = ~n11606 & ~n11622;
  assign n11624 = ~pi235 & n11623;
  assign n11625 = pi235 & ~n11623;
  assign n11626 = ~n11624 & ~n11625;
  assign n11627 = n6578 & n11626;
  assign n11628 = pi382 & ~n6578;
  assign n11629 = ~n11627 & ~n11628;
  assign n11630 = ~n1761 & ~n11629;
  assign n11631 = ~n11599 & ~n11630;
  assign n11632 = ~n1754 & ~n11631;
  assign n11633 = pi841 & n11623;
  assign n11634 = ~pi841 & ~n11623;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = n1754 & n11635;
  assign po531 = n11632 | n11636;
  assign n11638 = pi383 & n1761;
  assign n11639 = pi723 & ~n6579;
  assign n11640 = pi596 & n6579;
  assign n11641 = ~n11639 & ~n11640;
  assign n11642 = ~n2449 & ~n11641;
  assign n11643 = pi180 & n2449;
  assign n11644 = ~n11642 & ~n11643;
  assign n11645 = pi562 & n11644;
  assign n11646 = pi596 & n6592;
  assign n11647 = pi180 & n6594;
  assign n11648 = ~n6594 & ~n11644;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = ~n6592 & ~n11649;
  assign n11651 = ~n11646 & ~n11650;
  assign n11652 = n6591 & ~n11651;
  assign n11653 = pi180 & ~pi669;
  assign n11654 = ~n6591 & n11653;
  assign n11655 = n6603 & ~n11651;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = ~n11652 & n11656;
  assign n11658 = n2564 & ~n11657;
  assign n11659 = pi180 & ~n2564;
  assign n11660 = ~n11658 & ~n11659;
  assign n11661 = ~pi562 & n11660;
  assign n11662 = ~n11645 & ~n11661;
  assign n11663 = ~pi240 & n11662;
  assign n11664 = pi240 & ~n11662;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = n6578 & n11665;
  assign n11667 = pi383 & ~n6578;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = ~n1761 & ~n11668;
  assign n11670 = ~n11638 & ~n11669;
  assign n11671 = ~n1754 & ~n11670;
  assign n11672 = pi851 & n11662;
  assign n11673 = ~pi851 & ~n11662;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = n1754 & n11674;
  assign po532 = n11671 | n11675;
  assign n11677 = pi384 & n1761;
  assign n11678 = pi726 & ~n6579;
  assign n11679 = pi630 & n6579;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n2449 & ~n11680;
  assign n11682 = pi095 & n2449;
  assign n11683 = ~n11681 & ~n11682;
  assign n11684 = pi562 & n11683;
  assign n11685 = pi630 & n6592;
  assign n11686 = pi095 & n6594;
  assign n11687 = ~n6594 & ~n11683;
  assign n11688 = ~n11686 & ~n11687;
  assign n11689 = ~n6592 & ~n11688;
  assign n11690 = ~n11685 & ~n11689;
  assign n11691 = n6591 & ~n11690;
  assign n11692 = pi095 & ~pi669;
  assign n11693 = ~n6591 & n11692;
  assign n11694 = n6603 & ~n11690;
  assign n11695 = ~n11693 & ~n11694;
  assign n11696 = ~n11691 & n11695;
  assign n11697 = n2564 & ~n11696;
  assign n11698 = pi095 & ~n2564;
  assign n11699 = ~n11697 & ~n11698;
  assign n11700 = ~pi562 & n11699;
  assign n11701 = ~n11684 & ~n11700;
  assign n11702 = ~pi243 & n11701;
  assign n11703 = pi243 & ~n11701;
  assign n11704 = ~n11702 & ~n11703;
  assign n11705 = n6578 & n11704;
  assign n11706 = pi384 & ~n6578;
  assign n11707 = ~n11705 & ~n11706;
  assign n11708 = ~n1761 & ~n11707;
  assign n11709 = ~n11677 & ~n11708;
  assign n11710 = ~n1754 & ~n11709;
  assign n11711 = pi854 & n11701;
  assign n11712 = ~pi854 & ~n11701;
  assign n11713 = ~n11711 & ~n11712;
  assign n11714 = n1754 & n11713;
  assign po533 = n11710 | n11714;
  assign n11716 = pi385 & n1761;
  assign n11717 = pi729 & ~n6579;
  assign n11718 = pi618 & n6579;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = ~n2449 & ~n11719;
  assign n11721 = pi096 & n2449;
  assign n11722 = ~n11720 & ~n11721;
  assign n11723 = pi562 & n11722;
  assign n11724 = pi618 & n6592;
  assign n11725 = pi096 & n6594;
  assign n11726 = ~n6594 & ~n11722;
  assign n11727 = ~n11725 & ~n11726;
  assign n11728 = ~n6592 & ~n11727;
  assign n11729 = ~n11724 & ~n11728;
  assign n11730 = n6591 & ~n11729;
  assign n11731 = pi096 & ~pi669;
  assign n11732 = ~n6591 & n11731;
  assign n11733 = n6603 & ~n11729;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = ~n11730 & n11734;
  assign n11736 = n2564 & ~n11735;
  assign n11737 = pi096 & ~n2564;
  assign n11738 = ~n11736 & ~n11737;
  assign n11739 = ~pi562 & n11738;
  assign n11740 = ~n11723 & ~n11739;
  assign n11741 = ~pi236 & n11740;
  assign n11742 = pi236 & ~n11740;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = n6578 & n11743;
  assign n11745 = pi385 & ~n6578;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = ~n1761 & ~n11746;
  assign n11748 = ~n11716 & ~n11747;
  assign n11749 = ~n1754 & ~n11748;
  assign n11750 = pi857 & n11740;
  assign n11751 = ~pi857 & ~n11740;
  assign n11752 = ~n11750 & ~n11751;
  assign n11753 = n1754 & n11752;
  assign po534 = n11749 | n11753;
  assign n11755 = pi386 & n1761;
  assign n11756 = pi691 & ~n6579;
  assign n11757 = pi518 & n6579;
  assign n11758 = ~n11756 & ~n11757;
  assign n11759 = ~n2449 & ~n11758;
  assign n11760 = pi172 & n2449;
  assign n11761 = ~n11759 & ~n11760;
  assign n11762 = pi562 & n11761;
  assign n11763 = pi518 & n6592;
  assign n11764 = pi172 & n6594;
  assign n11765 = ~n6594 & ~n11761;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = ~n6592 & ~n11766;
  assign n11768 = ~n11763 & ~n11767;
  assign n11769 = n6591 & ~n11768;
  assign n11770 = pi172 & ~pi669;
  assign n11771 = ~n6591 & n11770;
  assign n11772 = n6603 & ~n11768;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = ~n11769 & n11773;
  assign n11775 = n2564 & ~n11774;
  assign n11776 = pi172 & ~n2564;
  assign n11777 = ~n11775 & ~n11776;
  assign n11778 = ~pi562 & n11777;
  assign n11779 = ~n11762 & ~n11778;
  assign n11780 = pi216 & n11779;
  assign n11781 = ~pi216 & ~n11779;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = n6578 & n11782;
  assign n11784 = pi386 & ~n6578;
  assign n11785 = ~n11783 & ~n11784;
  assign n11786 = ~n1761 & ~n11785;
  assign n11787 = ~n11755 & ~n11786;
  assign n11788 = ~n1754 & ~n11787;
  assign n11789 = pi819 & n11779;
  assign n11790 = ~pi819 & ~n11779;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = n1754 & n11791;
  assign po535 = n11788 | n11792;
  assign n11794 = pi387 & ~po814;
  assign n11795 = po814 & ~n5544;
  assign po536 = n11794 | n11795;
  assign n11797 = pi388 & ~po814;
  assign n11798 = po814 & ~n5644;
  assign po537 = n11797 | n11798;
  assign n11800 = pi389 & ~po814;
  assign n11801 = po814 & ~n5593;
  assign po538 = n11800 | n11801;
  assign n11803 = n5284 & ~n6577;
  assign n11804 = ~n5283 & ~n11803;
  assign n11805 = ~n1754 & ~n11804;
  assign n11806 = ~n2021 & ~n11805;
  assign po539 = n5288 | ~n11806;
  assign n11808 = pi391 & n1761;
  assign n11809 = pi792 & ~n6579;
  assign n11810 = pi629 & n6579;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = ~n2449 & ~n11811;
  assign n11813 = pi028 & n2449;
  assign n11814 = ~n11812 & ~n11813;
  assign n11815 = pi562 & n11814;
  assign n11816 = pi629 & n6592;
  assign n11817 = pi028 & n6594;
  assign n11818 = ~n6594 & ~n11814;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = ~n6592 & ~n11819;
  assign n11821 = ~n11816 & ~n11820;
  assign n11822 = n6591 & ~n11821;
  assign n11823 = pi028 & ~pi669;
  assign n11824 = ~n6591 & n11823;
  assign n11825 = n6603 & ~n11821;
  assign n11826 = ~n11824 & ~n11825;
  assign n11827 = ~n11822 & n11826;
  assign n11828 = n2564 & ~n11827;
  assign n11829 = pi028 & ~n2564;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = ~pi562 & n11830;
  assign n11832 = ~n11815 & ~n11831;
  assign n11833 = pi434 & n11832;
  assign n11834 = ~pi434 & ~n11832;
  assign n11835 = ~n11833 & ~n11834;
  assign n11836 = n6578 & n11835;
  assign n11837 = pi391 & ~n6578;
  assign n11838 = ~n11836 & ~n11837;
  assign n11839 = ~n1761 & ~n11838;
  assign n11840 = ~n11808 & ~n11839;
  assign n11841 = ~n1754 & ~n11840;
  assign n11842 = pi920 & n11832;
  assign n11843 = ~pi920 & ~n11832;
  assign n11844 = ~n11842 & ~n11843;
  assign n11845 = n1754 & n11844;
  assign po540 = n11841 | n11845;
  assign n11847 = pi392 & n1761;
  assign n11848 = pi763 & ~n6579;
  assign n11849 = pi600 & n6579;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = ~n2449 & ~n11850;
  assign n11852 = ~pi184 & n2449;
  assign n11853 = ~n11851 & ~n11852;
  assign n11854 = pi562 & n11853;
  assign n11855 = pi600 & n6592;
  assign n11856 = ~pi184 & n6594;
  assign n11857 = ~n6594 & ~n11853;
  assign n11858 = ~n11856 & ~n11857;
  assign n11859 = ~n6592 & ~n11858;
  assign n11860 = ~n11855 & ~n11859;
  assign n11861 = n6591 & ~n11860;
  assign n11862 = ~pi184 & ~pi669;
  assign n11863 = ~n6591 & n11862;
  assign n11864 = n6603 & ~n11860;
  assign n11865 = ~n11863 & ~n11864;
  assign n11866 = ~n11861 & n11865;
  assign n11867 = n2564 & ~n11866;
  assign n11868 = ~pi184 & ~n2564;
  assign n11869 = ~n11867 & ~n11868;
  assign n11870 = ~pi562 & n11869;
  assign n11871 = ~n11854 & ~n11870;
  assign n11872 = pi251 & n11871;
  assign n11873 = ~pi251 & ~n11871;
  assign n11874 = ~n11872 & ~n11873;
  assign n11875 = n6578 & n11874;
  assign n11876 = pi392 & ~n6578;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = ~n1761 & ~n11877;
  assign n11879 = ~n11847 & ~n11878;
  assign n11880 = ~n1754 & ~n11879;
  assign n11881 = pi891 & n11871;
  assign n11882 = ~pi891 & ~n11871;
  assign n11883 = ~n11881 & ~n11882;
  assign n11884 = n1754 & n11883;
  assign po541 = n11880 | n11884;
  assign n11886 = pi393 & n1761;
  assign n11887 = pi791 & ~n6579;
  assign n11888 = pi655 & n6579;
  assign n11889 = ~n11887 & ~n11888;
  assign n11890 = ~n2449 & ~n11889;
  assign n11891 = pi029 & n2449;
  assign n11892 = ~n11890 & ~n11891;
  assign n11893 = pi562 & n11892;
  assign n11894 = pi655 & n6592;
  assign n11895 = pi029 & n6594;
  assign n11896 = ~n6594 & ~n11892;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = ~n6592 & ~n11897;
  assign n11899 = ~n11894 & ~n11898;
  assign n11900 = n6591 & ~n11899;
  assign n11901 = pi029 & ~pi669;
  assign n11902 = ~n6591 & n11901;
  assign n11903 = n6603 & ~n11899;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n11900 & n11904;
  assign n11906 = n2564 & ~n11905;
  assign n11907 = pi029 & ~n2564;
  assign n11908 = ~n11906 & ~n11907;
  assign n11909 = ~pi562 & n11908;
  assign n11910 = ~n11893 & ~n11909;
  assign n11911 = pi436 & n11910;
  assign n11912 = ~pi436 & ~n11910;
  assign n11913 = ~n11911 & ~n11912;
  assign n11914 = n6578 & n11913;
  assign n11915 = pi393 & ~n6578;
  assign n11916 = ~n11914 & ~n11915;
  assign n11917 = ~n1761 & ~n11916;
  assign n11918 = ~n11886 & ~n11917;
  assign n11919 = ~n1754 & ~n11918;
  assign n11920 = pi919 & n11910;
  assign n11921 = ~pi919 & ~n11910;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = n1754 & n11922;
  assign po542 = n11919 | n11923;
  assign n11925 = pi394 & ~po814;
  assign n11926 = po814 & ~n5494;
  assign po543 = n11925 | n11926;
  assign n11928 = pi395 & n1761;
  assign n11929 = pi756 & ~n6579;
  assign n11930 = pi580 & n6579;
  assign n11931 = ~n11929 & ~n11930;
  assign n11932 = ~n2449 & ~n11931;
  assign n11933 = pi151 & n2449;
  assign n11934 = ~n11932 & ~n11933;
  assign n11935 = pi562 & n11934;
  assign n11936 = pi580 & n6592;
  assign n11937 = pi151 & n6594;
  assign n11938 = ~n6594 & ~n11934;
  assign n11939 = ~n11937 & ~n11938;
  assign n11940 = ~n6592 & ~n11939;
  assign n11941 = ~n11936 & ~n11940;
  assign n11942 = n6591 & ~n11941;
  assign n11943 = pi151 & ~pi669;
  assign n11944 = ~n6591 & n11943;
  assign n11945 = n6603 & ~n11941;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11942 & n11946;
  assign n11948 = n2564 & ~n11947;
  assign n11949 = pi151 & ~n2564;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = ~pi562 & n11950;
  assign n11952 = ~n11935 & ~n11951;
  assign n11953 = pi338 & n11952;
  assign n11954 = ~pi338 & ~n11952;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = n6578 & n11955;
  assign n11957 = pi395 & ~n6578;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = ~n1761 & ~n11958;
  assign n11960 = ~n11928 & ~n11959;
  assign n11961 = ~n1754 & ~n11960;
  assign n11962 = pi884 & n11952;
  assign n11963 = ~pi884 & ~n11952;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = n1754 & n11964;
  assign po544 = n11961 | n11965;
  assign n11967 = pi396 & ~po814;
  assign n11968 = po814 & ~n5695;
  assign po545 = n11967 | n11968;
  assign n11970 = pi397 & n1761;
  assign n11971 = pi788 & ~n6579;
  assign n11972 = pi657 & n6579;
  assign n11973 = ~n11971 & ~n11972;
  assign n11974 = ~n2449 & ~n11973;
  assign n11975 = pi143 & n2449;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = pi562 & n11976;
  assign n11978 = pi657 & n6592;
  assign n11979 = pi143 & n6594;
  assign n11980 = ~n6594 & ~n11976;
  assign n11981 = ~n11979 & ~n11980;
  assign n11982 = ~n6592 & ~n11981;
  assign n11983 = ~n11978 & ~n11982;
  assign n11984 = n6591 & ~n11983;
  assign n11985 = pi143 & ~pi669;
  assign n11986 = ~n6591 & n11985;
  assign n11987 = n6603 & ~n11983;
  assign n11988 = ~n11986 & ~n11987;
  assign n11989 = ~n11984 & n11988;
  assign n11990 = n2564 & ~n11989;
  assign n11991 = pi143 & ~n2564;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = ~pi562 & n11992;
  assign n11994 = ~n11977 & ~n11993;
  assign n11995 = pi433 & n11994;
  assign n11996 = ~pi433 & ~n11994;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 = n6578 & n11997;
  assign n11999 = pi397 & ~n6578;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = ~n1761 & ~n12000;
  assign n12002 = ~n11970 & ~n12001;
  assign n12003 = ~n1754 & ~n12002;
  assign n12004 = pi916 & n11994;
  assign n12005 = ~pi916 & ~n11994;
  assign n12006 = ~n12004 & ~n12005;
  assign n12007 = n1754 & n12006;
  assign po546 = n12003 | n12007;
  assign n12009 = pi398 & n1761;
  assign n12010 = pi728 & ~n6579;
  assign n12011 = pi640 & n6579;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = ~n2449 & ~n12012;
  assign n12014 = pi035 & n2449;
  assign n12015 = ~n12013 & ~n12014;
  assign n12016 = pi562 & n12015;
  assign n12017 = pi640 & n6592;
  assign n12018 = pi035 & n6594;
  assign n12019 = ~n6594 & ~n12015;
  assign n12020 = ~n12018 & ~n12019;
  assign n12021 = ~n6592 & ~n12020;
  assign n12022 = ~n12017 & ~n12021;
  assign n12023 = n6591 & ~n12022;
  assign n12024 = pi035 & ~pi669;
  assign n12025 = ~n6591 & n12024;
  assign n12026 = n6603 & ~n12022;
  assign n12027 = ~n12025 & ~n12026;
  assign n12028 = ~n12023 & n12027;
  assign n12029 = n2564 & ~n12028;
  assign n12030 = pi035 & ~n2564;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = ~pi562 & n12031;
  assign n12033 = ~n12016 & ~n12032;
  assign n12034 = ~pi244 & n12033;
  assign n12035 = pi244 & ~n12033;
  assign n12036 = ~n12034 & ~n12035;
  assign n12037 = n6578 & n12036;
  assign n12038 = pi398 & ~n6578;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = ~n1761 & ~n12039;
  assign n12041 = ~n12009 & ~n12040;
  assign n12042 = ~n1754 & ~n12041;
  assign n12043 = pi856 & n12033;
  assign n12044 = ~pi856 & ~n12033;
  assign n12045 = ~n12043 & ~n12044;
  assign n12046 = n1754 & n12045;
  assign po547 = n12042 | n12046;
  assign n12048 = pi399 & n1761;
  assign n12049 = pi745 & ~n6579;
  assign n12050 = pi589 & n6579;
  assign n12051 = ~n12049 & ~n12050;
  assign n12052 = ~n2449 & ~n12051;
  assign n12053 = pi102 & n2449;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = pi562 & n12054;
  assign n12056 = pi589 & n6592;
  assign n12057 = pi102 & n6594;
  assign n12058 = ~n6594 & ~n12054;
  assign n12059 = ~n12057 & ~n12058;
  assign n12060 = ~n6592 & ~n12059;
  assign n12061 = ~n12056 & ~n12060;
  assign n12062 = n6591 & ~n12061;
  assign n12063 = pi102 & ~pi669;
  assign n12064 = ~n6591 & n12063;
  assign n12065 = n6603 & ~n12061;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = ~n12062 & n12066;
  assign n12068 = n2564 & ~n12067;
  assign n12069 = pi102 & ~n2564;
  assign n12070 = ~n12068 & ~n12069;
  assign n12071 = ~pi562 & n12070;
  assign n12072 = ~n12055 & ~n12071;
  assign n12073 = pi295 & n12072;
  assign n12074 = ~pi295 & ~n12072;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = n6578 & n12075;
  assign n12077 = pi399 & ~n6578;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = ~n1761 & ~n12078;
  assign n12080 = ~n12048 & ~n12079;
  assign n12081 = ~n1754 & ~n12080;
  assign n12082 = pi873 & n12072;
  assign n12083 = ~pi873 & ~n12072;
  assign n12084 = ~n12082 & ~n12083;
  assign n12085 = n1754 & n12084;
  assign po548 = n12081 | n12085;
  assign n12087 = pi400 & n1761;
  assign n12088 = pi690 & ~n6579;
  assign n12089 = pi535 & n6579;
  assign n12090 = ~n12088 & ~n12089;
  assign n12091 = ~n2449 & ~n12090;
  assign n12092 = pi064 & n2449;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = pi562 & n12093;
  assign n12095 = pi535 & n6592;
  assign n12096 = pi064 & n6594;
  assign n12097 = ~n6594 & ~n12093;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = ~n6592 & ~n12098;
  assign n12100 = ~n12095 & ~n12099;
  assign n12101 = n6591 & ~n12100;
  assign n12102 = pi064 & ~pi669;
  assign n12103 = ~n6591 & n12102;
  assign n12104 = n6603 & ~n12100;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = ~n12101 & n12105;
  assign n12107 = n2564 & ~n12106;
  assign n12108 = pi064 & ~n2564;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~pi562 & n12109;
  assign n12111 = ~n12094 & ~n12110;
  assign n12112 = pi217 & n12111;
  assign n12113 = ~pi217 & ~n12111;
  assign n12114 = ~n12112 & ~n12113;
  assign n12115 = n6578 & n12114;
  assign n12116 = pi400 & ~n6578;
  assign n12117 = ~n12115 & ~n12116;
  assign n12118 = ~n1761 & ~n12117;
  assign n12119 = ~n12087 & ~n12118;
  assign n12120 = ~n1754 & ~n12119;
  assign n12121 = pi818 & n12111;
  assign n12122 = ~pi818 & ~n12111;
  assign n12123 = ~n12121 & ~n12122;
  assign n12124 = n1754 & n12123;
  assign po549 = n12120 | n12124;
  assign n12126 = pi401 & n1761;
  assign n12127 = pi742 & ~n6579;
  assign n12128 = pi627 & n6579;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~n2449 & ~n12129;
  assign n12131 = pi098 & n2449;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = pi562 & n12132;
  assign n12134 = pi627 & n6592;
  assign n12135 = pi098 & n6594;
  assign n12136 = ~n6594 & ~n12132;
  assign n12137 = ~n12135 & ~n12136;
  assign n12138 = ~n6592 & ~n12137;
  assign n12139 = ~n12134 & ~n12138;
  assign n12140 = n6591 & ~n12139;
  assign n12141 = pi098 & ~pi669;
  assign n12142 = ~n6591 & n12141;
  assign n12143 = n6603 & ~n12139;
  assign n12144 = ~n12142 & ~n12143;
  assign n12145 = ~n12140 & n12144;
  assign n12146 = n2564 & ~n12145;
  assign n12147 = pi098 & ~n2564;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = ~pi562 & n12148;
  assign n12150 = ~n12133 & ~n12149;
  assign n12151 = pi293 & n12150;
  assign n12152 = ~pi293 & ~n12150;
  assign n12153 = ~n12151 & ~n12152;
  assign n12154 = n6578 & n12153;
  assign n12155 = pi401 & ~n6578;
  assign n12156 = ~n12154 & ~n12155;
  assign n12157 = ~n1761 & ~n12156;
  assign n12158 = ~n12126 & ~n12157;
  assign n12159 = ~n1754 & ~n12158;
  assign n12160 = pi870 & n12150;
  assign n12161 = ~pi870 & ~n12150;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = n1754 & n12162;
  assign po550 = n12159 | n12163;
  assign n12165 = pi402 & n1761;
  assign n12166 = pi727 & ~n6579;
  assign n12167 = pi613 & n6579;
  assign n12168 = ~n12166 & ~n12167;
  assign n12169 = ~n2449 & ~n12168;
  assign n12170 = pi034 & n2449;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = pi562 & n12171;
  assign n12173 = pi613 & n6592;
  assign n12174 = pi034 & n6594;
  assign n12175 = ~n6594 & ~n12171;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = ~n6592 & ~n12176;
  assign n12178 = ~n12173 & ~n12177;
  assign n12179 = n6591 & ~n12178;
  assign n12180 = pi034 & ~pi669;
  assign n12181 = ~n6591 & n12180;
  assign n12182 = n6603 & ~n12178;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = ~n12179 & n12183;
  assign n12185 = n2564 & ~n12184;
  assign n12186 = pi034 & ~n2564;
  assign n12187 = ~n12185 & ~n12186;
  assign n12188 = ~pi562 & n12187;
  assign n12189 = ~n12172 & ~n12188;
  assign n12190 = ~pi246 & n12189;
  assign n12191 = pi246 & ~n12189;
  assign n12192 = ~n12190 & ~n12191;
  assign n12193 = n6578 & n12192;
  assign n12194 = pi402 & ~n6578;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = ~n1761 & ~n12195;
  assign n12197 = ~n12165 & ~n12196;
  assign n12198 = ~n1754 & ~n12197;
  assign n12199 = pi855 & n12189;
  assign n12200 = ~pi855 & ~n12189;
  assign n12201 = ~n12199 & ~n12200;
  assign n12202 = n1754 & n12201;
  assign po551 = n12198 | n12202;
  assign n12204 = pi403 & n1761;
  assign n12205 = pi787 & ~n6579;
  assign n12206 = pi651 & n6579;
  assign n12207 = ~n12205 & ~n12206;
  assign n12208 = ~n2449 & ~n12207;
  assign n12209 = pi181 & n2449;
  assign n12210 = ~n12208 & ~n12209;
  assign n12211 = pi562 & n12210;
  assign n12212 = pi651 & n6592;
  assign n12213 = pi181 & n6594;
  assign n12214 = ~n6594 & ~n12210;
  assign n12215 = ~n12213 & ~n12214;
  assign n12216 = ~n6592 & ~n12215;
  assign n12217 = ~n12212 & ~n12216;
  assign n12218 = n6591 & ~n12217;
  assign n12219 = pi181 & ~pi669;
  assign n12220 = ~n6591 & n12219;
  assign n12221 = n6603 & ~n12217;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = ~n12218 & n12222;
  assign n12224 = n2564 & ~n12223;
  assign n12225 = pi181 & ~n2564;
  assign n12226 = ~n12224 & ~n12225;
  assign n12227 = ~pi562 & n12226;
  assign n12228 = ~n12211 & ~n12227;
  assign n12229 = pi421 & n12228;
  assign n12230 = ~pi421 & ~n12228;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = n6578 & n12231;
  assign n12233 = pi403 & ~n6578;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = ~n1761 & ~n12234;
  assign n12236 = ~n12204 & ~n12235;
  assign n12237 = ~n1754 & ~n12236;
  assign n12238 = pi915 & n12228;
  assign n12239 = ~pi915 & ~n12228;
  assign n12240 = ~n12238 & ~n12239;
  assign n12241 = n1754 & n12240;
  assign po552 = n12237 | n12241;
  assign n12243 = pi404 & n1761;
  assign n12244 = pi693 & ~n6579;
  assign n12245 = pi511 & n6579;
  assign n12246 = ~n12244 & ~n12245;
  assign n12247 = ~n2449 & ~n12246;
  assign n12248 = pi090 & n2449;
  assign n12249 = ~n12247 & ~n12248;
  assign n12250 = pi562 & n12249;
  assign n12251 = pi511 & n6592;
  assign n12252 = pi090 & n6594;
  assign n12253 = ~n6594 & ~n12249;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = ~n6592 & ~n12254;
  assign n12256 = ~n12251 & ~n12255;
  assign n12257 = n6591 & ~n12256;
  assign n12258 = pi090 & ~pi669;
  assign n12259 = ~n6591 & n12258;
  assign n12260 = n6603 & ~n12256;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = ~n12257 & n12261;
  assign n12263 = n2564 & ~n12262;
  assign n12264 = pi090 & ~n2564;
  assign n12265 = ~n12263 & ~n12264;
  assign n12266 = ~pi562 & n12265;
  assign n12267 = ~n12250 & ~n12266;
  assign n12268 = pi218 & n12267;
  assign n12269 = ~pi218 & ~n12267;
  assign n12270 = ~n12268 & ~n12269;
  assign n12271 = n6578 & n12270;
  assign n12272 = pi404 & ~n6578;
  assign n12273 = ~n12271 & ~n12272;
  assign n12274 = ~n1761 & ~n12273;
  assign n12275 = ~n12243 & ~n12274;
  assign n12276 = ~n1754 & ~n12275;
  assign n12277 = pi821 & n12267;
  assign n12278 = ~pi821 & ~n12267;
  assign n12279 = ~n12277 & ~n12278;
  assign n12280 = n1754 & n12279;
  assign po553 = n12276 | n12280;
  assign n12282 = pi405 & n1761;
  assign n12283 = pi725 & ~n6579;
  assign n12284 = pi633 & n6579;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = ~n2449 & ~n12285;
  assign n12287 = pi094 & n2449;
  assign n12288 = ~n12286 & ~n12287;
  assign n12289 = pi562 & n12288;
  assign n12290 = pi633 & n6592;
  assign n12291 = pi094 & n6594;
  assign n12292 = ~n6594 & ~n12288;
  assign n12293 = ~n12291 & ~n12292;
  assign n12294 = ~n6592 & ~n12293;
  assign n12295 = ~n12290 & ~n12294;
  assign n12296 = n6591 & ~n12295;
  assign n12297 = pi094 & ~pi669;
  assign n12298 = ~n6591 & n12297;
  assign n12299 = n6603 & ~n12295;
  assign n12300 = ~n12298 & ~n12299;
  assign n12301 = ~n12296 & n12300;
  assign n12302 = n2564 & ~n12301;
  assign n12303 = pi094 & ~n2564;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = ~pi562 & n12304;
  assign n12306 = ~n12289 & ~n12305;
  assign n12307 = ~pi242 & n12306;
  assign n12308 = pi242 & ~n12306;
  assign n12309 = ~n12307 & ~n12308;
  assign n12310 = n6578 & n12309;
  assign n12311 = pi405 & ~n6578;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = ~n1761 & ~n12312;
  assign n12314 = ~n12282 & ~n12313;
  assign n12315 = ~n1754 & ~n12314;
  assign n12316 = pi853 & n12306;
  assign n12317 = ~pi853 & ~n12306;
  assign n12318 = ~n12316 & ~n12317;
  assign n12319 = n1754 & n12318;
  assign po554 = n12315 | n12319;
  assign n12321 = pi406 & n1761;
  assign n12322 = pi724 & ~n6579;
  assign n12323 = pi641 & n6579;
  assign n12324 = ~n12322 & ~n12323;
  assign n12325 = ~n2449 & ~n12324;
  assign n12326 = pi149 & n2449;
  assign n12327 = ~n12325 & ~n12326;
  assign n12328 = pi562 & n12327;
  assign n12329 = pi641 & n6592;
  assign n12330 = pi149 & n6594;
  assign n12331 = ~n6594 & ~n12327;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = ~n6592 & ~n12332;
  assign n12334 = ~n12329 & ~n12333;
  assign n12335 = n6591 & ~n12334;
  assign n12336 = pi149 & ~pi669;
  assign n12337 = ~n6591 & n12336;
  assign n12338 = n6603 & ~n12334;
  assign n12339 = ~n12337 & ~n12338;
  assign n12340 = ~n12335 & n12339;
  assign n12341 = n2564 & ~n12340;
  assign n12342 = pi149 & ~n2564;
  assign n12343 = ~n12341 & ~n12342;
  assign n12344 = ~pi562 & n12343;
  assign n12345 = ~n12328 & ~n12344;
  assign n12346 = ~pi241 & n12345;
  assign n12347 = pi241 & ~n12345;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = n6578 & n12348;
  assign n12350 = pi406 & ~n6578;
  assign n12351 = ~n12349 & ~n12350;
  assign n12352 = ~n1761 & ~n12351;
  assign n12353 = ~n12321 & ~n12352;
  assign n12354 = ~n1754 & ~n12353;
  assign n12355 = pi852 & n12345;
  assign n12356 = ~pi852 & ~n12345;
  assign n12357 = ~n12355 & ~n12356;
  assign n12358 = n1754 & n12357;
  assign po555 = n12354 | n12358;
  assign n12360 = pi407 & n1761;
  assign n12361 = pi692 & ~n6579;
  assign n12362 = pi519 & n6579;
  assign n12363 = ~n12361 & ~n12362;
  assign n12364 = ~n2449 & ~n12363;
  assign n12365 = pi147 & n2449;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = pi562 & n12366;
  assign n12368 = pi519 & n6592;
  assign n12369 = pi147 & n6594;
  assign n12370 = ~n6594 & ~n12366;
  assign n12371 = ~n12369 & ~n12370;
  assign n12372 = ~n6592 & ~n12371;
  assign n12373 = ~n12368 & ~n12372;
  assign n12374 = n6591 & ~n12373;
  assign n12375 = pi147 & ~pi669;
  assign n12376 = ~n6591 & n12375;
  assign n12377 = n6603 & ~n12373;
  assign n12378 = ~n12376 & ~n12377;
  assign n12379 = ~n12374 & n12378;
  assign n12380 = n2564 & ~n12379;
  assign n12381 = pi147 & ~n2564;
  assign n12382 = ~n12380 & ~n12381;
  assign n12383 = ~pi562 & n12382;
  assign n12384 = ~n12367 & ~n12383;
  assign n12385 = pi219 & n12384;
  assign n12386 = ~pi219 & ~n12384;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = n6578 & n12387;
  assign n12389 = pi407 & ~n6578;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391 = ~n1761 & ~n12390;
  assign n12392 = ~n12360 & ~n12391;
  assign n12393 = ~n1754 & ~n12392;
  assign n12394 = pi820 & n12384;
  assign n12395 = ~pi820 & ~n12384;
  assign n12396 = ~n12394 & ~n12395;
  assign n12397 = n1754 & n12396;
  assign po556 = n12393 | n12397;
  assign n12399 = pi408 & n1761;
  assign n12400 = pi722 & ~n6579;
  assign n12401 = pi583 & n6579;
  assign n12402 = ~n12400 & ~n12401;
  assign n12403 = ~n2449 & ~n12402;
  assign n12404 = pi068 & n2449;
  assign n12405 = ~n12403 & ~n12404;
  assign n12406 = pi562 & n12405;
  assign n12407 = pi583 & n6592;
  assign n12408 = pi068 & n6594;
  assign n12409 = ~n6594 & ~n12405;
  assign n12410 = ~n12408 & ~n12409;
  assign n12411 = ~n6592 & ~n12410;
  assign n12412 = ~n12407 & ~n12411;
  assign n12413 = n6591 & ~n12412;
  assign n12414 = pi068 & ~pi669;
  assign n12415 = ~n6591 & n12414;
  assign n12416 = n6603 & ~n12412;
  assign n12417 = ~n12415 & ~n12416;
  assign n12418 = ~n12413 & n12417;
  assign n12419 = n2564 & ~n12418;
  assign n12420 = pi068 & ~n2564;
  assign n12421 = ~n12419 & ~n12420;
  assign n12422 = ~pi562 & n12421;
  assign n12423 = ~n12406 & ~n12422;
  assign n12424 = ~pi245 & n12423;
  assign n12425 = pi245 & ~n12423;
  assign n12426 = ~n12424 & ~n12425;
  assign n12427 = n6578 & n12426;
  assign n12428 = pi408 & ~n6578;
  assign n12429 = ~n12427 & ~n12428;
  assign n12430 = ~n1761 & ~n12429;
  assign n12431 = ~n12399 & ~n12430;
  assign n12432 = ~n1754 & ~n12431;
  assign n12433 = pi850 & n12423;
  assign n12434 = ~pi850 & ~n12423;
  assign n12435 = ~n12433 & ~n12434;
  assign n12436 = n1754 & n12435;
  assign po557 = n12432 | n12436;
  assign n12438 = pi409 & ~po814;
  assign n12439 = po814 & ~n6027;
  assign po558 = n12438 | n12439;
  assign n12441 = ~pi410 & ~n10112;
  assign n12442 = ~n9605 & ~n12441;
  assign n12443 = n9610 & n10112;
  assign n12444 = ~pi410 & ~n12443;
  assign n12445 = ~n9696 & n10361;
  assign n12446 = n9696 & ~n10361;
  assign n12447 = ~n12445 & ~n12446;
  assign n12448 = n9873 & ~n10243;
  assign n12449 = ~n9873 & n10243;
  assign n12450 = ~n12448 & ~n12449;
  assign n12451 = ~n10186 & n12450;
  assign n12452 = n10186 & ~n12450;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12447 & n12453;
  assign n12455 = n12447 & ~n12453;
  assign n12456 = ~n12454 & ~n12455;
  assign n12457 = ~pi673 & ~n12456;
  assign n12458 = ~n9804 & n9826;
  assign n12459 = n9804 & ~n9826;
  assign n12460 = ~n12458 & ~n12459;
  assign n12461 = n10276 & ~n12460;
  assign n12462 = ~n10276 & n12460;
  assign n12463 = ~n12461 & ~n12462;
  assign n12464 = pi060 & ~n2449;
  assign n12465 = pi307 & n2449;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = n9619 & ~n12466;
  assign n12468 = pi310 & n2449;
  assign n12469 = pi058 & ~n2449;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = n9611 & ~n12470;
  assign n12472 = ~n12467 & ~n12471;
  assign n12473 = pi059 & ~n2449;
  assign n12474 = pi299 & n2449;
  assign n12475 = ~n12473 & ~n12474;
  assign n12476 = n9622 & ~n12475;
  assign n12477 = pi264 & n2449;
  assign n12478 = pi061 & ~n2449;
  assign n12479 = ~n12477 & ~n12478;
  assign n12480 = po815 & ~n12479;
  assign n12481 = ~n12476 & ~n12480;
  assign n12482 = n12472 & n12481;
  assign n12483 = pi376 & n2449;
  assign n12484 = pi067 & ~n2449;
  assign n12485 = ~n12483 & ~n12484;
  assign n12486 = n9611 & ~n12485;
  assign n12487 = pi092 & ~n2449;
  assign n12488 = pi374 & n2449;
  assign n12489 = ~n12487 & ~n12488;
  assign n12490 = n9622 & ~n12489;
  assign n12491 = pi266 & n2449;
  assign n12492 = ~pi062 & ~n2449;
  assign n12493 = ~n12491 & ~n12492;
  assign n12494 = po815 & ~n12493;
  assign n12495 = ~n12490 & ~n12494;
  assign n12496 = pi353 & n2449;
  assign n12497 = pi065 & ~n2449;
  assign n12498 = ~n12496 & ~n12497;
  assign n12499 = n9619 & ~n12498;
  assign n12500 = n12495 & ~n12499;
  assign n12501 = ~n12486 & n12500;
  assign n12502 = n12482 & n12501;
  assign n12503 = ~n12482 & ~n12501;
  assign n12504 = ~n12502 & ~n12503;
  assign n12505 = ~n10186 & ~n12504;
  assign n12506 = n10186 & n12504;
  assign n12507 = ~n12505 & ~n12506;
  assign n12508 = n10364 & n12507;
  assign n12509 = ~n10364 & ~n12507;
  assign n12510 = ~n12508 & ~n12509;
  assign n12511 = pi064 & ~n2449;
  assign n12512 = pi400 & n2449;
  assign n12513 = ~n12511 & ~n12512;
  assign n12514 = po815 & ~n12513;
  assign n12515 = pi352 & n2449;
  assign n12516 = pi063 & ~n2449;
  assign n12517 = ~n12515 & ~n12516;
  assign n12518 = n9611 & ~n12517;
  assign n12519 = ~n12514 & ~n12518;
  assign n12520 = pi068 & ~n2449;
  assign n12521 = pi408 & n2449;
  assign n12522 = ~n12520 & ~n12521;
  assign n12523 = n9622 & ~n12522;
  assign n12524 = pi366 & n2449;
  assign n12525 = pi066 & ~n2449;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = n9619 & ~n12526;
  assign n12528 = ~n12523 & ~n12527;
  assign n12529 = n12519 & n12528;
  assign n12530 = pi373 & n2449;
  assign n12531 = pi109 & ~n2449;
  assign n12532 = ~n12530 & ~n12531;
  assign n12533 = n9619 & ~n12532;
  assign n12534 = pi322 & n2449;
  assign n12535 = pi106 & ~n2449;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = n9611 & ~n12536;
  assign n12538 = pi108 & ~n2449;
  assign n12539 = pi330 & n2449;
  assign n12540 = ~n12538 & ~n12539;
  assign n12541 = n9622 & ~n12540;
  assign n12542 = pi107 & ~n2449;
  assign n12543 = pi306 & n2449;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = po815 & ~n12544;
  assign n12546 = ~n12541 & ~n12545;
  assign n12547 = ~n12537 & n12546;
  assign n12548 = ~n12533 & n12547;
  assign n12549 = n12529 & n12548;
  assign n12550 = ~n12529 & ~n12548;
  assign n12551 = ~n12549 & ~n12550;
  assign n12552 = n12456 & n12551;
  assign n12553 = ~n12456 & ~n12551;
  assign n12554 = ~n12552 & ~n12553;
  assign n12555 = ~n12510 & n12554;
  assign n12556 = n12510 & ~n12554;
  assign n12557 = ~n12555 & ~n12556;
  assign n12558 = ~n12463 & n12557;
  assign n12559 = n12463 & ~n12557;
  assign n12560 = ~n12558 & ~n12559;
  assign n12561 = pi673 & ~n12560;
  assign n12562 = ~n12457 & ~n12561;
  assign n12563 = n9610 & ~n12562;
  assign n12564 = ~n12444 & ~n12563;
  assign n12565 = ~n12442 & ~n12564;
  assign n12566 = ~pi410 & po815;
  assign po559 = n12565 | n12566;
  assign n12568 = n9718 & ~n10161;
  assign n12569 = ~n9718 & n10161;
  assign n12570 = ~n12568 & ~n12569;
  assign n12571 = n9892 & n10243;
  assign n12572 = ~n9892 & ~n10243;
  assign n12573 = ~n12571 & ~n12572;
  assign n12574 = ~n10326 & ~n12573;
  assign n12575 = n10326 & n12573;
  assign n12576 = ~n12574 & ~n12575;
  assign n12577 = ~n12570 & n12576;
  assign n12578 = n12570 & ~n12576;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = ~pi673 & ~n12579;
  assign n12581 = n9785 & ~n9845;
  assign n12582 = ~n9785 & n9845;
  assign n12583 = ~n12581 & ~n12582;
  assign n12584 = n10096 & ~n12583;
  assign n12585 = ~n10096 & n12583;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = n12482 & ~n12529;
  assign n12588 = ~n12482 & n12529;
  assign n12589 = ~n12587 & ~n12588;
  assign n12590 = ~n10326 & n12589;
  assign n12591 = n10326 & ~n12589;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n9759 & n12592;
  assign n12594 = n9759 & ~n12592;
  assign n12595 = ~n12593 & ~n12594;
  assign n12596 = ~n12501 & n12548;
  assign n12597 = n12501 & ~n12548;
  assign n12598 = ~n12596 & ~n12597;
  assign n12599 = n12579 & ~n12598;
  assign n12600 = ~n12579 & n12598;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = ~n12595 & n12601;
  assign n12603 = n12595 & ~n12601;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = ~n12586 & n12604;
  assign n12606 = n12586 & ~n12604;
  assign n12607 = ~n12605 & ~n12606;
  assign n12608 = pi673 & ~n12607;
  assign n12609 = ~n12580 & ~n12608;
  assign n12610 = n9610 & ~n12609;
  assign n12611 = ~pi411 & ~n9610;
  assign n12612 = ~n12610 & ~n12611;
  assign n12613 = n9605 & ~n12612;
  assign n12614 = ~pi411 & ~n10112;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = ~pi411 & po815;
  assign po560 = ~n12615 | n12616;
  assign n12618 = ~n9715 & ~n10323;
  assign n12619 = n9715 & n10323;
  assign n12620 = ~n12618 & ~n12619;
  assign n12621 = n9873 & n10224;
  assign n12622 = ~n9873 & ~n10224;
  assign n12623 = ~n12621 & ~n12622;
  assign n12624 = ~n9759 & ~n12623;
  assign n12625 = n9759 & n12623;
  assign n12626 = ~n12624 & ~n12625;
  assign n12627 = ~n12620 & n12626;
  assign n12628 = n12620 & ~n12626;
  assign n12629 = ~n12627 & ~n12628;
  assign n12630 = ~pi673 & ~n12629;
  assign n12631 = ~n9759 & n12598;
  assign n12632 = n9759 & ~n12598;
  assign n12633 = ~n12631 & ~n12632;
  assign n12634 = ~n10326 & n12633;
  assign n12635 = n10326 & ~n12633;
  assign n12636 = ~n12634 & ~n12635;
  assign n12637 = ~n12589 & n12629;
  assign n12638 = n12589 & ~n12629;
  assign n12639 = ~n12637 & ~n12638;
  assign n12640 = ~n12636 & n12639;
  assign n12641 = n12636 & ~n12639;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = ~n12586 & n12642;
  assign n12644 = n12586 & ~n12642;
  assign n12645 = ~n12643 & ~n12644;
  assign n12646 = pi673 & ~n12645;
  assign n12647 = ~n12630 & ~n12646;
  assign n12648 = n9610 & ~n12647;
  assign n12649 = ~pi412 & ~n9610;
  assign n12650 = ~n12648 & ~n12649;
  assign n12651 = n9605 & ~n12650;
  assign n12652 = ~pi412 & ~n10112;
  assign n12653 = ~n12651 & ~n12652;
  assign n12654 = ~pi412 & po815;
  assign po561 = ~n12653 | n12654;
  assign n12656 = pi413 & ~po814;
  assign n12657 = po814 & ~n5979;
  assign po562 = n12656 | n12657;
  assign n12659 = pi414 & ~po814;
  assign n12660 = po814 & ~n5737;
  assign po563 = n12659 | n12660;
  assign n12662 = pi415 & ~po814;
  assign n12663 = po814 & ~n5835;
  assign po564 = n12662 | n12663;
  assign n12665 = pi416 & ~po814;
  assign n12666 = po814 & ~n5883;
  assign po565 = n12665 | n12666;
  assign n12668 = pi417 & ~po814;
  assign n12669 = po814 & ~n5931;
  assign po566 = n12668 | n12669;
  assign n12671 = pi418 & ~po814;
  assign n12672 = po814 & ~n6123;
  assign po567 = n12671 | n12672;
  assign n12674 = pi419 & ~po814;
  assign n12675 = po814 & ~n6075;
  assign po568 = n12674 | n12675;
  assign n12677 = ~pi420 & ~n10112;
  assign n12678 = n10164 & ~n10320;
  assign n12679 = ~n10164 & n10320;
  assign n12680 = ~n12678 & ~n12679;
  assign n12681 = n9892 & ~n10224;
  assign n12682 = ~n9892 & n10224;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~n10364 & n12683;
  assign n12685 = n10364 & ~n12683;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = ~n12680 & ~n12686;
  assign n12688 = n12680 & n12686;
  assign n12689 = ~n12687 & ~n12688;
  assign n12690 = ~pi673 & ~n12689;
  assign n12691 = n10364 & ~n12551;
  assign n12692 = ~n10364 & n12551;
  assign n12693 = ~n12691 & ~n12692;
  assign n12694 = ~n10186 & n12693;
  assign n12695 = n10186 & ~n12693;
  assign n12696 = ~n12694 & ~n12695;
  assign n12697 = n12504 & n12689;
  assign n12698 = ~n12504 & ~n12689;
  assign n12699 = ~n12697 & ~n12698;
  assign n12700 = ~n12696 & n12699;
  assign n12701 = n12696 & ~n12699;
  assign n12702 = ~n12700 & ~n12701;
  assign n12703 = ~n12463 & n12702;
  assign n12704 = n12463 & ~n12702;
  assign n12705 = ~n12703 & ~n12704;
  assign n12706 = pi673 & ~n12705;
  assign n12707 = ~n12690 & ~n12706;
  assign n12708 = n9610 & ~n12707;
  assign n12709 = ~pi420 & ~n9610;
  assign n12710 = ~n12708 & ~n12709;
  assign n12711 = n9605 & ~n12710;
  assign n12712 = ~n12677 & ~n12711;
  assign n12713 = ~pi420 & po815;
  assign po569 = ~n12712 | n12713;
  assign n12715 = pi421 & ~po814;
  assign n12716 = po814 & ~n6177;
  assign po570 = n12715 | n12716;
  assign n12718 = n9622 & ~n10107;
  assign n12719 = ~n9605 & ~n9619;
  assign n12720 = ~pi422 & ~n12719;
  assign n12721 = ~n12718 & ~n12720;
  assign n12722 = ~pi422 & po815;
  assign po571 = ~n12721 | n12722;
  assign n12724 = n9622 & ~n10287;
  assign n12725 = ~pi423 & ~n12719;
  assign n12726 = ~n12724 & ~n12725;
  assign n12727 = ~pi423 & po815;
  assign po572 = ~n12726 | n12727;
  assign n12729 = n9622 & ~n10382;
  assign n12730 = ~pi424 & ~n12719;
  assign n12731 = ~n12729 & ~n12730;
  assign n12732 = ~pi424 & po815;
  assign po573 = ~n12731 | n12732;
  assign n12734 = n9619 & ~n10107;
  assign n12735 = ~n9605 & ~n9622;
  assign n12736 = ~pi425 & ~n12735;
  assign n12737 = ~n12734 & ~n12736;
  assign n12738 = ~pi425 & po815;
  assign po574 = ~n12737 | n12738;
  assign n12740 = n9622 & ~n10344;
  assign n12741 = ~pi426 & ~n12719;
  assign n12742 = ~n12740 & ~n12741;
  assign n12743 = ~pi426 & po815;
  assign po575 = ~n12742 | n12743;
  assign n12745 = n9619 & ~n10344;
  assign n12746 = ~pi427 & ~n12735;
  assign n12747 = ~n12745 & ~n12746;
  assign n12748 = ~pi427 & po815;
  assign po576 = ~n12747 | n12748;
  assign n12750 = n9619 & ~n10287;
  assign n12751 = ~pi428 & ~n12735;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = ~pi428 & po815;
  assign po577 = ~n12752 | n12753;
  assign n12755 = n9619 & ~n10382;
  assign n12756 = ~pi429 & ~n12735;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = ~pi429 & po815;
  assign po578 = ~n12757 | n12758;
  assign n12760 = pi430 & ~po814;
  assign n12761 = po814 & ~n6225;
  assign po579 = n12760 | n12761;
  assign n12763 = pi431 & ~po814;
  assign n12764 = po814 & ~n6273;
  assign po580 = n12763 | n12764;
  assign n12766 = pi432 & ~po814;
  assign n12767 = po814 & ~n6465;
  assign po581 = n12766 | n12767;
  assign n12769 = pi433 & ~po814;
  assign n12770 = po814 & ~n6321;
  assign po582 = n12769 | n12770;
  assign n12772 = pi434 & ~po814;
  assign n12773 = po814 & ~n6417;
  assign po583 = n12772 | n12773;
  assign n12775 = n1791 & n6577;
  assign po584 = n1754 | n12775;
  assign n12777 = pi436 & ~po814;
  assign n12778 = po814 & ~n6369;
  assign po585 = n12777 | n12778;
  assign n12780 = pi437 & ~po814;
  assign n12781 = po814 & ~n5796;
  assign po586 = n12780 | n12781;
  assign n12783 = ~n9785 & n10199;
  assign n12784 = n9785 & ~n10199;
  assign n12785 = ~n12783 & ~n12784;
  assign n12786 = ~n12507 & n12785;
  assign n12787 = n12507 & ~n12785;
  assign n12788 = ~n12786 & ~n12787;
  assign n12789 = ~pi673 & ~n12788;
  assign n12790 = n10279 & n12788;
  assign n12791 = ~n10279 & ~n12788;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = pi673 & ~n12792;
  assign n12794 = ~n12789 & ~n12793;
  assign n12795 = n9610 & ~n12794;
  assign n12796 = ~pi438 & ~n9610;
  assign n12797 = ~n12795 & ~n12796;
  assign n12798 = n9605 & ~n12797;
  assign n12799 = ~pi438 & ~n10112;
  assign n12800 = ~n12798 & ~n12799;
  assign n12801 = ~pi438 & po815;
  assign po587 = ~n12800 | n12801;
  assign n12803 = ~n9873 & n12683;
  assign n12804 = n9873 & ~n12683;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = ~n10196 & ~n12805;
  assign n12807 = n10196 & n12805;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = ~pi673 & ~n12808;
  assign n12810 = n12482 & ~n12548;
  assign n12811 = ~n12482 & n12548;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = ~n10186 & ~n10364;
  assign n12814 = n10186 & n10364;
  assign n12815 = ~n12813 & ~n12814;
  assign n12816 = ~n12812 & n12815;
  assign n12817 = n12812 & ~n12815;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = ~n10261 & n12808;
  assign n12820 = n10261 & ~n12808;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n12818 & n12821;
  assign n12823 = n12818 & ~n12821;
  assign n12824 = ~n12822 & ~n12823;
  assign n12825 = pi673 & ~n12824;
  assign n12826 = ~n12809 & ~n12825;
  assign n12827 = n9610 & ~n12826;
  assign n12828 = ~pi439 & ~n9610;
  assign n12829 = ~n12827 & ~n12828;
  assign n12830 = n9605 & ~n12829;
  assign n12831 = ~pi439 & ~n10112;
  assign n12832 = ~n12830 & ~n12831;
  assign n12833 = ~pi439 & po815;
  assign po588 = ~n12832 | n12833;
  assign n12835 = n9807 & ~n9826;
  assign n12836 = ~n9807 & n9826;
  assign n12837 = ~n12835 & ~n12836;
  assign n12838 = ~n12592 & n12837;
  assign n12839 = n12592 & ~n12837;
  assign n12840 = ~n12838 & ~n12839;
  assign n12841 = ~pi673 & ~n12840;
  assign n12842 = ~n10099 & n12840;
  assign n12843 = n10099 & ~n12840;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = pi673 & ~n12844;
  assign n12846 = ~n12841 & ~n12845;
  assign n12847 = n9610 & ~n12846;
  assign n12848 = ~pi440 & ~n9610;
  assign n12849 = ~n12847 & ~n12848;
  assign n12850 = n9605 & ~n12849;
  assign n12851 = ~pi440 & ~n10112;
  assign n12852 = ~n12850 & ~n12851;
  assign n12853 = ~pi440 & po815;
  assign po589 = ~n12852 | n12853;
  assign n12855 = ~n10243 & ~n12623;
  assign n12856 = n10243 & n12623;
  assign n12857 = ~n12855 & ~n12856;
  assign n12858 = ~n9848 & ~n12857;
  assign n12859 = n9848 & n12857;
  assign n12860 = ~n12858 & ~n12859;
  assign n12861 = ~pi673 & ~n12860;
  assign n12862 = ~n12501 & n12529;
  assign n12863 = n12501 & ~n12529;
  assign n12864 = ~n12862 & ~n12863;
  assign n12865 = n9759 & ~n10326;
  assign n12866 = ~n9759 & n10326;
  assign n12867 = ~n12865 & ~n12866;
  assign n12868 = ~n12864 & n12867;
  assign n12869 = n12864 & ~n12867;
  assign n12870 = ~n12868 & ~n12869;
  assign n12871 = ~n10005 & n12860;
  assign n12872 = n10005 & ~n12860;
  assign n12873 = ~n12871 & ~n12872;
  assign n12874 = ~n12870 & n12873;
  assign n12875 = n12870 & ~n12873;
  assign n12876 = ~n12874 & ~n12875;
  assign n12877 = pi673 & ~n12876;
  assign n12878 = ~n12861 & ~n12877;
  assign n12879 = n9610 & ~n12878;
  assign n12880 = ~pi441 & ~n9610;
  assign n12881 = ~n12879 & ~n12880;
  assign n12882 = n9605 & ~n12881;
  assign n12883 = ~pi441 & ~n10112;
  assign n12884 = ~n12882 & ~n12883;
  assign n12885 = ~pi441 & po815;
  assign po590 = ~n12884 | n12885;
  assign n12887 = ~n9845 & ~n10196;
  assign n12888 = n9845 & n10196;
  assign n12889 = ~n12887 & ~n12888;
  assign n12890 = ~n12693 & n12889;
  assign n12891 = n12693 & ~n12889;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = ~pi673 & ~n12892;
  assign n12894 = n10279 & n12892;
  assign n12895 = ~n10279 & ~n12892;
  assign n12896 = ~n12894 & ~n12895;
  assign n12897 = pi673 & ~n12896;
  assign n12898 = ~n12893 & ~n12897;
  assign n12899 = n9610 & ~n12898;
  assign n12900 = ~pi442 & ~n9610;
  assign n12901 = ~n12899 & ~n12900;
  assign n12902 = n9605 & ~n12901;
  assign n12903 = ~pi442 & ~n10112;
  assign n12904 = ~n12902 & ~n12903;
  assign n12905 = ~pi442 & po815;
  assign po591 = ~n12904 | n12905;
  assign n12907 = ~pi443 & ~n10112;
  assign n12908 = ~n9892 & n12450;
  assign n12909 = n9892 & ~n12450;
  assign n12910 = ~n12908 & ~n12909;
  assign n12911 = n10199 & ~n12910;
  assign n12912 = ~n10199 & n12910;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = ~pi673 & ~n12913;
  assign n12915 = n10261 & ~n12913;
  assign n12916 = ~n10261 & n12913;
  assign n12917 = ~n12915 & ~n12916;
  assign n12918 = ~n12818 & n12917;
  assign n12919 = n12818 & ~n12917;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = pi673 & ~n12920;
  assign n12922 = ~n12914 & ~n12921;
  assign n12923 = n9610 & ~n12922;
  assign n12924 = ~pi443 & ~n9610;
  assign n12925 = ~n12923 & ~n12924;
  assign n12926 = n9605 & ~n12925;
  assign n12927 = ~n12907 & ~n12926;
  assign n12928 = ~pi443 & po815;
  assign po592 = ~n12927 | n12928;
  assign n12930 = n9622 & ~n12647;
  assign n12931 = ~pi444 & ~n12719;
  assign n12932 = ~n12930 & ~n12931;
  assign n12933 = ~pi444 & po815;
  assign po593 = ~n12932 | n12933;
  assign n12935 = n9622 & ~n12562;
  assign n12936 = ~pi445 & ~n12719;
  assign n12937 = ~n12935 & ~n12936;
  assign n12938 = ~pi445 & po815;
  assign po594 = ~n12937 | n12938;
  assign n12940 = n9622 & ~n12609;
  assign n12941 = ~pi446 & ~n12719;
  assign n12942 = ~n12940 & ~n12941;
  assign n12943 = ~pi446 & po815;
  assign po595 = ~n12942 | n12943;
  assign n12945 = n9622 & ~n12707;
  assign n12946 = ~pi447 & ~n12719;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = ~pi447 & po815;
  assign po596 = ~n12947 | n12948;
  assign n12950 = n9619 & ~n12647;
  assign n12951 = ~pi448 & ~n12735;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = ~pi448 & po815;
  assign po597 = ~n12952 | n12953;
  assign n12955 = n9619 & ~n12562;
  assign n12956 = ~pi449 & ~n12735;
  assign n12957 = ~n12955 & ~n12956;
  assign n12958 = ~pi449 & po815;
  assign po598 = ~n12957 | n12958;
  assign n12960 = ~n9804 & ~n9848;
  assign n12961 = n9804 & n9848;
  assign n12962 = ~n12960 & ~n12961;
  assign n12963 = ~n12633 & n12962;
  assign n12964 = n12633 & ~n12962;
  assign n12965 = ~n12963 & ~n12964;
  assign n12966 = ~pi673 & ~n12965;
  assign n12967 = ~n10099 & n12965;
  assign n12968 = n10099 & ~n12965;
  assign n12969 = ~n12967 & ~n12968;
  assign n12970 = pi673 & ~n12969;
  assign n12971 = ~n12966 & ~n12970;
  assign n12972 = n9610 & ~n12971;
  assign n12973 = ~pi450 & ~n9610;
  assign n12974 = ~n12972 & ~n12973;
  assign n12975 = n9605 & ~n12974;
  assign n12976 = ~pi450 & ~n10112;
  assign n12977 = ~n12975 & ~n12976;
  assign n12978 = ~pi450 & po815;
  assign po599 = ~n12977 | n12978;
  assign n12980 = ~n10224 & ~n12573;
  assign n12981 = n10224 & n12573;
  assign n12982 = ~n12980 & ~n12981;
  assign n12983 = n9807 & ~n12982;
  assign n12984 = ~n9807 & n12982;
  assign n12985 = ~n12983 & ~n12984;
  assign n12986 = ~pi673 & ~n12985;
  assign n12987 = ~n10005 & n12985;
  assign n12988 = n10005 & ~n12985;
  assign n12989 = ~n12987 & ~n12988;
  assign n12990 = ~n12870 & n12989;
  assign n12991 = n12870 & ~n12989;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = pi673 & ~n12992;
  assign n12994 = ~n12986 & ~n12993;
  assign n12995 = n9610 & ~n12994;
  assign n12996 = ~pi451 & ~n9610;
  assign n12997 = ~n12995 & ~n12996;
  assign n12998 = n9605 & ~n12997;
  assign n12999 = ~pi451 & ~n10112;
  assign n13000 = ~n12998 & ~n12999;
  assign n13001 = ~pi451 & po815;
  assign po600 = ~n13000 | n13001;
  assign n13003 = n9619 & ~n12707;
  assign n13004 = ~pi452 & ~n12735;
  assign n13005 = ~n13003 & ~n13004;
  assign n13006 = ~pi452 & po815;
  assign po601 = ~n13005 | n13006;
  assign n13008 = n9619 & ~n12609;
  assign n13009 = ~pi453 & ~n12735;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~pi453 & po815;
  assign po602 = ~n13010 | n13011;
  assign n13013 = ~n12504 & ~n12529;
  assign n13014 = n12504 & n12529;
  assign n13015 = ~n13013 & ~n13014;
  assign n13016 = n10364 & n13015;
  assign n13017 = ~n10364 & ~n13015;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = ~pi673 & ~n13018;
  assign n13020 = ~n10276 & n13018;
  assign n13021 = n10276 & ~n13018;
  assign n13022 = ~n13020 & ~n13021;
  assign n13023 = pi673 & ~n13022;
  assign n13024 = ~n13019 & ~n13023;
  assign n13025 = n9610 & ~n13024;
  assign n13026 = ~pi454 & ~n9610;
  assign n13027 = ~n13025 & ~n13026;
  assign n13028 = n9605 & ~n13027;
  assign n13029 = ~pi454 & ~n10112;
  assign n13030 = ~n13028 & ~n13029;
  assign n13031 = ~pi454 & po815;
  assign po603 = ~n13030 | n13031;
  assign n13033 = ~n10046 & n10090;
  assign n13034 = n10046 & ~n10090;
  assign n13035 = ~n13033 & ~n13034;
  assign n13036 = ~n9674 & ~n13035;
  assign n13037 = n9674 & n13035;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = ~pi673 & ~n13038;
  assign n13040 = ~n9696 & n12576;
  assign n13041 = n9696 & ~n12576;
  assign n13042 = ~n13040 & ~n13041;
  assign n13043 = ~n12626 & n13042;
  assign n13044 = n12626 & ~n13042;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = n10005 & ~n10320;
  assign n13047 = ~n10005 & n10320;
  assign n13048 = ~n13046 & ~n13047;
  assign n13049 = ~n13038 & n13048;
  assign n13050 = n13038 & ~n13048;
  assign n13051 = ~n13049 & ~n13050;
  assign n13052 = ~n13045 & n13051;
  assign n13053 = n13045 & ~n13051;
  assign n13054 = ~n13052 & ~n13053;
  assign n13055 = pi673 & ~n13054;
  assign n13056 = ~n13039 & ~n13055;
  assign n13057 = n9610 & ~n13056;
  assign n13058 = ~pi455 & ~n9610;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = n9605 & ~n13059;
  assign n13061 = ~pi455 & ~n10112;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = ~pi455 & po815;
  assign po604 = ~n13062 | n13063;
  assign n13065 = ~n10027 & n10267;
  assign n13066 = n10027 & ~n10267;
  assign n13067 = ~n13065 & ~n13066;
  assign n13068 = n10139 & ~n13067;
  assign n13069 = ~n10139 & n13067;
  assign n13070 = ~n13068 & ~n13069;
  assign n13071 = ~pi673 & ~n13070;
  assign n13072 = ~n10161 & ~n12686;
  assign n13073 = n10161 & n12686;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = n12453 & ~n13074;
  assign n13076 = ~n12453 & n13074;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = ~n9715 & n10261;
  assign n13079 = n9715 & ~n10261;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = ~n13070 & n13080;
  assign n13082 = n13070 & ~n13080;
  assign n13083 = ~n13081 & ~n13082;
  assign n13084 = ~n13077 & n13083;
  assign n13085 = n13077 & ~n13083;
  assign n13086 = ~n13084 & ~n13085;
  assign n13087 = pi673 & ~n13086;
  assign n13088 = ~n13071 & ~n13087;
  assign n13089 = n9610 & ~n13088;
  assign n13090 = ~pi456 & ~n9610;
  assign n13091 = ~n13089 & ~n13090;
  assign n13092 = n9605 & ~n13091;
  assign n13093 = ~pi456 & ~n10112;
  assign n13094 = ~n13092 & ~n13093;
  assign n13095 = ~pi456 & po815;
  assign po605 = ~n13094 | n13095;
  assign n13097 = n9958 & ~n9996;
  assign n13098 = ~n9958 & n9996;
  assign n13099 = ~n13097 & ~n13098;
  assign n13100 = ~n10049 & n13099;
  assign n13101 = n10049 & ~n13099;
  assign n13102 = ~n13100 & ~n13101;
  assign n13103 = ~pi673 & ~n13102;
  assign n13104 = ~n9718 & n13102;
  assign n13105 = n9718 & ~n13102;
  assign n13106 = ~n13104 & ~n13105;
  assign n13107 = ~n9652 & n10136;
  assign n13108 = n9652 & ~n10136;
  assign n13109 = ~n13107 & ~n13108;
  assign n13110 = ~n9759 & n10329;
  assign n13111 = n9759 & ~n10329;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = ~n13109 & n13112;
  assign n13114 = n13109 & ~n13112;
  assign n13115 = ~n13113 & ~n13114;
  assign n13116 = ~n13106 & n13115;
  assign n13117 = n13106 & ~n13115;
  assign n13118 = ~n13116 & ~n13117;
  assign n13119 = pi673 & ~n13118;
  assign n13120 = ~n13103 & ~n13119;
  assign n13121 = n9610 & ~n13120;
  assign n13122 = ~pi457 & ~n9610;
  assign n13123 = ~n13121 & ~n13122;
  assign n13124 = n9605 & ~n13123;
  assign n13125 = ~pi457 & ~n10112;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = ~pi457 & po815;
  assign po606 = ~n13126 | n13127;
  assign n13129 = ~n12501 & ~n12551;
  assign n13130 = n12501 & n12551;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = ~n10186 & n13131;
  assign n13133 = n10186 & ~n13131;
  assign n13134 = ~n13132 & ~n13133;
  assign n13135 = ~pi673 & ~n13134;
  assign n13136 = ~n10276 & n13134;
  assign n13137 = n10276 & ~n13134;
  assign n13138 = ~n13136 & ~n13137;
  assign n13139 = pi673 & ~n13138;
  assign n13140 = ~n13135 & ~n13139;
  assign n13141 = n9610 & ~n13140;
  assign n13142 = ~pi458 & ~n9610;
  assign n13143 = ~n13141 & ~n13142;
  assign n13144 = n9605 & ~n13143;
  assign n13145 = ~pi458 & ~n10112;
  assign n13146 = ~n13144 & ~n13145;
  assign n13147 = ~pi458 & po815;
  assign po607 = ~n13146 | n13147;
  assign n13149 = ~n12482 & n12598;
  assign n13150 = n12482 & ~n12598;
  assign n13151 = ~n13149 & ~n13150;
  assign n13152 = ~n10326 & n13151;
  assign n13153 = n10326 & ~n13151;
  assign n13154 = ~n13152 & ~n13153;
  assign n13155 = ~pi673 & ~n13154;
  assign n13156 = ~n10096 & n13154;
  assign n13157 = n10096 & ~n13154;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = pi673 & ~n13158;
  assign n13160 = ~n13155 & ~n13159;
  assign n13161 = n9610 & ~n13160;
  assign n13162 = ~pi459 & ~n9610;
  assign n13163 = ~n13161 & ~n13162;
  assign n13164 = n9605 & ~n13163;
  assign n13165 = ~pi459 & ~n10112;
  assign n13166 = ~n13164 & ~n13165;
  assign n13167 = ~pi459 & po815;
  assign po608 = ~n13166 | n13167;
  assign n13169 = ~n12548 & n12589;
  assign n13170 = n12548 & ~n12589;
  assign n13171 = ~n13169 & ~n13170;
  assign n13172 = ~n9759 & n13171;
  assign n13173 = n9759 & ~n13171;
  assign n13174 = ~n13172 & ~n13173;
  assign n13175 = ~pi673 & ~n13174;
  assign n13176 = ~n10096 & n13174;
  assign n13177 = n10096 & ~n13174;
  assign n13178 = ~n13176 & ~n13177;
  assign n13179 = pi673 & ~n13178;
  assign n13180 = ~n13175 & ~n13179;
  assign n13181 = n9610 & ~n13180;
  assign n13182 = ~pi460 & ~n9610;
  assign n13183 = ~n13181 & ~n13182;
  assign n13184 = n9605 & ~n13183;
  assign n13185 = ~pi460 & ~n10112;
  assign n13186 = ~n13184 & ~n13185;
  assign n13187 = ~pi460 & po815;
  assign po609 = ~n13186 | n13187;
  assign n13189 = ~n9977 & n10252;
  assign n13190 = n9977 & ~n10252;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n10270 & n13191;
  assign n13193 = n10270 & ~n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = ~pi673 & ~n13194;
  assign n13196 = ~n10164 & n13194;
  assign n13197 = n10164 & ~n13194;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = ~n9633 & n9671;
  assign n13200 = n9633 & ~n9671;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = ~n10186 & n10367;
  assign n13203 = n10186 & ~n10367;
  assign n13204 = ~n13202 & ~n13203;
  assign n13205 = ~n13201 & n13204;
  assign n13206 = n13201 & ~n13204;
  assign n13207 = ~n13205 & ~n13206;
  assign n13208 = ~n13198 & n13207;
  assign n13209 = n13198 & ~n13207;
  assign n13210 = ~n13208 & ~n13209;
  assign n13211 = pi673 & ~n13210;
  assign n13212 = ~n13195 & ~n13211;
  assign n13213 = n9610 & ~n13212;
  assign n13214 = ~pi461 & ~n9610;
  assign n13215 = ~n13213 & ~n13214;
  assign n13216 = n9605 & ~n13215;
  assign n13217 = ~pi461 & ~n10112;
  assign n13218 = ~n13216 & ~n13217;
  assign n13219 = ~pi461 & po815;
  assign po610 = ~n13218 | n13219;
  assign n13221 = ~n9936 & n10255;
  assign n13222 = n9936 & ~n10255;
  assign n13223 = ~n13221 & ~n13222;
  assign n13224 = ~n10267 & n13223;
  assign n13225 = n10267 & ~n13223;
  assign n13226 = ~n13224 & ~n13225;
  assign n13227 = ~pi673 & ~n13226;
  assign n13228 = ~n10361 & n13226;
  assign n13229 = n10361 & ~n13226;
  assign n13230 = ~n13228 & ~n13229;
  assign n13231 = n10189 & n10364;
  assign n13232 = ~n10189 & ~n10364;
  assign n13233 = ~n13231 & ~n13232;
  assign n13234 = ~n13201 & n13233;
  assign n13235 = n13201 & ~n13233;
  assign n13236 = ~n13234 & ~n13235;
  assign n13237 = ~n13230 & n13236;
  assign n13238 = n13230 & ~n13236;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = pi673 & ~n13239;
  assign n13241 = ~n13227 & ~n13240;
  assign n13242 = n9610 & ~n13241;
  assign n13243 = ~pi462 & ~n9610;
  assign n13244 = ~n13242 & ~n13243;
  assign n13245 = n9605 & ~n13244;
  assign n13246 = ~pi462 & ~n10112;
  assign n13247 = ~n13245 & ~n13246;
  assign n13248 = ~pi462 & po815;
  assign po611 = ~n13247 | n13248;
  assign n13250 = ~n9955 & n9999;
  assign n13251 = n9955 & ~n9999;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = ~n10090 & n13252;
  assign n13254 = n10090 & ~n13252;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = ~pi673 & ~n13255;
  assign n13257 = n10323 & n13255;
  assign n13258 = ~n10323 & ~n13255;
  assign n13259 = ~n13257 & ~n13258;
  assign n13260 = n9762 & ~n10326;
  assign n13261 = ~n9762 & n10326;
  assign n13262 = ~n13260 & ~n13261;
  assign n13263 = ~n13109 & n13262;
  assign n13264 = n13109 & ~n13262;
  assign n13265 = ~n13263 & ~n13264;
  assign n13266 = ~n13259 & n13265;
  assign n13267 = n13259 & ~n13265;
  assign n13268 = ~n13266 & ~n13267;
  assign n13269 = pi673 & ~n13268;
  assign n13270 = ~n13256 & ~n13269;
  assign n13271 = n9610 & ~n13270;
  assign n13272 = ~pi463 & ~n9610;
  assign n13273 = ~n13271 & ~n13272;
  assign n13274 = n9605 & ~n13273;
  assign n13275 = ~pi463 & ~n10112;
  assign n13276 = ~n13274 & ~n13275;
  assign n13277 = ~pi463 & po815;
  assign po612 = ~n13276 | n13277;
  assign n13279 = ~n10068 & n10270;
  assign n13280 = n10068 & ~n10270;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = n10355 & ~n13281;
  assign n13283 = ~n10355 & n13281;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = ~pi673 & ~n13284;
  assign n13286 = ~n9715 & n12453;
  assign n13287 = n9715 & ~n12453;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = ~n12686 & ~n13288;
  assign n13290 = n12686 & n13288;
  assign n13291 = ~n13289 & ~n13290;
  assign n13292 = ~n10161 & n10261;
  assign n13293 = n10161 & ~n10261;
  assign n13294 = ~n13292 & ~n13293;
  assign n13295 = ~n13284 & n13294;
  assign n13296 = n13284 & ~n13294;
  assign n13297 = ~n13295 & ~n13296;
  assign n13298 = ~n13291 & n13297;
  assign n13299 = n13291 & ~n13297;
  assign n13300 = ~n13298 & ~n13299;
  assign n13301 = pi673 & ~n13300;
  assign n13302 = ~n13285 & ~n13301;
  assign n13303 = n9610 & ~n13302;
  assign n13304 = ~pi464 & ~n9610;
  assign n13305 = ~n13303 & ~n13304;
  assign n13306 = n9605 & ~n13305;
  assign n13307 = ~pi464 & ~n10112;
  assign n13308 = ~n13306 & ~n13307;
  assign n13309 = ~pi464 & po815;
  assign po613 = ~n13308 | n13309;
  assign n13311 = n10049 & ~n10087;
  assign n13312 = ~n10049 & n10087;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = ~n10298 & ~n13313;
  assign n13315 = n10298 & n13313;
  assign n13316 = ~n13314 & ~n13315;
  assign n13317 = ~pi673 & ~n13316;
  assign n13318 = ~n10320 & n12626;
  assign n13319 = n10320 & ~n12626;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n12576 & n13320;
  assign n13322 = n12576 & ~n13320;
  assign n13323 = ~n13321 & ~n13322;
  assign n13324 = ~n9696 & n10005;
  assign n13325 = n9696 & ~n10005;
  assign n13326 = ~n13324 & ~n13325;
  assign n13327 = ~n13316 & n13326;
  assign n13328 = n13316 & ~n13326;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = ~n13323 & n13329;
  assign n13331 = n13323 & ~n13329;
  assign n13332 = ~n13330 & ~n13331;
  assign n13333 = pi673 & ~n13332;
  assign n13334 = ~n13317 & ~n13333;
  assign n13335 = n9610 & ~n13334;
  assign n13336 = ~pi465 & ~n9610;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = n9605 & ~n13337;
  assign n13339 = ~pi465 & ~n10112;
  assign n13340 = ~n13338 & ~n13339;
  assign n13341 = ~pi465 & po815;
  assign po614 = ~n13340 | n13341;
  assign n13343 = ~n9622 & n12719;
  assign n13344 = pi466 & ~n13343;
  assign n13345 = po815 & ~n10287;
  assign po615 = n13344 | n13345;
  assign n13347 = pi467 & ~n13343;
  assign n13348 = po815 & ~n10344;
  assign po616 = n13347 | n13348;
  assign n13350 = pi468 & ~n13343;
  assign n13351 = po815 & ~n10382;
  assign po617 = n13350 | n13351;
  assign n13353 = pi469 & ~n13343;
  assign n13354 = po815 & ~n10107;
  assign po618 = n13353 | n13354;
  assign n13356 = n9622 & ~n12971;
  assign n13357 = ~pi470 & ~n12719;
  assign n13358 = ~n13356 & ~n13357;
  assign n13359 = ~pi470 & po815;
  assign po619 = ~n13358 | n13359;
  assign n13361 = n9622 & ~n12994;
  assign n13362 = ~pi471 & ~n12719;
  assign n13363 = ~n13361 & ~n13362;
  assign n13364 = ~pi471 & po815;
  assign po620 = ~n13363 | n13364;
  assign n13366 = n9622 & ~n12826;
  assign n13367 = ~pi472 & ~n12719;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = ~pi472 & po815;
  assign po621 = ~n13368 | n13369;
  assign n13371 = n9622 & ~n12794;
  assign n13372 = ~pi473 & ~n12719;
  assign n13373 = ~n13371 & ~n13372;
  assign n13374 = ~pi473 & po815;
  assign po622 = ~n13373 | n13374;
  assign n13376 = n9622 & ~n12846;
  assign n13377 = ~pi474 & ~n12719;
  assign n13378 = ~n13376 & ~n13377;
  assign n13379 = ~pi474 & po815;
  assign po623 = ~n13378 | n13379;
  assign n13381 = n9622 & ~n12878;
  assign n13382 = ~pi475 & ~n12719;
  assign n13383 = ~n13381 & ~n13382;
  assign n13384 = ~pi475 & po815;
  assign po624 = ~n13383 | n13384;
  assign n13386 = n9622 & ~n12898;
  assign n13387 = ~pi476 & ~n12719;
  assign n13388 = ~n13386 & ~n13387;
  assign n13389 = ~pi476 & po815;
  assign po625 = ~n13388 | n13389;
  assign n13391 = n9622 & ~n12922;
  assign n13392 = ~pi477 & ~n12719;
  assign n13393 = ~n13391 & ~n13392;
  assign n13394 = ~pi477 & po815;
  assign po626 = ~n13393 | n13394;
  assign n13396 = n9619 & ~n12971;
  assign n13397 = ~pi478 & ~n12735;
  assign n13398 = ~n13396 & ~n13397;
  assign n13399 = ~pi478 & po815;
  assign po627 = ~n13398 | n13399;
  assign n13401 = n9619 & ~n12994;
  assign n13402 = ~pi479 & ~n12735;
  assign n13403 = ~n13401 & ~n13402;
  assign n13404 = ~pi479 & po815;
  assign po628 = ~n13403 | n13404;
  assign n13406 = n9619 & ~n12826;
  assign n13407 = ~pi480 & ~n12735;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = ~pi480 & po815;
  assign po629 = ~n13408 | n13409;
  assign n13411 = n9619 & ~n12794;
  assign n13412 = ~pi481 & ~n12735;
  assign n13413 = ~n13411 & ~n13412;
  assign n13414 = ~pi481 & po815;
  assign po630 = ~n13413 | n13414;
  assign n13416 = n9619 & ~n12846;
  assign n13417 = ~pi482 & ~n12735;
  assign n13418 = ~n13416 & ~n13417;
  assign n13419 = ~pi482 & po815;
  assign po631 = ~n13418 | n13419;
  assign n13421 = n9619 & ~n12878;
  assign n13422 = ~pi483 & ~n12735;
  assign n13423 = ~n13421 & ~n13422;
  assign n13424 = ~pi483 & po815;
  assign po632 = ~n13423 | n13424;
  assign n13426 = n9619 & ~n12898;
  assign n13427 = ~pi484 & ~n12735;
  assign n13428 = ~n13426 & ~n13427;
  assign n13429 = ~pi484 & po815;
  assign po633 = ~n13428 | n13429;
  assign n13431 = n9619 & ~n12922;
  assign n13432 = ~pi485 & ~n12735;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = ~pi485 & po815;
  assign po634 = ~n13433 | n13434;
  assign n13436 = n9622 & ~n13088;
  assign n13437 = ~pi486 & ~n12719;
  assign n13438 = ~n13436 & ~n13437;
  assign n13439 = ~pi486 & po815;
  assign po635 = ~n13438 | n13439;
  assign n13441 = n9622 & ~n13212;
  assign n13442 = ~pi487 & ~n12719;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~pi487 & po815;
  assign po636 = ~n13443 | n13444;
  assign n13446 = n9619 & ~n13334;
  assign n13447 = ~pi488 & ~n12735;
  assign n13448 = ~n13446 & ~n13447;
  assign n13449 = ~pi488 & po815;
  assign po637 = ~n13448 | n13449;
  assign n13451 = n9622 & ~n13302;
  assign n13452 = ~pi489 & ~n12719;
  assign n13453 = ~n13451 & ~n13452;
  assign n13454 = ~pi489 & po815;
  assign po638 = ~n13453 | n13454;
  assign n13456 = n9622 & ~n13334;
  assign n13457 = ~pi490 & ~n12719;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = ~pi490 & po815;
  assign po639 = ~n13458 | n13459;
  assign n13461 = n9622 & ~n13056;
  assign n13462 = ~pi491 & ~n12719;
  assign n13463 = ~n13461 & ~n13462;
  assign n13464 = ~pi491 & po815;
  assign po640 = ~n13463 | n13464;
  assign n13466 = n9619 & ~n13302;
  assign n13467 = ~pi492 & ~n12735;
  assign n13468 = ~n13466 & ~n13467;
  assign n13469 = ~pi492 & po815;
  assign po641 = ~n13468 | n13469;
  assign n13471 = pi493 & ~n13343;
  assign n13472 = po815 & ~n12647;
  assign po642 = n13471 | n13472;
  assign n13474 = n9622 & ~n13270;
  assign n13475 = ~pi494 & ~n12719;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~pi494 & po815;
  assign po643 = ~n13476 | n13477;
  assign n13479 = n9622 & ~n13241;
  assign n13480 = ~pi495 & ~n12719;
  assign n13481 = ~n13479 & ~n13480;
  assign n13482 = ~pi495 & po815;
  assign po644 = ~n13481 | n13482;
  assign n13484 = n9622 & ~n13120;
  assign n13485 = ~pi496 & ~n12719;
  assign n13486 = ~n13484 & ~n13485;
  assign n13487 = ~pi496 & po815;
  assign po645 = ~n13486 | n13487;
  assign n13489 = n9619 & ~n13270;
  assign n13490 = ~pi497 & ~n12735;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = ~pi497 & po815;
  assign po646 = ~n13491 | n13492;
  assign n13494 = n9619 & ~n13241;
  assign n13495 = ~pi498 & ~n12735;
  assign n13496 = ~n13494 & ~n13495;
  assign n13497 = ~pi498 & po815;
  assign po647 = ~n13496 | n13497;
  assign n13499 = n9619 & ~n13120;
  assign n13500 = ~pi499 & ~n12735;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = ~pi499 & po815;
  assign po648 = ~n13501 | n13502;
  assign n13504 = n9619 & ~n13212;
  assign n13505 = ~pi500 & ~n12735;
  assign n13506 = ~n13504 & ~n13505;
  assign n13507 = ~pi500 & po815;
  assign po649 = ~n13506 | n13507;
  assign n13509 = n9622 & ~n13180;
  assign n13510 = ~pi501 & ~n12719;
  assign n13511 = ~n13509 & ~n13510;
  assign n13512 = ~pi501 & po815;
  assign po650 = ~n13511 | n13512;
  assign n13514 = n9622 & ~n13160;
  assign n13515 = ~pi502 & ~n12719;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = ~pi502 & po815;
  assign po651 = ~n13516 | n13517;
  assign n13519 = n9622 & ~n13024;
  assign n13520 = ~pi503 & ~n12719;
  assign n13521 = ~n13519 & ~n13520;
  assign n13522 = ~pi503 & po815;
  assign po652 = ~n13521 | n13522;
  assign n13524 = n9619 & ~n13180;
  assign n13525 = ~pi504 & ~n12735;
  assign n13526 = ~n13524 & ~n13525;
  assign n13527 = ~pi504 & po815;
  assign po653 = ~n13526 | n13527;
  assign n13529 = n9619 & ~n13024;
  assign n13530 = ~pi505 & ~n12735;
  assign n13531 = ~n13529 & ~n13530;
  assign n13532 = ~pi505 & po815;
  assign po654 = ~n13531 | n13532;
  assign n13534 = n9619 & ~n13160;
  assign n13535 = ~pi506 & ~n12735;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = ~pi506 & po815;
  assign po655 = ~n13536 | n13537;
  assign n13539 = n9619 & ~n13140;
  assign n13540 = ~pi507 & ~n12735;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = ~pi507 & po815;
  assign po656 = ~n13541 | n13542;
  assign n13544 = n9622 & ~n13140;
  assign n13545 = ~pi508 & ~n12719;
  assign n13546 = ~n13544 & ~n13545;
  assign n13547 = ~pi508 & po815;
  assign po657 = ~n13546 | n13547;
  assign n13549 = pi509 & ~n13343;
  assign n13550 = po815 & ~n12707;
  assign po658 = n13549 | n13550;
  assign n13552 = pi510 & ~n13343;
  assign n13553 = po815 & ~n12562;
  assign po659 = n13552 | n13553;
  assign n13555 = pi511 & ~n13343;
  assign n13556 = po815 & ~n12609;
  assign po660 = n13555 | n13556;
  assign n13558 = n9619 & ~n13056;
  assign n13559 = ~pi512 & ~n12735;
  assign n13560 = ~n13558 & ~n13559;
  assign n13561 = ~pi512 & po815;
  assign po661 = ~n13560 | n13561;
  assign n13563 = n9619 & ~n13088;
  assign n13564 = ~pi513 & ~n12735;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = ~pi513 & po815;
  assign po662 = ~n13565 | n13566;
  assign n13568 = ~n9737 & n10326;
  assign n13569 = n9737 & ~n10326;
  assign n13570 = ~n13568 & ~n13569;
  assign n13571 = ~n9958 & n13570;
  assign n13572 = n9958 & ~n13570;
  assign n13573 = ~n13571 & ~n13572;
  assign n13574 = ~pi673 & ~n13573;
  assign n13575 = ~n9674 & n10298;
  assign n13576 = n9674 & ~n10298;
  assign n13577 = ~n13575 & ~n13576;
  assign n13578 = n10027 & ~n10068;
  assign n13579 = ~n10027 & n10068;
  assign n13580 = ~n13578 & ~n13579;
  assign n13581 = n13573 & ~n13580;
  assign n13582 = ~n13573 & n13580;
  assign n13583 = ~n13581 & ~n13582;
  assign n13584 = ~n13577 & n13583;
  assign n13585 = n13577 & ~n13583;
  assign n13586 = ~n13584 & ~n13585;
  assign n13587 = pi673 & ~n13586;
  assign n13588 = ~n13574 & ~n13587;
  assign n13589 = n9610 & ~n13588;
  assign n13590 = ~pi514 & ~n9610;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = n9605 & ~n13591;
  assign n13593 = ~pi514 & ~n10112;
  assign n13594 = ~n13592 & ~n13593;
  assign n13595 = ~pi514 & po815;
  assign po663 = ~n13594 | n13595;
  assign n13597 = ~n9756 & ~n10364;
  assign n13598 = n9756 & n10364;
  assign n13599 = ~n13597 & ~n13598;
  assign n13600 = ~n10252 & n13599;
  assign n13601 = n10252 & ~n13599;
  assign n13602 = ~n13600 & ~n13601;
  assign n13603 = ~pi673 & ~n13602;
  assign n13604 = ~n10139 & n10355;
  assign n13605 = n10139 & ~n10355;
  assign n13606 = ~n13604 & ~n13605;
  assign n13607 = n10046 & ~n10087;
  assign n13608 = ~n10046 & n10087;
  assign n13609 = ~n13607 & ~n13608;
  assign n13610 = n13602 & ~n13609;
  assign n13611 = ~n13602 & n13609;
  assign n13612 = ~n13610 & ~n13611;
  assign n13613 = ~n13606 & n13612;
  assign n13614 = n13606 & ~n13612;
  assign n13615 = ~n13613 & ~n13614;
  assign n13616 = pi673 & ~n13615;
  assign n13617 = ~n13603 & ~n13616;
  assign n13618 = n9610 & ~n13617;
  assign n13619 = ~pi515 & ~n9610;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = n9605 & ~n13620;
  assign n13622 = ~pi515 & ~n10112;
  assign n13623 = ~n13621 & ~n13622;
  assign n13624 = ~pi515 & po815;
  assign po664 = ~n13623 | n13624;
  assign n13626 = ~n9914 & n10186;
  assign n13627 = n9914 & ~n10186;
  assign n13628 = ~n13626 & ~n13627;
  assign n13629 = ~n10255 & n13628;
  assign n13630 = n10255 & ~n13628;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~pi673 & ~n13631;
  assign n13633 = ~n13609 & n13631;
  assign n13634 = n13609 & ~n13631;
  assign n13635 = ~n13633 & ~n13634;
  assign n13636 = ~n13606 & n13635;
  assign n13637 = n13606 & ~n13635;
  assign n13638 = ~n13636 & ~n13637;
  assign n13639 = pi673 & ~n13638;
  assign n13640 = ~n13632 & ~n13639;
  assign n13641 = n9610 & ~n13640;
  assign n13642 = ~pi516 & ~n9610;
  assign n13643 = ~n13641 & ~n13642;
  assign n13644 = n9605 & ~n13643;
  assign n13645 = ~pi516 & ~n10112;
  assign n13646 = ~n13644 & ~n13645;
  assign n13647 = ~pi516 & po815;
  assign po665 = ~n13646 | n13647;
  assign n13649 = n9759 & ~n10183;
  assign n13650 = ~n9759 & n10183;
  assign n13651 = ~n13649 & ~n13650;
  assign n13652 = ~n9999 & n13651;
  assign n13653 = n9999 & ~n13651;
  assign n13654 = ~n13652 & ~n13653;
  assign n13655 = ~pi673 & ~n13654;
  assign n13656 = ~n13580 & n13654;
  assign n13657 = n13580 & ~n13654;
  assign n13658 = ~n13656 & ~n13657;
  assign n13659 = ~n13577 & n13658;
  assign n13660 = n13577 & ~n13658;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = pi673 & ~n13661;
  assign n13663 = ~n13655 & ~n13662;
  assign n13664 = n9610 & ~n13663;
  assign n13665 = ~pi517 & ~n9610;
  assign n13666 = ~n13664 & ~n13665;
  assign n13667 = n9605 & ~n13666;
  assign n13668 = ~pi517 & ~n10112;
  assign n13669 = ~n13667 & ~n13668;
  assign n13670 = ~pi517 & po815;
  assign po666 = ~n13669 | n13670;
  assign n13672 = pi518 & ~n13343;
  assign n13673 = po815 & ~n12846;
  assign po667 = n13672 | n13673;
  assign n13675 = pi519 & ~n13343;
  assign n13676 = po815 & ~n12878;
  assign po668 = n13675 | n13676;
  assign n13678 = pi520 & ~n13343;
  assign n13679 = po815 & ~n12971;
  assign po669 = n13678 | n13679;
  assign n13681 = pi521 & ~n13343;
  assign n13682 = po815 & ~n12898;
  assign po670 = n13681 | n13682;
  assign n13684 = pi522 & ~n13343;
  assign n13685 = po815 & ~n12922;
  assign po671 = n13684 | n13685;
  assign n13687 = pi523 & ~n13343;
  assign n13688 = po815 & ~n12794;
  assign po672 = n13687 | n13688;
  assign n13690 = pi524 & ~n13343;
  assign n13691 = po815 & ~n12994;
  assign po673 = n13690 | n13691;
  assign n13693 = pi525 & ~n13343;
  assign n13694 = po815 & ~n12826;
  assign po674 = n13693 | n13694;
  assign n13696 = n9619 & ~n13617;
  assign n13697 = ~pi526 & ~n12735;
  assign n13698 = ~n13696 & ~n13697;
  assign n13699 = ~pi526 & po815;
  assign po675 = ~n13698 | n13699;
  assign n13701 = pi527 & ~n13343;
  assign n13702 = po815 & ~n13140;
  assign po676 = n13701 | n13702;
  assign n13704 = n9622 & ~n13663;
  assign n13705 = ~pi528 & ~n12719;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = ~pi528 & po815;
  assign po677 = ~n13706 | n13707;
  assign n13709 = n9619 & ~n13588;
  assign n13710 = ~pi529 & ~n12735;
  assign n13711 = ~n13709 & ~n13710;
  assign n13712 = ~pi529 & po815;
  assign po678 = ~n13711 | n13712;
  assign n13714 = pi530 & ~n13343;
  assign n13715 = po815 & ~n13302;
  assign po679 = n13714 | n13715;
  assign n13717 = pi531 & ~n13343;
  assign n13718 = po815 & ~n13056;
  assign po680 = n13717 | n13718;
  assign n13720 = n9622 & ~n13640;
  assign n13721 = ~pi532 & ~n12719;
  assign n13722 = ~n13720 & ~n13721;
  assign n13723 = ~pi532 & po815;
  assign po681 = ~n13722 | n13723;
  assign n13725 = pi533 & ~n13343;
  assign n13726 = po815 & ~n13120;
  assign po682 = n13725 | n13726;
  assign n13728 = pi534 & ~n13343;
  assign n13729 = po815 & ~n13212;
  assign po683 = n13728 | n13729;
  assign n13731 = pi535 & ~n13343;
  assign n13732 = po815 & ~n13160;
  assign po684 = n13731 | n13732;
  assign n13734 = n9622 & ~n13617;
  assign n13735 = ~pi536 & ~n12719;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = ~pi536 & po815;
  assign po685 = ~n13736 | n13737;
  assign n13739 = n9622 & ~n13588;
  assign n13740 = ~pi537 & ~n12719;
  assign n13741 = ~n13739 & ~n13740;
  assign n13742 = ~pi537 & po815;
  assign po686 = ~n13741 | n13742;
  assign n13744 = pi538 & ~n13343;
  assign n13745 = po815 & ~n13270;
  assign po687 = n13744 | n13745;
  assign n13747 = pi539 & ~n13343;
  assign n13748 = po815 & ~n13241;
  assign po688 = n13747 | n13748;
  assign n13750 = pi540 & ~n13343;
  assign n13751 = po815 & ~n13180;
  assign po689 = n13750 | n13751;
  assign n13753 = pi541 & ~n13343;
  assign n13754 = po815 & ~n13024;
  assign po690 = n13753 | n13754;
  assign n13756 = n9619 & ~n13640;
  assign n13757 = ~pi542 & ~n12735;
  assign n13758 = ~n13756 & ~n13757;
  assign n13759 = ~pi542 & po815;
  assign po691 = ~n13758 | n13759;
  assign n13761 = pi543 & ~n13343;
  assign n13762 = po815 & ~n13088;
  assign po692 = n13761 | n13762;
  assign n13764 = pi544 & ~n13343;
  assign n13765 = po815 & ~n13334;
  assign po693 = n13764 | n13765;
  assign n13767 = n9619 & ~n13663;
  assign n13768 = ~pi545 & ~n12735;
  assign n13769 = ~n13767 & ~n13768;
  assign n13770 = ~pi545 & po815;
  assign po694 = ~n13769 | n13770;
  assign n13772 = pi546 & ~n13343;
  assign n13773 = po815 & ~n13588;
  assign po695 = n13772 | n13773;
  assign n13775 = pi547 & ~n13343;
  assign n13776 = po815 & ~n13663;
  assign po696 = n13775 | n13776;
  assign n13778 = pi548 & ~n13343;
  assign n13779 = po815 & ~n13640;
  assign po697 = n13778 | n13779;
  assign n13781 = pi549 & ~n13343;
  assign n13782 = po815 & ~n13617;
  assign po698 = n13781 | n13782;
  assign n13784 = n5295 & ~n6577;
  assign n13785 = ~n5294 & ~n13784;
  assign n13786 = n5290 & ~n13785;
  assign po699 = n5298 | n13786;
  assign n13788 = n5305 & ~n6577;
  assign n13789 = ~n5304 & ~n13788;
  assign n13790 = n5290 & ~n13789;
  assign po700 = n5308 | n13790;
  assign n13792 = n5314 & ~n6577;
  assign n13793 = ~n5313 & ~n13792;
  assign n13794 = n5290 & ~n13793;
  assign po701 = n5310 | n13794;
  assign n13796 = n2018 & ~n2019;
  assign n13797 = pi553 & n2019;
  assign n13798 = ~n13796 & ~n13797;
  assign po702 = n2023 | ~n13798;
  assign n13800 = n2019 & n2022;
  assign n13801 = pi554 & n13800;
  assign n13802 = ~n2019 & n2440;
  assign po703 = n13801 | n13802;
  assign n13804 = pi562 & ~pi672;
  assign n13805 = pi555 & n13804;
  assign n13806 = ~pi435 & n2565;
  assign n13807 = ~pi562 & n2564;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = pi555 & ~n6594;
  assign n13810 = pi555 & pi557;
  assign n13811 = ~n1751 & ~n13810;
  assign n13812 = n6594 & ~n13811;
  assign n13813 = ~n13809 & ~n13812;
  assign n13814 = ~n6592 & ~n13813;
  assign n13815 = ~pi555 & pi557;
  assign n13816 = pi555 & ~pi557;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = n6592 & ~n13817;
  assign n13819 = ~n13814 & ~n13818;
  assign n13820 = n6591 & ~n13819;
  assign n13821 = pi669 & ~n13819;
  assign n13822 = ~pi669 & ~n13817;
  assign n13823 = ~n13821 & ~n13822;
  assign n13824 = ~n6591 & ~n13823;
  assign n13825 = ~n13820 & ~n13824;
  assign n13826 = ~n13808 & ~n13825;
  assign n13827 = ~n13805 & ~n13826;
  assign po816 = pi562 & pi672;
  assign n13829 = pi673 & po816;
  assign po704 = ~n13827 | n13829;
  assign n13831 = pi556 & n13810;
  assign n13832 = ~pi556 & ~n13810;
  assign n13833 = ~n13831 & ~n13832;
  assign n13834 = n6592 & ~n13833;
  assign n13835 = pi556 & ~n1751;
  assign n13836 = ~n1752 & ~n13835;
  assign n13837 = n6594 & ~n13836;
  assign n13838 = pi556 & ~n6594;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = ~n6592 & n13839;
  assign n13841 = ~n13834 & ~n13840;
  assign n13842 = pi669 & ~n13841;
  assign n13843 = ~pi669 & ~n13833;
  assign n13844 = ~n13842 & ~n13843;
  assign n13845 = ~n6591 & n13844;
  assign n13846 = n6591 & n13841;
  assign n13847 = ~n13845 & ~n13846;
  assign n13848 = ~n13808 & ~n13847;
  assign n13849 = pi556 & pi562;
  assign n13850 = ~pi672 & n13849;
  assign po705 = n13848 | n13850;
  assign n13852 = pi557 & n6594;
  assign n13853 = ~pi557 & ~n6594;
  assign n13854 = ~n13852 & ~n13853;
  assign n13855 = ~n6592 & ~n13854;
  assign n13856 = pi557 & n6592;
  assign n13857 = ~n13855 & ~n13856;
  assign n13858 = pi669 & ~n13857;
  assign n13859 = pi557 & ~pi669;
  assign n13860 = ~n13858 & ~n13859;
  assign n13861 = ~n6591 & n13860;
  assign n13862 = n6591 & n13857;
  assign n13863 = ~n13861 & ~n13862;
  assign n13864 = ~n13808 & ~n13863;
  assign n13865 = pi557 & pi562;
  assign n13866 = ~pi672 & n13865;
  assign po706 = n13864 | n13866;
  assign n13868 = pi558 & n13804;
  assign n13869 = pi558 & n13831;
  assign n13870 = ~pi558 & ~n13831;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = n6592 & ~n13871;
  assign n13873 = pi558 & ~n1752;
  assign n13874 = ~n1753 & ~n13873;
  assign n13875 = n6594 & ~n13874;
  assign n13876 = pi558 & ~n6594;
  assign n13877 = ~n13875 & ~n13876;
  assign n13878 = ~n6592 & n13877;
  assign n13879 = ~n13872 & ~n13878;
  assign n13880 = n6591 & n13879;
  assign n13881 = pi669 & ~n13879;
  assign n13882 = ~pi669 & ~n13871;
  assign n13883 = ~n13881 & ~n13882;
  assign n13884 = ~n6591 & n13883;
  assign n13885 = ~n13880 & ~n13884;
  assign n13886 = ~n13808 & ~n13885;
  assign n13887 = ~n13868 & ~n13886;
  assign po707 = n13829 | ~n13887;
  assign n13889 = pi667 & ~n6594;
  assign n13890 = ~n6592 & n13889;
  assign n13891 = n6591 & ~n13890;
  assign n13892 = ~pi669 & ~n6591;
  assign n13893 = ~n13891 & ~n13892;
  assign n13894 = n13807 & ~n13893;
  assign n13895 = pi562 & ~pi667;
  assign n13896 = ~n13894 & ~n13895;
  assign n13897 = n13806 & ~n13893;
  assign po708 = ~n13896 | n13897;
  assign n13899 = ~pi560 & ~n9610;
  assign n13900 = n9605 & ~n13899;
  assign po709 = n9622 | n13900;
  assign n13902 = n9605 & ~n9610;
  assign n13903 = pi561 & n13902;
  assign n13904 = ~n9622 & ~n13903;
  assign po710 = n9619 | ~n13904;
  assign n13906 = pi435 & ~n2564;
  assign n13907 = ~pi562 & ~n13906;
  assign po711 = po816 | n13907;
  assign n13909 = ~pi563 & ~n2572;
  assign n13910 = n2558 & ~n13909;
  assign n13911 = ~pi563 & n2559;
  assign po712 = n13910 | n13911;
  assign po713 = pi435 & n2565;
  assign n13914 = pi565 & ~n2494;
  assign n13915 = ~n2495 & ~n13914;
  assign n13916 = n2559 & ~n13915;
  assign n13917 = pi565 & n2558;
  assign n13918 = ~n2572 & n13917;
  assign po714 = n13916 | n13918;
  assign n13920 = pi566 & n2558;
  assign n13921 = ~n2572 & n13920;
  assign n13922 = ~pi566 & ~n2460;
  assign n13923 = ~n2494 & ~n13922;
  assign n13924 = n2559 & n13923;
  assign po715 = n13921 | n13924;
  assign n13926 = pi567 & n2558;
  assign n13927 = ~n2572 & n13926;
  assign n13928 = ~n2454 & ~n2474;
  assign n13929 = n2559 & ~n13928;
  assign po716 = n13927 | n13929;
  assign n13931 = pi568 & n2558;
  assign n13932 = ~n2572 & n13931;
  assign n13933 = pi568 & n2517;
  assign n13934 = ~pi568 & ~n2517;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = n2559 & n13935;
  assign po717 = n13932 | n13936;
  assign n13938 = pi569 & ~n13343;
  assign po718 = n13147 | n13938;
  assign n13940 = pi570 & ~n13343;
  assign po719 = n13277 | n13940;
  assign n13942 = pi571 & ~n13343;
  assign po720 = n12801 | n13942;
  assign n13944 = pi572 & ~n13343;
  assign po721 = n10293 | n13944;
  assign n13946 = pi573 & ~n13343;
  assign po722 = n13248 | n13946;
  assign n13948 = pi574 & ~n13343;
  assign po723 = n13167 | n13948;
  assign n13950 = pi575 & ~n13343;
  assign po724 = n13454 | n13950;
  assign n13952 = pi576 & ~n13343;
  assign po725 = n12953 | n13952;
  assign n13954 = pi577 & ~n13343;
  assign po726 = n13492 | n13954;
  assign n13956 = pi578 & ~n13343;
  assign po727 = n13561 | n13956;
  assign n13958 = pi579 & ~n13343;
  assign po728 = n13001 | n13958;
  assign n13960 = pi580 & ~n13343;
  assign po729 = n13424 | n13960;
  assign n13962 = pi581 & ~n13343;
  assign po730 = n12654 | n13962;
  assign n13964 = pi582 & ~n13343;
  assign po731 = n13542 | n13964;
  assign n13966 = pi583 & ~n13343;
  assign po732 = n13517 | n13966;
  assign n13968 = pi584 & ~n13343;
  assign po733 = n13006 | n13968;
  assign n13970 = pi585 & ~n13343;
  assign po734 = n13449 | n13970;
  assign n13972 = pi586 & ~n13343;
  assign po735 = n13389 | n13972;
  assign n13974 = pi587 & ~n13343;
  assign po736 = n13359 | n13974;
  assign n13976 = pi588 & ~n13343;
  assign po737 = n13399 | n13976;
  assign n13978 = pi589 & ~n13343;
  assign po738 = n13712 | n13978;
  assign n13980 = pi590 & ~n13343;
  assign po739 = n13566 | n13980;
  assign n13982 = pi591 & ~n13343;
  assign po740 = n12833 | n13982;
  assign n13984 = pi592 & ~n13343;
  assign po741 = n13469 | n13984;
  assign n13986 = pi593 & ~n13343;
  assign po742 = n13497 | n13986;
  assign n13988 = pi594 & ~n13343;
  assign po743 = n12928 | n13988;
  assign n13990 = pi595 & ~n13343;
  assign po744 = n13527 | n13990;
  assign n13992 = pi596 & ~n13343;
  assign po745 = n13379 | n13992;
  assign n13994 = pi597 & ~n13343;
  assign po746 = n10350 | n13994;
  assign n13996 = pi598 & ~n13343;
  assign po747 = n13502 | n13996;
  assign n13998 = pi599 & ~n13343;
  assign po748 = n13532 | n13998;
  assign n14000 = pi600 & ~n13343;
  assign po749 = n13429 | n14000;
  assign n14002 = pi601 & ~n13343;
  assign po750 = n13219 | n14002;
  assign n14004 = pi602 & ~n13343;
  assign po751 = n13434 | n14004;
  assign n14006 = pi603 & ~n13343;
  assign po752 = n13409 | n14006;
  assign n14008 = pi604 & ~n13343;
  assign po753 = n13522 | n14008;
  assign n14010 = pi605 & ~n13343;
  assign po754 = n13737 | n14010;
  assign n14012 = pi606 & ~n13343;
  assign po755 = n12978 | n14012;
  assign n14014 = pi607 & ~n13343;
  assign po756 = n12938 | n14014;
  assign n14016 = pi608 & ~n13343;
  assign po757 = n12753 | n14016;
  assign n14018 = pi609 & ~n13343;
  assign po758 = n13459 | n14018;
  assign n14020 = pi610 & ~n13343;
  assign po759 = n12748 | n14020;
  assign n14022 = pi611 & ~n13343;
  assign po760 = n13595 | n14022;
  assign n14024 = pi612 & ~n13343;
  assign po761 = n13309 | n14024;
  assign n14026 = pi613 & ~n13343;
  assign po762 = n13464 | n14026;
  assign n14028 = pi614 & ~n13343;
  assign po763 = n13670 | n14028;
  assign n14030 = pi615 & ~n13343;
  assign po764 = n13095 | n14030;
  assign n14032 = pi616 & ~n13343;
  assign po765 = n12722 | n14032;
  assign n14034 = pi617 & ~n13343;
  assign po766 = n13742 | n14034;
  assign n14036 = pi618 & ~n13343;
  assign po767 = n13707 | n14036;
  assign n14038 = pi619 & ~n13343;
  assign po768 = n13444 | n14038;
  assign n14040 = pi620 & ~n13343;
  assign po769 = n13187 | n14040;
  assign n14042 = pi621 & ~n13343;
  assign po770 = n12616 | n14042;
  assign n14044 = pi622 & ~n13343;
  assign po771 = n13482 | n14044;
  assign n14046 = pi623 & ~n13343;
  assign po772 = n13537 | n14046;
  assign n14048 = pi624 & ~n13343;
  assign po773 = n12713 | n14048;
  assign n14050 = pi625 & ~n13343;
  assign po774 = n13011 | n14050;
  assign n14052 = pi626 & ~n13343;
  assign po775 = n13394 | n14052;
  assign n14054 = pi627 & ~n13343;
  assign po776 = n12738 | n14054;
  assign n14056 = pi628 & ~n13343;
  assign po777 = n13341 | n14056;
  assign n14058 = pi629 & ~n13343;
  assign po778 = n13127 | n14058;
  assign n14060 = pi630 & ~n13343;
  assign po779 = n12743 | n14060;
  assign n14062 = pi631 & ~n13343;
  assign po780 = n12948 | n14062;
  assign n14064 = pi632 & ~n13343;
  assign po781 = n13770 | n14064;
  assign n14066 = pi633 & ~n13343;
  assign po782 = n12943 | n14066;
  assign n14068 = pi634 & ~n13343;
  assign po783 = n13404 | n14068;
  assign n14070 = pi635 & ~n13343;
  assign po784 = n13419 | n14070;
  assign n14072 = pi636 & ~n13343;
  assign po785 = n12566 | n14072;
  assign n14074 = pi637 & ~n13343;
  assign po786 = n12727 | n14074;
  assign n14076 = pi638 & ~n13343;
  assign po787 = n13369 | n14076;
  assign n14078 = pi639 & ~n13343;
  assign po788 = n13507 | n14078;
  assign n14080 = pi640 & ~n13343;
  assign po789 = n13487 | n14080;
  assign n14082 = pi641 & ~n13343;
  assign po790 = n13384 | n14082;
  assign n14084 = pi642 & ~n13343;
  assign po791 = n10388 | n14084;
  assign n14086 = pi643 & ~n13343;
  assign po792 = n13512 | n14086;
  assign n14088 = pi644 & ~n13343;
  assign po793 = n12958 | n14088;
  assign n14090 = pi645 & ~n13343;
  assign po794 = n13439 | n14090;
  assign n14092 = pi646 & ~n13343;
  assign po795 = n13723 | n14092;
  assign n14094 = pi647 & ~n13343;
  assign po796 = n13031 | n14094;
  assign n14096 = pi648 & ~n13343;
  assign po797 = n13547 | n14096;
  assign n14098 = pi649 & ~n13343;
  assign po798 = n13624 | n14098;
  assign n14100 = pi650 & ~n13343;
  assign po799 = n13364 | n14100;
  assign n14102 = pi651 & ~n13343;
  assign po800 = n12853 | n14102;
  assign n14104 = pi652 & ~n13343;
  assign po801 = n13374 | n14104;
  assign n14106 = pi653 & ~n13343;
  assign po802 = n12905 | n14106;
  assign n14108 = pi654 & ~n13343;
  assign po803 = n12758 | n14108;
  assign n14110 = pi655 & ~n13343;
  assign po804 = n13063 | n14110;
  assign n14112 = pi656 & ~n13343;
  assign po805 = n12732 | n14112;
  assign n14114 = pi657 & ~n13343;
  assign po806 = n12885 | n14114;
  assign n14116 = pi658 & ~n13343;
  assign po807 = n13477 | n14116;
  assign n14118 = pi659 & ~n13343;
  assign po808 = n13414 | n14118;
  assign n14120 = pi660 & ~n13343;
  assign po809 = n13647 | n14120;
  assign n14122 = pi661 & ~n13343;
  assign po810 = n13759 | n14122;
  assign n14124 = pi662 & ~n13343;
  assign po811 = n13699 | n14124;
  assign n14126 = pi663 & ~n13343;
  assign po812 = n12933 | n14126;
  assign n14128 = pi664 & ~n13343;
  assign po813 = n10115 | n14128;
  assign n14130 = ~n2019 & n2411;
  assign po817 = n13796 | n14130;
  assign n14132 = ~pi563 & n2465;
  assign n14133 = ~pi567 & pi568;
  assign po818 = n14132 & n14133;
  assign po130 = 1'b1;
  assign po145 = ~po814;
  assign po000 = pi564;
  assign po001 = pi266;
  assign po002 = pi303;
  assign po003 = pi312;
  assign po004 = pi270;
  assign po005 = pi326;
  assign po006 = pi297;
  assign po007 = pi256;
  assign po008 = pi308;
  assign po009 = pi264;
  assign po010 = pi323;
  assign po011 = pi282;
  assign po012 = pi319;
  assign po013 = pi327;
  assign po014 = pi283;
  assign po015 = pi329;
  assign po016 = pi331;
  assign po017 = pi400;
  assign po018 = pi386;
  assign po019 = pi407;
  assign po020 = pi404;
  assign po021 = pi355;
  assign po022 = pi358;
  assign po023 = pi360;
  assign po024 = pi363;
  assign po025 = pi306;
  assign po026 = pi258;
  assign po027 = pi262;
  assign po028 = pi340;
  assign po029 = pi309;
  assign po030 = pi263;
  assign po031 = pi311;
  assign po032 = pi313;
  assign po033 = pi374;
  assign po034 = pi343;
  assign po035 = pi317;
  assign po036 = pi346;
  assign po037 = pi378;
  assign po038 = pi380;
  assign po039 = pi381;
  assign po040 = pi382;
  assign po041 = pi299;
  assign po042 = pi271;
  assign po043 = pi273;
  assign po044 = pi274;
  assign po045 = pi275;
  assign po046 = pi325;
  assign po047 = pi278;
  assign po048 = pi279;
  assign po049 = pi408;
  assign po050 = pi383;
  assign po051 = pi406;
  assign po052 = pi405;
  assign po053 = pi384;
  assign po054 = pi402;
  assign po055 = pi398;
  assign po056 = pi385;
  assign po057 = pi330;
  assign po058 = pi286;
  assign po059 = pi285;
  assign po060 = pi287;
  assign po061 = pi253;
  assign po062 = pi301;
  assign po063 = pi302;
  assign po064 = pi255;
  assign po065 = pi353;
  assign po066 = pi354;
  assign po067 = pi356;
  assign po068 = pi357;
  assign po069 = pi401;
  assign po070 = pi359;
  assign po071 = pi361;
  assign po072 = pi399;
  assign po073 = pi307;
  assign po074 = pi304;
  assign po075 = pi305;
  assign po076 = pi341;
  assign po077 = pi257;
  assign po078 = pi259;
  assign po079 = pi260;
  assign po080 = pi261;
  assign po081 = pi366;
  assign po082 = pi367;
  assign po083 = pi395;
  assign po084 = pi368;
  assign po085 = pi371;
  assign po086 = pi369;
  assign po087 = pi370;
  assign po088 = pi372;
  assign po089 = pi373;
  assign po090 = pi392;
  assign po091 = pi314;
  assign po092 = pi315;
  assign po093 = pi316;
  assign po094 = pi318;
  assign po095 = pi320;
  assign po096 = pi321;
  assign po097 = pi376;
  assign po098 = pi377;
  assign po099 = pi345;
  assign po100 = pi379;
  assign po101 = pi342;
  assign po102 = pi351;
  assign po103 = pi362;
  assign po104 = pi344;
  assign po105 = pi310;
  assign po106 = pi265;
  assign po107 = pi267;
  assign po108 = pi268;
  assign po109 = pi276;
  assign po110 = pi328;
  assign po111 = pi284;
  assign po112 = pi254;
  assign po113 = pi352;
  assign po114 = pi403;
  assign po115 = pi397;
  assign po116 = pi364;
  assign po117 = pi365;
  assign po118 = pi393;
  assign po119 = pi391;
  assign po120 = pi375;
  assign po121 = pi322;
  assign po122 = pi324;
  assign po123 = pi269;
  assign po124 = pi272;
  assign po125 = pi300;
  assign po126 = pi277;
  assign po127 = pi280;
  assign po128 = pi281;
  assign po129 = pi671;
  assign po131 = pi670;
  assign po146 = pi012;
  assign po148 = pi013;
  assign po150 = pi014;
  assign po152 = pi015;
  assign po154 = pi016;
  assign po156 = pi017;
  assign po182 = pi042;
  assign po184 = pi043;
  assign po186 = pi044;
  assign po188 = pi045;
  assign po192 = pi048;
  assign po194 = pi049;
  assign po202 = pi056;
  assign po204 = pi057;
  assign po314 = pi166;
  assign po316 = pi167;
endmodule


