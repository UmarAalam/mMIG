//Written by the Majority Logic Package Thu Apr 30 23:14:44 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325;
assign w0 = pi00 & pi32;
assign w1 = pi64 & w0;
assign w2 = ~pi64 & ~w0;
assign w3 = ~w1 & ~w2;
assign w4 = pi00 & pi33;
assign w5 = pi01 & pi32;
assign w6 = pi65 & w5;
assign w7 = ~pi65 & ~w5;
assign w8 = ~w6 & ~w7;
assign w9 = w4 & w8;
assign w10 = ~w4 & ~w8;
assign w11 = ~w9 & ~w10;
assign w12 = w1 & w11;
assign w13 = ~w1 & ~w11;
assign w14 = ~w12 & ~w13;
assign w15 = (~w9 & ~w11) | (~w9 & w8577) | (~w11 & w8577);
assign w16 = pi01 & pi33;
assign w17 = pi00 & pi34;
assign w18 = ~w16 & ~w17;
assign w19 = pi01 & pi34;
assign w20 = w4 & w19;
assign w21 = ~w18 & ~w20;
assign w22 = pi02 & pi32;
assign w23 = pi66 & w22;
assign w24 = ~pi66 & ~w22;
assign w25 = ~w23 & ~w24;
assign w26 = w21 & w25;
assign w27 = ~w21 & ~w25;
assign w28 = ~w26 & ~w27;
assign w29 = w6 & w28;
assign w30 = ~w6 & ~w28;
assign w31 = ~w29 & ~w30;
assign w32 = ~w15 & w31;
assign w33 = w15 & ~w31;
assign w34 = ~w32 & ~w33;
assign w35 = (~w29 & ~w31) | (~w29 & w8578) | (~w31 & w8578);
assign w36 = ~w20 & ~w26;
assign w37 = pi00 & pi35;
assign w38 = w23 & w37;
assign w39 = ~w23 & ~w37;
assign w40 = ~w38 & ~w39;
assign w41 = pi03 & pi32;
assign w42 = pi67 & w41;
assign w43 = ~pi67 & ~w41;
assign w44 = ~w42 & ~w43;
assign w45 = pi02 & pi33;
assign w46 = ~w19 & ~w45;
assign w47 = pi02 & pi34;
assign w48 = w16 & w47;
assign w49 = ~w46 & ~w48;
assign w50 = w44 & ~w49;
assign w51 = ~w44 & w49;
assign w52 = ~w50 & ~w51;
assign w53 = w40 & ~w52;
assign w54 = ~w40 & w52;
assign w55 = ~w53 & ~w54;
assign w56 = ~w36 & w55;
assign w57 = w36 & ~w55;
assign w58 = ~w56 & ~w57;
assign w59 = w35 & ~w58;
assign w60 = ~w35 & w58;
assign w61 = ~w59 & ~w60;
assign w62 = ~w38 & ~w53;
assign w63 = pi00 & pi36;
assign w64 = w44 & ~w46;
assign w65 = w42 & ~w48;
assign w66 = w43 & w48;
assign w67 = ~w65 & ~w66;
assign w68 = ~w64 & w67;
assign w69 = w63 & ~w68;
assign w70 = ~w63 & w68;
assign w71 = ~w69 & ~w70;
assign w72 = pi01 & pi35;
assign w73 = ~w47 & ~w72;
assign w74 = pi02 & pi35;
assign w75 = w19 & w74;
assign w76 = ~w73 & ~w75;
assign w77 = pi03 & pi33;
assign w78 = pi04 & pi32;
assign w79 = pi68 & w78;
assign w80 = ~pi68 & ~w78;
assign w81 = ~w79 & ~w80;
assign w82 = w77 & ~w81;
assign w83 = ~w77 & w81;
assign w84 = ~w82 & ~w83;
assign w85 = w76 & ~w84;
assign w86 = ~w76 & w84;
assign w87 = ~w85 & ~w86;
assign w88 = w71 & w87;
assign w89 = ~w71 & ~w87;
assign w90 = ~w88 & ~w89;
assign w91 = w62 & ~w90;
assign w92 = ~w62 & w90;
assign w93 = ~w91 & ~w92;
assign w94 = (~w56 & ~w58) | (~w56 & w8579) | (~w58 & w8579);
assign w95 = ~w93 & w94;
assign w96 = w93 & ~w94;
assign w97 = ~w95 & ~w96;
assign w98 = ~w69 & ~w88;
assign w99 = w42 & w48;
assign w100 = pi05 & pi32;
assign w101 = pi69 & w100;
assign w102 = ~pi69 & ~w100;
assign w103 = ~w101 & ~w102;
assign w104 = pi04 & pi33;
assign w105 = pi00 & pi37;
assign w106 = ~w104 & ~w105;
assign w107 = ~w103 & w106;
assign w108 = ~w102 & w104;
assign w109 = ~w101 & ~w105;
assign w110 = w108 & w109;
assign w111 = ~w107 & ~w110;
assign w112 = ~w104 & w105;
assign w113 = w103 & ~w112;
assign w114 = pi04 & pi37;
assign w115 = w4 & w114;
assign w116 = ~w103 & ~w115;
assign w117 = ~w113 & ~w116;
assign w118 = w111 & ~w117;
assign w119 = pi01 & pi36;
assign w120 = pi03 & pi34;
assign w121 = ~w74 & ~w120;
assign w122 = pi03 & pi35;
assign w123 = w47 & w122;
assign w124 = ~w121 & ~w123;
assign w125 = w119 & ~w124;
assign w126 = ~w119 & w124;
assign w127 = ~w125 & ~w126;
assign w128 = ~w118 & w127;
assign w129 = w118 & ~w127;
assign w130 = ~w128 & ~w129;
assign w131 = w99 & w130;
assign w132 = ~w99 & ~w130;
assign w133 = ~w131 & ~w132;
assign w134 = ~w75 & ~w85;
assign w135 = ~w77 & ~w79;
assign w136 = ~w80 & ~w135;
assign w137 = ~w134 & w136;
assign w138 = w134 & ~w136;
assign w139 = ~w137 & ~w138;
assign w140 = w133 & w139;
assign w141 = ~w133 & ~w139;
assign w142 = ~w140 & ~w141;
assign w143 = w98 & ~w142;
assign w144 = ~w98 & w142;
assign w145 = ~w143 & ~w144;
assign w146 = ~w92 & w94;
assign w147 = ~w91 & ~w146;
assign w148 = w145 & ~w147;
assign w149 = ~w145 & w147;
assign w150 = ~w148 & ~w149;
assign w151 = w111 & ~w127;
assign w152 = ~w117 & ~w151;
assign w153 = ~w101 & ~w108;
assign w154 = w119 & ~w121;
assign w155 = ~w123 & ~w154;
assign w156 = ~w153 & ~w155;
assign w157 = w153 & w155;
assign w158 = ~w156 & ~w157;
assign w159 = ~w152 & w158;
assign w160 = w152 & ~w158;
assign w161 = ~w159 & ~w160;
assign w162 = w137 & w161;
assign w163 = ~w137 & ~w161;
assign w164 = ~w162 & ~w163;
assign w165 = pi06 & pi32;
assign w166 = pi70 & w165;
assign w167 = ~pi70 & ~w165;
assign w168 = ~w166 & ~w167;
assign w169 = pi05 & pi33;
assign w170 = pi04 & pi34;
assign w171 = ~w169 & ~w170;
assign w172 = pi05 & pi34;
assign w173 = w104 & w172;
assign w174 = ~w171 & ~w173;
assign w175 = w122 & ~w174;
assign w176 = ~w122 & w174;
assign w177 = ~w175 & ~w176;
assign w178 = ~w168 & w177;
assign w179 = w168 & ~w177;
assign w180 = ~w178 & ~w179;
assign w181 = pi00 & pi38;
assign w182 = pi01 & pi37;
assign w183 = pi02 & pi36;
assign w184 = ~w182 & ~w183;
assign w185 = pi02 & pi37;
assign w186 = w119 & w185;
assign w187 = ~w184 & ~w186;
assign w188 = w181 & ~w187;
assign w189 = ~w181 & w187;
assign w190 = ~w188 & ~w189;
assign w191 = w180 & w190;
assign w192 = ~w180 & ~w190;
assign w193 = ~w191 & ~w192;
assign w194 = w164 & ~w193;
assign w195 = ~w164 & w193;
assign w196 = ~w194 & ~w195;
assign w197 = ~w131 & ~w140;
assign w198 = ~w196 & w197;
assign w199 = w196 & ~w197;
assign w200 = ~w198 & ~w199;
assign w201 = ~w144 & ~w147;
assign w202 = ~w143 & ~w201;
assign w203 = ~w200 & w202;
assign w204 = w200 & ~w202;
assign w205 = ~w203 & ~w204;
assign w206 = ~w198 & ~w204;
assign w207 = (~w162 & ~w164) | (~w162 & w8665) | (~w164 & w8665);
assign w208 = w181 & ~w184;
assign w209 = ~w186 & ~w208;
assign w210 = w122 & ~w171;
assign w211 = ~w173 & ~w210;
assign w212 = ~w209 & ~w211;
assign w213 = w209 & w211;
assign w214 = ~w212 & ~w213;
assign w215 = (~w178 & ~w180) | (~w178 & w8666) | (~w180 & w8666);
assign w216 = w214 & w215;
assign w217 = ~w214 & ~w215;
assign w218 = ~w216 & ~w217;
assign w219 = (~w156 & w152) | (~w156 & w8667) | (w152 & w8667);
assign w220 = pi07 & pi32;
assign w221 = pi71 & w220;
assign w222 = ~pi71 & ~w220;
assign w223 = ~w221 & ~w222;
assign w224 = pi06 & pi33;
assign w225 = ~w172 & ~w224;
assign w226 = pi06 & pi34;
assign w227 = w169 & w226;
assign w228 = ~w225 & ~w227;
assign w229 = w223 & ~w228;
assign w230 = ~w223 & w228;
assign w231 = ~w229 & ~w230;
assign w232 = pi00 & pi39;
assign w233 = pi01 & pi38;
assign w234 = ~w232 & ~w233;
assign w235 = pi01 & pi39;
assign w236 = w181 & w235;
assign w237 = ~w234 & ~w236;
assign w238 = w166 & ~w237;
assign w239 = ~w166 & w237;
assign w240 = ~w238 & ~w239;
assign w241 = w231 & w240;
assign w242 = ~w231 & ~w240;
assign w243 = ~w241 & ~w242;
assign w244 = pi03 & pi36;
assign w245 = pi04 & pi35;
assign w246 = ~w244 & ~w245;
assign w247 = pi04 & pi36;
assign w248 = w122 & w247;
assign w249 = ~w246 & ~w248;
assign w250 = w185 & ~w249;
assign w251 = ~w185 & w249;
assign w252 = ~w250 & ~w251;
assign w253 = w243 & ~w252;
assign w254 = ~w243 & w252;
assign w255 = ~w253 & ~w254;
assign w256 = ~w219 & w255;
assign w257 = w219 & ~w255;
assign w258 = ~w256 & ~w257;
assign w259 = w218 & ~w258;
assign w260 = ~w218 & w258;
assign w261 = ~w259 & ~w260;
assign w262 = ~w207 & ~w261;
assign w263 = w207 & w261;
assign w264 = ~w262 & ~w263;
assign w265 = w206 & w264;
assign w266 = ~w206 & ~w264;
assign w267 = ~w265 & ~w266;
assign w268 = ~w198 & ~w263;
assign w269 = (~w262 & w204) | (~w262 & w8580) | (w204 & w8580);
assign w270 = ~w212 & ~w216;
assign w271 = pi05 & pi35;
assign w272 = ~w226 & ~w271;
assign w273 = pi06 & pi35;
assign w274 = w172 & w273;
assign w275 = ~w272 & ~w274;
assign w276 = pi07 & pi33;
assign w277 = pi08 & pi32;
assign w278 = pi72 & w277;
assign w279 = ~pi72 & ~w277;
assign w280 = ~w278 & ~w279;
assign w281 = w276 & w280;
assign w282 = ~w276 & ~w280;
assign w283 = ~w281 & ~w282;
assign w284 = w275 & w283;
assign w285 = ~w275 & ~w283;
assign w286 = ~w284 & ~w285;
assign w287 = pi02 & pi38;
assign w288 = pi03 & pi37;
assign w289 = ~w247 & ~w288;
assign w290 = w114 & w244;
assign w291 = ~w289 & ~w290;
assign w292 = w287 & ~w291;
assign w293 = ~w287 & w291;
assign w294 = ~w292 & ~w293;
assign w295 = ~w286 & w294;
assign w296 = w286 & ~w294;
assign w297 = ~w295 & ~w296;
assign w298 = pi00 & pi40;
assign w299 = ~w235 & ~w298;
assign w300 = pi01 & pi40;
assign w301 = w232 & w300;
assign w302 = ~w299 & ~w301;
assign w303 = w221 & w227;
assign w304 = ~w221 & ~w227;
assign w305 = ~w303 & ~w304;
assign w306 = w223 & ~w225;
assign w307 = ~w305 & ~w306;
assign w308 = w302 & ~w307;
assign w309 = ~w302 & w307;
assign w310 = ~w308 & ~w309;
assign w311 = w297 & ~w310;
assign w312 = ~w297 & w310;
assign w313 = ~w311 & ~w312;
assign w314 = (~w242 & ~w243) | (~w242 & w8668) | (~w243 & w8668);
assign w315 = w166 & ~w234;
assign w316 = ~w236 & ~w315;
assign w317 = w185 & ~w246;
assign w318 = ~w248 & ~w317;
assign w319 = ~w316 & ~w318;
assign w320 = w316 & w318;
assign w321 = ~w319 & ~w320;
assign w322 = ~w314 & w321;
assign w323 = w314 & ~w321;
assign w324 = ~w322 & ~w323;
assign w325 = w313 & ~w324;
assign w326 = ~w313 & w324;
assign w327 = ~w325 & ~w326;
assign w328 = w270 & ~w327;
assign w329 = ~w270 & w327;
assign w330 = ~w328 & ~w329;
assign w331 = ~w257 & ~w260;
assign w332 = w330 & w331;
assign w333 = ~w330 & ~w331;
assign w334 = ~w332 & ~w333;
assign w335 = ~w269 & w334;
assign w336 = w269 & ~w334;
assign w337 = ~w335 & ~w336;
assign w338 = pi00 & pi41;
assign w339 = w303 & w338;
assign w340 = ~w303 & ~w338;
assign w341 = ~w339 & ~w340;
assign w342 = ~w278 & ~w281;
assign w343 = (~w274 & ~w283) | (~w274 & w8581) | (~w283 & w8581);
assign w344 = ~w342 & ~w343;
assign w345 = w342 & w343;
assign w346 = ~w344 & ~w345;
assign w347 = w341 & w346;
assign w348 = ~w341 & ~w346;
assign w349 = ~w347 & ~w348;
assign w350 = pi03 & pi38;
assign w351 = pi02 & pi39;
assign w352 = ~w350 & ~w351;
assign w353 = pi03 & pi39;
assign w354 = w287 & w353;
assign w355 = ~w352 & ~w354;
assign w356 = w300 & ~w355;
assign w357 = ~w300 & w355;
assign w358 = ~w356 & ~w357;
assign w359 = pi08 & pi33;
assign w360 = pi09 & pi32;
assign w361 = pi73 & w360;
assign w362 = ~pi73 & ~w360;
assign w363 = ~w361 & ~w362;
assign w364 = w359 & w363;
assign w365 = ~w359 & ~w363;
assign w366 = ~w364 & ~w365;
assign w367 = ~w114 & ~w366;
assign w368 = w114 & w366;
assign w369 = ~w367 & ~w368;
assign w370 = pi05 & pi36;
assign w371 = pi07 & pi34;
assign w372 = ~w273 & ~w371;
assign w373 = pi07 & pi35;
assign w374 = w226 & w373;
assign w375 = ~w372 & ~w374;
assign w376 = w370 & ~w375;
assign w377 = ~w370 & w375;
assign w378 = ~w376 & ~w377;
assign w379 = w369 & ~w378;
assign w380 = ~w369 & w378;
assign w381 = ~w379 & ~w380;
assign w382 = ~w358 & w381;
assign w383 = w358 & ~w381;
assign w384 = ~w382 & ~w383;
assign w385 = w349 & w384;
assign w386 = ~w349 & ~w384;
assign w387 = ~w385 & ~w386;
assign w388 = ~w319 & ~w322;
assign w389 = (~w295 & ~w297) | (~w295 & w8582) | (~w297 & w8582);
assign w390 = ~w301 & ~w308;
assign w391 = w287 & ~w289;
assign w392 = ~w290 & ~w391;
assign w393 = ~w390 & ~w392;
assign w394 = w390 & w392;
assign w395 = ~w393 & ~w394;
assign w396 = w389 & w395;
assign w397 = ~w389 & ~w395;
assign w398 = ~w396 & ~w397;
assign w399 = ~w388 & w398;
assign w400 = w388 & ~w398;
assign w401 = ~w399 & ~w400;
assign w402 = w387 & w401;
assign w403 = ~w387 & ~w401;
assign w404 = ~w402 & ~w403;
assign w405 = ~w326 & ~w329;
assign w406 = ~w404 & w405;
assign w407 = w404 & ~w405;
assign w408 = ~w406 & ~w407;
assign w409 = ~w332 & ~w335;
assign w410 = w408 & w409;
assign w411 = ~w408 & ~w409;
assign w412 = ~w410 & ~w411;
assign w413 = ~w332 & ~w407;
assign w414 = ~w335 & w413;
assign w415 = ~w406 & ~w414;
assign w416 = ~w399 & ~w402;
assign w417 = ~w393 & ~w396;
assign w418 = (~w382 & ~w384) | (~w382 & w8583) | (~w384 & w8583);
assign w419 = (~w339 & ~w346) | (~w339 & w8669) | (~w346 & w8669);
assign w420 = w300 & ~w352;
assign w421 = ~w354 & ~w420;
assign w422 = ~w419 & ~w421;
assign w423 = w419 & w421;
assign w424 = ~w422 & ~w423;
assign w425 = ~w418 & w424;
assign w426 = w418 & ~w424;
assign w427 = ~w425 & ~w426;
assign w428 = ~w417 & w427;
assign w429 = w417 & ~w427;
assign w430 = ~w428 & ~w429;
assign w431 = pi04 & pi38;
assign w432 = ~w353 & ~w431;
assign w433 = pi04 & pi39;
assign w434 = w350 & w433;
assign w435 = ~w432 & ~w434;
assign w436 = pi00 & pi42;
assign w437 = pi01 & pi41;
assign w438 = pi02 & pi40;
assign w439 = ~w437 & ~w438;
assign w440 = pi02 & pi41;
assign w441 = w300 & w440;
assign w442 = ~w439 & ~w441;
assign w443 = w436 & ~w442;
assign w444 = ~w436 & w442;
assign w445 = ~w443 & ~w444;
assign w446 = w435 & ~w445;
assign w447 = ~w435 & w445;
assign w448 = ~w446 & ~w447;
assign w449 = pi05 & pi37;
assign w450 = pi09 & pi33;
assign w451 = pi10 & pi32;
assign w452 = pi74 & w451;
assign w453 = ~pi74 & ~w451;
assign w454 = ~w452 & ~w453;
assign w455 = w450 & w454;
assign w456 = ~w450 & ~w454;
assign w457 = ~w455 & ~w456;
assign w458 = w449 & w457;
assign w459 = ~w449 & ~w457;
assign w460 = ~w458 & ~w459;
assign w461 = pi06 & pi36;
assign w462 = pi08 & pi34;
assign w463 = ~w373 & ~w462;
assign w464 = pi08 & pi35;
assign w465 = w371 & w464;
assign w466 = ~w463 & ~w465;
assign w467 = w461 & ~w466;
assign w468 = ~w461 & w466;
assign w469 = ~w467 & ~w468;
assign w470 = w460 & ~w469;
assign w471 = ~w460 & w469;
assign w472 = ~w470 & ~w471;
assign w473 = (~w361 & ~w363) | (~w361 & w8670) | (~w363 & w8670);
assign w474 = w370 & ~w372;
assign w475 = ~w374 & ~w474;
assign w476 = ~w473 & ~w475;
assign w477 = w473 & w475;
assign w478 = ~w476 & ~w477;
assign w479 = ~w368 & w378;
assign w480 = ~w367 & ~w479;
assign w481 = ~w479 & w8671;
assign w482 = (~w478 & w479) | (~w478 & w8672) | (w479 & w8672);
assign w483 = ~w481 & ~w482;
assign w484 = w344 & w483;
assign w485 = ~w344 & ~w483;
assign w486 = ~w484 & ~w485;
assign w487 = w472 & w486;
assign w488 = ~w472 & ~w486;
assign w489 = ~w487 & ~w488;
assign w490 = w448 & w489;
assign w491 = ~w448 & ~w489;
assign w492 = ~w490 & ~w491;
assign w493 = w430 & w492;
assign w494 = ~w430 & ~w492;
assign w495 = ~w493 & ~w494;
assign w496 = ~w416 & w495;
assign w497 = w416 & ~w495;
assign w498 = ~w496 & ~w497;
assign w499 = ~w415 & ~w498;
assign w500 = w415 & w498;
assign w501 = ~w499 & ~w500;
assign w502 = ~w496 & ~w500;
assign w503 = ~w428 & ~w493;
assign w504 = ~w422 & ~w425;
assign w505 = pi06 & pi37;
assign w506 = pi10 & pi33;
assign w507 = pi11 & pi32;
assign w508 = pi75 & w507;
assign w509 = ~pi75 & ~w507;
assign w510 = ~w508 & ~w509;
assign w511 = w506 & w510;
assign w512 = ~w506 & ~w510;
assign w513 = ~w511 & ~w512;
assign w514 = w505 & w513;
assign w515 = ~w505 & ~w513;
assign w516 = ~w514 & ~w515;
assign w517 = pi07 & pi36;
assign w518 = pi09 & pi34;
assign w519 = ~w464 & ~w518;
assign w520 = pi09 & pi35;
assign w521 = w462 & w520;
assign w522 = ~w519 & ~w521;
assign w523 = w517 & ~w522;
assign w524 = ~w517 & w522;
assign w525 = ~w523 & ~w524;
assign w526 = w516 & ~w525;
assign w527 = ~w516 & w525;
assign w528 = ~w526 & ~w527;
assign w529 = (~w458 & ~w460) | (~w458 & w8673) | (~w460 & w8673);
assign w530 = (~w452 & ~w454) | (~w452 & w8674) | (~w454 & w8674);
assign w531 = w461 & ~w463;
assign w532 = ~w465 & ~w531;
assign w533 = ~w530 & ~w532;
assign w534 = w530 & w532;
assign w535 = ~w533 & ~w534;
assign w536 = ~w434 & w535;
assign w537 = w434 & ~w535;
assign w538 = ~w536 & ~w537;
assign w539 = w529 & ~w538;
assign w540 = ~w529 & w538;
assign w541 = ~w539 & ~w540;
assign w542 = w528 & ~w541;
assign w543 = ~w528 & w541;
assign w544 = ~w542 & ~w543;
assign w545 = pi00 & pi43;
assign w546 = pi01 & pi42;
assign w547 = ~w545 & ~w546;
assign w548 = pi01 & pi43;
assign w549 = w436 & w548;
assign w550 = ~w547 & ~w549;
assign w551 = (w480 & w8675) | (w480 & w8676) | (w8675 & w8676);
assign w552 = ~w550 & w9294;
assign w553 = ~w551 & ~w552;
assign w554 = pi03 & pi40;
assign w555 = pi05 & pi38;
assign w556 = ~w433 & ~w555;
assign w557 = pi05 & pi39;
assign w558 = w431 & w557;
assign w559 = ~w556 & ~w558;
assign w560 = w554 & w559;
assign w561 = ~w554 & ~w559;
assign w562 = ~w560 & ~w561;
assign w563 = w440 & w562;
assign w564 = ~w440 & ~w562;
assign w565 = ~w563 & ~w564;
assign w566 = w553 & w565;
assign w567 = ~w553 & ~w565;
assign w568 = ~w566 & ~w567;
assign w569 = w544 & w568;
assign w570 = ~w544 & ~w568;
assign w571 = ~w569 & ~w570;
assign w572 = w504 & ~w571;
assign w573 = ~w504 & w571;
assign w574 = ~w572 & ~w573;
assign w575 = (~w446 & ~w489) | (~w446 & w8585) | (~w489 & w8585);
assign w576 = (~w484 & ~w486) | (~w484 & w8586) | (~w486 & w8586);
assign w577 = w436 & ~w439;
assign w578 = ~w441 & ~w577;
assign w579 = ~w576 & ~w578;
assign w580 = w576 & w578;
assign w581 = ~w579 & ~w580;
assign w582 = ~w575 & w581;
assign w583 = w575 & ~w581;
assign w584 = ~w582 & ~w583;
assign w585 = w574 & ~w584;
assign w586 = ~w574 & w584;
assign w587 = ~w585 & ~w586;
assign w588 = ~w503 & ~w587;
assign w589 = w503 & w587;
assign w590 = ~w588 & ~w589;
assign w591 = w502 & w590;
assign w592 = ~w502 & ~w590;
assign w593 = ~w591 & ~w592;
assign w594 = ~w496 & ~w588;
assign w595 = (~w589 & w500) | (~w589 & w8677) | (w500 & w8677);
assign w596 = ~w579 & ~w582;
assign w597 = pi07 & pi37;
assign w598 = pi11 & pi33;
assign w599 = pi12 & pi32;
assign w600 = pi76 & w599;
assign w601 = ~pi76 & ~w599;
assign w602 = ~w600 & ~w601;
assign w603 = w598 & w602;
assign w604 = ~w598 & ~w602;
assign w605 = ~w603 & ~w604;
assign w606 = w597 & w605;
assign w607 = ~w597 & ~w605;
assign w608 = ~w606 & ~w607;
assign w609 = pi08 & pi36;
assign w610 = pi10 & pi34;
assign w611 = ~w520 & ~w610;
assign w612 = pi10 & pi35;
assign w613 = w518 & w612;
assign w614 = ~w611 & ~w613;
assign w615 = w609 & ~w614;
assign w616 = ~w609 & w614;
assign w617 = ~w615 & ~w616;
assign w618 = w608 & ~w617;
assign w619 = ~w608 & w617;
assign w620 = ~w618 & ~w619;
assign w621 = (~w514 & ~w516) | (~w514 & w8678) | (~w516 & w8678);
assign w622 = w562 & w8587;
assign w623 = w440 & w554;
assign w624 = w558 & ~w623;
assign w625 = ~w560 & ~w624;
assign w626 = ~w622 & w625;
assign w627 = (~w508 & ~w510) | (~w508 & w8679) | (~w510 & w8679);
assign w628 = w517 & ~w519;
assign w629 = ~w521 & ~w628;
assign w630 = ~w627 & ~w629;
assign w631 = w627 & w629;
assign w632 = ~w630 & ~w631;
assign w633 = w626 & ~w632;
assign w634 = ~w626 & w632;
assign w635 = ~w633 & ~w634;
assign w636 = w621 & ~w635;
assign w637 = ~w621 & w635;
assign w638 = ~w636 & ~w637;
assign w639 = w620 & w638;
assign w640 = ~w620 & ~w638;
assign w641 = ~w639 & ~w640;
assign w642 = ~w529 & ~w534;
assign w643 = ~w533 & ~w642;
assign w644 = pi00 & pi44;
assign w645 = ~w548 & ~w644;
assign w646 = pi01 & pi44;
assign w647 = w545 & w646;
assign w648 = ~w645 & ~w647;
assign w649 = pi03 & pi41;
assign w650 = pi02 & pi42;
assign w651 = ~w649 & ~w650;
assign w652 = pi03 & pi42;
assign w653 = w440 & w652;
assign w654 = ~w651 & ~w653;
assign w655 = pi04 & pi40;
assign w656 = pi06 & pi38;
assign w657 = ~w557 & ~w656;
assign w658 = pi06 & pi39;
assign w659 = w555 & w658;
assign w660 = ~w657 & ~w659;
assign w661 = w655 & ~w660;
assign w662 = ~w655 & w660;
assign w663 = ~w661 & ~w662;
assign w664 = w654 & ~w663;
assign w665 = ~w654 & w663;
assign w666 = ~w664 & ~w665;
assign w667 = w648 & ~w666;
assign w668 = ~w648 & w666;
assign w669 = ~w667 & ~w668;
assign w670 = w643 & w669;
assign w671 = ~w643 & ~w669;
assign w672 = ~w670 & ~w671;
assign w673 = w641 & w672;
assign w674 = ~w641 & ~w672;
assign w675 = ~w673 & ~w674;
assign w676 = ~w596 & w675;
assign w677 = w596 & ~w675;
assign w678 = ~w676 & ~w677;
assign w679 = ~w566 & ~w569;
assign w680 = ~w549 & ~w551;
assign w681 = w434 & w541;
assign w682 = ~w542 & ~w681;
assign w683 = ~w680 & ~w682;
assign w684 = w680 & w682;
assign w685 = ~w683 & ~w684;
assign w686 = w679 & ~w685;
assign w687 = ~w679 & w685;
assign w688 = ~w686 & ~w687;
assign w689 = w678 & ~w688;
assign w690 = ~w678 & w688;
assign w691 = ~w689 & ~w690;
assign w692 = ~w572 & ~w585;
assign w693 = w691 & ~w692;
assign w694 = ~w691 & w692;
assign w695 = ~w693 & ~w694;
assign w696 = w595 & ~w695;
assign w697 = ~w595 & w695;
assign w698 = ~w696 & ~w697;
assign w699 = ~w595 & ~w694;
assign w700 = ~w693 & ~w699;
assign w701 = ~w677 & ~w689;
assign w702 = pi05 & pi40;
assign w703 = pi07 & pi38;
assign w704 = ~w658 & ~w703;
assign w705 = pi07 & pi39;
assign w706 = w656 & w705;
assign w707 = ~w704 & ~w706;
assign w708 = w702 & ~w707;
assign w709 = ~w702 & w707;
assign w710 = ~w708 & ~w709;
assign w711 = w646 & ~w710;
assign w712 = ~w646 & w710;
assign w713 = ~w711 & ~w712;
assign w714 = pi02 & pi43;
assign w715 = pi04 & pi41;
assign w716 = ~w652 & ~w715;
assign w717 = pi04 & pi42;
assign w718 = w649 & w717;
assign w719 = ~w716 & ~w718;
assign w720 = w714 & ~w719;
assign w721 = ~w714 & w719;
assign w722 = ~w720 & ~w721;
assign w723 = w713 & ~w722;
assign w724 = ~w713 & w722;
assign w725 = ~w723 & ~w724;
assign w726 = pi00 & pi45;
assign w727 = w558 & w623;
assign w728 = w726 & w727;
assign w729 = ~w726 & ~w727;
assign w730 = ~w728 & ~w729;
assign w731 = (~w630 & w621) | (~w630 & w9234) | (w621 & w9234);
assign w732 = ~w730 & w731;
assign w733 = w730 & ~w731;
assign w734 = ~w732 & ~w733;
assign w735 = w725 & w734;
assign w736 = ~w725 & ~w734;
assign w737 = ~w735 & ~w736;
assign w738 = (~w606 & ~w608) | (~w606 & w8680) | (~w608 & w8680);
assign w739 = ~w600 & ~w603;
assign w740 = w609 & ~w611;
assign w741 = ~w613 & ~w740;
assign w742 = ~w739 & ~w741;
assign w743 = w739 & w741;
assign w744 = ~w742 & ~w743;
assign w745 = ~w738 & w744;
assign w746 = w738 & ~w744;
assign w747 = ~w745 & ~w746;
assign w748 = pi08 & pi37;
assign w749 = pi12 & pi33;
assign w750 = pi13 & pi32;
assign w751 = pi77 & w750;
assign w752 = ~pi77 & ~w750;
assign w753 = ~w751 & ~w752;
assign w754 = w749 & w753;
assign w755 = ~w749 & ~w753;
assign w756 = ~w754 & ~w755;
assign w757 = w748 & w756;
assign w758 = ~w748 & ~w756;
assign w759 = ~w757 & ~w758;
assign w760 = pi09 & pi36;
assign w761 = pi11 & pi34;
assign w762 = ~w612 & ~w761;
assign w763 = pi11 & pi35;
assign w764 = w610 & w763;
assign w765 = ~w762 & ~w764;
assign w766 = w760 & ~w765;
assign w767 = ~w760 & w765;
assign w768 = ~w766 & ~w767;
assign w769 = w759 & ~w768;
assign w770 = ~w759 & w768;
assign w771 = ~w769 & ~w770;
assign w772 = (~w653 & w663) | (~w653 & w9235) | (w663 & w9235);
assign w773 = w655 & ~w657;
assign w774 = ~w659 & ~w773;
assign w775 = ~w772 & ~w774;
assign w776 = w772 & w774;
assign w777 = ~w775 & ~w776;
assign w778 = ~w771 & ~w777;
assign w779 = w771 & w777;
assign w780 = ~w778 & ~w779;
assign w781 = w747 & ~w780;
assign w782 = ~w747 & w780;
assign w783 = ~w781 & ~w782;
assign w784 = w737 & ~w783;
assign w785 = ~w737 & w783;
assign w786 = ~w784 & ~w785;
assign w787 = w666 & ~w672;
assign w788 = ~w673 & ~w787;
assign w789 = ~w626 & ~w638;
assign w790 = ~w639 & ~w789;
assign w791 = ~w643 & ~w645;
assign w792 = ~w647 & ~w791;
assign w793 = ~w790 & ~w792;
assign w794 = w790 & w792;
assign w795 = ~w793 & ~w794;
assign w796 = ~w788 & w795;
assign w797 = w788 & ~w795;
assign w798 = ~w796 & ~w797;
assign w799 = ~w683 & ~w687;
assign w800 = ~w798 & w799;
assign w801 = w798 & ~w799;
assign w802 = ~w800 & ~w801;
assign w803 = w786 & ~w802;
assign w804 = ~w786 & w802;
assign w805 = ~w803 & ~w804;
assign w806 = w701 & ~w805;
assign w807 = ~w701 & w805;
assign w808 = ~w806 & ~w807;
assign w809 = ~w700 & ~w808;
assign w810 = ~w693 & w808;
assign w811 = ~w699 & w810;
assign w812 = ~w809 & ~w811;
assign w813 = ~w806 & ~w811;
assign w814 = pi08 & pi38;
assign w815 = pi09 & pi37;
assign w816 = pi10 & pi36;
assign w817 = ~w815 & ~w816;
assign w818 = pi10 & pi37;
assign w819 = w760 & w818;
assign w820 = ~w817 & ~w819;
assign w821 = w814 & ~w820;
assign w822 = ~w814 & w820;
assign w823 = ~w821 & ~w822;
assign w824 = pi12 & pi34;
assign w825 = pi13 & pi33;
assign w826 = ~w824 & ~w825;
assign w827 = pi13 & pi34;
assign w828 = w749 & w827;
assign w829 = ~w826 & ~w828;
assign w830 = ~w705 & w763;
assign w831 = w705 & ~w763;
assign w832 = ~w830 & ~w831;
assign w833 = w829 & w832;
assign w834 = ~w829 & ~w832;
assign w835 = ~w833 & ~w834;
assign w836 = ~w823 & ~w835;
assign w837 = w823 & w835;
assign w838 = ~w836 & ~w837;
assign w839 = (~w757 & ~w759) | (~w757 & w8588) | (~w759 & w8588);
assign w840 = (~w751 & ~w753) | (~w751 & w9236) | (~w753 & w9236);
assign w841 = w760 & ~w762;
assign w842 = ~w764 & ~w841;
assign w843 = ~w840 & ~w842;
assign w844 = w840 & w842;
assign w845 = ~w843 & ~w844;
assign w846 = ~w839 & w845;
assign w847 = w839 & ~w845;
assign w848 = ~w846 & ~w847;
assign w849 = (~w711 & ~w713) | (~w711 & w8681) | (~w713 & w8681);
assign w850 = w714 & ~w716;
assign w851 = ~w718 & ~w850;
assign w852 = w702 & ~w704;
assign w853 = ~w706 & ~w852;
assign w854 = ~w851 & ~w853;
assign w855 = w851 & w853;
assign w856 = ~w854 & ~w855;
assign w857 = w849 & ~w856;
assign w858 = ~w849 & w856;
assign w859 = ~w857 & ~w858;
assign w860 = w848 & w859;
assign w861 = ~w848 & ~w859;
assign w862 = ~w860 & ~w861;
assign w863 = w838 & w862;
assign w864 = ~w838 & ~w862;
assign w865 = ~w863 & ~w864;
assign w866 = pi00 & pi46;
assign w867 = pi05 & pi41;
assign w868 = pi06 & pi40;
assign w869 = ~w867 & ~w868;
assign w870 = pi06 & pi41;
assign w871 = w702 & w870;
assign w872 = ~w869 & ~w871;
assign w873 = w717 & ~w872;
assign w874 = ~w717 & w872;
assign w875 = ~w873 & ~w874;
assign w876 = w866 & ~w875;
assign w877 = ~w866 & w875;
assign w878 = ~w876 & ~w877;
assign w879 = pi01 & pi45;
assign w880 = pi02 & pi44;
assign w881 = pi03 & pi43;
assign w882 = ~w880 & ~w881;
assign w883 = pi03 & pi44;
assign w884 = w714 & w883;
assign w885 = ~w882 & ~w884;
assign w886 = w879 & ~w885;
assign w887 = ~w879 & w885;
assign w888 = ~w886 & ~w887;
assign w889 = w878 & ~w888;
assign w890 = ~w878 & w888;
assign w891 = ~w889 & ~w890;
assign w892 = (~w742 & w738) | (~w742 & w9237) | (w738 & w9237);
assign w893 = pi14 & pi32;
assign w894 = pi78 & w893;
assign w895 = ~pi78 & ~w893;
assign w896 = ~w894 & ~w895;
assign w897 = ~w775 & ~w896;
assign w898 = w775 & w896;
assign w899 = ~w897 & ~w898;
assign w900 = w892 & ~w899;
assign w901 = ~w892 & w899;
assign w902 = ~w900 & ~w901;
assign w903 = w891 & w902;
assign w904 = ~w891 & ~w902;
assign w905 = ~w903 & ~w904;
assign w906 = w865 & w905;
assign w907 = ~w865 & ~w905;
assign w908 = ~w906 & ~w907;
assign w909 = ~w793 & ~w796;
assign w910 = ~w735 & ~w784;
assign w911 = ~w778 & ~w782;
assign w912 = ~w728 & ~w733;
assign w913 = w911 & ~w912;
assign w914 = ~w911 & w912;
assign w915 = ~w913 & ~w914;
assign w916 = ~w910 & w915;
assign w917 = w910 & ~w915;
assign w918 = ~w916 & ~w917;
assign w919 = ~w909 & w918;
assign w920 = w909 & ~w918;
assign w921 = ~w919 & ~w920;
assign w922 = w908 & w921;
assign w923 = ~w908 & ~w921;
assign w924 = ~w922 & ~w923;
assign w925 = ~w800 & ~w804;
assign w926 = w924 & w925;
assign w927 = ~w924 & ~w925;
assign w928 = ~w926 & ~w927;
assign w929 = w813 & ~w928;
assign w930 = ~w813 & w928;
assign w931 = ~w929 & ~w930;
assign w932 = ~w806 & ~w926;
assign w933 = (~w927 & w811) | (~w927 & w8682) | (w811 & w8682);
assign w934 = ~w919 & ~w922;
assign w935 = ~w913 & ~w916;
assign w936 = (~w903 & ~w865) | (~w903 & w9238) | (~w865 & w9238);
assign w937 = (~w860 & ~w862) | (~w860 & w9239) | (~w862 & w9239);
assign w938 = ~w898 & ~w901;
assign w939 = ~w937 & ~w938;
assign w940 = w937 & w938;
assign w941 = ~w939 & ~w940;
assign w942 = ~w936 & w941;
assign w943 = w936 & ~w941;
assign w944 = ~w942 & ~w943;
assign w945 = w935 & ~w944;
assign w946 = ~w935 & w944;
assign w947 = ~w945 & ~w946;
assign w948 = pi04 & pi43;
assign w949 = pi05 & pi42;
assign w950 = ~w948 & ~w949;
assign w951 = pi05 & pi43;
assign w952 = w717 & w951;
assign w953 = ~w950 & ~w952;
assign w954 = w883 & ~w953;
assign w955 = ~w883 & w953;
assign w956 = ~w954 & ~w955;
assign w957 = w894 & ~w956;
assign w958 = ~w894 & w956;
assign w959 = ~w957 & ~w958;
assign w960 = pi00 & pi47;
assign w961 = pi01 & pi46;
assign w962 = pi02 & pi45;
assign w963 = ~w961 & ~w962;
assign w964 = pi02 & pi46;
assign w965 = w879 & w964;
assign w966 = ~w963 & ~w965;
assign w967 = w960 & ~w966;
assign w968 = ~w960 & w966;
assign w969 = ~w967 & ~w968;
assign w970 = w959 & ~w969;
assign w971 = ~w959 & w969;
assign w972 = ~w970 & ~w971;
assign w973 = pi15 & pi32;
assign w974 = ~pi79 & ~w973;
assign w975 = pi79 & w973;
assign w976 = ~w974 & ~w975;
assign w977 = pi14 & pi33;
assign w978 = ~w827 & ~w977;
assign w979 = w827 & w977;
assign w980 = ~w978 & ~w979;
assign w981 = w976 & ~w980;
assign w982 = ~w976 & w980;
assign w983 = ~w981 & ~w982;
assign w984 = ~w844 & w983;
assign w985 = (w984 & ~w839) | (w984 & w8683) | (~w839 & w8683);
assign w986 = ~w843 & ~w983;
assign w987 = (w986 & w839) | (w986 & w8684) | (w839 & w8684);
assign w988 = ~w985 & ~w987;
assign w989 = (~w854 & w849) | (~w854 & w9240) | (w849 & w9240);
assign w990 = ~w988 & w989;
assign w991 = w988 & ~w989;
assign w992 = ~w990 & ~w991;
assign w993 = w972 & ~w992;
assign w994 = ~w972 & w992;
assign w995 = ~w993 & ~w994;
assign w996 = pi11 & pi36;
assign w997 = pi12 & pi35;
assign w998 = ~w996 & ~w997;
assign w999 = pi12 & pi36;
assign w1000 = w763 & w999;
assign w1001 = ~w998 & ~w1000;
assign w1002 = w818 & ~w1001;
assign w1003 = ~w818 & w1001;
assign w1004 = ~w1002 & ~w1003;
assign w1005 = w870 & ~w1004;
assign w1006 = ~w870 & w1004;
assign w1007 = ~w1005 & ~w1006;
assign w1008 = pi07 & pi40;
assign w1009 = pi08 & pi39;
assign w1010 = pi09 & pi38;
assign w1011 = ~w1009 & ~w1010;
assign w1012 = pi09 & pi39;
assign w1013 = w814 & w1012;
assign w1014 = ~w1011 & ~w1013;
assign w1015 = w1008 & ~w1014;
assign w1016 = ~w1008 & w1014;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = w1007 & ~w1017;
assign w1019 = ~w1007 & w1017;
assign w1020 = ~w1018 & ~w1019;
assign w1021 = (~w876 & ~w878) | (~w876 & w8685) | (~w878 & w8685);
assign w1022 = w879 & ~w882;
assign w1023 = ~w884 & ~w1022;
assign w1024 = w717 & ~w869;
assign w1025 = ~w871 & ~w1024;
assign w1026 = ~w1023 & ~w1025;
assign w1027 = w1023 & w1025;
assign w1028 = ~w1026 & ~w1027;
assign w1029 = ~w1021 & w1028;
assign w1030 = w1021 & ~w1028;
assign w1031 = ~w1029 & ~w1030;
assign w1032 = w763 & ~w826;
assign w1033 = ~w828 & ~w1032;
assign w1034 = w814 & ~w817;
assign w1035 = ~w819 & ~w1034;
assign w1036 = ~w1033 & ~w1035;
assign w1037 = w1033 & w1035;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = w705 & w835;
assign w1040 = ~w836 & ~w1039;
assign w1041 = w1038 & ~w1040;
assign w1042 = ~w1038 & w1040;
assign w1043 = ~w1041 & ~w1042;
assign w1044 = w1031 & w1043;
assign w1045 = ~w1031 & ~w1043;
assign w1046 = ~w1044 & ~w1045;
assign w1047 = w1020 & ~w1046;
assign w1048 = ~w1020 & w1046;
assign w1049 = ~w1047 & ~w1048;
assign w1050 = ~w995 & w1049;
assign w1051 = w995 & ~w1049;
assign w1052 = ~w1050 & ~w1051;
assign w1053 = w947 & ~w1052;
assign w1054 = ~w947 & w1052;
assign w1055 = ~w1053 & ~w1054;
assign w1056 = ~w934 & ~w1055;
assign w1057 = w934 & w1055;
assign w1058 = ~w1056 & ~w1057;
assign w1059 = w933 & ~w1058;
assign w1060 = ~w933 & w1058;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = (~w1026 & w1021) | (~w1026 & w9241) | (w1021 & w9241);
assign w1063 = pi14 & pi34;
assign w1064 = pi13 & pi35;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = pi14 & pi35;
assign w1067 = w827 & w1066;
assign w1068 = ~w1065 & ~w1067;
assign w1069 = pi15 & pi33;
assign w1070 = pi16 & pi32;
assign w1071 = pi80 & w1070;
assign w1072 = ~pi80 & ~w1070;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = w1069 & ~w1073;
assign w1075 = ~w1069 & w1073;
assign w1076 = ~w1074 & ~w1075;
assign w1077 = w1068 & ~w1076;
assign w1078 = ~w1068 & w1076;
assign w1079 = ~w1077 & ~w1078;
assign w1080 = (~w1036 & w1040) | (~w1036 & w8686) | (w1040 & w8686);
assign w1081 = w1079 & ~w1080;
assign w1082 = ~w1079 & w1080;
assign w1083 = ~w1081 & ~w1082;
assign w1084 = ~w1062 & w1083;
assign w1085 = w1062 & ~w1083;
assign w1086 = ~w1084 & ~w1085;
assign w1087 = pi03 & pi45;
assign w1088 = pi04 & pi44;
assign w1089 = ~w951 & ~w1088;
assign w1090 = pi05 & pi44;
assign w1091 = w948 & w1090;
assign w1092 = ~w1089 & ~w1091;
assign w1093 = w1087 & ~w1092;
assign w1094 = ~w1087 & w1092;
assign w1095 = ~w1093 & ~w1094;
assign w1096 = w976 & ~w978;
assign w1097 = w975 & ~w979;
assign w1098 = w974 & w979;
assign w1099 = ~w1097 & ~w1098;
assign w1100 = ~w1096 & w1099;
assign w1101 = ~w1095 & ~w1100;
assign w1102 = w1095 & w1100;
assign w1103 = ~w1101 & ~w1102;
assign w1104 = pi00 & pi48;
assign w1105 = pi01 & pi47;
assign w1106 = ~w964 & ~w1105;
assign w1107 = pi02 & pi47;
assign w1108 = w961 & w1107;
assign w1109 = ~w1106 & ~w1108;
assign w1110 = w1104 & ~w1109;
assign w1111 = ~w1104 & w1109;
assign w1112 = ~w1110 & ~w1111;
assign w1113 = w1103 & w1112;
assign w1114 = ~w1103 & ~w1112;
assign w1115 = ~w1113 & ~w1114;
assign w1116 = w1086 & ~w1115;
assign w1117 = ~w1086 & w1115;
assign w1118 = ~w1116 & ~w1117;
assign w1119 = pi06 & pi42;
assign w1120 = pi11 & pi37;
assign w1121 = ~w999 & ~w1120;
assign w1122 = pi12 & pi37;
assign w1123 = w996 & w1122;
assign w1124 = ~w1121 & ~w1123;
assign w1125 = pi10 & pi38;
assign w1126 = ~w1124 & w1125;
assign w1127 = w1124 & ~w1125;
assign w1128 = ~w1126 & ~w1127;
assign w1129 = w1119 & ~w1128;
assign w1130 = ~w1119 & w1128;
assign w1131 = ~w1129 & ~w1130;
assign w1132 = pi07 & pi41;
assign w1133 = pi08 & pi40;
assign w1134 = ~w1012 & ~w1133;
assign w1135 = pi09 & pi40;
assign w1136 = w1009 & w1135;
assign w1137 = ~w1134 & ~w1136;
assign w1138 = w1132 & ~w1137;
assign w1139 = ~w1132 & w1137;
assign w1140 = ~w1138 & ~w1139;
assign w1141 = w1131 & ~w1140;
assign w1142 = ~w1131 & w1140;
assign w1143 = ~w1141 & ~w1142;
assign w1144 = (~w957 & ~w959) | (~w957 & w8687) | (~w959 & w8687);
assign w1145 = w960 & ~w963;
assign w1146 = ~w965 & ~w1145;
assign w1147 = w883 & ~w950;
assign w1148 = ~w952 & ~w1147;
assign w1149 = ~w1146 & ~w1148;
assign w1150 = w1146 & w1148;
assign w1151 = ~w1149 & ~w1150;
assign w1152 = ~w1144 & w1151;
assign w1153 = w1144 & ~w1151;
assign w1154 = ~w1152 & ~w1153;
assign w1155 = w818 & ~w998;
assign w1156 = ~w1000 & ~w1155;
assign w1157 = w1008 & ~w1011;
assign w1158 = ~w1013 & ~w1157;
assign w1159 = ~w1156 & ~w1158;
assign w1160 = w1156 & w1158;
assign w1161 = ~w1159 & ~w1160;
assign w1162 = (~w1005 & ~w1007) | (~w1005 & w8688) | (~w1007 & w8688);
assign w1163 = w1161 & ~w1162;
assign w1164 = ~w1161 & w1162;
assign w1165 = ~w1163 & ~w1164;
assign w1166 = ~w1154 & ~w1165;
assign w1167 = w1154 & w1165;
assign w1168 = ~w1166 & ~w1167;
assign w1169 = w1143 & ~w1168;
assign w1170 = ~w1143 & w1168;
assign w1171 = ~w1169 & ~w1170;
assign w1172 = w1118 & ~w1171;
assign w1173 = ~w1118 & w1171;
assign w1174 = ~w1172 & ~w1173;
assign w1175 = ~w939 & ~w942;
assign w1176 = ~w993 & ~w1051;
assign w1177 = w983 & ~w985;
assign w1178 = ~w990 & ~w1177;
assign w1179 = (~w1045 & ~w1046) | (~w1045 & w9242) | (~w1046 & w9242);
assign w1180 = w1178 & w1179;
assign w1181 = ~w1178 & ~w1179;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = w1176 & ~w1182;
assign w1184 = ~w1176 & w1182;
assign w1185 = ~w1183 & ~w1184;
assign w1186 = w1175 & ~w1185;
assign w1187 = ~w1175 & w1185;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = w1174 & ~w1188;
assign w1190 = ~w1174 & w1188;
assign w1191 = ~w1189 & ~w1190;
assign w1192 = ~w945 & ~w1053;
assign w1193 = ~w1191 & w1192;
assign w1194 = w1191 & ~w1192;
assign w1195 = ~w1193 & ~w1194;
assign w1196 = ~w1056 & ~w933;
assign w1197 = ~w1057 & ~w1196;
assign w1198 = ~w1195 & ~w1197;
assign w1199 = w1195 & w1197;
assign w1200 = ~w1198 & ~w1199;
assign w1201 = ~w1193 & ~w1199;
assign w1202 = pi11 & pi38;
assign w1203 = pi10 & pi39;
assign w1204 = ~w1202 & ~w1203;
assign w1205 = pi11 & pi39;
assign w1206 = w1125 & w1205;
assign w1207 = ~w1204 & ~w1206;
assign w1208 = w1135 & ~w1207;
assign w1209 = ~w1135 & w1207;
assign w1210 = ~w1208 & ~w1209;
assign w1211 = w1090 & ~w1210;
assign w1212 = ~w1090 & w1210;
assign w1213 = ~w1211 & ~w1212;
assign w1214 = pi06 & pi43;
assign w1215 = pi07 & pi42;
assign w1216 = pi08 & pi41;
assign w1217 = ~w1215 & ~w1216;
assign w1218 = pi08 & pi42;
assign w1219 = w1132 & w1218;
assign w1220 = ~w1217 & ~w1219;
assign w1221 = w1214 & ~w1220;
assign w1222 = ~w1214 & w1220;
assign w1223 = ~w1221 & ~w1222;
assign w1224 = w1213 & ~w1223;
assign w1225 = ~w1213 & w1223;
assign w1226 = ~w1224 & ~w1225;
assign w1227 = ~w1121 & w1125;
assign w1228 = ~w1123 & ~w1227;
assign w1229 = w1132 & ~w1134;
assign w1230 = ~w1136 & ~w1229;
assign w1231 = ~w1228 & ~w1230;
assign w1232 = w1228 & w1230;
assign w1233 = ~w1231 & ~w1232;
assign w1234 = (~w1129 & ~w1131) | (~w1129 & w8689) | (~w1131 & w8689);
assign w1235 = w1233 & ~w1234;
assign w1236 = ~w1233 & w1234;
assign w1237 = ~w1235 & ~w1236;
assign w1238 = w1104 & ~w1106;
assign w1239 = ~w1108 & ~w1238;
assign w1240 = w1087 & ~w1089;
assign w1241 = ~w1091 & ~w1240;
assign w1242 = ~w1239 & ~w1241;
assign w1243 = w1239 & w1241;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = ~w1102 & ~w1113;
assign w1246 = w1244 & w1245;
assign w1247 = ~w1244 & ~w1245;
assign w1248 = ~w1246 & ~w1247;
assign w1249 = w1237 & w1248;
assign w1250 = ~w1237 & ~w1248;
assign w1251 = ~w1249 & ~w1250;
assign w1252 = w1226 & w1251;
assign w1253 = ~w1226 & ~w1251;
assign w1254 = ~w1252 & ~w1253;
assign w1255 = ~w1149 & ~w1152;
assign w1256 = pi13 & pi36;
assign w1257 = pi15 & pi34;
assign w1258 = ~w1066 & ~w1257;
assign w1259 = pi15 & pi35;
assign w1260 = w1063 & w1259;
assign w1261 = ~w1258 & ~w1260;
assign w1262 = w1256 & ~w1261;
assign w1263 = ~w1256 & w1261;
assign w1264 = ~w1262 & ~w1263;
assign w1265 = pi17 & pi32;
assign w1266 = pi81 & w1265;
assign w1267 = ~pi81 & ~w1265;
assign w1268 = ~w1266 & ~w1267;
assign w1269 = pi16 & pi33;
assign w1270 = ~w1122 & w1269;
assign w1271 = w1122 & ~w1269;
assign w1272 = ~w1270 & ~w1271;
assign w1273 = w1268 & w1272;
assign w1274 = ~w1268 & ~w1272;
assign w1275 = ~w1273 & ~w1274;
assign w1276 = ~w1264 & ~w1275;
assign w1277 = w1264 & w1275;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = (~w1159 & w1162) | (~w1159 & w9243) | (w1162 & w9243);
assign w1280 = ~w1278 & w1279;
assign w1281 = w1278 & ~w1279;
assign w1282 = ~w1280 & ~w1281;
assign w1283 = w1255 & w1282;
assign w1284 = ~w1255 & ~w1282;
assign w1285 = ~w1283 & ~w1284;
assign w1286 = ~w1069 & ~w1071;
assign w1287 = ~w1072 & ~w1286;
assign w1288 = (w1076 & w8690) | (w1076 & w8691) | (w8690 & w8691);
assign w1289 = (~w1076 & w8692) | (~w1076 & w8693) | (w8692 & w8693);
assign w1290 = ~w1288 & ~w1289;
assign w1291 = pi03 & pi46;
assign w1292 = pi04 & pi45;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = pi04 & pi46;
assign w1295 = w1087 & w1294;
assign w1296 = ~w1293 & ~w1295;
assign w1297 = w1107 & ~w1296;
assign w1298 = ~w1107 & w1296;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = w1290 & ~w1299;
assign w1301 = ~w1290 & w1299;
assign w1302 = ~w1300 & ~w1301;
assign w1303 = pi00 & pi49;
assign w1304 = pi01 & pi48;
assign w1305 = ~w1303 & ~w1304;
assign w1306 = pi01 & pi49;
assign w1307 = w1104 & w1306;
assign w1308 = ~w1305 & ~w1307;
assign w1309 = w975 & w979;
assign w1310 = ~w1308 & w1309;
assign w1311 = w1308 & ~w1309;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = w1302 & w1312;
assign w1314 = ~w1302 & ~w1312;
assign w1315 = ~w1313 & ~w1314;
assign w1316 = ~w1285 & ~w1315;
assign w1317 = w1285 & w1315;
assign w1318 = ~w1316 & ~w1317;
assign w1319 = w1254 & w1318;
assign w1320 = ~w1254 & ~w1318;
assign w1321 = ~w1319 & ~w1320;
assign w1322 = (~w1180 & w1176) | (~w1180 & w9244) | (w1176 & w9244);
assign w1323 = w1321 & ~w1322;
assign w1324 = ~w1321 & w1322;
assign w1325 = ~w1323 & ~w1324;
assign w1326 = ~w1116 & ~w1172;
assign w1327 = ~w1081 & ~w1084;
assign w1328 = (~w1166 & ~w1168) | (~w1166 & w9245) | (~w1168 & w9245);
assign w1329 = ~w1327 & w1328;
assign w1330 = w1327 & ~w1328;
assign w1331 = ~w1329 & ~w1330;
assign w1332 = w1326 & w1331;
assign w1333 = ~w1326 & ~w1331;
assign w1334 = ~w1332 & ~w1333;
assign w1335 = w1325 & ~w1334;
assign w1336 = ~w1325 & w1334;
assign w1337 = ~w1335 & ~w1336;
assign w1338 = (~w1186 & ~w1188) | (~w1186 & w9246) | (~w1188 & w9246);
assign w1339 = ~w1337 & ~w1338;
assign w1340 = w1337 & w1338;
assign w1341 = ~w1339 & ~w1340;
assign w1342 = w1201 & w1341;
assign w1343 = ~w1201 & ~w1341;
assign w1344 = ~w1342 & ~w1343;
assign w1345 = ~w1323 & ~w1335;
assign w1346 = ~w1316 & ~w1319;
assign w1347 = ~w1280 & ~w1283;
assign w1348 = ~w1249 & ~w1252;
assign w1349 = w1347 & ~w1348;
assign w1350 = ~w1347 & w1348;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = ~w1346 & w1351;
assign w1353 = w1346 & ~w1351;
assign w1354 = ~w1352 & ~w1353;
assign w1355 = ~w1242 & ~w1246;
assign w1356 = pi12 & pi38;
assign w1357 = ~w1205 & ~w1356;
assign w1358 = pi12 & pi39;
assign w1359 = w1202 & w1358;
assign w1360 = ~w1357 & ~w1359;
assign w1361 = (~w1231 & w1234) | (~w1231 & w9247) | (w1234 & w9247);
assign w1362 = ~w1360 & w1361;
assign w1363 = w1360 & ~w1361;
assign w1364 = ~w1362 & ~w1363;
assign w1365 = w1355 & w1364;
assign w1366 = ~w1355 & ~w1364;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = pi14 & pi36;
assign w1369 = pi16 & pi34;
assign w1370 = ~w1259 & ~w1369;
assign w1371 = pi16 & pi35;
assign w1372 = w1257 & w1371;
assign w1373 = ~w1370 & ~w1372;
assign w1374 = w1368 & ~w1373;
assign w1375 = ~w1368 & w1373;
assign w1376 = ~w1374 & ~w1375;
assign w1377 = pi18 & pi32;
assign w1378 = pi82 & w1377;
assign w1379 = ~pi82 & ~w1377;
assign w1380 = ~w1378 & ~w1379;
assign w1381 = pi13 & pi37;
assign w1382 = pi17 & pi33;
assign w1383 = ~w1381 & w1382;
assign w1384 = w1381 & ~w1382;
assign w1385 = ~w1383 & ~w1384;
assign w1386 = w1380 & w1385;
assign w1387 = ~w1380 & ~w1385;
assign w1388 = ~w1386 & ~w1387;
assign w1389 = w1376 & w1388;
assign w1390 = ~w1376 & ~w1388;
assign w1391 = ~w1389 & ~w1390;
assign w1392 = pi02 & pi48;
assign w1393 = pi03 & pi47;
assign w1394 = ~w1392 & ~w1393;
assign w1395 = pi03 & pi48;
assign w1396 = w1107 & w1395;
assign w1397 = ~w1394 & ~w1396;
assign w1398 = w1306 & ~w1397;
assign w1399 = ~w1306 & w1397;
assign w1400 = ~w1398 & ~w1399;
assign w1401 = w1391 & ~w1400;
assign w1402 = ~w1391 & w1400;
assign w1403 = ~w1401 & ~w1402;
assign w1404 = w1256 & ~w1258;
assign w1405 = ~w1260 & ~w1404;
assign w1406 = ~w1266 & ~w1269;
assign w1407 = ~w1267 & ~w1406;
assign w1408 = ~w1405 & w1407;
assign w1409 = w1405 & ~w1407;
assign w1410 = ~w1408 & ~w1409;
assign w1411 = w1122 & w1275;
assign w1412 = ~w1276 & ~w1411;
assign w1413 = w1410 & ~w1412;
assign w1414 = ~w1410 & w1412;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = pi00 & pi50;
assign w1417 = ~w1289 & ~w1416;
assign w1418 = w1289 & w1416;
assign w1419 = ~w1417 & ~w1418;
assign w1420 = ~w1415 & w1419;
assign w1421 = w1415 & ~w1419;
assign w1422 = ~w1420 & ~w1421;
assign w1423 = w1403 & ~w1422;
assign w1424 = ~w1403 & w1422;
assign w1425 = ~w1423 & ~w1424;
assign w1426 = w1367 & ~w1425;
assign w1427 = ~w1367 & w1425;
assign w1428 = ~w1426 & ~w1427;
assign w1429 = (~w1211 & ~w1213) | (~w1211 & w9248) | (~w1213 & w9248);
assign w1430 = w1214 & ~w1217;
assign w1431 = ~w1219 & ~w1430;
assign w1432 = w1135 & ~w1204;
assign w1433 = ~w1206 & ~w1432;
assign w1434 = ~w1431 & ~w1433;
assign w1435 = w1431 & w1433;
assign w1436 = ~w1434 & ~w1435;
assign w1437 = ~w1429 & w1436;
assign w1438 = w1429 & ~w1436;
assign w1439 = ~w1437 & ~w1438;
assign w1440 = pi09 & pi41;
assign w1441 = pi10 & pi40;
assign w1442 = ~w1440 & ~w1441;
assign w1443 = pi10 & pi41;
assign w1444 = w1135 & w1443;
assign w1445 = ~w1442 & ~w1444;
assign w1446 = w1218 & ~w1445;
assign w1447 = ~w1218 & w1445;
assign w1448 = ~w1446 & ~w1447;
assign w1449 = w1294 & ~w1448;
assign w1450 = ~w1294 & w1448;
assign w1451 = ~w1449 & ~w1450;
assign w1452 = pi05 & pi45;
assign w1453 = pi06 & pi44;
assign w1454 = pi07 & pi43;
assign w1455 = ~w1453 & ~w1454;
assign w1456 = pi07 & pi44;
assign w1457 = w1214 & w1456;
assign w1458 = ~w1455 & ~w1457;
assign w1459 = w1452 & ~w1458;
assign w1460 = ~w1452 & w1458;
assign w1461 = ~w1459 & ~w1460;
assign w1462 = w1451 & ~w1461;
assign w1463 = ~w1451 & w1461;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = w1439 & w1464;
assign w1466 = ~w1439 & ~w1464;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = w1107 & ~w1293;
assign w1469 = ~w1295 & ~w1468;
assign w1470 = ~w1305 & w1309;
assign w1471 = ~w1307 & ~w1470;
assign w1472 = ~w1469 & ~w1471;
assign w1473 = w1469 & w1471;
assign w1474 = ~w1472 & ~w1473;
assign w1475 = (~w1301 & ~w1302) | (~w1301 & w9249) | (~w1302 & w9249);
assign w1476 = w1474 & w1475;
assign w1477 = ~w1474 & ~w1475;
assign w1478 = ~w1476 & ~w1477;
assign w1479 = w1467 & ~w1478;
assign w1480 = ~w1467 & w1478;
assign w1481 = ~w1479 & ~w1480;
assign w1482 = w1428 & w1481;
assign w1483 = ~w1428 & ~w1481;
assign w1484 = ~w1482 & ~w1483;
assign w1485 = (~w1330 & ~w1326) | (~w1330 & w9250) | (~w1326 & w9250);
assign w1486 = ~w1484 & w1485;
assign w1487 = w1484 & ~w1485;
assign w1488 = ~w1486 & ~w1487;
assign w1489 = w1354 & ~w1488;
assign w1490 = ~w1354 & w1488;
assign w1491 = ~w1489 & ~w1490;
assign w1492 = ~w1345 & ~w1491;
assign w1493 = w1345 & w1491;
assign w1494 = ~w1492 & ~w1493;
assign w1495 = ~w1339 & ~w1342;
assign w1496 = w1494 & w1495;
assign w1497 = ~w1494 & ~w1495;
assign w1498 = ~w1496 & ~w1497;
assign w1499 = ~w1492 & ~w1496;
assign w1500 = pi14 & pi37;
assign w1501 = pi18 & pi33;
assign w1502 = pi19 & pi32;
assign w1503 = pi83 & w1502;
assign w1504 = ~pi83 & ~w1502;
assign w1505 = ~w1503 & ~w1504;
assign w1506 = w1501 & w1505;
assign w1507 = ~w1501 & ~w1505;
assign w1508 = ~w1506 & ~w1507;
assign w1509 = w1500 & w1508;
assign w1510 = ~w1500 & ~w1508;
assign w1511 = ~w1509 & ~w1510;
assign w1512 = pi15 & pi36;
assign w1513 = pi17 & pi34;
assign w1514 = ~w1371 & ~w1513;
assign w1515 = pi17 & pi35;
assign w1516 = w1369 & w1515;
assign w1517 = ~w1514 & ~w1516;
assign w1518 = w1512 & ~w1517;
assign w1519 = ~w1512 & w1517;
assign w1520 = ~w1518 & ~w1519;
assign w1521 = w1511 & ~w1520;
assign w1522 = ~w1511 & w1520;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = pi00 & pi51;
assign w1525 = pi01 & pi50;
assign w1526 = pi02 & pi49;
assign w1527 = ~w1525 & ~w1526;
assign w1528 = pi02 & pi50;
assign w1529 = w1306 & w1528;
assign w1530 = ~w1527 & ~w1529;
assign w1531 = w1524 & ~w1530;
assign w1532 = ~w1524 & w1530;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = w1523 & ~w1533;
assign w1535 = ~w1523 & w1533;
assign w1536 = ~w1534 & ~w1535;
assign w1537 = w1368 & ~w1370;
assign w1538 = ~w1372 & ~w1537;
assign w1539 = ~w1378 & ~w1382;
assign w1540 = ~w1379 & ~w1539;
assign w1541 = ~w1538 & w1540;
assign w1542 = w1538 & ~w1540;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = w1381 & w1388;
assign w1545 = ~w1390 & ~w1544;
assign w1546 = w1543 & ~w1545;
assign w1547 = ~w1543 & w1545;
assign w1548 = ~w1546 & ~w1547;
assign w1549 = (~w1408 & w1412) | (~w1408 & w8590) | (w1412 & w8590);
assign w1550 = w1359 & ~w1549;
assign w1551 = ~w1359 & w1549;
assign w1552 = ~w1550 & ~w1551;
assign w1553 = w1548 & w1552;
assign w1554 = ~w1548 & ~w1552;
assign w1555 = ~w1553 & ~w1554;
assign w1556 = w1536 & w1555;
assign w1557 = ~w1536 & ~w1555;
assign w1558 = ~w1556 & ~w1557;
assign w1559 = ~w1434 & ~w1437;
assign w1560 = pi11 & pi40;
assign w1561 = pi13 & pi38;
assign w1562 = ~w1358 & ~w1561;
assign w1563 = pi13 & pi39;
assign w1564 = w1356 & w1563;
assign w1565 = ~w1562 & ~w1564;
assign w1566 = w1560 & w1565;
assign w1567 = ~w1560 & ~w1565;
assign w1568 = ~w1566 & ~w1567;
assign w1569 = w1443 & w1568;
assign w1570 = ~w1443 & ~w1568;
assign w1571 = ~w1569 & ~w1570;
assign w1572 = ~w1559 & w1571;
assign w1573 = w1559 & ~w1571;
assign w1574 = ~w1572 & ~w1573;
assign w1575 = ~w1472 & ~w1476;
assign w1576 = w1574 & ~w1575;
assign w1577 = ~w1574 & w1575;
assign w1578 = ~w1576 & ~w1577;
assign w1579 = w1558 & w1578;
assign w1580 = ~w1558 & ~w1578;
assign w1581 = ~w1579 & ~w1580;
assign w1582 = ~w1449 & ~w1462;
assign w1583 = w1452 & ~w1455;
assign w1584 = ~w1457 & ~w1583;
assign w1585 = w1218 & ~w1442;
assign w1586 = ~w1444 & ~w1585;
assign w1587 = ~w1584 & ~w1586;
assign w1588 = w1584 & w1586;
assign w1589 = ~w1587 & ~w1588;
assign w1590 = ~w1582 & w1589;
assign w1591 = w1582 & ~w1589;
assign w1592 = ~w1590 & ~w1591;
assign w1593 = pi08 & pi43;
assign w1594 = pi09 & pi42;
assign w1595 = ~w1593 & ~w1594;
assign w1596 = pi09 & pi43;
assign w1597 = w1218 & w1596;
assign w1598 = ~w1595 & ~w1597;
assign w1599 = w1456 & ~w1598;
assign w1600 = ~w1456 & w1598;
assign w1601 = ~w1599 & ~w1600;
assign w1602 = w1395 & ~w1601;
assign w1603 = ~w1395 & w1601;
assign w1604 = ~w1602 & ~w1603;
assign w1605 = pi04 & pi47;
assign w1606 = pi05 & pi46;
assign w1607 = pi06 & pi45;
assign w1608 = ~w1606 & ~w1607;
assign w1609 = pi06 & pi46;
assign w1610 = w1452 & w1609;
assign w1611 = ~w1608 & ~w1610;
assign w1612 = w1605 & ~w1611;
assign w1613 = ~w1605 & w1611;
assign w1614 = ~w1612 & ~w1613;
assign w1615 = w1604 & ~w1614;
assign w1616 = ~w1604 & w1614;
assign w1617 = ~w1615 & ~w1616;
assign w1618 = w1592 & w1617;
assign w1619 = ~w1592 & ~w1617;
assign w1620 = ~w1618 & ~w1619;
assign w1621 = (~w1401 & w1422) | (~w1401 & w8694) | (w1422 & w8694);
assign w1622 = w1306 & ~w1394;
assign w1623 = ~w1396 & ~w1622;
assign w1624 = (~w1623 & w1289) | (~w1623 & w9251) | (w1289 & w9251);
assign w1625 = (w1624 & w1415) | (w1624 & w8695) | (w1415 & w8695);
assign w1626 = ~w1418 & w1623;
assign w1627 = ~w1625 & ~w1626;
assign w1628 = w1415 & w9252;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = ~w1621 & ~w1629;
assign w1631 = w1621 & w1629;
assign w1632 = ~w1630 & ~w1631;
assign w1633 = w1620 & ~w1632;
assign w1634 = ~w1620 & w1632;
assign w1635 = ~w1633 & ~w1634;
assign w1636 = w1581 & ~w1635;
assign w1637 = ~w1581 & w1635;
assign w1638 = ~w1636 & ~w1637;
assign w1639 = ~w1349 & ~w1352;
assign w1640 = ~w1426 & ~w1482;
assign w1641 = ~w1362 & ~w1365;
assign w1642 = ~w1466 & ~w1479;
assign w1643 = w1641 & w1642;
assign w1644 = ~w1641 & ~w1642;
assign w1645 = ~w1643 & ~w1644;
assign w1646 = w1640 & w1645;
assign w1647 = ~w1640 & ~w1645;
assign w1648 = ~w1646 & ~w1647;
assign w1649 = ~w1639 & w1648;
assign w1650 = w1639 & ~w1648;
assign w1651 = ~w1649 & ~w1650;
assign w1652 = w1638 & w1651;
assign w1653 = ~w1638 & ~w1651;
assign w1654 = ~w1652 & ~w1653;
assign w1655 = ~w1487 & ~w1490;
assign w1656 = ~w1654 & ~w1655;
assign w1657 = w1654 & w1655;
assign w1658 = ~w1656 & ~w1657;
assign w1659 = w1499 & ~w1658;
assign w1660 = ~w1499 & w1658;
assign w1661 = ~w1659 & ~w1660;
assign w1662 = ~w1057 & w1195;
assign w1663 = w1341 & w1494;
assign w1664 = w1662 & w1663;
assign w1665 = w1658 & w1664;
assign w1666 = ~w1196 & w1665;
assign w1667 = ~w1193 & ~w1340;
assign w1668 = ~w1339 & ~w1493;
assign w1669 = ~w1667 & w1668;
assign w1670 = ~w1492 & ~w1657;
assign w1671 = ~w1669 & w1670;
assign w1672 = ~w1656 & ~w1671;
assign w1673 = ~w1666 & ~w1672;
assign w1674 = ~w1649 & ~w1652;
assign w1675 = ~w1643 & ~w1646;
assign w1676 = ~w1579 & ~w1636;
assign w1677 = ~w1572 & ~w1576;
assign w1678 = ~w1619 & ~w1633;
assign w1679 = ~w1677 & w1678;
assign w1680 = w1677 & ~w1678;
assign w1681 = ~w1679 & ~w1680;
assign w1682 = ~w1676 & w1681;
assign w1683 = w1676 & ~w1681;
assign w1684 = ~w1682 & ~w1683;
assign w1685 = ~w1675 & w1684;
assign w1686 = w1675 & ~w1684;
assign w1687 = ~w1685 & ~w1686;
assign w1688 = ~w1587 & ~w1590;
assign w1689 = pi11 & pi41;
assign w1690 = pi10 & pi42;
assign w1691 = ~w1689 & ~w1690;
assign w1692 = pi11 & pi42;
assign w1693 = w1443 & w1692;
assign w1694 = ~w1691 & ~w1693;
assign w1695 = pi12 & pi40;
assign w1696 = pi14 & pi38;
assign w1697 = ~w1563 & ~w1696;
assign w1698 = pi14 & pi39;
assign w1699 = w1561 & w1698;
assign w1700 = ~w1697 & ~w1699;
assign w1701 = w1695 & ~w1700;
assign w1702 = ~w1695 & w1700;
assign w1703 = ~w1701 & ~w1702;
assign w1704 = w1694 & ~w1703;
assign w1705 = ~w1694 & w1703;
assign w1706 = ~w1704 & ~w1705;
assign w1707 = ~w1688 & w1706;
assign w1708 = w1688 & ~w1706;
assign w1709 = ~w1707 & ~w1708;
assign w1710 = ~w1625 & ~w1630;
assign w1711 = w1709 & ~w1710;
assign w1712 = ~w1709 & w1710;
assign w1713 = ~w1711 & ~w1712;
assign w1714 = pi15 & pi37;
assign w1715 = pi19 & pi33;
assign w1716 = pi20 & pi32;
assign w1717 = pi84 & w1716;
assign w1718 = ~pi84 & ~w1716;
assign w1719 = ~w1717 & ~w1718;
assign w1720 = w1715 & w1719;
assign w1721 = ~w1715 & ~w1719;
assign w1722 = ~w1720 & ~w1721;
assign w1723 = w1714 & w1722;
assign w1724 = ~w1714 & ~w1722;
assign w1725 = ~w1723 & ~w1724;
assign w1726 = pi16 & pi36;
assign w1727 = pi18 & pi34;
assign w1728 = ~w1515 & ~w1727;
assign w1729 = pi18 & pi35;
assign w1730 = w1513 & w1729;
assign w1731 = ~w1728 & ~w1730;
assign w1732 = w1726 & ~w1731;
assign w1733 = ~w1726 & w1731;
assign w1734 = ~w1732 & ~w1733;
assign w1735 = w1725 & ~w1734;
assign w1736 = ~w1725 & w1734;
assign w1737 = ~w1735 & ~w1736;
assign w1738 = pi00 & pi52;
assign w1739 = pi01 & pi51;
assign w1740 = ~w1528 & ~w1739;
assign w1741 = pi02 & pi51;
assign w1742 = w1525 & w1741;
assign w1743 = ~w1740 & ~w1742;
assign w1744 = w1738 & ~w1743;
assign w1745 = ~w1738 & w1743;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = w1737 & ~w1746;
assign w1748 = ~w1737 & w1746;
assign w1749 = ~w1747 & ~w1748;
assign w1750 = (~w1509 & ~w1511) | (~w1509 & w8591) | (~w1511 & w8591);
assign w1751 = (~w1503 & ~w1505) | (~w1503 & w9253) | (~w1505 & w9253);
assign w1752 = w1512 & ~w1514;
assign w1753 = ~w1516 & ~w1752;
assign w1754 = ~w1751 & ~w1753;
assign w1755 = w1751 & w1753;
assign w1756 = ~w1754 & ~w1755;
assign w1757 = ~w1750 & w1756;
assign w1758 = w1750 & ~w1756;
assign w1759 = ~w1757 & ~w1758;
assign w1760 = (~w1541 & w1545) | (~w1541 & w8592) | (w1545 & w8592);
assign w1761 = (~w1564 & ~w1568) | (~w1564 & w8593) | (~w1568 & w8593);
assign w1762 = w1568 & w8594;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = ~w1566 & ~w1763;
assign w1765 = w1760 & w1764;
assign w1766 = ~w1760 & ~w1764;
assign w1767 = ~w1765 & ~w1766;
assign w1768 = w1759 & ~w1767;
assign w1769 = ~w1759 & w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = w1749 & ~w1770;
assign w1772 = ~w1749 & w1770;
assign w1773 = ~w1771 & ~w1772;
assign w1774 = w1713 & w1773;
assign w1775 = ~w1713 & ~w1773;
assign w1776 = ~w1774 & ~w1775;
assign w1777 = (~w1534 & ~w1555) | (~w1534 & w8696) | (~w1555 & w8696);
assign w1778 = (~w1550 & ~w1552) | (~w1550 & w8697) | (~w1552 & w8697);
assign w1779 = w1524 & ~w1527;
assign w1780 = ~w1529 & ~w1779;
assign w1781 = ~w1778 & ~w1780;
assign w1782 = w1778 & w1780;
assign w1783 = ~w1781 & ~w1782;
assign w1784 = ~w1777 & w1783;
assign w1785 = w1777 & ~w1783;
assign w1786 = ~w1784 & ~w1785;
assign w1787 = pi03 & pi49;
assign w1788 = pi07 & pi45;
assign w1789 = pi08 & pi44;
assign w1790 = ~w1596 & ~w1789;
assign w1791 = pi09 & pi44;
assign w1792 = w1593 & w1791;
assign w1793 = ~w1790 & ~w1792;
assign w1794 = w1788 & ~w1793;
assign w1795 = ~w1788 & w1793;
assign w1796 = ~w1794 & ~w1795;
assign w1797 = w1787 & ~w1796;
assign w1798 = ~w1787 & w1796;
assign w1799 = ~w1797 & ~w1798;
assign w1800 = pi04 & pi48;
assign w1801 = pi05 & pi47;
assign w1802 = ~w1609 & ~w1801;
assign w1803 = pi06 & pi47;
assign w1804 = w1606 & w1803;
assign w1805 = ~w1802 & ~w1804;
assign w1806 = w1800 & ~w1805;
assign w1807 = ~w1800 & w1805;
assign w1808 = ~w1806 & ~w1807;
assign w1809 = w1799 & ~w1808;
assign w1810 = ~w1799 & w1808;
assign w1811 = ~w1809 & ~w1810;
assign w1812 = ~w1602 & ~w1615;
assign w1813 = w1605 & ~w1608;
assign w1814 = ~w1610 & ~w1813;
assign w1815 = w1456 & ~w1595;
assign w1816 = ~w1597 & ~w1815;
assign w1817 = ~w1814 & ~w1816;
assign w1818 = w1814 & w1816;
assign w1819 = ~w1817 & ~w1818;
assign w1820 = ~w1812 & w1819;
assign w1821 = w1812 & ~w1819;
assign w1822 = ~w1820 & ~w1821;
assign w1823 = w1811 & w1822;
assign w1824 = ~w1811 & ~w1822;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = ~w1786 & ~w1825;
assign w1827 = w1786 & w1825;
assign w1828 = ~w1826 & ~w1827;
assign w1829 = w1776 & w1828;
assign w1830 = ~w1776 & ~w1828;
assign w1831 = ~w1829 & ~w1830;
assign w1832 = w1687 & w1831;
assign w1833 = ~w1687 & ~w1831;
assign w1834 = ~w1832 & ~w1833;
assign w1835 = ~w1674 & w1834;
assign w1836 = w1674 & ~w1834;
assign w1837 = ~w1835 & ~w1836;
assign w1838 = ~w1673 & w1837;
assign w1839 = w1673 & ~w1837;
assign w1840 = ~w1838 & ~w1839;
assign w1841 = ~w1685 & ~w1832;
assign w1842 = pi16 & pi37;
assign w1843 = pi20 & pi33;
assign w1844 = pi21 & pi32;
assign w1845 = pi85 & w1844;
assign w1846 = ~pi85 & ~w1844;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = w1843 & w1847;
assign w1849 = ~w1843 & ~w1847;
assign w1850 = ~w1848 & ~w1849;
assign w1851 = w1842 & w1850;
assign w1852 = ~w1842 & ~w1850;
assign w1853 = ~w1851 & ~w1852;
assign w1854 = pi17 & pi36;
assign w1855 = pi19 & pi34;
assign w1856 = ~w1729 & ~w1855;
assign w1857 = pi19 & pi35;
assign w1858 = w1727 & w1857;
assign w1859 = ~w1856 & ~w1858;
assign w1860 = w1854 & ~w1859;
assign w1861 = ~w1854 & w1859;
assign w1862 = ~w1860 & ~w1861;
assign w1863 = w1853 & ~w1862;
assign w1864 = ~w1853 & w1862;
assign w1865 = ~w1863 & ~w1864;
assign w1866 = pi00 & pi53;
assign w1867 = pi01 & pi52;
assign w1868 = ~w1866 & ~w1867;
assign w1869 = pi01 & pi53;
assign w1870 = w1738 & w1869;
assign w1871 = ~w1868 & ~w1870;
assign w1872 = w1871 & w9295;
assign w1873 = (w1750 & w9254) | (w1750 & w9255) | (w9254 & w9255);
assign w1874 = ~w1872 & ~w1873;
assign w1875 = w1865 & w1874;
assign w1876 = ~w1865 & ~w1874;
assign w1877 = ~w1875 & ~w1876;
assign w1878 = (~w1693 & w1703) | (~w1693 & w8699) | (w1703 & w8699);
assign w1879 = w1695 & ~w1697;
assign w1880 = ~w1699 & ~w1879;
assign w1881 = ~w1878 & ~w1880;
assign w1882 = w1878 & w1880;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = (~w1723 & ~w1725) | (~w1723 & w8595) | (~w1725 & w8595);
assign w1885 = (~w1717 & ~w1719) | (~w1717 & w8596) | (~w1719 & w8596);
assign w1886 = w1726 & ~w1728;
assign w1887 = ~w1730 & ~w1886;
assign w1888 = ~w1885 & ~w1887;
assign w1889 = w1885 & w1887;
assign w1890 = ~w1888 & ~w1889;
assign w1891 = w1884 & ~w1890;
assign w1892 = ~w1884 & w1890;
assign w1893 = ~w1891 & ~w1892;
assign w1894 = w1762 & w1893;
assign w1895 = ~w1762 & ~w1893;
assign w1896 = ~w1894 & ~w1895;
assign w1897 = w1883 & ~w1896;
assign w1898 = ~w1883 & w1896;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = w1877 & ~w1899;
assign w1901 = ~w1877 & w1899;
assign w1902 = ~w1900 & ~w1901;
assign w1903 = ~w1817 & ~w1820;
assign w1904 = pi13 & pi40;
assign w1905 = pi15 & pi38;
assign w1906 = ~w1698 & ~w1905;
assign w1907 = pi15 & pi39;
assign w1908 = w1696 & w1907;
assign w1909 = ~w1906 & ~w1908;
assign w1910 = w1904 & ~w1909;
assign w1911 = ~w1904 & w1909;
assign w1912 = ~w1910 & ~w1911;
assign w1913 = w1791 & ~w1912;
assign w1914 = ~w1791 & w1912;
assign w1915 = ~w1913 & ~w1914;
assign w1916 = pi10 & pi43;
assign w1917 = pi12 & pi41;
assign w1918 = ~w1692 & ~w1917;
assign w1919 = pi12 & pi42;
assign w1920 = w1689 & w1919;
assign w1921 = ~w1918 & ~w1920;
assign w1922 = w1916 & ~w1921;
assign w1923 = ~w1916 & w1921;
assign w1924 = ~w1922 & ~w1923;
assign w1925 = w1915 & ~w1924;
assign w1926 = ~w1915 & w1924;
assign w1927 = ~w1925 & ~w1926;
assign w1928 = ~w1903 & w1927;
assign w1929 = w1903 & ~w1927;
assign w1930 = ~w1928 & ~w1929;
assign w1931 = (w1930 & w1784) | (w1930 & w9256) | (w1784 & w9256);
assign w1932 = ~w1784 & w9257;
assign w1933 = ~w1931 & ~w1932;
assign w1934 = w1902 & w1933;
assign w1935 = ~w1902 & ~w1933;
assign w1936 = ~w1934 & ~w1935;
assign w1937 = pi08 & pi45;
assign w1938 = pi07 & pi46;
assign w1939 = ~w1937 & ~w1938;
assign w1940 = pi08 & pi46;
assign w1941 = w1788 & w1940;
assign w1942 = ~w1939 & ~w1941;
assign w1943 = w1803 & ~w1942;
assign w1944 = ~w1803 & w1942;
assign w1945 = ~w1943 & ~w1944;
assign w1946 = w1741 & ~w1945;
assign w1947 = ~w1741 & w1945;
assign w1948 = ~w1946 & ~w1947;
assign w1949 = pi03 & pi50;
assign w1950 = pi04 & pi49;
assign w1951 = pi05 & pi48;
assign w1952 = ~w1950 & ~w1951;
assign w1953 = pi05 & pi49;
assign w1954 = w1800 & w1953;
assign w1955 = ~w1952 & ~w1954;
assign w1956 = w1949 & ~w1955;
assign w1957 = ~w1949 & w1955;
assign w1958 = ~w1956 & ~w1957;
assign w1959 = w1948 & ~w1958;
assign w1960 = ~w1948 & w1958;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = ~w1797 & ~w1809;
assign w1963 = w1800 & ~w1802;
assign w1964 = ~w1804 & ~w1963;
assign w1965 = w1788 & ~w1790;
assign w1966 = ~w1792 & ~w1965;
assign w1967 = ~w1964 & ~w1966;
assign w1968 = w1964 & w1966;
assign w1969 = ~w1967 & ~w1968;
assign w1970 = ~w1962 & w1969;
assign w1971 = w1962 & ~w1969;
assign w1972 = ~w1970 & ~w1971;
assign w1973 = (~w1747 & w1770) | (~w1747 & w8700) | (w1770 & w8700);
assign w1974 = w1738 & ~w1740;
assign w1975 = ~w1742 & ~w1974;
assign w1976 = ~w1769 & w8701;
assign w1977 = (w1975 & w1769) | (w1975 & w8702) | (w1769 & w8702);
assign w1978 = ~w1976 & ~w1977;
assign w1979 = ~w1973 & w1978;
assign w1980 = w1973 & ~w1978;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = w1972 & w1981;
assign w1983 = ~w1972 & ~w1981;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = w1961 & ~w1984;
assign w1986 = ~w1961 & w1984;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = w1936 & ~w1987;
assign w1989 = ~w1936 & w1987;
assign w1990 = ~w1988 & ~w1989;
assign w1991 = ~w1679 & ~w1682;
assign w1992 = ~w1707 & ~w1711;
assign w1993 = (~w1823 & ~w1786) | (~w1823 & w9258) | (~w1786 & w9258);
assign w1994 = ~w1992 & ~w1993;
assign w1995 = w1992 & w1993;
assign w1996 = ~w1994 & ~w1995;
assign w1997 = ~w1774 & ~w1828;
assign w1998 = ~w1775 & ~w1997;
assign w1999 = w1996 & w1998;
assign w2000 = ~w1996 & ~w1998;
assign w2001 = ~w1999 & ~w2000;
assign w2002 = ~w1991 & w2001;
assign w2003 = w1991 & ~w2001;
assign w2004 = ~w2002 & ~w2003;
assign w2005 = w1990 & w2004;
assign w2006 = ~w1990 & ~w2004;
assign w2007 = ~w2005 & ~w2006;
assign w2008 = w1841 & ~w2007;
assign w2009 = ~w1841 & w2007;
assign w2010 = ~w2008 & ~w2009;
assign w2011 = ~w1835 & ~w1838;
assign w2012 = w2010 & w2011;
assign w2013 = ~w2010 & ~w2011;
assign w2014 = ~w2012 & ~w2013;
assign w2015 = (~w2002 & ~w2004) | (~w2002 & w9259) | (~w2004 & w9259);
assign w2016 = (~w1934 & w1987) | (~w1934 & w9260) | (w1987 & w9260);
assign w2017 = ~w1928 & ~w1931;
assign w2018 = (~w1983 & ~w1984) | (~w1983 & w9261) | (~w1984 & w9261);
assign w2019 = ~w2017 & w2018;
assign w2020 = w2017 & ~w2018;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = ~w2016 & w2021;
assign w2023 = w2016 & ~w2021;
assign w2024 = ~w2022 & ~w2023;
assign w2025 = (~w1994 & ~w1998) | (~w1994 & w9262) | (~w1998 & w9262);
assign w2026 = pi00 & pi54;
assign w2027 = (~w1889 & w1735) | (~w1889 & w8597) | (w1735 & w8597);
assign w2028 = (w1735 & w8703) | (w1735 & w8704) | (w8703 & w8704);
assign w2029 = ~w1723 & w8598;
assign w2030 = w1889 & w2026;
assign w2031 = (~w2030 & w1735) | (~w2030 & w8599) | (w1735 & w8599);
assign w2032 = w1881 & w2031;
assign w2033 = ~w2028 & w2032;
assign w2034 = ~w1881 & ~w2031;
assign w2035 = ~w1881 & ~w2026;
assign w2036 = w2027 & w2035;
assign w2037 = ~w2034 & ~w2036;
assign w2038 = ~w2033 & w2037;
assign w2039 = pi10 & pi44;
assign w2040 = pi14 & pi40;
assign w2041 = pi16 & pi38;
assign w2042 = ~w1907 & ~w2041;
assign w2043 = pi16 & pi39;
assign w2044 = w1905 & w2043;
assign w2045 = ~w2042 & ~w2044;
assign w2046 = w2040 & ~w2045;
assign w2047 = ~w2040 & w2045;
assign w2048 = ~w2046 & ~w2047;
assign w2049 = w2039 & ~w2048;
assign w2050 = ~w2039 & w2048;
assign w2051 = ~w2049 & ~w2050;
assign w2052 = pi11 & pi43;
assign w2053 = pi13 & pi41;
assign w2054 = ~w1919 & ~w2053;
assign w2055 = pi13 & pi42;
assign w2056 = w1917 & w2055;
assign w2057 = ~w2054 & ~w2056;
assign w2058 = w2052 & ~w2057;
assign w2059 = ~w2052 & w2057;
assign w2060 = ~w2058 & ~w2059;
assign w2061 = w2051 & ~w2060;
assign w2062 = ~w2051 & w2060;
assign w2063 = ~w2061 & ~w2062;
assign w2064 = ~w2038 & w2063;
assign w2065 = w2038 & ~w2063;
assign w2066 = ~w2064 & ~w2065;
assign w2067 = pi17 & pi37;
assign w2068 = pi21 & pi33;
assign w2069 = pi22 & pi32;
assign w2070 = pi86 & w2069;
assign w2071 = ~pi86 & ~w2069;
assign w2072 = ~w2070 & ~w2071;
assign w2073 = w2068 & w2072;
assign w2074 = ~w2068 & ~w2072;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = w2067 & w2075;
assign w2077 = ~w2067 & ~w2075;
assign w2078 = ~w2076 & ~w2077;
assign w2079 = pi18 & pi36;
assign w2080 = pi20 & pi34;
assign w2081 = ~w1857 & ~w2080;
assign w2082 = pi20 & pi35;
assign w2083 = w1855 & w2082;
assign w2084 = ~w2081 & ~w2083;
assign w2085 = w2079 & ~w2084;
assign w2086 = ~w2079 & w2084;
assign w2087 = ~w2085 & ~w2086;
assign w2088 = w2078 & ~w2087;
assign w2089 = ~w2078 & w2087;
assign w2090 = ~w2088 & ~w2089;
assign w2091 = (~w1913 & ~w1915) | (~w1913 & w8600) | (~w1915 & w8600);
assign w2092 = w1916 & ~w1918;
assign w2093 = ~w1920 & ~w2092;
assign w2094 = w1904 & ~w1906;
assign w2095 = ~w1908 & ~w2094;
assign w2096 = w2093 & w2095;
assign w2097 = ~w2093 & ~w2095;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = w2091 & ~w2098;
assign w2100 = ~w2091 & w2098;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = (~w1851 & ~w1853) | (~w1851 & w8601) | (~w1853 & w8601);
assign w2103 = ~w1845 & ~w1848;
assign w2104 = w1854 & ~w1856;
assign w2105 = ~w1858 & ~w2104;
assign w2106 = ~w2103 & ~w2105;
assign w2107 = w2103 & w2105;
assign w2108 = ~w2106 & ~w2107;
assign w2109 = w2102 & ~w2108;
assign w2110 = ~w2102 & w2108;
assign w2111 = ~w2109 & ~w2110;
assign w2112 = ~w2101 & ~w2111;
assign w2113 = w2101 & w2111;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = w2090 & ~w2114;
assign w2116 = ~w2090 & w2114;
assign w2117 = ~w2115 & ~w2116;
assign w2118 = w2066 & ~w2117;
assign w2119 = ~w2066 & w2117;
assign w2120 = ~w2118 & ~w2119;
assign w2121 = pi09 & pi45;
assign w2122 = ~w1940 & ~w2121;
assign w2123 = pi09 & pi46;
assign w2124 = w1937 & w2123;
assign w2125 = ~w2122 & ~w2124;
assign w2126 = ~w1967 & ~w1970;
assign w2127 = w2125 & ~w2126;
assign w2128 = ~w2125 & w2126;
assign w2129 = ~w2127 & ~w2128;
assign w2130 = (w2129 & w1979) | (w2129 & w9263) | (w1979 & w9263);
assign w2131 = ~w1979 & w9264;
assign w2132 = ~w2130 & ~w2131;
assign w2133 = w2120 & w2132;
assign w2134 = ~w2120 & ~w2132;
assign w2135 = ~w2133 & ~w2134;
assign w2136 = (~w1875 & w1899) | (~w1875 & w8705) | (w1899 & w8705);
assign w2137 = ~w1870 & ~w1872;
assign w2138 = ~w2137 & w9296;
assign w2139 = (w1896 & w9265) | (w1896 & w9266) | (w9265 & w9266);
assign w2140 = ~w2138 & ~w2139;
assign w2141 = ~w2136 & w2140;
assign w2142 = w2136 & ~w2140;
assign w2143 = ~w2141 & ~w2142;
assign w2144 = ~w1946 & ~w1959;
assign w2145 = w1949 & ~w1952;
assign w2146 = ~w1954 & ~w2145;
assign w2147 = w1803 & ~w1939;
assign w2148 = ~w1941 & ~w2147;
assign w2149 = ~w2146 & ~w2148;
assign w2150 = w2146 & w2148;
assign w2151 = ~w2149 & ~w2150;
assign w2152 = ~w2144 & w2151;
assign w2153 = w2144 & ~w2151;
assign w2154 = ~w2152 & ~w2153;
assign w2155 = pi06 & pi48;
assign w2156 = pi07 & pi47;
assign w2157 = ~w2155 & ~w2156;
assign w2158 = pi07 & pi48;
assign w2159 = w1803 & w2158;
assign w2160 = ~w2157 & ~w2159;
assign w2161 = w1953 & ~w2160;
assign w2162 = ~w1953 & w2160;
assign w2163 = ~w2161 & ~w2162;
assign w2164 = w1869 & ~w2163;
assign w2165 = ~w1869 & w2163;
assign w2166 = ~w2164 & ~w2165;
assign w2167 = pi02 & pi52;
assign w2168 = pi03 & pi51;
assign w2169 = pi04 & pi50;
assign w2170 = ~w2168 & ~w2169;
assign w2171 = pi04 & pi51;
assign w2172 = w1949 & w2171;
assign w2173 = ~w2170 & ~w2172;
assign w2174 = w2167 & ~w2173;
assign w2175 = ~w2167 & w2173;
assign w2176 = ~w2174 & ~w2175;
assign w2177 = w2166 & ~w2176;
assign w2178 = ~w2166 & w2176;
assign w2179 = ~w2177 & ~w2178;
assign w2180 = w2154 & w2179;
assign w2181 = ~w2154 & ~w2179;
assign w2182 = ~w2180 & ~w2181;
assign w2183 = w2143 & ~w2182;
assign w2184 = ~w2143 & w2182;
assign w2185 = ~w2183 & ~w2184;
assign w2186 = w2135 & ~w2185;
assign w2187 = ~w2135 & w2185;
assign w2188 = ~w2186 & ~w2187;
assign w2189 = ~w2025 & w2188;
assign w2190 = w2025 & ~w2188;
assign w2191 = ~w2189 & ~w2190;
assign w2192 = w2024 & w2191;
assign w2193 = ~w2024 & ~w2191;
assign w2194 = ~w2192 & ~w2193;
assign w2195 = ~w2015 & w2194;
assign w2196 = w2015 & ~w2194;
assign w2197 = ~w2195 & ~w2196;
assign w2198 = ~w2008 & ~w2012;
assign w2199 = ~w2197 & ~w2198;
assign w2200 = ~w2008 & w2197;
assign w2201 = ~w1835 & ~w2009;
assign w2202 = w2200 & ~w2201;
assign w2203 = w2197 & w9267;
assign w2204 = ~w1673 & w2203;
assign w2205 = ~w2202 & ~w2204;
assign w2206 = ~w2199 & w2205;
assign w2207 = ~w2195 & w2205;
assign w2208 = ~w2149 & ~w2152;
assign w2209 = pi08 & pi47;
assign w2210 = pi10 & pi45;
assign w2211 = ~w2123 & ~w2210;
assign w2212 = pi10 & pi46;
assign w2213 = w2121 & w2212;
assign w2214 = ~w2211 & ~w2213;
assign w2215 = w2209 & w2214;
assign w2216 = ~w2209 & ~w2214;
assign w2217 = ~w2215 & ~w2216;
assign w2218 = w2158 & w2217;
assign w2219 = ~w2158 & ~w2217;
assign w2220 = ~w2218 & ~w2219;
assign w2221 = ~w2208 & w2220;
assign w2222 = w2208 & ~w2220;
assign w2223 = ~w2221 & ~w2222;
assign w2224 = ~w2138 & w2223;
assign w2225 = ~w2141 & w2224;
assign w2226 = w2136 & ~w2138;
assign w2227 = ~w2139 & ~w2223;
assign w2228 = ~w2226 & w2227;
assign w2229 = ~w2225 & ~w2228;
assign w2230 = pi18 & pi37;
assign w2231 = pi22 & pi33;
assign w2232 = pi23 & pi32;
assign w2233 = pi87 & w2232;
assign w2234 = ~pi87 & ~w2232;
assign w2235 = ~w2233 & ~w2234;
assign w2236 = w2231 & w2235;
assign w2237 = ~w2231 & ~w2235;
assign w2238 = ~w2236 & ~w2237;
assign w2239 = w2230 & w2238;
assign w2240 = ~w2230 & ~w2238;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = pi19 & pi36;
assign w2243 = pi21 & pi34;
assign w2244 = ~w2082 & ~w2243;
assign w2245 = pi21 & pi35;
assign w2246 = w2080 & w2245;
assign w2247 = ~w2244 & ~w2246;
assign w2248 = w2242 & ~w2247;
assign w2249 = ~w2242 & w2247;
assign w2250 = ~w2248 & ~w2249;
assign w2251 = w2241 & ~w2250;
assign w2252 = ~w2241 & w2250;
assign w2253 = ~w2251 & ~w2252;
assign w2254 = (~w2049 & ~w2051) | (~w2049 & w8602) | (~w2051 & w8602);
assign w2255 = w2052 & ~w2054;
assign w2256 = ~w2056 & ~w2255;
assign w2257 = w2040 & ~w2042;
assign w2258 = ~w2044 & ~w2257;
assign w2259 = ~w2256 & ~w2258;
assign w2260 = w2256 & w2258;
assign w2261 = ~w2259 & ~w2260;
assign w2262 = w2254 & ~w2261;
assign w2263 = ~w2254 & w2261;
assign w2264 = ~w2262 & ~w2263;
assign w2265 = w2124 & w2264;
assign w2266 = ~w2124 & ~w2264;
assign w2267 = ~w2265 & ~w2266;
assign w2268 = w2253 & w2267;
assign w2269 = ~w2253 & ~w2267;
assign w2270 = ~w2268 & ~w2269;
assign w2271 = pi11 & pi44;
assign w2272 = pi15 & pi40;
assign w2273 = pi17 & pi38;
assign w2274 = ~w2043 & ~w2273;
assign w2275 = pi17 & pi39;
assign w2276 = w2041 & w2275;
assign w2277 = ~w2274 & ~w2276;
assign w2278 = w2272 & ~w2277;
assign w2279 = ~w2272 & w2277;
assign w2280 = ~w2278 & ~w2279;
assign w2281 = w2271 & ~w2280;
assign w2282 = ~w2271 & w2280;
assign w2283 = ~w2281 & ~w2282;
assign w2284 = pi12 & pi43;
assign w2285 = pi14 & pi41;
assign w2286 = ~w2055 & ~w2285;
assign w2287 = pi14 & pi42;
assign w2288 = w2053 & w2287;
assign w2289 = ~w2286 & ~w2288;
assign w2290 = w2284 & ~w2289;
assign w2291 = ~w2284 & w2289;
assign w2292 = ~w2290 & ~w2291;
assign w2293 = w2283 & ~w2292;
assign w2294 = ~w2283 & w2292;
assign w2295 = ~w2293 & ~w2294;
assign w2296 = (~w2097 & w2091) | (~w2097 & w8707) | (w2091 & w8707);
assign w2297 = (~w2106 & w2102) | (~w2106 & w8708) | (w2102 & w8708);
assign w2298 = ~w2296 & ~w2297;
assign w2299 = w2296 & w2297;
assign w2300 = ~w2298 & ~w2299;
assign w2301 = (~w2076 & ~w2078) | (~w2076 & w8603) | (~w2078 & w8603);
assign w2302 = ~w2070 & ~w2073;
assign w2303 = w2079 & ~w2081;
assign w2304 = ~w2083 & ~w2303;
assign w2305 = ~w2302 & ~w2304;
assign w2306 = w2302 & w2304;
assign w2307 = ~w2305 & ~w2306;
assign w2308 = w2301 & ~w2307;
assign w2309 = ~w2301 & w2307;
assign w2310 = ~w2308 & ~w2309;
assign w2311 = w2300 & w2310;
assign w2312 = ~w2300 & ~w2310;
assign w2313 = ~w2311 & ~w2312;
assign w2314 = ~w2295 & ~w2313;
assign w2315 = w2295 & w2313;
assign w2316 = ~w2314 & ~w2315;
assign w2317 = w2270 & ~w2316;
assign w2318 = ~w2270 & w2316;
assign w2319 = ~w2317 & ~w2318;
assign w2320 = ~w2229 & ~w2319;
assign w2321 = w2229 & w2319;
assign w2322 = ~w2320 & ~w2321;
assign w2323 = ~w2064 & ~w2118;
assign w2324 = (~w2112 & ~w2114) | (~w2112 & w8709) | (~w2114 & w8709);
assign w2325 = w1881 & ~w2031;
assign w2326 = w2027 & ~w2035;
assign w2327 = ~w2325 & ~w2326;
assign w2328 = w2324 & ~w2327;
assign w2329 = ~w2324 & w2327;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = ~w2323 & w2330;
assign w2332 = w2323 & ~w2330;
assign w2333 = ~w2331 & ~w2332;
assign w2334 = pi00 & pi55;
assign w2335 = pi05 & pi50;
assign w2336 = pi06 & pi49;
assign w2337 = ~w2335 & ~w2336;
assign w2338 = pi06 & pi50;
assign w2339 = w1953 & w2338;
assign w2340 = ~w2337 & ~w2339;
assign w2341 = w2171 & ~w2340;
assign w2342 = ~w2171 & w2340;
assign w2343 = ~w2341 & ~w2342;
assign w2344 = w2334 & ~w2343;
assign w2345 = ~w2334 & w2343;
assign w2346 = ~w2344 & ~w2345;
assign w2347 = pi01 & pi54;
assign w2348 = pi02 & pi53;
assign w2349 = pi03 & pi52;
assign w2350 = ~w2348 & ~w2349;
assign w2351 = pi03 & pi53;
assign w2352 = w2167 & w2351;
assign w2353 = ~w2350 & ~w2352;
assign w2354 = w2347 & ~w2353;
assign w2355 = ~w2347 & w2353;
assign w2356 = ~w2354 & ~w2355;
assign w2357 = w2346 & ~w2356;
assign w2358 = ~w2346 & w2356;
assign w2359 = ~w2357 & ~w2358;
assign w2360 = ~w2164 & ~w2177;
assign w2361 = w2167 & ~w2170;
assign w2362 = ~w2172 & ~w2361;
assign w2363 = w1953 & ~w2157;
assign w2364 = ~w2159 & ~w2363;
assign w2365 = ~w2362 & ~w2364;
assign w2366 = w2362 & w2364;
assign w2367 = ~w2365 & ~w2366;
assign w2368 = ~w2360 & w2367;
assign w2369 = w2360 & ~w2367;
assign w2370 = ~w2368 & ~w2369;
assign w2371 = w2359 & w2370;
assign w2372 = ~w2359 & ~w2370;
assign w2373 = ~w2371 & ~w2372;
assign w2374 = w2333 & ~w2373;
assign w2375 = ~w2333 & w2373;
assign w2376 = ~w2374 & ~w2375;
assign w2377 = w2322 & ~w2376;
assign w2378 = ~w2322 & w2376;
assign w2379 = ~w2377 & ~w2378;
assign w2380 = ~w2019 & ~w2022;
assign w2381 = ~w2133 & ~w2186;
assign w2382 = ~w2127 & ~w2130;
assign w2383 = ~w2181 & ~w2184;
assign w2384 = ~w2382 & w2383;
assign w2385 = w2382 & ~w2383;
assign w2386 = ~w2384 & ~w2385;
assign w2387 = w2381 & ~w2386;
assign w2388 = ~w2381 & w2386;
assign w2389 = ~w2387 & ~w2388;
assign w2390 = ~w2380 & w2389;
assign w2391 = w2380 & ~w2389;
assign w2392 = ~w2390 & ~w2391;
assign w2393 = w2379 & w2392;
assign w2394 = ~w2379 & ~w2392;
assign w2395 = ~w2393 & ~w2394;
assign w2396 = ~w2189 & ~w2192;
assign w2397 = w2395 & ~w2396;
assign w2398 = ~w2395 & w2396;
assign w2399 = ~w2397 & ~w2398;
assign w2400 = w2207 & w2399;
assign w2401 = ~w2207 & ~w2399;
assign w2402 = ~w2400 & ~w2401;
assign w2403 = ~w2195 & ~w2397;
assign w2404 = ~w2204 & w9268;
assign w2405 = ~w2398 & ~w2404;
assign w2406 = ~w2390 & ~w2393;
assign w2407 = ~w2365 & ~w2368;
assign w2408 = pi08 & pi48;
assign w2409 = pi07 & pi49;
assign w2410 = ~w2408 & ~w2409;
assign w2411 = pi08 & pi49;
assign w2412 = w2158 & w2411;
assign w2413 = ~w2410 & ~w2412;
assign w2414 = pi09 & pi47;
assign w2415 = pi11 & pi45;
assign w2416 = ~w2212 & ~w2415;
assign w2417 = pi11 & pi46;
assign w2418 = w2210 & w2417;
assign w2419 = ~w2416 & ~w2418;
assign w2420 = w2414 & ~w2419;
assign w2421 = ~w2414 & w2419;
assign w2422 = ~w2420 & ~w2421;
assign w2423 = w2413 & ~w2422;
assign w2424 = ~w2413 & w2422;
assign w2425 = ~w2423 & ~w2424;
assign w2426 = ~w2407 & w2425;
assign w2427 = w2407 & ~w2425;
assign w2428 = ~w2426 & ~w2427;
assign w2429 = ~w2328 & w2428;
assign w2430 = (w2429 & w2323) | (w2429 & w8710) | (w2323 & w8710);
assign w2431 = ~w2118 & w8711;
assign w2432 = ~w2329 & ~w2428;
assign w2433 = ~w2431 & w2432;
assign w2434 = ~w2430 & ~w2433;
assign w2435 = pi19 & pi37;
assign w2436 = pi23 & pi33;
assign w2437 = pi24 & pi32;
assign w2438 = pi88 & w2437;
assign w2439 = ~pi88 & ~w2437;
assign w2440 = ~w2438 & ~w2439;
assign w2441 = w2436 & w2440;
assign w2442 = ~w2436 & ~w2440;
assign w2443 = ~w2441 & ~w2442;
assign w2444 = w2435 & w2443;
assign w2445 = ~w2435 & ~w2443;
assign w2446 = ~w2444 & ~w2445;
assign w2447 = pi20 & pi36;
assign w2448 = pi22 & pi34;
assign w2449 = ~w2245 & ~w2448;
assign w2450 = pi22 & pi35;
assign w2451 = w2243 & w2450;
assign w2452 = ~w2449 & ~w2451;
assign w2453 = w2447 & ~w2452;
assign w2454 = ~w2447 & w2452;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = w2446 & ~w2455;
assign w2457 = ~w2446 & w2455;
assign w2458 = ~w2456 & ~w2457;
assign w2459 = (~w2281 & ~w2283) | (~w2281 & w8604) | (~w2283 & w8604);
assign w2460 = w2284 & ~w2286;
assign w2461 = ~w2288 & ~w2460;
assign w2462 = w2272 & ~w2274;
assign w2463 = ~w2276 & ~w2462;
assign w2464 = ~w2461 & ~w2463;
assign w2465 = w2461 & w2463;
assign w2466 = ~w2464 & ~w2465;
assign w2467 = ~w2459 & w2466;
assign w2468 = w2459 & ~w2466;
assign w2469 = ~w2467 & ~w2468;
assign w2470 = ~w2213 & ~w2218;
assign w2471 = w2213 & w2218;
assign w2472 = ~w2470 & ~w2471;
assign w2473 = ~w2215 & ~w2472;
assign w2474 = w2469 & ~w2473;
assign w2475 = ~w2469 & w2473;
assign w2476 = ~w2474 & ~w2475;
assign w2477 = w2458 & w2476;
assign w2478 = ~w2458 & ~w2476;
assign w2479 = ~w2477 & ~w2478;
assign w2480 = pi12 & pi44;
assign w2481 = pi16 & pi40;
assign w2482 = pi18 & pi38;
assign w2483 = ~w2275 & ~w2482;
assign w2484 = pi18 & pi39;
assign w2485 = w2273 & w2484;
assign w2486 = ~w2483 & ~w2485;
assign w2487 = w2481 & ~w2486;
assign w2488 = ~w2481 & w2486;
assign w2489 = ~w2487 & ~w2488;
assign w2490 = w2480 & ~w2489;
assign w2491 = ~w2480 & w2489;
assign w2492 = ~w2490 & ~w2491;
assign w2493 = pi13 & pi43;
assign w2494 = pi15 & pi41;
assign w2495 = ~w2287 & ~w2494;
assign w2496 = pi15 & pi42;
assign w2497 = w2285 & w2496;
assign w2498 = ~w2495 & ~w2497;
assign w2499 = w2493 & ~w2498;
assign w2500 = ~w2493 & w2498;
assign w2501 = ~w2499 & ~w2500;
assign w2502 = w2492 & ~w2501;
assign w2503 = ~w2492 & w2501;
assign w2504 = ~w2502 & ~w2503;
assign w2505 = (~w2239 & ~w2241) | (~w2239 & w8605) | (~w2241 & w8605);
assign w2506 = ~w2233 & ~w2236;
assign w2507 = w2242 & ~w2244;
assign w2508 = ~w2246 & ~w2507;
assign w2509 = ~w2506 & ~w2508;
assign w2510 = w2506 & w2508;
assign w2511 = ~w2509 & ~w2510;
assign w2512 = ~w2505 & w2511;
assign w2513 = w2505 & ~w2511;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = (~w2259 & w2254) | (~w2259 & w8712) | (w2254 & w8712);
assign w2516 = (~w2305 & w2301) | (~w2305 & w8713) | (w2301 & w8713);
assign w2517 = ~w2515 & ~w2516;
assign w2518 = w2515 & w2516;
assign w2519 = ~w2517 & ~w2518;
assign w2520 = w2514 & w2519;
assign w2521 = ~w2514 & ~w2519;
assign w2522 = ~w2520 & ~w2521;
assign w2523 = ~w2504 & ~w2522;
assign w2524 = w2504 & w2522;
assign w2525 = ~w2523 & ~w2524;
assign w2526 = w2479 & ~w2525;
assign w2527 = ~w2479 & w2525;
assign w2528 = ~w2526 & ~w2527;
assign w2529 = ~w2434 & ~w2528;
assign w2530 = w2434 & w2528;
assign w2531 = ~w2529 & ~w2530;
assign w2532 = ~w2265 & ~w2268;
assign w2533 = ~w2298 & ~w2311;
assign w2534 = ~w2532 & ~w2533;
assign w2535 = w2532 & w2533;
assign w2536 = ~w2534 & ~w2535;
assign w2537 = w2270 & ~w2314;
assign w2538 = ~w2315 & ~w2537;
assign w2539 = w2536 & ~w2538;
assign w2540 = ~w2536 & w2538;
assign w2541 = ~w2539 & ~w2540;
assign w2542 = ~w2344 & ~w2357;
assign w2543 = w2347 & ~w2350;
assign w2544 = ~w2352 & ~w2543;
assign w2545 = w2171 & ~w2337;
assign w2546 = ~w2339 & ~w2545;
assign w2547 = ~w2544 & ~w2546;
assign w2548 = w2544 & w2546;
assign w2549 = ~w2547 & ~w2548;
assign w2550 = ~w2542 & w2549;
assign w2551 = w2542 & ~w2549;
assign w2552 = ~w2550 & ~w2551;
assign w2553 = pi00 & pi56;
assign w2554 = pi04 & pi52;
assign w2555 = pi05 & pi51;
assign w2556 = ~w2338 & ~w2555;
assign w2557 = pi06 & pi51;
assign w2558 = w2335 & w2557;
assign w2559 = ~w2556 & ~w2558;
assign w2560 = w2554 & ~w2559;
assign w2561 = ~w2554 & w2559;
assign w2562 = ~w2560 & ~w2561;
assign w2563 = w2553 & ~w2562;
assign w2564 = ~w2553 & w2562;
assign w2565 = ~w2563 & ~w2564;
assign w2566 = pi01 & pi55;
assign w2567 = pi02 & pi54;
assign w2568 = ~w2351 & ~w2567;
assign w2569 = pi03 & pi54;
assign w2570 = w2348 & w2569;
assign w2571 = ~w2568 & ~w2570;
assign w2572 = w2566 & ~w2571;
assign w2573 = ~w2566 & w2571;
assign w2574 = ~w2572 & ~w2573;
assign w2575 = w2565 & ~w2574;
assign w2576 = ~w2565 & w2574;
assign w2577 = ~w2575 & ~w2576;
assign w2578 = w2552 & w2577;
assign w2579 = ~w2552 & ~w2577;
assign w2580 = ~w2578 & ~w2579;
assign w2581 = w2541 & w2580;
assign w2582 = ~w2541 & ~w2580;
assign w2583 = ~w2581 & ~w2582;
assign w2584 = w2531 & w2583;
assign w2585 = ~w2531 & ~w2583;
assign w2586 = ~w2584 & ~w2585;
assign w2587 = ~w2320 & ~w2377;
assign w2588 = ~w2372 & ~w2375;
assign w2589 = ~w2222 & ~w2225;
assign w2590 = w2588 & w2589;
assign w2591 = ~w2588 & ~w2589;
assign w2592 = ~w2590 & ~w2591;
assign w2593 = ~w2587 & w2592;
assign w2594 = w2587 & ~w2592;
assign w2595 = ~w2593 & ~w2594;
assign w2596 = ~w2384 & ~w2388;
assign w2597 = w2595 & ~w2596;
assign w2598 = ~w2595 & w2596;
assign w2599 = ~w2597 & ~w2598;
assign w2600 = w2586 & w2599;
assign w2601 = ~w2586 & ~w2599;
assign w2602 = ~w2600 & ~w2601;
assign w2603 = ~w2406 & w2602;
assign w2604 = w2406 & ~w2602;
assign w2605 = ~w2603 & ~w2604;
assign w2606 = w2405 & w2605;
assign w2607 = ~w2405 & ~w2605;
assign w2608 = ~w2606 & ~w2607;
assign w2609 = ~w2597 & ~w2600;
assign w2610 = ~w2474 & ~w2477;
assign w2611 = ~w2517 & ~w2520;
assign w2612 = ~w2610 & ~w2611;
assign w2613 = w2610 & w2611;
assign w2614 = ~w2612 & ~w2613;
assign w2615 = w2479 & ~w2523;
assign w2616 = ~w2524 & ~w2615;
assign w2617 = w2614 & ~w2616;
assign w2618 = ~w2614 & w2616;
assign w2619 = ~w2617 & ~w2618;
assign w2620 = (~w2509 & w2505) | (~w2509 & w8714) | (w2505 & w8714);
assign w2621 = pi05 & pi52;
assign w2622 = pi04 & pi53;
assign w2623 = ~w2621 & ~w2622;
assign w2624 = pi05 & pi53;
assign w2625 = w2554 & w2624;
assign w2626 = ~w2623 & ~w2625;
assign w2627 = w2569 & ~w2626;
assign w2628 = ~w2569 & w2626;
assign w2629 = ~w2627 & ~w2628;
assign w2630 = ~w2620 & ~w2629;
assign w2631 = w2620 & w2629;
assign w2632 = ~w2630 & ~w2631;
assign w2633 = pi00 & pi57;
assign w2634 = pi01 & pi56;
assign w2635 = pi02 & pi55;
assign w2636 = ~w2634 & ~w2635;
assign w2637 = pi02 & pi56;
assign w2638 = w2566 & w2637;
assign w2639 = ~w2636 & ~w2638;
assign w2640 = w2633 & ~w2639;
assign w2641 = ~w2633 & w2639;
assign w2642 = ~w2640 & ~w2641;
assign w2643 = w2632 & ~w2642;
assign w2644 = ~w2632 & w2642;
assign w2645 = ~w2643 & ~w2644;
assign w2646 = ~w2563 & ~w2575;
assign w2647 = w2566 & ~w2568;
assign w2648 = ~w2570 & ~w2647;
assign w2649 = w2554 & ~w2556;
assign w2650 = ~w2558 & ~w2649;
assign w2651 = ~w2648 & ~w2650;
assign w2652 = w2648 & w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = ~w2646 & w2653;
assign w2655 = w2646 & ~w2653;
assign w2656 = ~w2654 & ~w2655;
assign w2657 = w2645 & w2656;
assign w2658 = ~w2645 & ~w2656;
assign w2659 = ~w2657 & ~w2658;
assign w2660 = w2619 & ~w2659;
assign w2661 = ~w2619 & w2659;
assign w2662 = ~w2660 & ~w2661;
assign w2663 = ~w2534 & ~w2539;
assign w2664 = ~w2547 & ~w2550;
assign w2665 = pi10 & pi47;
assign w2666 = pi12 & pi45;
assign w2667 = ~w2417 & ~w2666;
assign w2668 = pi12 & pi46;
assign w2669 = w2415 & w2668;
assign w2670 = ~w2667 & ~w2669;
assign w2671 = w2665 & ~w2670;
assign w2672 = ~w2665 & w2670;
assign w2673 = ~w2671 & ~w2672;
assign w2674 = w2557 & ~w2673;
assign w2675 = ~w2557 & w2673;
assign w2676 = ~w2674 & ~w2675;
assign w2677 = pi07 & pi50;
assign w2678 = pi09 & pi48;
assign w2679 = ~w2411 & ~w2678;
assign w2680 = pi09 & pi49;
assign w2681 = w2408 & w2680;
assign w2682 = ~w2679 & ~w2681;
assign w2683 = w2677 & ~w2682;
assign w2684 = ~w2677 & w2682;
assign w2685 = ~w2683 & ~w2684;
assign w2686 = w2676 & ~w2685;
assign w2687 = ~w2676 & w2685;
assign w2688 = ~w2686 & ~w2687;
assign w2689 = ~w2664 & w2688;
assign w2690 = w2664 & ~w2688;
assign w2691 = ~w2689 & ~w2690;
assign w2692 = pi13 & pi44;
assign w2693 = pi17 & pi40;
assign w2694 = pi19 & pi38;
assign w2695 = ~w2484 & ~w2694;
assign w2696 = pi19 & pi39;
assign w2697 = w2482 & w2696;
assign w2698 = ~w2695 & ~w2697;
assign w2699 = w2693 & ~w2698;
assign w2700 = ~w2693 & w2698;
assign w2701 = ~w2699 & ~w2700;
assign w2702 = w2692 & ~w2701;
assign w2703 = ~w2692 & w2701;
assign w2704 = ~w2702 & ~w2703;
assign w2705 = pi14 & pi43;
assign w2706 = pi16 & pi41;
assign w2707 = ~w2496 & ~w2706;
assign w2708 = pi16 & pi42;
assign w2709 = w2494 & w2708;
assign w2710 = ~w2707 & ~w2709;
assign w2711 = w2705 & ~w2710;
assign w2712 = ~w2705 & w2710;
assign w2713 = ~w2711 & ~w2712;
assign w2714 = w2704 & ~w2713;
assign w2715 = ~w2704 & w2713;
assign w2716 = ~w2714 & ~w2715;
assign w2717 = ~w2464 & w2471;
assign w2718 = ~w2467 & w2717;
assign w2719 = (~w2465 & w2293) | (~w2465 & w8606) | (w2293 & w8606);
assign w2720 = (w2293 & w8715) | (w2293 & w8716) | (w8715 & w8716);
assign w2721 = ~w2718 & ~w2720;
assign w2722 = (~w2444 & ~w2446) | (~w2444 & w8717) | (~w2446 & w8717);
assign w2723 = ~w2438 & ~w2441;
assign w2724 = w2447 & ~w2449;
assign w2725 = ~w2451 & ~w2724;
assign w2726 = ~w2723 & ~w2725;
assign w2727 = w2723 & w2725;
assign w2728 = ~w2726 & ~w2727;
assign w2729 = ~w2722 & w2728;
assign w2730 = w2722 & ~w2728;
assign w2731 = ~w2729 & ~w2730;
assign w2732 = ~w2721 & w2731;
assign w2733 = w2721 & ~w2731;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = w2716 & w2734;
assign w2736 = ~w2716 & ~w2734;
assign w2737 = ~w2735 & ~w2736;
assign w2738 = pi20 & pi37;
assign w2739 = pi24 & pi33;
assign w2740 = pi25 & pi32;
assign w2741 = pi89 & w2740;
assign w2742 = ~pi89 & ~w2740;
assign w2743 = ~w2741 & ~w2742;
assign w2744 = w2739 & w2743;
assign w2745 = ~w2739 & ~w2743;
assign w2746 = ~w2744 & ~w2745;
assign w2747 = w2738 & w2746;
assign w2748 = ~w2738 & ~w2746;
assign w2749 = ~w2747 & ~w2748;
assign w2750 = pi21 & pi36;
assign w2751 = pi23 & pi34;
assign w2752 = ~w2450 & ~w2751;
assign w2753 = pi23 & pi35;
assign w2754 = w2448 & w2753;
assign w2755 = ~w2752 & ~w2754;
assign w2756 = w2750 & ~w2755;
assign w2757 = ~w2750 & w2755;
assign w2758 = ~w2756 & ~w2757;
assign w2759 = w2749 & ~w2758;
assign w2760 = ~w2749 & w2758;
assign w2761 = ~w2759 & ~w2760;
assign w2762 = (~w2412 & w2422) | (~w2412 & w8607) | (w2422 & w8607);
assign w2763 = w2414 & ~w2416;
assign w2764 = ~w2418 & ~w2763;
assign w2765 = ~w2764 & ~w2762;
assign w2766 = w2762 & w2764;
assign w2767 = ~w2765 & ~w2766;
assign w2768 = w2761 & w2767;
assign w2769 = ~w2761 & ~w2767;
assign w2770 = ~w2768 & ~w2769;
assign w2771 = (~w2490 & ~w2492) | (~w2490 & w9125) | (~w2492 & w9125);
assign w2772 = w2493 & ~w2495;
assign w2773 = ~w2497 & ~w2772;
assign w2774 = w2481 & ~w2483;
assign w2775 = ~w2485 & ~w2774;
assign w2776 = ~w2773 & ~w2775;
assign w2777 = w2773 & w2775;
assign w2778 = ~w2776 & ~w2777;
assign w2779 = ~w2771 & w2778;
assign w2780 = w2771 & ~w2778;
assign w2781 = ~w2779 & ~w2780;
assign w2782 = w2770 & ~w2781;
assign w2783 = ~w2770 & w2781;
assign w2784 = ~w2782 & ~w2783;
assign w2785 = w2737 & w2784;
assign w2786 = ~w2737 & ~w2784;
assign w2787 = ~w2785 & ~w2786;
assign w2788 = w2691 & ~w2787;
assign w2789 = ~w2691 & w2787;
assign w2790 = ~w2788 & ~w2789;
assign w2791 = w2663 & w2790;
assign w2792 = ~w2663 & ~w2790;
assign w2793 = ~w2791 & ~w2792;
assign w2794 = ~w2662 & ~w2793;
assign w2795 = w2662 & w2793;
assign w2796 = ~w2794 & ~w2795;
assign w2797 = ~w2590 & ~w2593;
assign w2798 = ~w2529 & ~w2584;
assign w2799 = ~w2427 & ~w2430;
assign w2800 = ~w2578 & ~w2581;
assign w2801 = w2799 & ~w2800;
assign w2802 = ~w2799 & w2800;
assign w2803 = ~w2801 & ~w2802;
assign w2804 = ~w2798 & w2803;
assign w2805 = w2798 & ~w2803;
assign w2806 = ~w2804 & ~w2805;
assign w2807 = ~w2797 & w2806;
assign w2808 = w2797 & ~w2806;
assign w2809 = ~w2807 & ~w2808;
assign w2810 = w2796 & w2809;
assign w2811 = ~w2796 & ~w2809;
assign w2812 = ~w2810 & ~w2811;
assign w2813 = w2609 & ~w2812;
assign w2814 = ~w2609 & w2812;
assign w2815 = ~w2813 & ~w2814;
assign w2816 = ~w2603 & ~w2606;
assign w2817 = w2815 & ~w2816;
assign w2818 = ~w2815 & w2816;
assign w2819 = ~w2817 & ~w2818;
assign w2820 = ~w2807 & ~w2810;
assign w2821 = w2471 & w2719;
assign w2822 = ~w2732 & ~w2821;
assign w2823 = ~w2769 & ~w2782;
assign w2824 = ~w2822 & w2823;
assign w2825 = w2822 & ~w2823;
assign w2826 = ~w2824 & ~w2825;
assign w2827 = ~w2736 & ~w2784;
assign w2828 = ~w2735 & ~w2827;
assign w2829 = w2826 & ~w2828;
assign w2830 = ~w2826 & w2828;
assign w2831 = ~w2829 & ~w2830;
assign w2832 = ~w2630 & ~w2643;
assign w2833 = w2633 & ~w2636;
assign w2834 = ~w2638 & ~w2833;
assign w2835 = w2569 & ~w2623;
assign w2836 = ~w2625 & ~w2835;
assign w2837 = ~w2834 & ~w2836;
assign w2838 = w2834 & w2836;
assign w2839 = ~w2837 & ~w2838;
assign w2840 = ~w2832 & w2839;
assign w2841 = w2832 & ~w2839;
assign w2842 = ~w2840 & ~w2841;
assign w2843 = ~w2776 & ~w2779;
assign w2844 = pi03 & pi55;
assign w2845 = pi04 & pi54;
assign w2846 = ~w2844 & ~w2845;
assign w2847 = pi04 & pi55;
assign w2848 = w2569 & w2847;
assign w2849 = ~w2846 & ~w2848;
assign w2850 = w2637 & ~w2849;
assign w2851 = ~w2637 & w2849;
assign w2852 = ~w2850 & ~w2851;
assign w2853 = ~w2843 & ~w2852;
assign w2854 = w2843 & w2852;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = pi00 & pi58;
assign w2857 = pi01 & pi57;
assign w2858 = ~w2856 & ~w2857;
assign w2859 = pi01 & pi58;
assign w2860 = w2633 & w2859;
assign w2861 = ~w2858 & ~w2860;
assign w2862 = ~w2726 & ~w2729;
assign w2863 = w2861 & ~w2862;
assign w2864 = ~w2861 & w2862;
assign w2865 = ~w2863 & ~w2864;
assign w2866 = w2855 & w2865;
assign w2867 = ~w2855 & ~w2865;
assign w2868 = ~w2866 & ~w2867;
assign w2869 = w2842 & w2868;
assign w2870 = ~w2842 & ~w2868;
assign w2871 = ~w2869 & ~w2870;
assign w2872 = w2831 & w2871;
assign w2873 = ~w2831 & ~w2871;
assign w2874 = ~w2872 & ~w2873;
assign w2875 = ~w2612 & ~w2617;
assign w2876 = pi06 & pi52;
assign w2877 = ~w2624 & ~w2876;
assign w2878 = pi06 & pi53;
assign w2879 = w2621 & w2878;
assign w2880 = ~w2877 & ~w2879;
assign w2881 = ~w2651 & ~w2654;
assign w2882 = w2880 & ~w2881;
assign w2883 = ~w2880 & w2881;
assign w2884 = ~w2882 & ~w2883;
assign w2885 = pi07 & pi51;
assign w2886 = pi11 & pi47;
assign w2887 = pi13 & pi45;
assign w2888 = ~w2668 & ~w2887;
assign w2889 = pi13 & pi46;
assign w2890 = w2666 & w2889;
assign w2891 = ~w2888 & ~w2890;
assign w2892 = w2886 & ~w2891;
assign w2893 = ~w2886 & w2891;
assign w2894 = ~w2892 & ~w2893;
assign w2895 = w2885 & ~w2894;
assign w2896 = ~w2885 & w2894;
assign w2897 = ~w2895 & ~w2896;
assign w2898 = pi08 & pi50;
assign w2899 = pi10 & pi48;
assign w2900 = ~w2680 & ~w2899;
assign w2901 = pi10 & pi49;
assign w2902 = w2678 & w2901;
assign w2903 = ~w2900 & ~w2902;
assign w2904 = w2898 & ~w2903;
assign w2905 = ~w2898 & w2903;
assign w2906 = ~w2904 & ~w2905;
assign w2907 = w2897 & ~w2906;
assign w2908 = ~w2897 & w2906;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = (~w2702 & ~w2704) | (~w2702 & w8718) | (~w2704 & w8718);
assign w2911 = w2705 & ~w2707;
assign w2912 = ~w2709 & ~w2911;
assign w2913 = w2693 & ~w2695;
assign w2914 = ~w2697 & ~w2913;
assign w2915 = ~w2912 & ~w2914;
assign w2916 = w2912 & w2914;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = ~w2910 & w2917;
assign w2919 = w2910 & ~w2917;
assign w2920 = ~w2918 & ~w2919;
assign w2921 = (~w2747 & ~w2749) | (~w2747 & w8608) | (~w2749 & w8608);
assign w2922 = (~w2741 & ~w2743) | (~w2741 & w8719) | (~w2743 & w8719);
assign w2923 = w2750 & ~w2752;
assign w2924 = ~w2754 & ~w2923;
assign w2925 = ~w2922 & ~w2924;
assign w2926 = w2922 & w2924;
assign w2927 = ~w2925 & ~w2926;
assign w2928 = w2765 & ~w2927;
assign w2929 = ~w2765 & w2927;
assign w2930 = ~w2928 & ~w2929;
assign w2931 = w2921 & ~w2930;
assign w2932 = ~w2921 & w2930;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = w2920 & ~w2933;
assign w2935 = ~w2920 & w2933;
assign w2936 = ~w2934 & ~w2935;
assign w2937 = ~w2909 & ~w2936;
assign w2938 = w2909 & w2936;
assign w2939 = ~w2937 & ~w2938;
assign w2940 = pi14 & pi44;
assign w2941 = pi18 & pi40;
assign w2942 = pi20 & pi38;
assign w2943 = ~w2696 & ~w2942;
assign w2944 = pi20 & pi39;
assign w2945 = w2694 & w2944;
assign w2946 = ~w2943 & ~w2945;
assign w2947 = w2941 & ~w2946;
assign w2948 = ~w2941 & w2946;
assign w2949 = ~w2947 & ~w2948;
assign w2950 = w2940 & ~w2949;
assign w2951 = ~w2940 & w2949;
assign w2952 = ~w2950 & ~w2951;
assign w2953 = pi15 & pi43;
assign w2954 = pi17 & pi41;
assign w2955 = ~w2708 & ~w2954;
assign w2956 = pi17 & pi42;
assign w2957 = w2706 & w2956;
assign w2958 = ~w2955 & ~w2957;
assign w2959 = w2953 & ~w2958;
assign w2960 = ~w2953 & w2958;
assign w2961 = ~w2959 & ~w2960;
assign w2962 = w2952 & ~w2961;
assign w2963 = ~w2952 & w2961;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = pi21 & pi37;
assign w2966 = pi25 & pi33;
assign w2967 = pi26 & pi32;
assign w2968 = pi90 & w2967;
assign w2969 = ~pi90 & ~w2967;
assign w2970 = ~w2968 & ~w2969;
assign w2971 = w2966 & w2970;
assign w2972 = ~w2966 & ~w2970;
assign w2973 = ~w2971 & ~w2972;
assign w2974 = w2965 & w2973;
assign w2975 = ~w2965 & ~w2973;
assign w2976 = ~w2974 & ~w2975;
assign w2977 = pi22 & pi36;
assign w2978 = pi24 & pi34;
assign w2979 = ~w2753 & ~w2978;
assign w2980 = pi24 & pi35;
assign w2981 = w2751 & w2980;
assign w2982 = ~w2979 & ~w2981;
assign w2983 = w2977 & ~w2982;
assign w2984 = ~w2977 & w2982;
assign w2985 = ~w2983 & ~w2984;
assign w2986 = w2976 & ~w2985;
assign w2987 = ~w2976 & w2985;
assign w2988 = ~w2986 & ~w2987;
assign w2989 = (~w2674 & ~w2676) | (~w2674 & w8720) | (~w2676 & w8720);
assign w2990 = w2677 & ~w2679;
assign w2991 = ~w2681 & ~w2990;
assign w2992 = w2665 & ~w2667;
assign w2993 = ~w2669 & ~w2992;
assign w2994 = ~w2991 & ~w2993;
assign w2995 = w2991 & w2993;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = ~w2989 & w2996;
assign w2998 = w2989 & ~w2996;
assign w2999 = ~w2997 & ~w2998;
assign w3000 = w2988 & w2999;
assign w3001 = ~w2988 & ~w2999;
assign w3002 = ~w3000 & ~w3001;
assign w3003 = w2964 & w3002;
assign w3004 = ~w2964 & ~w3002;
assign w3005 = ~w3003 & ~w3004;
assign w3006 = w2939 & ~w3005;
assign w3007 = ~w2939 & w3005;
assign w3008 = ~w3006 & ~w3007;
assign w3009 = w2884 & ~w3008;
assign w3010 = ~w2884 & w3008;
assign w3011 = ~w3009 & ~w3010;
assign w3012 = w2875 & w3011;
assign w3013 = ~w2875 & ~w3011;
assign w3014 = ~w3012 & ~w3013;
assign w3015 = w2874 & ~w3014;
assign w3016 = ~w2874 & w3014;
assign w3017 = ~w3015 & ~w3016;
assign w3018 = ~w2801 & ~w2804;
assign w3019 = ~w2787 & w2793;
assign w3020 = ~w2794 & ~w3019;
assign w3021 = ~w2658 & ~w2661;
assign w3022 = ~w2663 & ~w2690;
assign w3023 = ~w2689 & ~w3022;
assign w3024 = w3021 & ~w3023;
assign w3025 = ~w3021 & w3023;
assign w3026 = ~w3024 & ~w3025;
assign w3027 = ~w3020 & w3026;
assign w3028 = w3020 & ~w3026;
assign w3029 = ~w3027 & ~w3028;
assign w3030 = ~w3018 & w3029;
assign w3031 = w3018 & ~w3029;
assign w3032 = ~w3030 & ~w3031;
assign w3033 = w3017 & w3032;
assign w3034 = ~w3017 & ~w3032;
assign w3035 = ~w3033 & ~w3034;
assign w3036 = ~w2820 & w3035;
assign w3037 = w2820 & ~w3035;
assign w3038 = ~w3036 & ~w3037;
assign w3039 = ~w2814 & ~w2817;
assign w3040 = w3038 & ~w3039;
assign w3041 = ~w3038 & w3039;
assign w3042 = ~w3040 & ~w3041;
assign w3043 = ~w3036 & ~w3040;
assign w3044 = (~w3030 & ~w3032) | (~w3030 & w8721) | (~w3032 & w8721);
assign w3045 = pi22 & pi37;
assign w3046 = pi26 & pi33;
assign w3047 = pi27 & pi32;
assign w3048 = pi91 & w3047;
assign w3049 = ~pi91 & ~w3047;
assign w3050 = ~w3048 & ~w3049;
assign w3051 = w3046 & w3050;
assign w3052 = ~w3046 & ~w3050;
assign w3053 = ~w3051 & ~w3052;
assign w3054 = w3045 & w3053;
assign w3055 = ~w3045 & ~w3053;
assign w3056 = ~w3054 & ~w3055;
assign w3057 = pi23 & pi36;
assign w3058 = pi25 & pi34;
assign w3059 = ~w2980 & ~w3058;
assign w3060 = pi25 & pi35;
assign w3061 = w2978 & w3060;
assign w3062 = ~w3059 & ~w3061;
assign w3063 = w3057 & ~w3062;
assign w3064 = ~w3057 & w3062;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = w3056 & ~w3065;
assign w3067 = ~w3056 & w3065;
assign w3068 = ~w3066 & ~w3067;
assign w3069 = w2879 & w3068;
assign w3070 = ~w2879 & ~w3068;
assign w3071 = ~w3069 & ~w3070;
assign w3072 = pi15 & pi44;
assign w3073 = pi19 & pi40;
assign w3074 = pi21 & pi38;
assign w3075 = ~w2944 & ~w3074;
assign w3076 = pi21 & pi39;
assign w3077 = w2942 & w3076;
assign w3078 = ~w3075 & ~w3077;
assign w3079 = w3073 & ~w3078;
assign w3080 = ~w3073 & w3078;
assign w3081 = ~w3079 & ~w3080;
assign w3082 = w3072 & ~w3081;
assign w3083 = ~w3072 & w3081;
assign w3084 = ~w3082 & ~w3083;
assign w3085 = pi16 & pi43;
assign w3086 = pi18 & pi41;
assign w3087 = ~w2956 & ~w3086;
assign w3088 = pi18 & pi42;
assign w3089 = w2954 & w3088;
assign w3090 = ~w3087 & ~w3089;
assign w3091 = w3085 & ~w3090;
assign w3092 = ~w3085 & w3090;
assign w3093 = ~w3091 & ~w3092;
assign w3094 = w3084 & ~w3093;
assign w3095 = ~w3084 & w3093;
assign w3096 = ~w3094 & ~w3095;
assign w3097 = w3071 & w3096;
assign w3098 = ~w3071 & ~w3096;
assign w3099 = ~w3097 & ~w3098;
assign w3100 = (~w2895 & ~w2897) | (~w2895 & w8918) | (~w2897 & w8918);
assign w3101 = w2898 & ~w2900;
assign w3102 = ~w2902 & ~w3101;
assign w3103 = w2886 & ~w2888;
assign w3104 = ~w2890 & ~w3103;
assign w3105 = ~w3102 & ~w3104;
assign w3106 = w3102 & w3104;
assign w3107 = ~w3105 & ~w3106;
assign w3108 = ~w3100 & w3107;
assign w3109 = w3100 & ~w3107;
assign w3110 = ~w3108 & ~w3109;
assign w3111 = (~w2950 & ~w2952) | (~w2950 & w8609) | (~w2952 & w8609);
assign w3112 = w2953 & ~w2955;
assign w3113 = ~w2957 & ~w3112;
assign w3114 = w2941 & ~w2943;
assign w3115 = ~w2945 & ~w3114;
assign w3116 = ~w3113 & ~w3115;
assign w3117 = w3113 & w3115;
assign w3118 = ~w3116 & ~w3117;
assign w3119 = ~w3111 & w3118;
assign w3120 = w3111 & ~w3118;
assign w3121 = ~w3119 & ~w3120;
assign w3122 = (~w2974 & ~w2976) | (~w2974 & w8610) | (~w2976 & w8610);
assign w3123 = (~w2968 & ~w2970) | (~w2968 & w8919) | (~w2970 & w8919);
assign w3124 = w2977 & ~w2979;
assign w3125 = ~w2981 & ~w3124;
assign w3126 = ~w3123 & ~w3125;
assign w3127 = w3123 & w3125;
assign w3128 = ~w3126 & ~w3127;
assign w3129 = ~w3122 & w3128;
assign w3130 = w3122 & ~w3128;
assign w3131 = ~w3129 & ~w3130;
assign w3132 = w3121 & w3131;
assign w3133 = ~w3121 & ~w3131;
assign w3134 = ~w3132 & ~w3133;
assign w3135 = w3110 & w3134;
assign w3136 = ~w3110 & ~w3134;
assign w3137 = ~w3135 & ~w3136;
assign w3138 = pi08 & pi51;
assign w3139 = pi12 & pi47;
assign w3140 = pi14 & pi45;
assign w3141 = ~w2889 & ~w3140;
assign w3142 = pi14 & pi46;
assign w3143 = w2887 & w3142;
assign w3144 = ~w3141 & ~w3143;
assign w3145 = w3139 & ~w3144;
assign w3146 = ~w3139 & w3144;
assign w3147 = ~w3145 & ~w3146;
assign w3148 = w3138 & ~w3147;
assign w3149 = ~w3138 & w3147;
assign w3150 = ~w3148 & ~w3149;
assign w3151 = pi09 & pi50;
assign w3152 = pi11 & pi48;
assign w3153 = ~w2901 & ~w3152;
assign w3154 = pi11 & pi49;
assign w3155 = w2899 & w3154;
assign w3156 = ~w3153 & ~w3155;
assign w3157 = w3151 & ~w3156;
assign w3158 = ~w3151 & w3156;
assign w3159 = ~w3157 & ~w3158;
assign w3160 = w3150 & ~w3159;
assign w3161 = ~w3150 & w3159;
assign w3162 = ~w3160 & ~w3161;
assign w3163 = w3137 & w3162;
assign w3164 = ~w3137 & ~w3162;
assign w3165 = ~w3163 & ~w3164;
assign w3166 = w3099 & w3165;
assign w3167 = ~w3099 & ~w3165;
assign w3168 = ~w3166 & ~w3167;
assign w3169 = (~w2824 & w2828) | (~w2824 & w8722) | (w2828 & w8722);
assign w3170 = ~w2837 & ~w2840;
assign w3171 = pi05 & pi54;
assign w3172 = pi07 & pi52;
assign w3173 = ~w2878 & ~w3172;
assign w3174 = pi07 & pi53;
assign w3175 = w2876 & w3174;
assign w3176 = ~w3173 & ~w3175;
assign w3177 = w3171 & w3176;
assign w3178 = ~w3171 & ~w3176;
assign w3179 = ~w3177 & ~w3178;
assign w3180 = w2847 & w3179;
assign w3181 = ~w2847 & ~w3179;
assign w3182 = ~w3180 & ~w3181;
assign w3183 = ~w3170 & w3182;
assign w3184 = w3170 & ~w3182;
assign w3185 = ~w3183 & ~w3184;
assign w3186 = ~w3169 & w3185;
assign w3187 = w3169 & ~w3185;
assign w3188 = ~w3186 & ~w3187;
assign w3189 = w3168 & w3188;
assign w3190 = ~w3168 & ~w3188;
assign w3191 = ~w3189 & ~w3190;
assign w3192 = ~w2853 & ~w2866;
assign w3193 = ~w2860 & ~w2863;
assign w3194 = w2637 & ~w2846;
assign w3195 = ~w2848 & ~w3194;
assign w3196 = ~w3193 & ~w3195;
assign w3197 = w3193 & w3195;
assign w3198 = ~w3196 & ~w3197;
assign w3199 = ~w3192 & w3198;
assign w3200 = w3192 & ~w3198;
assign w3201 = ~w3199 & ~w3200;
assign w3202 = (~w2994 & w2989) | (~w2994 & w9126) | (w2989 & w9126);
assign w3203 = pi02 & pi57;
assign w3204 = pi03 & pi56;
assign w3205 = ~w3203 & ~w3204;
assign w3206 = pi03 & pi57;
assign w3207 = w2637 & w3206;
assign w3208 = ~w3205 & ~w3207;
assign w3209 = w2859 & ~w3208;
assign w3210 = ~w2859 & w3208;
assign w3211 = ~w3209 & ~w3210;
assign w3212 = w3202 & w3211;
assign w3213 = ~w3202 & ~w3211;
assign w3214 = ~w3212 & ~w3213;
assign w3215 = (~w2915 & w2910) | (~w2915 & w9127) | (w2910 & w9127);
assign w3216 = pi00 & pi59;
assign w3217 = w3216 & w9297;
assign w3218 = (w2921 & w8920) | (w2921 & w8921) | (w8920 & w8921);
assign w3219 = ~w3217 & ~w3218;
assign w3220 = ~w3215 & w3219;
assign w3221 = w3215 & ~w3219;
assign w3222 = ~w3220 & ~w3221;
assign w3223 = w3214 & ~w3222;
assign w3224 = ~w3214 & w3222;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = w3201 & ~w3225;
assign w3227 = ~w3201 & w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = ~w2937 & ~w3006;
assign w3230 = w2765 & w2933;
assign w3231 = ~w2934 & ~w3230;
assign w3232 = ~w3000 & ~w3003;
assign w3233 = ~w3231 & ~w3232;
assign w3234 = w3231 & w3232;
assign w3235 = ~w3233 & ~w3234;
assign w3236 = w3229 & w3235;
assign w3237 = ~w3229 & ~w3235;
assign w3238 = ~w3236 & ~w3237;
assign w3239 = w3228 & ~w3238;
assign w3240 = ~w3228 & w3238;
assign w3241 = ~w3239 & ~w3240;
assign w3242 = w3191 & ~w3241;
assign w3243 = ~w3191 & w3241;
assign w3244 = ~w3242 & ~w3243;
assign w3245 = (~w3024 & w3020) | (~w3024 & w8724) | (w3020 & w8724);
assign w3246 = ~w3008 & w3014;
assign w3247 = ~w3015 & ~w3246;
assign w3248 = ~w2869 & ~w2872;
assign w3249 = w2875 & ~w2882;
assign w3250 = ~w2883 & ~w3249;
assign w3251 = ~w3248 & w3250;
assign w3252 = w3248 & ~w3250;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = ~w3247 & w3253;
assign w3255 = w3247 & ~w3253;
assign w3256 = ~w3254 & ~w3255;
assign w3257 = ~w3245 & w3256;
assign w3258 = w3245 & ~w3256;
assign w3259 = ~w3257 & ~w3258;
assign w3260 = w3244 & w3259;
assign w3261 = ~w3244 & ~w3259;
assign w3262 = ~w3260 & ~w3261;
assign w3263 = ~w3044 & w3262;
assign w3264 = w3044 & ~w3262;
assign w3265 = ~w3263 & ~w3264;
assign w3266 = w3043 & w3265;
assign w3267 = ~w3043 & ~w3265;
assign w3268 = ~w3266 & ~w3267;
assign w3269 = ~w2603 & ~w2814;
assign w3270 = ~w2813 & ~w3037;
assign w3271 = ~w3269 & w3270;
assign w3272 = (~w3264 & w3271) | (~w3264 & w8725) | (w3271 & w8725);
assign w3273 = w2605 & w2815;
assign w3274 = w3038 & w3265;
assign w3275 = w3273 & w3274;
assign w3276 = w2405 & w3275;
assign w3277 = ~w3272 & ~w3276;
assign w3278 = ~w3257 & ~w3260;
assign w3279 = (~w3105 & w3100) | (~w3105 & w9128) | (w3100 & w9128);
assign w3280 = pi01 & pi59;
assign w3281 = pi02 & pi58;
assign w3282 = ~w3206 & ~w3281;
assign w3283 = pi03 & pi58;
assign w3284 = w3203 & w3283;
assign w3285 = ~w3282 & ~w3284;
assign w3286 = w3280 & ~w3285;
assign w3287 = ~w3280 & w3285;
assign w3288 = ~w3286 & ~w3287;
assign w3289 = w3279 & w3288;
assign w3290 = ~w3279 & ~w3288;
assign w3291 = ~w3289 & ~w3290;
assign w3292 = (~w3116 & w3111) | (~w3116 & w9129) | (w3111 & w9129);
assign w3293 = pi00 & pi60;
assign w3294 = (~w3122 & w8922) | (~w3122 & w8923) | (w8922 & w8923);
assign w3295 = (w3122 & w8924) | (w3122 & w8925) | (w8924 & w8925);
assign w3296 = ~w3294 & ~w3295;
assign w3297 = ~w3292 & w3296;
assign w3298 = w3292 & ~w3296;
assign w3299 = ~w3297 & ~w3298;
assign w3300 = w3291 & ~w3299;
assign w3301 = ~w3291 & w3299;
assign w3302 = ~w3300 & ~w3301;
assign w3303 = (~w3212 & w3222) | (~w3212 & w9130) | (w3222 & w9130);
assign w3304 = (~w3217 & ~w3219) | (~w3217 & w9131) | (~w3219 & w9131);
assign w3305 = w2859 & ~w3205;
assign w3306 = ~w3207 & ~w3305;
assign w3307 = ~w3304 & ~w3306;
assign w3308 = w3304 & w3306;
assign w3309 = ~w3307 & ~w3308;
assign w3310 = w3303 & w3309;
assign w3311 = ~w3303 & ~w3309;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = (~w3163 & ~w3165) | (~w3163 & w8726) | (~w3165 & w8726);
assign w3314 = ~w3069 & ~w3097;
assign w3315 = (~w3132 & ~w3134) | (~w3132 & w9132) | (~w3134 & w9132);
assign w3316 = ~w3314 & ~w3315;
assign w3317 = w3314 & w3315;
assign w3318 = ~w3316 & ~w3317;
assign w3319 = (w3165 & w9133) | (w3165 & w9134) | (w9133 & w9134);
assign w3320 = ~w3318 & w3313;
assign w3321 = ~w3319 & ~w3320;
assign w3322 = w3312 & w3321;
assign w3323 = ~w3312 & ~w3321;
assign w3324 = ~w3322 & ~w3323;
assign w3325 = ~w3302 & w3324;
assign w3326 = w3302 & ~w3324;
assign w3327 = ~w3325 & ~w3326;
assign w3328 = pi16 & pi44;
assign w3329 = pi20 & pi40;
assign w3330 = pi22 & pi38;
assign w3331 = ~w3076 & ~w3330;
assign w3332 = pi22 & pi39;
assign w3333 = w3074 & w3332;
assign w3334 = ~w3331 & ~w3333;
assign w3335 = w3329 & ~w3334;
assign w3336 = ~w3329 & w3334;
assign w3337 = ~w3335 & ~w3336;
assign w3338 = w3328 & ~w3337;
assign w3339 = ~w3328 & w3337;
assign w3340 = ~w3338 & ~w3339;
assign w3341 = pi17 & pi43;
assign w3342 = pi19 & pi41;
assign w3343 = ~w3088 & ~w3342;
assign w3344 = pi19 & pi42;
assign w3345 = w3086 & w3344;
assign w3346 = ~w3343 & ~w3345;
assign w3347 = w3341 & ~w3346;
assign w3348 = ~w3341 & w3346;
assign w3349 = ~w3347 & ~w3348;
assign w3350 = w3340 & ~w3349;
assign w3351 = ~w3340 & w3349;
assign w3352 = ~w3350 & ~w3351;
assign w3353 = pi23 & pi37;
assign w3354 = pi27 & pi33;
assign w3355 = pi28 & pi32;
assign w3356 = pi92 & w3355;
assign w3357 = ~pi92 & ~w3355;
assign w3358 = ~w3356 & ~w3357;
assign w3359 = w3354 & w3358;
assign w3360 = ~w3354 & ~w3358;
assign w3361 = ~w3359 & ~w3360;
assign w3362 = w3353 & w3361;
assign w3363 = ~w3353 & ~w3361;
assign w3364 = ~w3362 & ~w3363;
assign w3365 = pi24 & pi36;
assign w3366 = pi26 & pi34;
assign w3367 = ~w3060 & ~w3366;
assign w3368 = pi26 & pi35;
assign w3369 = w3058 & w3368;
assign w3370 = ~w3367 & ~w3369;
assign w3371 = w3365 & ~w3370;
assign w3372 = ~w3365 & w3370;
assign w3373 = ~w3371 & ~w3372;
assign w3374 = w3364 & ~w3373;
assign w3375 = ~w3364 & w3373;
assign w3376 = ~w3374 & ~w3375;
assign w3377 = ~w3175 & ~w3180;
assign w3378 = w3175 & w3180;
assign w3379 = ~w3377 & ~w3378;
assign w3380 = ~w3177 & ~w3379;
assign w3381 = w3376 & ~w3380;
assign w3382 = ~w3376 & w3380;
assign w3383 = ~w3381 & ~w3382;
assign w3384 = w3352 & w3383;
assign w3385 = ~w3352 & ~w3383;
assign w3386 = ~w3384 & ~w3385;
assign w3387 = (~w3148 & ~w3150) | (~w3148 & w8926) | (~w3150 & w8926);
assign w3388 = w3151 & ~w3153;
assign w3389 = ~w3155 & ~w3388;
assign w3390 = w3139 & ~w3141;
assign w3391 = ~w3143 & ~w3390;
assign w3392 = ~w3389 & ~w3391;
assign w3393 = w3389 & w3391;
assign w3394 = ~w3392 & ~w3393;
assign w3395 = ~w3387 & w3394;
assign w3396 = w3387 & ~w3394;
assign w3397 = ~w3395 & ~w3396;
assign w3398 = (~w3082 & ~w3084) | (~w3082 & w8611) | (~w3084 & w8611);
assign w3399 = w3085 & ~w3087;
assign w3400 = ~w3089 & ~w3399;
assign w3401 = w3073 & ~w3075;
assign w3402 = ~w3077 & ~w3401;
assign w3403 = ~w3400 & ~w3402;
assign w3404 = w3400 & w3402;
assign w3405 = ~w3403 & ~w3404;
assign w3406 = ~w3398 & w3405;
assign w3407 = w3398 & ~w3405;
assign w3408 = ~w3406 & ~w3407;
assign w3409 = (~w3054 & ~w3056) | (~w3054 & w8612) | (~w3056 & w8612);
assign w3410 = (~w3048 & ~w3050) | (~w3048 & w8927) | (~w3050 & w8927);
assign w3411 = w3057 & ~w3059;
assign w3412 = ~w3061 & ~w3411;
assign w3413 = ~w3410 & ~w3412;
assign w3414 = w3410 & w3412;
assign w3415 = ~w3413 & ~w3414;
assign w3416 = ~w3409 & w3415;
assign w3417 = w3409 & ~w3415;
assign w3418 = ~w3416 & ~w3417;
assign w3419 = w3408 & w3418;
assign w3420 = ~w3408 & ~w3418;
assign w3421 = ~w3419 & ~w3420;
assign w3422 = w3397 & w3421;
assign w3423 = ~w3397 & ~w3421;
assign w3424 = ~w3422 & ~w3423;
assign w3425 = pi09 & pi51;
assign w3426 = pi13 & pi47;
assign w3427 = pi15 & pi45;
assign w3428 = ~w3142 & ~w3427;
assign w3429 = pi15 & pi46;
assign w3430 = w3140 & w3429;
assign w3431 = ~w3428 & ~w3430;
assign w3432 = w3426 & ~w3431;
assign w3433 = ~w3426 & w3431;
assign w3434 = ~w3432 & ~w3433;
assign w3435 = w3425 & ~w3434;
assign w3436 = ~w3425 & w3434;
assign w3437 = ~w3435 & ~w3436;
assign w3438 = pi10 & pi50;
assign w3439 = pi12 & pi48;
assign w3440 = ~w3154 & ~w3439;
assign w3441 = pi12 & pi49;
assign w3442 = w3152 & w3441;
assign w3443 = ~w3440 & ~w3442;
assign w3444 = w3438 & ~w3443;
assign w3445 = ~w3438 & w3443;
assign w3446 = ~w3444 & ~w3445;
assign w3447 = w3437 & ~w3446;
assign w3448 = ~w3437 & w3446;
assign w3449 = ~w3447 & ~w3448;
assign w3450 = w3424 & w3449;
assign w3451 = ~w3424 & ~w3449;
assign w3452 = ~w3450 & ~w3451;
assign w3453 = w3386 & w3452;
assign w3454 = ~w3386 & ~w3452;
assign w3455 = ~w3453 & ~w3454;
assign w3456 = ~w3196 & ~w3199;
assign w3457 = pi05 & pi55;
assign w3458 = pi04 & pi56;
assign w3459 = ~w3457 & ~w3458;
assign w3460 = pi05 & pi56;
assign w3461 = w2847 & w3460;
assign w3462 = ~w3459 & ~w3461;
assign w3463 = pi06 & pi54;
assign w3464 = pi08 & pi52;
assign w3465 = ~w3174 & ~w3464;
assign w3466 = pi08 & pi53;
assign w3467 = w3172 & w3466;
assign w3468 = ~w3465 & ~w3467;
assign w3469 = w3463 & ~w3468;
assign w3470 = ~w3463 & w3468;
assign w3471 = ~w3469 & ~w3470;
assign w3472 = w3462 & ~w3471;
assign w3473 = ~w3462 & w3471;
assign w3474 = ~w3472 & ~w3473;
assign w3475 = ~w3456 & w3474;
assign w3476 = w3456 & ~w3474;
assign w3477 = ~w3475 & ~w3476;
assign w3478 = ~w3233 & ~w3236;
assign w3479 = w3477 & ~w3478;
assign w3480 = ~w3477 & w3478;
assign w3481 = ~w3479 & ~w3480;
assign w3482 = w3455 & w3481;
assign w3483 = ~w3455 & ~w3481;
assign w3484 = ~w3482 & ~w3483;
assign w3485 = w3327 & w3484;
assign w3486 = ~w3327 & ~w3484;
assign w3487 = ~w3485 & ~w3486;
assign w3488 = ~w3251 & ~w3254;
assign w3489 = ~w3183 & ~w3186;
assign w3490 = ~w3227 & ~w3239;
assign w3491 = ~w3489 & w3490;
assign w3492 = w3489 & ~w3490;
assign w3493 = ~w3491 & ~w3492;
assign w3494 = ~w3189 & ~w3242;
assign w3495 = w3493 & ~w3494;
assign w3496 = ~w3493 & w3494;
assign w3497 = ~w3495 & ~w3496;
assign w3498 = ~w3488 & w3497;
assign w3499 = w3488 & ~w3497;
assign w3500 = ~w3498 & ~w3499;
assign w3501 = w3487 & w3500;
assign w3502 = ~w3487 & ~w3500;
assign w3503 = ~w3501 & ~w3502;
assign w3504 = ~w3278 & w3503;
assign w3505 = w3278 & ~w3503;
assign w3506 = ~w3504 & ~w3505;
assign w3507 = ~w3277 & w3506;
assign w3508 = w3277 & ~w3506;
assign w3509 = ~w3507 & ~w3508;
assign w3510 = ~w3498 & ~w3501;
assign w3511 = ~w3482 & ~w3485;
assign w3512 = ~w3475 & ~w3479;
assign w3513 = ~w3322 & ~w3325;
assign w3514 = ~w3512 & ~w3513;
assign w3515 = w3512 & w3513;
assign w3516 = ~w3514 & ~w3515;
assign w3517 = ~w3511 & w3516;
assign w3518 = w3511 & ~w3516;
assign w3519 = ~w3517 & ~w3518;
assign w3520 = ~w3491 & ~w3495;
assign w3521 = (~w3289 & w3299) | (~w3289 & w9135) | (w3299 & w9135);
assign w3522 = (~w3294 & ~w3296) | (~w3294 & w9136) | (~w3296 & w9136);
assign w3523 = w3280 & ~w3282;
assign w3524 = ~w3284 & ~w3523;
assign w3525 = ~w3522 & ~w3524;
assign w3526 = w3522 & w3524;
assign w3527 = ~w3525 & ~w3526;
assign w3528 = w3521 & w3527;
assign w3529 = ~w3521 & ~w3527;
assign w3530 = ~w3528 & ~w3529;
assign w3531 = (~w3450 & ~w3452) | (~w3450 & w8727) | (~w3452 & w8727);
assign w3532 = ~w3381 & ~w3384;
assign w3533 = (~w3419 & ~w3421) | (~w3419 & w9137) | (~w3421 & w9137);
assign w3534 = ~w3532 & ~w3533;
assign w3535 = w3532 & w3533;
assign w3536 = ~w3534 & ~w3535;
assign w3537 = (w3452 & w9138) | (w3452 & w9139) | (w9138 & w9139);
assign w3538 = ~w3536 & w3531;
assign w3539 = ~w3537 & ~w3538;
assign w3540 = w3530 & w3539;
assign w3541 = ~w3530 & ~w3539;
assign w3542 = ~w3540 & ~w3541;
assign w3543 = pi00 & pi61;
assign w3544 = pi02 & pi59;
assign w3545 = pi01 & pi60;
assign w3546 = ~w3544 & ~w3545;
assign w3547 = pi02 & pi60;
assign w3548 = w3280 & w3547;
assign w3549 = ~w3546 & ~w3548;
assign w3550 = w3543 & ~w3549;
assign w3551 = ~w3543 & w3549;
assign w3552 = ~w3550 & ~w3551;
assign w3553 = w3378 & ~w3552;
assign w3554 = ~w3378 & w3552;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = (~w3392 & w3387) | (~w3392 & w9140) | (w3387 & w9140);
assign w3557 = (~w3413 & w3409) | (~w3413 & w8728) | (w3409 & w8728);
assign w3558 = (~w3403 & w3398) | (~w3403 & w8729) | (w3398 & w8729);
assign w3559 = ~w3557 & ~w3558;
assign w3560 = w3557 & w3558;
assign w3561 = ~w3559 & ~w3560;
assign w3562 = ~w3556 & w3561;
assign w3563 = w3556 & ~w3561;
assign w3564 = ~w3562 & ~w3563;
assign w3565 = w3555 & w3564;
assign w3566 = ~w3555 & ~w3564;
assign w3567 = ~w3565 & ~w3566;
assign w3568 = w3542 & w3567;
assign w3569 = ~w3542 & ~w3567;
assign w3570 = ~w3568 & ~w3569;
assign w3571 = pi17 & pi44;
assign w3572 = pi21 & pi40;
assign w3573 = pi23 & pi38;
assign w3574 = ~w3332 & ~w3573;
assign w3575 = pi23 & pi39;
assign w3576 = w3330 & w3575;
assign w3577 = ~w3574 & ~w3576;
assign w3578 = w3572 & ~w3577;
assign w3579 = ~w3572 & w3577;
assign w3580 = ~w3578 & ~w3579;
assign w3581 = w3571 & ~w3580;
assign w3582 = ~w3571 & w3580;
assign w3583 = ~w3581 & ~w3582;
assign w3584 = pi18 & pi43;
assign w3585 = pi20 & pi41;
assign w3586 = ~w3344 & ~w3585;
assign w3587 = pi20 & pi42;
assign w3588 = w3342 & w3587;
assign w3589 = ~w3586 & ~w3588;
assign w3590 = w3584 & ~w3589;
assign w3591 = ~w3584 & w3589;
assign w3592 = ~w3590 & ~w3591;
assign w3593 = w3583 & ~w3592;
assign w3594 = ~w3583 & w3592;
assign w3595 = ~w3593 & ~w3594;
assign w3596 = pi24 & pi37;
assign w3597 = pi28 & pi33;
assign w3598 = pi29 & pi32;
assign w3599 = pi93 & w3598;
assign w3600 = ~pi93 & ~w3598;
assign w3601 = ~w3599 & ~w3600;
assign w3602 = w3597 & w3601;
assign w3603 = ~w3597 & ~w3601;
assign w3604 = ~w3602 & ~w3603;
assign w3605 = w3596 & w3604;
assign w3606 = ~w3596 & ~w3604;
assign w3607 = ~w3605 & ~w3606;
assign w3608 = pi25 & pi36;
assign w3609 = pi27 & pi34;
assign w3610 = ~w3368 & ~w3609;
assign w3611 = pi27 & pi35;
assign w3612 = w3366 & w3611;
assign w3613 = ~w3610 & ~w3612;
assign w3614 = w3608 & ~w3613;
assign w3615 = ~w3608 & w3613;
assign w3616 = ~w3614 & ~w3615;
assign w3617 = w3607 & ~w3616;
assign w3618 = ~w3607 & w3616;
assign w3619 = ~w3617 & ~w3618;
assign w3620 = ~w3461 & ~w3472;
assign w3621 = w3463 & ~w3465;
assign w3622 = ~w3467 & ~w3621;
assign w3623 = ~w3620 & ~w3622;
assign w3624 = w3620 & w3622;
assign w3625 = ~w3623 & ~w3624;
assign w3626 = ~w3619 & ~w3625;
assign w3627 = w3619 & w3625;
assign w3628 = ~w3626 & ~w3627;
assign w3629 = ~w3595 & w3628;
assign w3630 = w3595 & ~w3628;
assign w3631 = ~w3629 & ~w3630;
assign w3632 = (~w3435 & ~w3437) | (~w3435 & w8928) | (~w3437 & w8928);
assign w3633 = w3438 & ~w3440;
assign w3634 = ~w3442 & ~w3633;
assign w3635 = w3426 & ~w3428;
assign w3636 = ~w3430 & ~w3635;
assign w3637 = ~w3634 & ~w3636;
assign w3638 = w3634 & w3636;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = ~w3632 & w3639;
assign w3641 = w3632 & ~w3639;
assign w3642 = ~w3640 & ~w3641;
assign w3643 = (~w3338 & ~w3340) | (~w3338 & w8613) | (~w3340 & w8613);
assign w3644 = w3341 & ~w3343;
assign w3645 = ~w3345 & ~w3644;
assign w3646 = w3329 & ~w3331;
assign w3647 = ~w3333 & ~w3646;
assign w3648 = ~w3645 & ~w3647;
assign w3649 = w3645 & w3647;
assign w3650 = ~w3648 & ~w3649;
assign w3651 = ~w3643 & w3650;
assign w3652 = w3643 & ~w3650;
assign w3653 = ~w3651 & ~w3652;
assign w3654 = (~w3362 & ~w3364) | (~w3362 & w8614) | (~w3364 & w8614);
assign w3655 = (~w3356 & ~w3358) | (~w3356 & w8929) | (~w3358 & w8929);
assign w3656 = w3365 & ~w3367;
assign w3657 = ~w3369 & ~w3656;
assign w3658 = ~w3655 & ~w3657;
assign w3659 = w3655 & w3657;
assign w3660 = ~w3658 & ~w3659;
assign w3661 = ~w3654 & w3660;
assign w3662 = w3654 & ~w3660;
assign w3663 = ~w3661 & ~w3662;
assign w3664 = w3653 & w3663;
assign w3665 = ~w3653 & ~w3663;
assign w3666 = ~w3664 & ~w3665;
assign w3667 = w3642 & w3666;
assign w3668 = ~w3642 & ~w3666;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = pi10 & pi51;
assign w3671 = pi14 & pi47;
assign w3672 = pi16 & pi45;
assign w3673 = ~w3429 & ~w3672;
assign w3674 = pi16 & pi46;
assign w3675 = w3427 & w3674;
assign w3676 = ~w3673 & ~w3675;
assign w3677 = w3671 & ~w3676;
assign w3678 = ~w3671 & w3676;
assign w3679 = ~w3677 & ~w3678;
assign w3680 = w3670 & ~w3679;
assign w3681 = ~w3670 & w3679;
assign w3682 = ~w3680 & ~w3681;
assign w3683 = pi11 & pi50;
assign w3684 = pi13 & pi48;
assign w3685 = ~w3441 & ~w3684;
assign w3686 = pi13 & pi49;
assign w3687 = w3439 & w3686;
assign w3688 = ~w3685 & ~w3687;
assign w3689 = w3683 & ~w3688;
assign w3690 = ~w3683 & w3688;
assign w3691 = ~w3689 & ~w3690;
assign w3692 = w3682 & ~w3691;
assign w3693 = ~w3682 & w3691;
assign w3694 = ~w3692 & ~w3693;
assign w3695 = w3669 & w3694;
assign w3696 = ~w3669 & ~w3694;
assign w3697 = ~w3695 & ~w3696;
assign w3698 = ~w3631 & w3697;
assign w3699 = w3631 & ~w3697;
assign w3700 = ~w3698 & ~w3699;
assign w3701 = (~w3316 & w3313) | (~w3316 & w8930) | (w3313 & w8930);
assign w3702 = ~w3307 & ~w3310;
assign w3703 = pi07 & pi54;
assign w3704 = pi09 & pi52;
assign w3705 = ~w3466 & ~w3704;
assign w3706 = pi09 & pi53;
assign w3707 = w3464 & w3706;
assign w3708 = ~w3705 & ~w3707;
assign w3709 = w3703 & ~w3708;
assign w3710 = ~w3703 & w3708;
assign w3711 = ~w3709 & ~w3710;
assign w3712 = w3283 & ~w3711;
assign w3713 = ~w3283 & w3711;
assign w3714 = ~w3712 & ~w3713;
assign w3715 = pi04 & pi57;
assign w3716 = pi06 & pi55;
assign w3717 = ~w3460 & ~w3716;
assign w3718 = pi06 & pi56;
assign w3719 = w3457 & w3718;
assign w3720 = ~w3717 & ~w3719;
assign w3721 = w3715 & ~w3720;
assign w3722 = ~w3715 & w3720;
assign w3723 = ~w3721 & ~w3722;
assign w3724 = w3714 & ~w3723;
assign w3725 = ~w3714 & w3723;
assign w3726 = ~w3724 & ~w3725;
assign w3727 = w3702 & ~w3726;
assign w3728 = ~w3702 & w3726;
assign w3729 = ~w3727 & ~w3728;
assign w3730 = w3701 & w3729;
assign w3731 = ~w3701 & ~w3729;
assign w3732 = ~w3730 & ~w3731;
assign w3733 = w3700 & ~w3732;
assign w3734 = ~w3700 & w3732;
assign w3735 = ~w3733 & ~w3734;
assign w3736 = w3570 & w3735;
assign w3737 = ~w3570 & ~w3735;
assign w3738 = ~w3736 & ~w3737;
assign w3739 = ~w3520 & w3738;
assign w3740 = w3520 & ~w3738;
assign w3741 = ~w3739 & ~w3740;
assign w3742 = w3519 & w3741;
assign w3743 = ~w3519 & ~w3741;
assign w3744 = ~w3742 & ~w3743;
assign w3745 = w3510 & ~w3744;
assign w3746 = ~w3510 & w3744;
assign w3747 = ~w3745 & ~w3746;
assign w3748 = ~w3504 & ~w3507;
assign w3749 = ~w3747 & w3748;
assign w3750 = w3747 & ~w3748;
assign w3751 = ~w3749 & ~w3750;
assign w3752 = w3506 & w3747;
assign w3753 = w3272 & w3752;
assign w3754 = w3275 & w9269;
assign w3755 = ~w3753 & ~w3754;
assign w3756 = ~w3504 & ~w3746;
assign w3757 = ~w3745 & ~w3756;
assign w3758 = w3755 & ~w3757;
assign w3759 = pi11 & pi51;
assign w3760 = pi15 & pi47;
assign w3761 = pi17 & pi45;
assign w3762 = ~w3674 & ~w3761;
assign w3763 = pi17 & pi46;
assign w3764 = w3672 & w3763;
assign w3765 = ~w3762 & ~w3764;
assign w3766 = w3760 & ~w3765;
assign w3767 = ~w3760 & w3765;
assign w3768 = ~w3766 & ~w3767;
assign w3769 = w3759 & ~w3768;
assign w3770 = ~w3759 & w3768;
assign w3771 = ~w3769 & ~w3770;
assign w3772 = pi12 & pi50;
assign w3773 = pi14 & pi48;
assign w3774 = ~w3686 & ~w3773;
assign w3775 = pi14 & pi49;
assign w3776 = w3684 & w3775;
assign w3777 = ~w3774 & ~w3776;
assign w3778 = w3772 & ~w3777;
assign w3779 = ~w3772 & w3777;
assign w3780 = ~w3778 & ~w3779;
assign w3781 = w3771 & ~w3780;
assign w3782 = ~w3771 & w3780;
assign w3783 = ~w3781 & ~w3782;
assign w3784 = pi18 & pi44;
assign w3785 = pi22 & pi40;
assign w3786 = pi24 & pi38;
assign w3787 = ~w3575 & ~w3786;
assign w3788 = pi24 & pi39;
assign w3789 = w3573 & w3788;
assign w3790 = ~w3787 & ~w3789;
assign w3791 = w3785 & ~w3790;
assign w3792 = ~w3785 & w3790;
assign w3793 = ~w3791 & ~w3792;
assign w3794 = w3784 & ~w3793;
assign w3795 = ~w3784 & w3793;
assign w3796 = ~w3794 & ~w3795;
assign w3797 = pi19 & pi43;
assign w3798 = pi21 & pi41;
assign w3799 = ~w3587 & ~w3798;
assign w3800 = pi21 & pi42;
assign w3801 = w3585 & w3800;
assign w3802 = ~w3799 & ~w3801;
assign w3803 = w3797 & ~w3802;
assign w3804 = ~w3797 & w3802;
assign w3805 = ~w3803 & ~w3804;
assign w3806 = w3796 & ~w3805;
assign w3807 = ~w3796 & w3805;
assign w3808 = ~w3806 & ~w3807;
assign w3809 = pi25 & pi37;
assign w3810 = pi29 & pi33;
assign w3811 = pi30 & pi32;
assign w3812 = pi94 & w3811;
assign w3813 = ~pi94 & ~w3811;
assign w3814 = ~w3812 & ~w3813;
assign w3815 = w3810 & w3814;
assign w3816 = ~w3810 & ~w3814;
assign w3817 = ~w3815 & ~w3816;
assign w3818 = w3809 & w3817;
assign w3819 = ~w3809 & ~w3817;
assign w3820 = ~w3818 & ~w3819;
assign w3821 = pi26 & pi36;
assign w3822 = pi28 & pi34;
assign w3823 = ~w3611 & ~w3822;
assign w3824 = pi28 & pi35;
assign w3825 = w3609 & w3824;
assign w3826 = ~w3823 & ~w3825;
assign w3827 = w3821 & ~w3826;
assign w3828 = ~w3821 & w3826;
assign w3829 = ~w3827 & ~w3828;
assign w3830 = w3820 & ~w3829;
assign w3831 = ~w3820 & w3829;
assign w3832 = ~w3830 & ~w3831;
assign w3833 = w3808 & w3832;
assign w3834 = ~w3808 & ~w3832;
assign w3835 = ~w3833 & ~w3834;
assign w3836 = w3783 & w3835;
assign w3837 = ~w3783 & ~w3835;
assign w3838 = ~w3836 & ~w3837;
assign w3839 = (~w3712 & ~w3714) | (~w3712 & w8615) | (~w3714 & w8615);
assign w3840 = w3715 & ~w3717;
assign w3841 = ~w3719 & ~w3840;
assign w3842 = w3703 & ~w3705;
assign w3843 = ~w3707 & ~w3842;
assign w3844 = ~w3841 & ~w3843;
assign w3845 = w3841 & w3843;
assign w3846 = ~w3844 & ~w3845;
assign w3847 = ~w3839 & w3846;
assign w3848 = w3839 & ~w3846;
assign w3849 = ~w3847 & ~w3848;
assign w3850 = (~w3680 & ~w3682) | (~w3680 & w8616) | (~w3682 & w8616);
assign w3851 = w3683 & ~w3685;
assign w3852 = ~w3687 & ~w3851;
assign w3853 = w3671 & ~w3673;
assign w3854 = ~w3675 & ~w3853;
assign w3855 = ~w3852 & ~w3854;
assign w3856 = w3852 & w3854;
assign w3857 = ~w3855 & ~w3856;
assign w3858 = ~w3850 & w3857;
assign w3859 = w3850 & ~w3857;
assign w3860 = ~w3858 & ~w3859;
assign w3861 = (~w3581 & ~w3583) | (~w3581 & w8617) | (~w3583 & w8617);
assign w3862 = w3584 & ~w3586;
assign w3863 = ~w3588 & ~w3862;
assign w3864 = w3572 & ~w3574;
assign w3865 = ~w3576 & ~w3864;
assign w3866 = ~w3863 & ~w3865;
assign w3867 = w3863 & w3865;
assign w3868 = ~w3866 & ~w3867;
assign w3869 = ~w3861 & w3868;
assign w3870 = w3861 & ~w3868;
assign w3871 = ~w3869 & ~w3870;
assign w3872 = w3860 & w3871;
assign w3873 = ~w3860 & ~w3871;
assign w3874 = ~w3872 & ~w3873;
assign w3875 = w3849 & w3874;
assign w3876 = ~w3849 & ~w3874;
assign w3877 = ~w3875 & ~w3876;
assign w3878 = pi04 & pi58;
assign w3879 = pi08 & pi54;
assign w3880 = pi10 & pi52;
assign w3881 = ~w3706 & ~w3880;
assign w3882 = pi10 & pi53;
assign w3883 = w3704 & w3882;
assign w3884 = ~w3881 & ~w3883;
assign w3885 = w3879 & ~w3884;
assign w3886 = ~w3879 & w3884;
assign w3887 = ~w3885 & ~w3886;
assign w3888 = w3878 & ~w3887;
assign w3889 = ~w3878 & w3887;
assign w3890 = ~w3888 & ~w3889;
assign w3891 = pi05 & pi57;
assign w3892 = pi07 & pi55;
assign w3893 = ~w3718 & ~w3892;
assign w3894 = pi07 & pi56;
assign w3895 = w3716 & w3894;
assign w3896 = ~w3893 & ~w3895;
assign w3897 = w3891 & ~w3896;
assign w3898 = ~w3891 & w3896;
assign w3899 = ~w3897 & ~w3898;
assign w3900 = w3890 & ~w3899;
assign w3901 = ~w3890 & w3899;
assign w3902 = ~w3900 & ~w3901;
assign w3903 = w3877 & w3902;
assign w3904 = ~w3877 & ~w3902;
assign w3905 = ~w3903 & ~w3904;
assign w3906 = w3838 & w3905;
assign w3907 = ~w3838 & ~w3905;
assign w3908 = ~w3906 & ~w3907;
assign w3909 = (~w3534 & w3531) | (~w3534 & w8931) | (w3531 & w8931);
assign w3910 = pi03 & pi59;
assign w3911 = ~w3547 & ~w3910;
assign w3912 = pi03 & pi60;
assign w3913 = w3544 & w3912;
assign w3914 = ~w3911 & ~w3913;
assign w3915 = ~w3525 & ~w3528;
assign w3916 = w3914 & ~w3915;
assign w3917 = ~w3914 & w3915;
assign w3918 = ~w3916 & ~w3917;
assign w3919 = w3909 & w3918;
assign w3920 = ~w3909 & ~w3918;
assign w3921 = ~w3919 & ~w3920;
assign w3922 = w3908 & ~w3921;
assign w3923 = ~w3908 & w3921;
assign w3924 = ~w3922 & ~w3923;
assign w3925 = (~w3605 & ~w3607) | (~w3605 & w8618) | (~w3607 & w8618);
assign w3926 = (~w3599 & ~w3601) | (~w3599 & w8932) | (~w3601 & w8932);
assign w3927 = w3608 & ~w3610;
assign w3928 = ~w3612 & ~w3927;
assign w3929 = ~w3926 & ~w3928;
assign w3930 = w3926 & w3928;
assign w3931 = ~w3929 & ~w3930;
assign w3932 = ~w3925 & w3931;
assign w3933 = w3925 & ~w3931;
assign w3934 = ~w3932 & ~w3933;
assign w3935 = pi01 & pi61;
assign w3936 = pi00 & pi62;
assign w3937 = ~w3935 & ~w3936;
assign w3938 = pi01 & pi62;
assign w3939 = w3543 & w3938;
assign w3940 = ~w3937 & ~w3939;
assign w3941 = (~w3654 & w8933) | (~w3654 & w8934) | (w8933 & w8934);
assign w3942 = (w3654 & w8935) | (w3654 & w8936) | (w8935 & w8936);
assign w3943 = ~w3941 & ~w3942;
assign w3944 = w3934 & w3943;
assign w3945 = ~w3934 & ~w3943;
assign w3946 = ~w3944 & ~w3945;
assign w3947 = (~w3637 & w3632) | (~w3637 & w9141) | (w3632 & w9141);
assign w3948 = (~w3648 & w3643) | (~w3648 & w8730) | (w3643 & w8730);
assign w3949 = w3623 & ~w3948;
assign w3950 = ~w3623 & w3948;
assign w3951 = ~w3949 & ~w3950;
assign w3952 = ~w3947 & ~w3951;
assign w3953 = w3947 & w3951;
assign w3954 = ~w3952 & ~w3953;
assign w3955 = w3946 & ~w3954;
assign w3956 = ~w3946 & w3954;
assign w3957 = ~w3955 & ~w3956;
assign w3958 = (~w3553 & ~w3564) | (~w3553 & w8937) | (~w3564 & w8937);
assign w3959 = (~w3559 & ~w3561) | (~w3559 & w8938) | (~w3561 & w8938);
assign w3960 = w3543 & ~w3546;
assign w3961 = ~w3548 & ~w3960;
assign w3962 = ~w3959 & ~w3961;
assign w3963 = w3959 & w3961;
assign w3964 = ~w3962 & ~w3963;
assign w3965 = ~w3958 & w3964;
assign w3966 = w3958 & ~w3964;
assign w3967 = ~w3965 & ~w3966;
assign w3968 = (~w3695 & ~w3697) | (~w3695 & w8731) | (~w3697 & w8731);
assign w3969 = ~w3626 & ~w3629;
assign w3970 = (~w3664 & ~w3666) | (~w3664 & w9142) | (~w3666 & w9142);
assign w3971 = w3969 & ~w3970;
assign w3972 = ~w3969 & w3970;
assign w3973 = ~w3971 & ~w3972;
assign w3974 = w3973 & w3968;
assign w3975 = (w3697 & w9143) | (w3697 & w9144) | (w9143 & w9144);
assign w3976 = ~w3974 & ~w3975;
assign w3977 = w3967 & ~w3976;
assign w3978 = ~w3967 & w3976;
assign w3979 = ~w3977 & ~w3978;
assign w3980 = w3957 & ~w3979;
assign w3981 = ~w3957 & w3979;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = w3924 & ~w3982;
assign w3984 = ~w3924 & w3982;
assign w3985 = ~w3983 & ~w3984;
assign w3986 = ~w3514 & ~w3517;
assign w3987 = (~w3733 & ~w3570) | (~w3733 & w8939) | (~w3570 & w8939);
assign w3988 = ~w3727 & ~w3730;
assign w3989 = (~w3540 & ~w3542) | (~w3540 & w8940) | (~w3542 & w8940);
assign w3990 = w3988 & ~w3989;
assign w3991 = ~w3988 & w3989;
assign w3992 = ~w3990 & ~w3991;
assign w3993 = ~w3987 & w3992;
assign w3994 = w3987 & ~w3992;
assign w3995 = ~w3993 & ~w3994;
assign w3996 = ~w3986 & w3995;
assign w3997 = w3986 & ~w3995;
assign w3998 = ~w3996 & ~w3997;
assign w3999 = w3985 & w3998;
assign w4000 = ~w3985 & ~w3998;
assign w4001 = ~w3999 & ~w4000;
assign w4002 = ~w3739 & ~w3742;
assign w4003 = w4001 & ~w4002;
assign w4004 = ~w4001 & w4002;
assign w4005 = ~w4003 & ~w4004;
assign w4006 = ~w3758 & w4005;
assign w4007 = w3758 & ~w4005;
assign w4008 = ~w4006 & ~w4007;
assign w4009 = ~w3757 & ~w4003;
assign w4010 = ~w3754 & w8732;
assign w4011 = ~w4004 & ~w4010;
assign w4012 = ~w3996 & ~w3999;
assign w4013 = pi12 & pi51;
assign w4014 = pi16 & pi47;
assign w4015 = pi18 & pi45;
assign w4016 = ~w3763 & ~w4015;
assign w4017 = pi18 & pi46;
assign w4018 = w3761 & w4017;
assign w4019 = ~w4016 & ~w4018;
assign w4020 = w4014 & ~w4019;
assign w4021 = ~w4014 & w4019;
assign w4022 = ~w4020 & ~w4021;
assign w4023 = w4013 & ~w4022;
assign w4024 = ~w4013 & w4022;
assign w4025 = ~w4023 & ~w4024;
assign w4026 = pi13 & pi50;
assign w4027 = pi15 & pi48;
assign w4028 = ~w3775 & ~w4027;
assign w4029 = pi15 & pi49;
assign w4030 = w3773 & w4029;
assign w4031 = ~w4028 & ~w4030;
assign w4032 = w4026 & ~w4031;
assign w4033 = ~w4026 & w4031;
assign w4034 = ~w4032 & ~w4033;
assign w4035 = w4025 & ~w4034;
assign w4036 = ~w4025 & w4034;
assign w4037 = ~w4035 & ~w4036;
assign w4038 = pi19 & pi44;
assign w4039 = pi23 & pi40;
assign w4040 = pi25 & pi38;
assign w4041 = ~w3788 & ~w4040;
assign w4042 = pi25 & pi39;
assign w4043 = w3786 & w4042;
assign w4044 = ~w4041 & ~w4043;
assign w4045 = w4039 & ~w4044;
assign w4046 = ~w4039 & w4044;
assign w4047 = ~w4045 & ~w4046;
assign w4048 = w4038 & ~w4047;
assign w4049 = ~w4038 & w4047;
assign w4050 = ~w4048 & ~w4049;
assign w4051 = pi20 & pi43;
assign w4052 = pi22 & pi41;
assign w4053 = ~w3800 & ~w4052;
assign w4054 = pi22 & pi42;
assign w4055 = w3798 & w4054;
assign w4056 = ~w4053 & ~w4055;
assign w4057 = w4051 & ~w4056;
assign w4058 = ~w4051 & w4056;
assign w4059 = ~w4057 & ~w4058;
assign w4060 = w4050 & ~w4059;
assign w4061 = ~w4050 & w4059;
assign w4062 = ~w4060 & ~w4061;
assign w4063 = pi26 & pi37;
assign w4064 = pi30 & pi33;
assign w4065 = pi31 & pi32;
assign w4066 = ~pi95 & ~w4065;
assign w4067 = pi95 & w4065;
assign w4068 = ~w4066 & ~w4067;
assign w4069 = w4064 & w4068;
assign w4070 = ~w4064 & ~w4068;
assign w4071 = ~w4069 & ~w4070;
assign w4072 = w4063 & w4071;
assign w4073 = ~w4063 & ~w4071;
assign w4074 = ~w4072 & ~w4073;
assign w4075 = pi27 & pi36;
assign w4076 = pi29 & pi34;
assign w4077 = ~w3824 & ~w4076;
assign w4078 = pi29 & pi35;
assign w4079 = w3822 & w4078;
assign w4080 = ~w4077 & ~w4079;
assign w4081 = w4075 & ~w4080;
assign w4082 = ~w4075 & w4080;
assign w4083 = ~w4081 & ~w4082;
assign w4084 = w4074 & ~w4083;
assign w4085 = ~w4074 & w4083;
assign w4086 = ~w4084 & ~w4085;
assign w4087 = w4062 & w4086;
assign w4088 = ~w4062 & ~w4086;
assign w4089 = ~w4087 & ~w4088;
assign w4090 = w4037 & w4089;
assign w4091 = ~w4037 & ~w4089;
assign w4092 = ~w4090 & ~w4091;
assign w4093 = pi05 & pi58;
assign w4094 = pi09 & pi54;
assign w4095 = pi11 & pi52;
assign w4096 = ~w3882 & ~w4095;
assign w4097 = pi11 & pi53;
assign w4098 = w3880 & w4097;
assign w4099 = ~w4096 & ~w4098;
assign w4100 = w4094 & ~w4099;
assign w4101 = ~w4094 & w4099;
assign w4102 = ~w4100 & ~w4101;
assign w4103 = w4093 & ~w4102;
assign w4104 = ~w4093 & w4102;
assign w4105 = ~w4103 & ~w4104;
assign w4106 = pi06 & pi57;
assign w4107 = pi08 & pi55;
assign w4108 = ~w3894 & ~w4107;
assign w4109 = pi08 & pi56;
assign w4110 = w3892 & w4109;
assign w4111 = ~w4108 & ~w4110;
assign w4112 = w4106 & ~w4111;
assign w4113 = ~w4106 & w4111;
assign w4114 = ~w4112 & ~w4113;
assign w4115 = w4105 & ~w4114;
assign w4116 = ~w4105 & w4114;
assign w4117 = ~w4115 & ~w4116;
assign w4118 = (~w3888 & ~w3890) | (~w3888 & w8619) | (~w3890 & w8619);
assign w4119 = w3891 & ~w3893;
assign w4120 = ~w3895 & ~w4119;
assign w4121 = w3879 & ~w3881;
assign w4122 = ~w3883 & ~w4121;
assign w4123 = ~w4120 & ~w4122;
assign w4124 = w4120 & w4122;
assign w4125 = ~w4123 & ~w4124;
assign w4126 = ~w4118 & w4125;
assign w4127 = w4118 & ~w4125;
assign w4128 = ~w4126 & ~w4127;
assign w4129 = (~w3769 & ~w3771) | (~w3769 & w8620) | (~w3771 & w8620);
assign w4130 = w3772 & ~w3774;
assign w4131 = ~w3776 & ~w4130;
assign w4132 = w3760 & ~w3762;
assign w4133 = ~w3764 & ~w4132;
assign w4134 = ~w4131 & ~w4133;
assign w4135 = w4131 & w4133;
assign w4136 = ~w4134 & ~w4135;
assign w4137 = ~w4129 & w4136;
assign w4138 = w4129 & ~w4136;
assign w4139 = ~w4137 & ~w4138;
assign w4140 = w4128 & w4139;
assign w4141 = ~w4128 & ~w4139;
assign w4142 = ~w4140 & ~w4141;
assign w4143 = w3913 & ~w4142;
assign w4144 = ~w3913 & w4142;
assign w4145 = ~w4143 & ~w4144;
assign w4146 = ~w4117 & w4145;
assign w4147 = w4117 & ~w4145;
assign w4148 = ~w4146 & ~w4147;
assign w4149 = ~w4092 & w4148;
assign w4150 = w4092 & ~w4148;
assign w4151 = ~w4149 & ~w4150;
assign w4152 = pi00 & pi63;
assign w4153 = w3938 & ~w4152;
assign w4154 = ~w3938 & w4152;
assign w4155 = ~w4153 & ~w4154;
assign w4156 = pi02 & pi61;
assign w4157 = pi04 & pi59;
assign w4158 = ~w3912 & ~w4157;
assign w4159 = pi04 & pi60;
assign w4160 = w3910 & w4159;
assign w4161 = ~w4158 & ~w4160;
assign w4162 = w4156 & ~w4161;
assign w4163 = ~w4156 & w4161;
assign w4164 = ~w4162 & ~w4163;
assign w4165 = w4155 & ~w4164;
assign w4166 = ~w4155 & w4164;
assign w4167 = ~w4165 & ~w4166;
assign w4168 = (w4167 & w3965) | (w4167 & w9145) | (w3965 & w9145);
assign w4169 = ~w3965 & w9146;
assign w4170 = ~w4168 & ~w4169;
assign w4171 = (~w3972 & ~w3968) | (~w3972 & w8941) | (~w3968 & w8941);
assign w4172 = w4170 & w4171;
assign w4173 = ~w4170 & ~w4171;
assign w4174 = ~w4172 & ~w4173;
assign w4175 = w4151 & ~w4174;
assign w4176 = ~w4151 & w4174;
assign w4177 = ~w4175 & ~w4176;
assign w4178 = (~w3818 & ~w3820) | (~w3818 & w8733) | (~w3820 & w8733);
assign w4179 = ~w3812 & ~w3815;
assign w4180 = w3821 & ~w3823;
assign w4181 = ~w3825 & ~w4180;
assign w4182 = ~w4179 & ~w4181;
assign w4183 = w4179 & w4181;
assign w4184 = ~w4182 & ~w4183;
assign w4185 = ~w4178 & w4184;
assign w4186 = w4178 & ~w4184;
assign w4187 = ~w4185 & ~w4186;
assign w4188 = (~w3855 & w3850) | (~w3855 & w8734) | (w3850 & w8734);
assign w4189 = (~w3844 & w3839) | (~w3844 & w8735) | (w3839 & w8735);
assign w4190 = ~w4188 & ~w4189;
assign w4191 = w4188 & w4189;
assign w4192 = ~w4190 & ~w4191;
assign w4193 = w4187 & w4192;
assign w4194 = ~w4187 & ~w4192;
assign w4195 = ~w4193 & ~w4194;
assign w4196 = (~w3794 & ~w3796) | (~w3794 & w8736) | (~w3796 & w8736);
assign w4197 = w3797 & ~w3799;
assign w4198 = ~w3801 & ~w4197;
assign w4199 = w3785 & ~w3787;
assign w4200 = ~w3789 & ~w4199;
assign w4201 = ~w4198 & ~w4200;
assign w4202 = w4198 & w4200;
assign w4203 = ~w4201 & ~w4202;
assign w4204 = ~w4196 & w4203;
assign w4205 = w4196 & ~w4203;
assign w4206 = ~w4204 & ~w4205;
assign w4207 = (~w3866 & w3861) | (~w3866 & w8737) | (w3861 & w8737);
assign w4208 = (~w3929 & w3925) | (~w3929 & w8738) | (w3925 & w8738);
assign w4209 = w4207 & w4208;
assign w4210 = ~w4207 & ~w4208;
assign w4211 = ~w4209 & ~w4210;
assign w4212 = w4206 & ~w4211;
assign w4213 = ~w4206 & w4211;
assign w4214 = ~w4212 & ~w4213;
assign w4215 = w4195 & w4214;
assign w4216 = ~w4195 & ~w4214;
assign w4217 = ~w4215 & ~w4216;
assign w4218 = (~w3944 & w3954) | (~w3944 & w8942) | (w3954 & w8942);
assign w4219 = ~w3939 & ~w3941;
assign w4220 = (~w3950 & ~w3951) | (~w3950 & w8943) | (~w3951 & w8943);
assign w4221 = ~w4219 & w4220;
assign w4222 = w4219 & ~w4220;
assign w4223 = ~w4221 & ~w4222;
assign w4224 = ~w4218 & w4223;
assign w4225 = w4218 & ~w4223;
assign w4226 = ~w4224 & ~w4225;
assign w4227 = (~w3903 & ~w3905) | (~w3903 & w8739) | (~w3905 & w8739);
assign w4228 = ~w3833 & ~w3836;
assign w4229 = (~w3872 & ~w3874) | (~w3872 & w9147) | (~w3874 & w9147);
assign w4230 = ~w4228 & ~w4229;
assign w4231 = w4228 & w4229;
assign w4232 = ~w4230 & ~w4231;
assign w4233 = ~w4232 & w4227;
assign w4234 = (w3905 & w9148) | (w3905 & w9149) | (w9148 & w9149);
assign w4235 = ~w4233 & ~w4234;
assign w4236 = w4226 & w4235;
assign w4237 = ~w4226 & ~w4235;
assign w4238 = ~w4236 & ~w4237;
assign w4239 = w4217 & ~w4238;
assign w4240 = ~w4217 & w4238;
assign w4241 = ~w4239 & ~w4240;
assign w4242 = ~w4177 & ~w4241;
assign w4243 = w4177 & w4241;
assign w4244 = ~w4242 & ~w4243;
assign w4245 = (~w3990 & w3987) | (~w3990 & w9150) | (w3987 & w9150);
assign w4246 = (~w3922 & w3982) | (~w3922 & w8944) | (w3982 & w8944);
assign w4247 = ~w3917 & ~w3919;
assign w4248 = (~w3978 & ~w3979) | (~w3978 & w8945) | (~w3979 & w8945);
assign w4249 = w4247 & w4248;
assign w4250 = ~w4247 & ~w4248;
assign w4251 = ~w4249 & ~w4250;
assign w4252 = w4246 & ~w4251;
assign w4253 = ~w4246 & w4251;
assign w4254 = ~w4252 & ~w4253;
assign w4255 = w4245 & ~w4254;
assign w4256 = ~w4245 & w4254;
assign w4257 = ~w4255 & ~w4256;
assign w4258 = w4244 & w4257;
assign w4259 = ~w4244 & ~w4257;
assign w4260 = ~w4258 & ~w4259;
assign w4261 = ~w4012 & ~w4260;
assign w4262 = w4012 & w4260;
assign w4263 = ~w4261 & ~w4262;
assign w4264 = w4011 & ~w4263;
assign w4265 = ~w4003 & w4263;
assign w4266 = ~w4006 & w4265;
assign w4267 = ~w4264 & ~w4266;
assign w4268 = pi19 & pi45;
assign w4269 = pi23 & pi41;
assign w4270 = pi24 & pi40;
assign w4271 = ~w4042 & ~w4270;
assign w4272 = pi25 & pi40;
assign w4273 = w3788 & w4272;
assign w4274 = ~w4271 & ~w4273;
assign w4275 = w4269 & ~w4274;
assign w4276 = ~w4269 & w4274;
assign w4277 = ~w4275 & ~w4276;
assign w4278 = w4268 & ~w4277;
assign w4279 = ~w4268 & w4277;
assign w4280 = ~w4278 & ~w4279;
assign w4281 = pi20 & pi44;
assign w4282 = pi21 & pi43;
assign w4283 = ~w4054 & ~w4282;
assign w4284 = pi22 & pi43;
assign w4285 = w3800 & w4284;
assign w4286 = ~w4283 & ~w4285;
assign w4287 = w4281 & ~w4286;
assign w4288 = ~w4281 & w4286;
assign w4289 = ~w4287 & ~w4288;
assign w4290 = w4280 & ~w4289;
assign w4291 = ~w4280 & w4289;
assign w4292 = ~w4290 & ~w4291;
assign w4293 = pi26 & pi38;
assign w4294 = pi30 & pi34;
assign w4295 = pi31 & pi33;
assign w4296 = ~w4294 & w4295;
assign w4297 = w4294 & ~w4295;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = w4293 & ~w4298;
assign w4300 = ~w4293 & w4298;
assign w4301 = ~w4299 & ~w4300;
assign w4302 = pi27 & pi37;
assign w4303 = pi28 & pi36;
assign w4304 = ~w4078 & ~w4303;
assign w4305 = pi29 & pi36;
assign w4306 = w3824 & w4305;
assign w4307 = ~w4304 & ~w4306;
assign w4308 = w4302 & ~w4307;
assign w4309 = ~w4302 & w4307;
assign w4310 = ~w4308 & ~w4309;
assign w4311 = w4301 & ~w4310;
assign w4312 = ~w4301 & w4310;
assign w4313 = ~w4311 & ~w4312;
assign w4314 = w4292 & w4313;
assign w4315 = ~w4292 & ~w4313;
assign w4316 = ~w4314 & ~w4315;
assign w4317 = pi12 & pi52;
assign w4318 = pi16 & pi48;
assign w4319 = pi17 & pi47;
assign w4320 = ~w4017 & ~w4319;
assign w4321 = pi18 & pi47;
assign w4322 = w3763 & w4321;
assign w4323 = ~w4320 & ~w4322;
assign w4324 = w4318 & ~w4323;
assign w4325 = ~w4318 & w4323;
assign w4326 = ~w4324 & ~w4325;
assign w4327 = w4317 & ~w4326;
assign w4328 = ~w4317 & w4326;
assign w4329 = ~w4327 & ~w4328;
assign w4330 = pi13 & pi51;
assign w4331 = pi14 & pi50;
assign w4332 = ~w4029 & ~w4331;
assign w4333 = pi15 & pi50;
assign w4334 = w3775 & w4333;
assign w4335 = ~w4332 & ~w4334;
assign w4336 = w4330 & ~w4335;
assign w4337 = ~w4330 & w4335;
assign w4338 = ~w4336 & ~w4337;
assign w4339 = w4329 & ~w4338;
assign w4340 = ~w4329 & w4338;
assign w4341 = ~w4339 & ~w4340;
assign w4342 = w4316 & w4341;
assign w4343 = ~w4316 & ~w4341;
assign w4344 = ~w4342 & ~w4343;
assign w4345 = pi05 & pi59;
assign w4346 = pi09 & pi55;
assign w4347 = pi10 & pi54;
assign w4348 = ~w4097 & ~w4347;
assign w4349 = pi11 & pi54;
assign w4350 = w3882 & w4349;
assign w4351 = ~w4348 & ~w4350;
assign w4352 = w4346 & ~w4351;
assign w4353 = ~w4346 & w4351;
assign w4354 = ~w4352 & ~w4353;
assign w4355 = w4345 & ~w4354;
assign w4356 = ~w4345 & w4354;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = pi06 & pi58;
assign w4359 = pi07 & pi57;
assign w4360 = ~w4109 & ~w4359;
assign w4361 = pi08 & pi57;
assign w4362 = w3894 & w4361;
assign w4363 = ~w4360 & ~w4362;
assign w4364 = w4358 & ~w4363;
assign w4365 = ~w4358 & w4363;
assign w4366 = ~w4364 & ~w4365;
assign w4367 = w4357 & ~w4366;
assign w4368 = ~w4357 & w4366;
assign w4369 = ~w4367 & ~w4368;
assign w4370 = (~w4103 & ~w4105) | (~w4103 & w8621) | (~w4105 & w8621);
assign w4371 = w4106 & ~w4108;
assign w4372 = ~w4110 & ~w4371;
assign w4373 = w4094 & ~w4096;
assign w4374 = ~w4098 & ~w4373;
assign w4375 = ~w4372 & ~w4374;
assign w4376 = w4372 & w4374;
assign w4377 = ~w4375 & ~w4376;
assign w4378 = ~w4370 & w4377;
assign w4379 = w4370 & ~w4377;
assign w4380 = ~w4378 & ~w4379;
assign w4381 = (~w4023 & ~w4025) | (~w4023 & w8622) | (~w4025 & w8622);
assign w4382 = w4026 & ~w4028;
assign w4383 = ~w4030 & ~w4382;
assign w4384 = w4014 & ~w4016;
assign w4385 = ~w4018 & ~w4384;
assign w4386 = ~w4383 & ~w4385;
assign w4387 = w4383 & w4385;
assign w4388 = ~w4386 & ~w4387;
assign w4389 = ~w4381 & w4388;
assign w4390 = w4381 & ~w4388;
assign w4391 = ~w4389 & ~w4390;
assign w4392 = w4380 & w4391;
assign w4393 = ~w4380 & ~w4391;
assign w4394 = ~w4392 & ~w4393;
assign w4395 = ~w4153 & ~w4165;
assign w4396 = w4156 & ~w4158;
assign w4397 = ~w4160 & ~w4396;
assign w4398 = ~w4395 & ~w4397;
assign w4399 = w4395 & w4397;
assign w4400 = ~w4398 & ~w4399;
assign w4401 = w4394 & w4400;
assign w4402 = ~w4394 & ~w4400;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = w4369 & w4403;
assign w4405 = ~w4369 & ~w4403;
assign w4406 = ~w4404 & ~w4405;
assign w4407 = w4344 & w4406;
assign w4408 = ~w4344 & ~w4406;
assign w4409 = ~w4407 & ~w4408;
assign w4410 = pi01 & pi63;
assign w4411 = pi02 & pi62;
assign w4412 = pi03 & pi61;
assign w4413 = ~w4159 & ~w4412;
assign w4414 = pi04 & pi61;
assign w4415 = w3912 & w4414;
assign w4416 = ~w4413 & ~w4415;
assign w4417 = w4411 & w4416;
assign w4418 = ~w4411 & ~w4416;
assign w4419 = ~w4417 & ~w4418;
assign w4420 = ~w4410 & w4419;
assign w4421 = w4410 & ~w4419;
assign w4422 = ~w4420 & ~w4421;
assign w4423 = (w4422 & w4224) | (w4422 & w9151) | (w4224 & w9151);
assign w4424 = ~w4224 & w9152;
assign w4425 = ~w4423 & ~w4424;
assign w4426 = (~w4230 & w4227) | (~w4230 & w8946) | (w4227 & w8946);
assign w4427 = w4425 & ~w4426;
assign w4428 = ~w4425 & w4426;
assign w4429 = ~w4427 & ~w4428;
assign w4430 = ~w4409 & ~w4429;
assign w4431 = w4409 & w4429;
assign w4432 = ~w4430 & ~w4431;
assign w4433 = (~w4072 & ~w4074) | (~w4072 & w8623) | (~w4074 & w8623);
assign w4434 = (~w4066 & ~w4068) | (~w4066 & w8947) | (~w4068 & w8947);
assign w4435 = w4075 & ~w4077;
assign w4436 = ~w4079 & ~w4435;
assign w4437 = ~w4434 & ~w4436;
assign w4438 = w4434 & w4436;
assign w4439 = ~w4437 & ~w4438;
assign w4440 = ~w4433 & w4439;
assign w4441 = w4433 & ~w4439;
assign w4442 = ~w4440 & ~w4441;
assign w4443 = (~w4134 & w4129) | (~w4134 & w9153) | (w4129 & w9153);
assign w4444 = (~w4123 & w4118) | (~w4123 & w9154) | (w4118 & w9154);
assign w4445 = ~w4443 & ~w4444;
assign w4446 = w4443 & w4444;
assign w4447 = ~w4445 & ~w4446;
assign w4448 = w4442 & w4447;
assign w4449 = ~w4442 & ~w4447;
assign w4450 = ~w4448 & ~w4449;
assign w4451 = (~w4048 & ~w4050) | (~w4048 & w8624) | (~w4050 & w8624);
assign w4452 = w4051 & ~w4053;
assign w4453 = ~w4055 & ~w4452;
assign w4454 = w4039 & ~w4041;
assign w4455 = ~w4043 & ~w4454;
assign w4456 = ~w4453 & ~w4455;
assign w4457 = w4453 & w4455;
assign w4458 = ~w4456 & ~w4457;
assign w4459 = ~w4451 & w4458;
assign w4460 = w4451 & ~w4458;
assign w4461 = ~w4459 & ~w4460;
assign w4462 = (~w4201 & w4196) | (~w4201 & w9155) | (w4196 & w9155);
assign w4463 = (~w4182 & w4178) | (~w4182 & w9156) | (w4178 & w9156);
assign w4464 = w4462 & w4463;
assign w4465 = ~w4462 & ~w4463;
assign w4466 = ~w4464 & ~w4465;
assign w4467 = w4461 & ~w4466;
assign w4468 = ~w4461 & w4466;
assign w4469 = ~w4467 & ~w4468;
assign w4470 = w4450 & w4469;
assign w4471 = ~w4450 & ~w4469;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = ~w4212 & ~w4215;
assign w4474 = (~w4190 & ~w4192) | (~w4190 & w8948) | (~w4192 & w8948);
assign w4475 = ~w4209 & ~w4474;
assign w4476 = w4209 & w4474;
assign w4477 = ~w4475 & ~w4476;
assign w4478 = ~w4473 & w4477;
assign w4479 = w4473 & ~w4477;
assign w4480 = ~w4478 & ~w4479;
assign w4481 = (~w4146 & ~w4148) | (~w4146 & w8740) | (~w4148 & w8740);
assign w4482 = (~w4087 & ~w4089) | (~w4087 & w9157) | (~w4089 & w9157);
assign w4483 = ~w3913 & ~w4140;
assign w4484 = ~w4141 & ~w4483;
assign w4485 = ~w4482 & w4484;
assign w4486 = w4482 & ~w4484;
assign w4487 = ~w4485 & ~w4486;
assign w4488 = (~w4148 & w8949) | (~w4148 & w8950) | (w8949 & w8950);
assign w4489 = (w4148 & w8951) | (w4148 & w8952) | (w8951 & w8952);
assign w4490 = ~w4488 & ~w4489;
assign w4491 = ~w4480 & ~w4490;
assign w4492 = w4480 & w4490;
assign w4493 = ~w4491 & ~w4492;
assign w4494 = w4472 & ~w4493;
assign w4495 = ~w4472 & w4493;
assign w4496 = ~w4494 & ~w4495;
assign w4497 = w4432 & w4496;
assign w4498 = ~w4432 & ~w4496;
assign w4499 = ~w4497 & ~w4498;
assign w4500 = (~w4175 & ~w4241) | (~w4175 & w8953) | (~w4241 & w8953);
assign w4501 = ~w4168 & ~w4172;
assign w4502 = (~w4237 & ~w4238) | (~w4237 & w8954) | (~w4238 & w8954);
assign w4503 = ~w4501 & w4502;
assign w4504 = w4501 & ~w4502;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = w4500 & w4505;
assign w4507 = ~w4500 & ~w4505;
assign w4508 = ~w4506 & ~w4507;
assign w4509 = (~w4249 & w4246) | (~w4249 & w9158) | (w4246 & w9158);
assign w4510 = w4508 & ~w4509;
assign w4511 = ~w4508 & w4509;
assign w4512 = ~w4510 & ~w4511;
assign w4513 = ~w4499 & w4512;
assign w4514 = w4499 & ~w4512;
assign w4515 = ~w4513 & ~w4514;
assign w4516 = (~w4255 & ~w4257) | (~w4255 & w9159) | (~w4257 & w9159);
assign w4517 = w4515 & w4516;
assign w4518 = ~w4515 & ~w4516;
assign w4519 = ~w4517 & ~w4518;
assign w4520 = (w8732 & w9270) | (w8732 & w9271) | (w9270 & w9271);
assign w4521 = ~w4262 & w9298;
assign w4522 = (~w4010 & w8955) | (~w4010 & w8956) | (w8955 & w8956);
assign w4523 = ~w4519 & ~w4521;
assign w4524 = ~w4522 & ~w4523;
assign w4525 = (w4010 & w9040) | (w4010 & w9041) | (w9040 & w9041);
assign w4526 = (~w4510 & ~w4512) | (~w4510 & w8786) | (~w4512 & w8786);
assign w4527 = pi16 & pi49;
assign w4528 = pi17 & pi48;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = pi17 & pi49;
assign w4531 = w4318 & w4530;
assign w4532 = ~w4529 & ~w4531;
assign w4533 = w4333 & ~w4532;
assign w4534 = ~w4333 & w4532;
assign w4535 = ~w4533 & ~w4534;
assign w4536 = w4349 & ~w4535;
assign w4537 = ~w4349 & w4535;
assign w4538 = ~w4536 & ~w4537;
assign w4539 = pi12 & pi53;
assign w4540 = pi13 & pi52;
assign w4541 = pi14 & pi51;
assign w4542 = ~w4540 & ~w4541;
assign w4543 = pi14 & pi52;
assign w4544 = w4330 & w4543;
assign w4545 = ~w4542 & ~w4544;
assign w4546 = w4539 & ~w4545;
assign w4547 = ~w4539 & w4545;
assign w4548 = ~w4546 & ~w4547;
assign w4549 = w4538 & ~w4548;
assign w4550 = ~w4538 & w4548;
assign w4551 = ~w4549 & ~w4550;
assign w4552 = pi23 & pi42;
assign w4553 = pi24 & pi41;
assign w4554 = ~w4552 & ~w4553;
assign w4555 = pi24 & pi42;
assign w4556 = w4269 & w4555;
assign w4557 = ~w4554 & ~w4556;
assign w4558 = w4284 & ~w4557;
assign w4559 = ~w4284 & w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = w4321 & ~w4560;
assign w4562 = ~w4321 & w4560;
assign w4563 = ~w4561 & ~w4562;
assign w4564 = pi19 & pi46;
assign w4565 = pi20 & pi45;
assign w4566 = pi21 & pi44;
assign w4567 = ~w4565 & ~w4566;
assign w4568 = pi21 & pi45;
assign w4569 = w4281 & w4568;
assign w4570 = ~w4567 & ~w4569;
assign w4571 = w4564 & ~w4570;
assign w4572 = ~w4564 & w4570;
assign w4573 = ~w4571 & ~w4572;
assign w4574 = w4563 & ~w4573;
assign w4575 = ~w4563 & w4573;
assign w4576 = ~w4574 & ~w4575;
assign w4577 = pi31 & pi34;
assign w4578 = pi30 & pi35;
assign w4579 = ~w4577 & w4578;
assign w4580 = w4577 & ~w4578;
assign w4581 = ~w4579 & ~w4580;
assign w4582 = w4305 & w4581;
assign w4583 = ~w4305 & ~w4581;
assign w4584 = ~w4582 & ~w4583;
assign w4585 = w4272 & w4584;
assign w4586 = ~w4272 & ~w4584;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = pi26 & pi39;
assign w4589 = pi27 & pi38;
assign w4590 = pi28 & pi37;
assign w4591 = ~w4589 & ~w4590;
assign w4592 = pi28 & pi38;
assign w4593 = w4302 & w4592;
assign w4594 = ~w4591 & ~w4593;
assign w4595 = w4588 & ~w4594;
assign w4596 = ~w4588 & w4594;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = w4587 & ~w4597;
assign w4599 = ~w4587 & w4597;
assign w4600 = ~w4598 & ~w4599;
assign w4601 = w4576 & w4600;
assign w4602 = ~w4576 & ~w4600;
assign w4603 = ~w4601 & ~w4602;
assign w4604 = w4551 & w4603;
assign w4605 = ~w4551 & ~w4603;
assign w4606 = ~w4604 & ~w4605;
assign w4607 = pi09 & pi56;
assign w4608 = pi10 & pi55;
assign w4609 = ~w4607 & ~w4608;
assign w4610 = pi10 & pi56;
assign w4611 = w4346 & w4610;
assign w4612 = ~w4609 & ~w4611;
assign w4613 = w4361 & ~w4612;
assign w4614 = ~w4361 & w4612;
assign w4615 = ~w4613 & ~w4614;
assign w4616 = w4414 & ~w4615;
assign w4617 = ~w4414 & w4615;
assign w4618 = ~w4616 & ~w4617;
assign w4619 = pi05 & pi60;
assign w4620 = pi06 & pi59;
assign w4621 = pi07 & pi58;
assign w4622 = ~w4620 & ~w4621;
assign w4623 = pi07 & pi59;
assign w4624 = w4358 & w4623;
assign w4625 = ~w4622 & ~w4624;
assign w4626 = w4619 & ~w4625;
assign w4627 = ~w4619 & w4625;
assign w4628 = ~w4626 & ~w4627;
assign w4629 = w4618 & ~w4628;
assign w4630 = ~w4618 & w4628;
assign w4631 = ~w4629 & ~w4630;
assign w4632 = w4415 & w4420;
assign w4633 = ~w4415 & ~w4420;
assign w4634 = ~w4632 & ~w4633;
assign w4635 = ~w4417 & ~w4634;
assign w4636 = (~w4355 & ~w4357) | (~w4355 & w8741) | (~w4357 & w8741);
assign w4637 = w4358 & ~w4360;
assign w4638 = ~w4362 & ~w4637;
assign w4639 = w4346 & ~w4348;
assign w4640 = ~w4350 & ~w4639;
assign w4641 = ~w4638 & ~w4640;
assign w4642 = w4638 & w4640;
assign w4643 = ~w4641 & ~w4642;
assign w4644 = ~w4636 & w4643;
assign w4645 = w4636 & ~w4643;
assign w4646 = ~w4644 & ~w4645;
assign w4647 = (~w4327 & ~w4329) | (~w4327 & w8742) | (~w4329 & w8742);
assign w4648 = w4330 & ~w4332;
assign w4649 = ~w4334 & ~w4648;
assign w4650 = w4318 & ~w4320;
assign w4651 = ~w4322 & ~w4650;
assign w4652 = ~w4649 & ~w4651;
assign w4653 = w4649 & w4651;
assign w4654 = ~w4652 & ~w4653;
assign w4655 = ~w4647 & w4654;
assign w4656 = w4647 & ~w4654;
assign w4657 = ~w4655 & ~w4656;
assign w4658 = w4646 & w4657;
assign w4659 = ~w4646 & ~w4657;
assign w4660 = ~w4658 & ~w4659;
assign w4661 = ~w4635 & w4660;
assign w4662 = w4635 & ~w4660;
assign w4663 = ~w4661 & ~w4662;
assign w4664 = ~w4631 & ~w4663;
assign w4665 = w4631 & w4663;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = ~w4606 & w4666;
assign w4668 = w4606 & ~w4666;
assign w4669 = ~w4667 & ~w4668;
assign w4670 = pi02 & pi63;
assign w4671 = pi03 & pi62;
assign w4672 = w4670 & ~w4671;
assign w4673 = ~w4670 & w4671;
assign w4674 = ~w4672 & ~w4673;
assign w4675 = (~w4674 & w8787) | (~w4674 & w4478) | (w8787 & w4478);
assign w4676 = (w8788 & w4473) | (w8788 & w8957) | (w4473 & w8957);
assign w4677 = ~w4675 & ~w4676;
assign w4678 = (~w4485 & ~w4481) | (~w4485 & w8789) | (~w4481 & w8789);
assign w4679 = w4677 & ~w4678;
assign w4680 = ~w4677 & w4678;
assign w4681 = ~w4679 & ~w4680;
assign w4682 = ~w4669 & w4681;
assign w4683 = w4669 & ~w4681;
assign w4684 = ~w4682 & ~w4683;
assign w4685 = ~w4299 & ~w4311;
assign w4686 = w4302 & ~w4304;
assign w4687 = ~w4306 & ~w4686;
assign w4688 = ~w4296 & ~w4687;
assign w4689 = w4296 & w4687;
assign w4690 = ~w4688 & ~w4689;
assign w4691 = ~w4685 & w4690;
assign w4692 = w4685 & ~w4690;
assign w4693 = ~w4691 & ~w4692;
assign w4694 = (~w4375 & w4370) | (~w4375 & w8958) | (w4370 & w8958);
assign w4695 = w4398 & ~w4694;
assign w4696 = ~w4398 & w4694;
assign w4697 = ~w4695 & ~w4696;
assign w4698 = w4693 & w4697;
assign w4699 = ~w4693 & ~w4697;
assign w4700 = ~w4698 & ~w4699;
assign w4701 = (~w4278 & ~w4280) | (~w4278 & w8625) | (~w4280 & w8625);
assign w4702 = w4281 & ~w4283;
assign w4703 = ~w4285 & ~w4702;
assign w4704 = w4269 & ~w4271;
assign w4705 = ~w4273 & ~w4704;
assign w4706 = ~w4703 & ~w4705;
assign w4707 = w4703 & w4705;
assign w4708 = ~w4706 & ~w4707;
assign w4709 = ~w4701 & w4708;
assign w4710 = w4701 & ~w4708;
assign w4711 = ~w4709 & ~w4710;
assign w4712 = ~w4386 & ~w4389;
assign w4713 = (~w4437 & w4433) | (~w4437 & w8743) | (w4433 & w8743);
assign w4714 = (~w4456 & w4451) | (~w4456 & w8744) | (w4451 & w8744);
assign w4715 = ~w4713 & ~w4714;
assign w4716 = w4713 & w4714;
assign w4717 = ~w4715 & ~w4716;
assign w4718 = ~w4712 & w4717;
assign w4719 = w4712 & ~w4717;
assign w4720 = ~w4718 & ~w4719;
assign w4721 = w4711 & w4720;
assign w4722 = ~w4711 & ~w4720;
assign w4723 = ~w4721 & ~w4722;
assign w4724 = w4700 & w4723;
assign w4725 = ~w4700 & ~w4723;
assign w4726 = ~w4724 & ~w4725;
assign w4727 = ~w4467 & ~w4470;
assign w4728 = (~w4445 & ~w4447) | (~w4445 & w8790) | (~w4447 & w8790);
assign w4729 = ~w4464 & ~w4728;
assign w4730 = w4464 & w4728;
assign w4731 = ~w4729 & ~w4730;
assign w4732 = ~w4727 & w4731;
assign w4733 = w4727 & ~w4731;
assign w4734 = ~w4732 & ~w4733;
assign w4735 = (~w4404 & ~w4406) | (~w4404 & w8745) | (~w4406 & w8745);
assign w4736 = ~w4314 & ~w4342;
assign w4737 = ~w4392 & ~w4401;
assign w4738 = ~w4736 & ~w4737;
assign w4739 = w4736 & w4737;
assign w4740 = ~w4738 & ~w4739;
assign w4741 = ~w4735 & w4740;
assign w4742 = w4735 & ~w4740;
assign w4743 = ~w4741 & ~w4742;
assign w4744 = w4734 & w4743;
assign w4745 = ~w4734 & ~w4743;
assign w4746 = ~w4744 & ~w4745;
assign w4747 = w4726 & ~w4746;
assign w4748 = ~w4726 & w4746;
assign w4749 = ~w4747 & ~w4748;
assign w4750 = w4684 & ~w4749;
assign w4751 = ~w4684 & w4749;
assign w4752 = ~w4750 & ~w4751;
assign w4753 = (~w4503 & ~w4500) | (~w4503 & w9160) | (~w4500 & w9160);
assign w4754 = ~w4430 & ~w4497;
assign w4755 = ~w4423 & ~w4427;
assign w4756 = (~w4491 & ~w4493) | (~w4491 & w8791) | (~w4493 & w8791);
assign w4757 = ~w4755 & w4756;
assign w4758 = w4755 & ~w4756;
assign w4759 = ~w4757 & ~w4758;
assign w4760 = w4754 & w4759;
assign w4761 = ~w4754 & ~w4759;
assign w4762 = ~w4760 & ~w4761;
assign w4763 = ~w4753 & w4762;
assign w4764 = w4753 & ~w4762;
assign w4765 = ~w4763 & ~w4764;
assign w4766 = w4752 & w4765;
assign w4767 = ~w4752 & ~w4765;
assign w4768 = ~w4766 & ~w4767;
assign w4769 = w4526 & ~w4768;
assign w4770 = ~w4526 & w4768;
assign w4771 = ~w4769 & ~w4770;
assign w4772 = w4525 & ~w4771;
assign w4773 = ~w4525 & w4771;
assign w4774 = ~w4772 & ~w4773;
assign w4775 = (~w4763 & ~w4765) | (~w4763 & w8792) | (~w4765 & w8792);
assign w4776 = pi11 & pi55;
assign w4777 = pi15 & pi51;
assign w4778 = pi16 & pi50;
assign w4779 = ~w4530 & ~w4778;
assign w4780 = pi17 & pi50;
assign w4781 = w4527 & w4780;
assign w4782 = ~w4779 & ~w4781;
assign w4783 = w4777 & ~w4782;
assign w4784 = ~w4777 & w4782;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = w4776 & ~w4785;
assign w4787 = ~w4776 & w4785;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = pi12 & pi54;
assign w4790 = pi13 & pi53;
assign w4791 = ~w4543 & ~w4790;
assign w4792 = pi14 & pi53;
assign w4793 = w4540 & w4792;
assign w4794 = ~w4791 & ~w4793;
assign w4795 = w4789 & ~w4794;
assign w4796 = ~w4789 & w4794;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = w4788 & ~w4797;
assign w4799 = ~w4788 & w4797;
assign w4800 = ~w4798 & ~w4799;
assign w4801 = pi18 & pi48;
assign w4802 = pi22 & pi44;
assign w4803 = pi23 & pi43;
assign w4804 = ~w4555 & ~w4803;
assign w4805 = pi24 & pi43;
assign w4806 = w4552 & w4805;
assign w4807 = ~w4804 & ~w4806;
assign w4808 = w4802 & ~w4807;
assign w4809 = ~w4802 & w4807;
assign w4810 = ~w4808 & ~w4809;
assign w4811 = w4801 & ~w4810;
assign w4812 = ~w4801 & w4810;
assign w4813 = ~w4811 & ~w4812;
assign w4814 = pi19 & pi47;
assign w4815 = pi20 & pi46;
assign w4816 = ~w4568 & ~w4815;
assign w4817 = pi21 & pi46;
assign w4818 = w4565 & w4817;
assign w4819 = ~w4816 & ~w4818;
assign w4820 = w4814 & ~w4819;
assign w4821 = ~w4814 & w4819;
assign w4822 = ~w4820 & ~w4821;
assign w4823 = w4813 & ~w4822;
assign w4824 = ~w4813 & w4822;
assign w4825 = ~w4823 & ~w4824;
assign w4826 = pi25 & pi41;
assign w4827 = pi29 & pi37;
assign w4828 = pi31 & pi35;
assign w4829 = pi30 & pi36;
assign w4830 = ~w4828 & w4829;
assign w4831 = w4828 & ~w4829;
assign w4832 = ~w4830 & ~w4831;
assign w4833 = w4827 & w4832;
assign w4834 = ~w4827 & ~w4832;
assign w4835 = ~w4833 & ~w4834;
assign w4836 = w4826 & w4835;
assign w4837 = ~w4826 & ~w4835;
assign w4838 = ~w4836 & ~w4837;
assign w4839 = pi26 & pi40;
assign w4840 = pi27 & pi39;
assign w4841 = ~w4592 & ~w4840;
assign w4842 = pi28 & pi39;
assign w4843 = w4589 & w4842;
assign w4844 = ~w4841 & ~w4843;
assign w4845 = w4839 & ~w4844;
assign w4846 = ~w4839 & w4844;
assign w4847 = ~w4845 & ~w4846;
assign w4848 = w4838 & ~w4847;
assign w4849 = ~w4838 & w4847;
assign w4850 = ~w4848 & ~w4849;
assign w4851 = w4825 & w4850;
assign w4852 = ~w4825 & ~w4850;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = w4800 & w4853;
assign w4855 = ~w4800 & ~w4853;
assign w4856 = ~w4854 & ~w4855;
assign w4857 = (~w4616 & ~w4618) | (~w4616 & w8746) | (~w4618 & w8746);
assign w4858 = w4619 & ~w4622;
assign w4859 = ~w4624 & ~w4858;
assign w4860 = w4361 & ~w4609;
assign w4861 = ~w4611 & ~w4860;
assign w4862 = ~w4859 & ~w4861;
assign w4863 = w4859 & w4861;
assign w4864 = ~w4862 & ~w4863;
assign w4865 = ~w4857 & w4864;
assign w4866 = w4857 & ~w4864;
assign w4867 = ~w4865 & ~w4866;
assign w4868 = (~w4536 & ~w4538) | (~w4536 & w8626) | (~w4538 & w8626);
assign w4869 = w4539 & ~w4542;
assign w4870 = ~w4544 & ~w4869;
assign w4871 = w4333 & ~w4529;
assign w4872 = ~w4531 & ~w4871;
assign w4873 = ~w4870 & ~w4872;
assign w4874 = w4870 & w4872;
assign w4875 = ~w4873 & ~w4874;
assign w4876 = ~w4868 & w4875;
assign w4877 = w4868 & ~w4875;
assign w4878 = ~w4876 & ~w4877;
assign w4879 = w4867 & w4878;
assign w4880 = ~w4867 & ~w4878;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = ~w4672 & w4881;
assign w4883 = w4672 & ~w4881;
assign w4884 = ~w4882 & ~w4883;
assign w4885 = pi04 & pi62;
assign w4886 = pi08 & pi58;
assign w4887 = pi09 & pi57;
assign w4888 = ~w4610 & ~w4887;
assign w4889 = pi10 & pi57;
assign w4890 = w4607 & w4889;
assign w4891 = ~w4888 & ~w4890;
assign w4892 = w4886 & ~w4891;
assign w4893 = ~w4886 & w4891;
assign w4894 = ~w4892 & ~w4893;
assign w4895 = w4885 & ~w4894;
assign w4896 = ~w4885 & w4894;
assign w4897 = ~w4895 & ~w4896;
assign w4898 = pi05 & pi61;
assign w4899 = pi06 & pi60;
assign w4900 = ~w4623 & ~w4899;
assign w4901 = pi07 & pi60;
assign w4902 = w4620 & w4901;
assign w4903 = ~w4900 & ~w4902;
assign w4904 = w4898 & ~w4903;
assign w4905 = ~w4898 & w4903;
assign w4906 = ~w4904 & ~w4905;
assign w4907 = w4897 & ~w4906;
assign w4908 = ~w4897 & w4906;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = w4884 & w4909;
assign w4911 = ~w4884 & ~w4909;
assign w4912 = ~w4910 & ~w4911;
assign w4913 = w4856 & w4912;
assign w4914 = ~w4856 & ~w4912;
assign w4915 = ~w4913 & ~w4914;
assign w4916 = (~w4738 & w4735) | (~w4738 & w9042) | (w4735 & w9042);
assign w4917 = pi03 & pi63;
assign w4918 = (~w4729 & w4727) | (~w4729 & w8793) | (w4727 & w8793);
assign w4919 = w4917 & ~w4918;
assign w4920 = ~w4917 & w4918;
assign w4921 = ~w4919 & ~w4920;
assign w4922 = ~w4916 & w4921;
assign w4923 = w4916 & ~w4921;
assign w4924 = ~w4922 & ~w4923;
assign w4925 = w4915 & w4924;
assign w4926 = ~w4915 & ~w4924;
assign w4927 = ~w4925 & ~w4926;
assign w4928 = (~w4585 & ~w4587) | (~w4585 & w8627) | (~w4587 & w8627);
assign w4929 = (~w4579 & ~w4581) | (~w4579 & w8794) | (~w4581 & w8794);
assign w4930 = w4588 & ~w4591;
assign w4931 = ~w4593 & ~w4930;
assign w4932 = ~w4929 & ~w4931;
assign w4933 = w4929 & w4931;
assign w4934 = ~w4932 & ~w4933;
assign w4935 = ~w4928 & w4934;
assign w4936 = w4928 & ~w4934;
assign w4937 = ~w4935 & ~w4936;
assign w4938 = (~w4641 & w4636) | (~w4641 & w9043) | (w4636 & w9043);
assign w4939 = w4632 & ~w4938;
assign w4940 = ~w4632 & w4938;
assign w4941 = ~w4939 & ~w4940;
assign w4942 = w4937 & w4941;
assign w4943 = ~w4937 & ~w4941;
assign w4944 = ~w4942 & ~w4943;
assign w4945 = (~w4561 & ~w4563) | (~w4561 & w8628) | (~w4563 & w8628);
assign w4946 = w4564 & ~w4567;
assign w4947 = ~w4569 & ~w4946;
assign w4948 = w4284 & ~w4554;
assign w4949 = ~w4556 & ~w4948;
assign w4950 = ~w4947 & ~w4949;
assign w4951 = w4947 & w4949;
assign w4952 = ~w4950 & ~w4951;
assign w4953 = ~w4945 & w4952;
assign w4954 = w4945 & ~w4952;
assign w4955 = ~w4953 & ~w4954;
assign w4956 = ~w4652 & ~w4655;
assign w4957 = (~w4688 & w4685) | (~w4688 & w8795) | (w4685 & w8795);
assign w4958 = (~w4706 & w4701) | (~w4706 & w8747) | (w4701 & w8747);
assign w4959 = ~w4957 & ~w4958;
assign w4960 = w4957 & w4958;
assign w4961 = ~w4959 & ~w4960;
assign w4962 = ~w4956 & w4961;
assign w4963 = w4956 & ~w4961;
assign w4964 = ~w4962 & ~w4963;
assign w4965 = w4955 & w4964;
assign w4966 = ~w4955 & ~w4964;
assign w4967 = ~w4965 & ~w4966;
assign w4968 = w4944 & w4967;
assign w4969 = ~w4944 & ~w4967;
assign w4970 = ~w4968 & ~w4969;
assign w4971 = (~w4721 & ~w4723) | (~w4721 & w8796) | (~w4723 & w8796);
assign w4972 = (~w4695 & ~w4697) | (~w4695 & w9044) | (~w4697 & w9044);
assign w4973 = (~w4715 & ~w4717) | (~w4715 & w9045) | (~w4717 & w9045);
assign w4974 = ~w4972 & ~w4973;
assign w4975 = w4972 & w4973;
assign w4976 = ~w4974 & ~w4975;
assign w4977 = ~w4971 & w4976;
assign w4978 = w4971 & ~w4976;
assign w4979 = ~w4977 & ~w4978;
assign w4980 = (~w4664 & ~w4666) | (~w4664 & w8797) | (~w4666 & w8797);
assign w4981 = ~w4601 & ~w4604;
assign w4982 = ~w4658 & ~w4661;
assign w4983 = ~w4981 & ~w4982;
assign w4984 = w4981 & w4982;
assign w4985 = ~w4983 & ~w4984;
assign w4986 = w4980 & w4985;
assign w4987 = ~w4980 & ~w4985;
assign w4988 = ~w4986 & ~w4987;
assign w4989 = ~w4979 & ~w4988;
assign w4990 = w4979 & w4988;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = w4970 & w4991;
assign w4993 = ~w4970 & ~w4991;
assign w4994 = ~w4992 & ~w4993;
assign w4995 = w4927 & w4994;
assign w4996 = ~w4927 & ~w4994;
assign w4997 = ~w4995 & ~w4996;
assign w4998 = (~w4757 & ~w4754) | (~w4757 & w8798) | (~w4754 & w8798);
assign w4999 = (~w4682 & w4749) | (~w4682 & w8799) | (w4749 & w8799);
assign w5000 = (~w4675 & w4678) | (~w4675 & w9046) | (w4678 & w9046);
assign w5001 = ~w5000 & w9299;
assign w5002 = (w4746 & w8959) | (w4746 & w8960) | (w8959 & w8960);
assign w5003 = ~w5001 & ~w5002;
assign w5004 = ~w4999 & w5003;
assign w5005 = w4999 & ~w5003;
assign w5006 = ~w5004 & ~w5005;
assign w5007 = ~w4998 & w5006;
assign w5008 = w4998 & ~w5006;
assign w5009 = ~w5007 & ~w5008;
assign w5010 = w4997 & w5009;
assign w5011 = ~w4997 & ~w5009;
assign w5012 = ~w5010 & ~w5011;
assign w5013 = ~w4775 & w5012;
assign w5014 = w4775 & ~w5012;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = (~w4769 & w9047) | (~w4769 & ~w4525) | (w9047 & ~w4525);
assign w5017 = (~w4010 & w9272) | (~w4010 & w9273) | (w9272 & w9273);
assign w5018 = ~w5015 & ~w5016;
assign w5019 = ~w5017 & ~w5018;
assign w5020 = ~w5013 & ~w5017;
assign w5021 = (~w5007 & ~w5009) | (~w5007 & w8961) | (~w5009 & w8961);
assign w5022 = (~w5001 & w4999) | (~w5001 & w8962) | (w4999 & w8962);
assign w5023 = ~w4862 & ~w4865;
assign w5024 = (~w4950 & w4945) | (~w4950 & w8748) | (w4945 & w8748);
assign w5025 = (~w4873 & w4868) | (~w4873 & w8749) | (w4868 & w8749);
assign w5026 = ~w5024 & ~w5025;
assign w5027 = w5024 & w5025;
assign w5028 = ~w5026 & ~w5027;
assign w5029 = ~w5023 & w5028;
assign w5030 = w5023 & ~w5028;
assign w5031 = ~w5029 & ~w5030;
assign w5032 = (~w4836 & ~w4838) | (~w4836 & w8629) | (~w4838 & w8629);
assign w5033 = ~w4830 & ~w4833;
assign w5034 = w4839 & ~w4841;
assign w5035 = ~w4843 & ~w5034;
assign w5036 = ~w5033 & ~w5035;
assign w5037 = w5033 & w5035;
assign w5038 = ~w5036 & ~w5037;
assign w5039 = ~w5032 & w5038;
assign w5040 = w5032 & ~w5038;
assign w5041 = ~w5039 & ~w5040;
assign w5042 = pi04 & pi63;
assign w5043 = (w4928 & w8801) | (w4928 & w8802) | (w8801 & w8802);
assign w5044 = ~w5042 & w9300;
assign w5045 = ~w5043 & ~w5044;
assign w5046 = w5041 & ~w5045;
assign w5047 = ~w5041 & w5045;
assign w5048 = ~w5046 & ~w5047;
assign w5049 = w5031 & w5048;
assign w5050 = ~w5031 & ~w5048;
assign w5051 = ~w5049 & ~w5050;
assign w5052 = (~w4910 & ~w4912) | (~w4910 & w8803) | (~w4912 & w8803);
assign w5053 = ~w4851 & ~w4854;
assign w5054 = ~w4879 & ~w4882;
assign w5055 = ~w5053 & ~w5054;
assign w5056 = w5053 & w5054;
assign w5057 = ~w5055 & ~w5056;
assign w5058 = ~w5052 & w5057;
assign w5059 = w5052 & ~w5057;
assign w5060 = ~w5058 & ~w5059;
assign w5061 = (~w4965 & ~w4967) | (~w4965 & w8804) | (~w4967 & w8804);
assign w5062 = ~w4939 & ~w4942;
assign w5063 = ~w4959 & ~w4962;
assign w5064 = ~w5062 & ~w5063;
assign w5065 = w5062 & w5063;
assign w5066 = ~w5064 & ~w5065;
assign w5067 = ~w5061 & w5066;
assign w5068 = w5061 & ~w5066;
assign w5069 = ~w5067 & ~w5068;
assign w5070 = w5060 & w5069;
assign w5071 = ~w5060 & ~w5069;
assign w5072 = ~w5070 & ~w5071;
assign w5073 = w5051 & w5072;
assign w5074 = ~w5051 & ~w5072;
assign w5075 = ~w5073 & ~w5074;
assign w5076 = pi25 & pi42;
assign w5077 = pi29 & pi38;
assign w5078 = pi31 & pi36;
assign w5079 = pi30 & pi37;
assign w5080 = ~w5078 & w5079;
assign w5081 = w5078 & ~w5079;
assign w5082 = ~w5080 & ~w5081;
assign w5083 = w5077 & w5082;
assign w5084 = ~w5077 & ~w5082;
assign w5085 = ~w5083 & ~w5084;
assign w5086 = w5076 & w5085;
assign w5087 = ~w5076 & ~w5085;
assign w5088 = ~w5086 & ~w5087;
assign w5089 = pi26 & pi41;
assign w5090 = pi27 & pi40;
assign w5091 = ~w4842 & ~w5090;
assign w5092 = pi28 & pi40;
assign w5093 = w4840 & w5092;
assign w5094 = ~w5091 & ~w5093;
assign w5095 = w5089 & ~w5094;
assign w5096 = ~w5089 & w5094;
assign w5097 = ~w5095 & ~w5096;
assign w5098 = w5088 & ~w5097;
assign w5099 = ~w5088 & w5097;
assign w5100 = ~w5098 & ~w5099;
assign w5101 = ~w4917 & w5100;
assign w5102 = w4917 & ~w5100;
assign w5103 = ~w5101 & ~w5102;
assign w5104 = pi18 & pi49;
assign w5105 = pi22 & pi45;
assign w5106 = pi23 & pi44;
assign w5107 = ~w4805 & ~w5106;
assign w5108 = pi24 & pi44;
assign w5109 = w4803 & w5108;
assign w5110 = ~w5107 & ~w5109;
assign w5111 = w5105 & ~w5110;
assign w5112 = ~w5105 & w5110;
assign w5113 = ~w5111 & ~w5112;
assign w5114 = w5104 & ~w5113;
assign w5115 = ~w5104 & w5113;
assign w5116 = ~w5114 & ~w5115;
assign w5117 = pi19 & pi48;
assign w5118 = pi20 & pi47;
assign w5119 = ~w4817 & ~w5118;
assign w5120 = pi21 & pi47;
assign w5121 = w4815 & w5120;
assign w5122 = ~w5119 & ~w5121;
assign w5123 = w5117 & ~w5122;
assign w5124 = ~w5117 & w5122;
assign w5125 = ~w5123 & ~w5124;
assign w5126 = w5116 & ~w5125;
assign w5127 = ~w5116 & w5125;
assign w5128 = ~w5126 & ~w5127;
assign w5129 = w5103 & w5128;
assign w5130 = ~w5103 & ~w5128;
assign w5131 = ~w5129 & ~w5130;
assign w5132 = pi11 & pi56;
assign w5133 = pi15 & pi52;
assign w5134 = pi16 & pi51;
assign w5135 = ~w4780 & ~w5134;
assign w5136 = pi17 & pi51;
assign w5137 = w4778 & w5136;
assign w5138 = ~w5135 & ~w5137;
assign w5139 = w5133 & ~w5138;
assign w5140 = ~w5133 & w5138;
assign w5141 = ~w5139 & ~w5140;
assign w5142 = w5132 & ~w5141;
assign w5143 = ~w5132 & w5141;
assign w5144 = ~w5142 & ~w5143;
assign w5145 = pi12 & pi55;
assign w5146 = pi13 & pi54;
assign w5147 = ~w4792 & ~w5146;
assign w5148 = pi14 & pi54;
assign w5149 = w4790 & w5148;
assign w5150 = ~w5147 & ~w5149;
assign w5151 = w5145 & ~w5150;
assign w5152 = ~w5145 & w5150;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = w5144 & ~w5153;
assign w5155 = ~w5144 & w5153;
assign w5156 = ~w5154 & ~w5155;
assign w5157 = ~w4895 & ~w4907;
assign w5158 = w4898 & ~w4900;
assign w5159 = ~w4902 & ~w5158;
assign w5160 = w4886 & ~w4888;
assign w5161 = ~w4890 & ~w5160;
assign w5162 = ~w5159 & ~w5161;
assign w5163 = w5159 & w5161;
assign w5164 = ~w5162 & ~w5163;
assign w5165 = ~w5157 & w5164;
assign w5166 = w5157 & ~w5164;
assign w5167 = ~w5165 & ~w5166;
assign w5168 = (~w4786 & ~w4788) | (~w4786 & w8630) | (~w4788 & w8630);
assign w5169 = w4789 & ~w4791;
assign w5170 = ~w4793 & ~w5169;
assign w5171 = w4777 & ~w4779;
assign w5172 = ~w4781 & ~w5171;
assign w5173 = ~w5170 & ~w5172;
assign w5174 = w5170 & w5172;
assign w5175 = ~w5173 & ~w5174;
assign w5176 = ~w5168 & w5175;
assign w5177 = w5168 & ~w5175;
assign w5178 = ~w5176 & ~w5177;
assign w5179 = (~w4811 & ~w4813) | (~w4811 & w8631) | (~w4813 & w8631);
assign w5180 = w4814 & ~w4816;
assign w5181 = ~w4818 & ~w5180;
assign w5182 = w4802 & ~w4804;
assign w5183 = ~w4806 & ~w5182;
assign w5184 = ~w5181 & ~w5183;
assign w5185 = w5181 & w5183;
assign w5186 = ~w5184 & ~w5185;
assign w5187 = ~w5179 & w5186;
assign w5188 = w5179 & ~w5186;
assign w5189 = ~w5187 & ~w5188;
assign w5190 = w5178 & w5189;
assign w5191 = ~w5178 & ~w5189;
assign w5192 = ~w5190 & ~w5191;
assign w5193 = w5167 & w5192;
assign w5194 = ~w5167 & ~w5192;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = ~w5156 & ~w5195;
assign w5197 = w5156 & w5195;
assign w5198 = ~w5196 & ~w5197;
assign w5199 = ~w5131 & w5198;
assign w5200 = w5131 & ~w5198;
assign w5201 = ~w5199 & ~w5200;
assign w5202 = (~w4983 & ~w4980) | (~w4983 & w9048) | (~w4980 & w9048);
assign w5203 = pi08 & pi59;
assign w5204 = pi09 & pi58;
assign w5205 = ~w4889 & ~w5204;
assign w5206 = pi10 & pi58;
assign w5207 = w4887 & w5206;
assign w5208 = ~w5205 & ~w5207;
assign w5209 = w5203 & ~w5208;
assign w5210 = ~w5203 & w5208;
assign w5211 = ~w5209 & ~w5210;
assign w5212 = pi05 & pi62;
assign w5213 = pi06 & pi61;
assign w5214 = ~w4901 & ~w5213;
assign w5215 = pi07 & pi61;
assign w5216 = w4899 & w5215;
assign w5217 = ~w5214 & ~w5216;
assign w5218 = w5212 & ~w5217;
assign w5219 = ~w5212 & w5217;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = ~w5211 & ~w5220;
assign w5222 = w5211 & w5220;
assign w5223 = ~w5221 & ~w5222;
assign w5224 = (w4971 & w9049) | (w4971 & w9050) | (w9049 & w9050);
assign w5225 = w5223 & w9301;
assign w5226 = ~w5224 & ~w5225;
assign w5227 = w5202 & w5226;
assign w5228 = ~w5202 & ~w5226;
assign w5229 = ~w5227 & ~w5228;
assign w5230 = ~w5201 & ~w5229;
assign w5231 = w5201 & w5229;
assign w5232 = ~w5230 & ~w5231;
assign w5233 = w5075 & w5232;
assign w5234 = ~w5075 & ~w5232;
assign w5235 = ~w5233 & ~w5234;
assign w5236 = ~w5022 & w5235;
assign w5237 = w5022 & ~w5235;
assign w5238 = ~w5236 & ~w5237;
assign w5239 = (~w4925 & ~w4994) | (~w4925 & w9163) | (~w4994 & w9163);
assign w5240 = ~w4919 & ~w4922;
assign w5241 = (~w4990 & ~w4991) | (~w4990 & w9051) | (~w4991 & w9051);
assign w5242 = ~w5240 & ~w5241;
assign w5243 = w5240 & w5241;
assign w5244 = ~w5242 & ~w5243;
assign w5245 = w5239 & ~w5244;
assign w5246 = ~w5239 & w5244;
assign w5247 = ~w5245 & ~w5246;
assign w5248 = w5238 & ~w5247;
assign w5249 = ~w5238 & w5247;
assign w5250 = ~w5248 & ~w5249;
assign w5251 = ~w5021 & ~w5250;
assign w5252 = w5021 & w5250;
assign w5253 = ~w5251 & ~w5252;
assign w5254 = w5020 & ~w5253;
assign w5255 = ~w5020 & w5253;
assign w5256 = ~w5254 & ~w5255;
assign w5257 = ~w5014 & w5253;
assign w5258 = ~w4770 & ~w5013;
assign w5259 = w4519 & ~w4769;
assign w5260 = w5259 & w8805;
assign w5261 = w4517 & ~w4769;
assign w5262 = w5258 & ~w5261;
assign w5263 = (~w5251 & w5262) | (~w5251 & w8806) | (w5262 & w8806);
assign w5264 = (w4010 & w8964) | (w4010 & w8965) | (w8964 & w8965);
assign w5265 = pi05 & pi63;
assign w5266 = pi06 & pi62;
assign w5267 = w5265 & ~w5266;
assign w5268 = ~w5265 & w5266;
assign w5269 = ~w5267 & ~w5268;
assign w5270 = (~w5269 & w5165) | (~w5269 & w8966) | (w5165 & w8966);
assign w5271 = ~w5165 & w8967;
assign w5272 = ~w5270 & ~w5271;
assign w5273 = ~w5173 & ~w5176;
assign w5274 = (~w5036 & w5032) | (~w5036 & w8807) | (w5032 & w8807);
assign w5275 = (~w5184 & w5179) | (~w5184 & w8808) | (w5179 & w8808);
assign w5276 = ~w5274 & ~w5275;
assign w5277 = w5274 & w5275;
assign w5278 = ~w5276 & ~w5277;
assign w5279 = ~w5273 & w5278;
assign w5280 = w5273 & ~w5278;
assign w5281 = ~w5279 & ~w5280;
assign w5282 = w5272 & w5281;
assign w5283 = ~w5272 & ~w5281;
assign w5284 = ~w5282 & ~w5283;
assign w5285 = (~w5046 & ~w5031) | (~w5046 & w8809) | (~w5031 & w8809);
assign w5286 = (~w5026 & ~w5028) | (~w5026 & w8810) | (~w5028 & w8810);
assign w5287 = ~w5043 & ~w5286;
assign w5288 = w5043 & w5286;
assign w5289 = ~w5287 & ~w5288;
assign w5290 = ~w5285 & w5289;
assign w5291 = w5285 & ~w5289;
assign w5292 = ~w5290 & ~w5291;
assign w5293 = (~w5196 & ~w5198) | (~w5196 & w8751) | (~w5198 & w8751);
assign w5294 = ~w5101 & ~w5129;
assign w5295 = (~w5190 & ~w5192) | (~w5190 & w8968) | (~w5192 & w8968);
assign w5296 = ~w5294 & ~w5295;
assign w5297 = w5294 & w5295;
assign w5298 = ~w5296 & ~w5297;
assign w5299 = w5298 & w5293;
assign w5300 = (w5198 & w9274) | (w5198 & w9275) | (w9274 & w9275);
assign w5301 = ~w5299 & ~w5300;
assign w5302 = w5292 & w5301;
assign w5303 = ~w5292 & ~w5301;
assign w5304 = ~w5302 & ~w5303;
assign w5305 = w5284 & w5304;
assign w5306 = ~w5284 & ~w5304;
assign w5307 = ~w5305 & ~w5306;
assign w5308 = pi18 & pi50;
assign w5309 = pi22 & pi46;
assign w5310 = pi23 & pi45;
assign w5311 = ~w5108 & ~w5310;
assign w5312 = pi24 & pi45;
assign w5313 = w5106 & w5312;
assign w5314 = ~w5311 & ~w5313;
assign w5315 = w5309 & ~w5314;
assign w5316 = ~w5309 & w5314;
assign w5317 = ~w5315 & ~w5316;
assign w5318 = w5308 & ~w5317;
assign w5319 = ~w5308 & w5317;
assign w5320 = ~w5318 & ~w5319;
assign w5321 = pi19 & pi49;
assign w5322 = pi20 & pi48;
assign w5323 = ~w5120 & ~w5322;
assign w5324 = pi21 & pi48;
assign w5325 = w5118 & w5324;
assign w5326 = ~w5323 & ~w5325;
assign w5327 = w5321 & ~w5326;
assign w5328 = ~w5321 & w5326;
assign w5329 = ~w5327 & ~w5328;
assign w5330 = w5320 & ~w5329;
assign w5331 = ~w5320 & w5329;
assign w5332 = ~w5330 & ~w5331;
assign w5333 = w5212 & ~w5214;
assign w5334 = ~w5216 & ~w5333;
assign w5335 = w5203 & ~w5205;
assign w5336 = ~w5207 & ~w5335;
assign w5337 = ~w5334 & ~w5336;
assign w5338 = w5334 & w5336;
assign w5339 = ~w5337 & ~w5338;
assign w5340 = w5221 & w5339;
assign w5341 = ~w5221 & ~w5339;
assign w5342 = ~w5340 & ~w5341;
assign w5343 = pi25 & pi43;
assign w5344 = pi29 & pi39;
assign w5345 = pi31 & pi37;
assign w5346 = pi30 & pi38;
assign w5347 = ~w5345 & w5346;
assign w5348 = w5345 & ~w5346;
assign w5349 = ~w5347 & ~w5348;
assign w5350 = w5344 & w5349;
assign w5351 = ~w5344 & ~w5349;
assign w5352 = ~w5350 & ~w5351;
assign w5353 = w5343 & w5352;
assign w5354 = ~w5343 & ~w5352;
assign w5355 = ~w5353 & ~w5354;
assign w5356 = pi26 & pi42;
assign w5357 = pi27 & pi41;
assign w5358 = ~w5092 & ~w5357;
assign w5359 = pi28 & pi41;
assign w5360 = w5090 & w5359;
assign w5361 = ~w5358 & ~w5360;
assign w5362 = w5356 & ~w5361;
assign w5363 = ~w5356 & w5361;
assign w5364 = ~w5362 & ~w5363;
assign w5365 = w5355 & ~w5364;
assign w5366 = ~w5355 & w5364;
assign w5367 = ~w5365 & ~w5366;
assign w5368 = w5342 & w5367;
assign w5369 = ~w5342 & ~w5367;
assign w5370 = ~w5368 & ~w5369;
assign w5371 = w5332 & w5370;
assign w5372 = ~w5332 & ~w5370;
assign w5373 = ~w5371 & ~w5372;
assign w5374 = (~w5142 & ~w5144) | (~w5142 & w8811) | (~w5144 & w8811);
assign w5375 = w5145 & ~w5147;
assign w5376 = ~w5149 & ~w5375;
assign w5377 = w5133 & ~w5135;
assign w5378 = ~w5137 & ~w5377;
assign w5379 = ~w5376 & ~w5378;
assign w5380 = w5376 & w5378;
assign w5381 = ~w5379 & ~w5380;
assign w5382 = ~w5374 & w5381;
assign w5383 = w5374 & ~w5381;
assign w5384 = ~w5382 & ~w5383;
assign w5385 = (~w5114 & ~w5116) | (~w5114 & w8632) | (~w5116 & w8632);
assign w5386 = w5117 & ~w5119;
assign w5387 = ~w5121 & ~w5386;
assign w5388 = w5105 & ~w5107;
assign w5389 = ~w5109 & ~w5388;
assign w5390 = ~w5387 & ~w5389;
assign w5391 = w5387 & w5389;
assign w5392 = ~w5390 & ~w5391;
assign w5393 = ~w5385 & w5392;
assign w5394 = w5385 & ~w5392;
assign w5395 = ~w5393 & ~w5394;
assign w5396 = (~w5086 & ~w5088) | (~w5086 & w8633) | (~w5088 & w8633);
assign w5397 = (~w5080 & ~w5082) | (~w5080 & w8969) | (~w5082 & w8969);
assign w5398 = w5089 & ~w5091;
assign w5399 = ~w5093 & ~w5398;
assign w5400 = ~w5397 & ~w5399;
assign w5401 = w5397 & w5399;
assign w5402 = ~w5400 & ~w5401;
assign w5403 = ~w5396 & w5402;
assign w5404 = w5396 & ~w5402;
assign w5405 = ~w5403 & ~w5404;
assign w5406 = w5395 & w5405;
assign w5407 = ~w5395 & ~w5405;
assign w5408 = ~w5406 & ~w5407;
assign w5409 = w5384 & w5408;
assign w5410 = ~w5384 & ~w5408;
assign w5411 = ~w5409 & ~w5410;
assign w5412 = pi11 & pi57;
assign w5413 = pi15 & pi53;
assign w5414 = pi16 & pi52;
assign w5415 = ~w5136 & ~w5414;
assign w5416 = pi17 & pi52;
assign w5417 = w5134 & w5416;
assign w5418 = ~w5415 & ~w5417;
assign w5419 = w5413 & ~w5418;
assign w5420 = ~w5413 & w5418;
assign w5421 = ~w5419 & ~w5420;
assign w5422 = w5412 & ~w5421;
assign w5423 = ~w5412 & w5421;
assign w5424 = ~w5422 & ~w5423;
assign w5425 = pi12 & pi56;
assign w5426 = pi13 & pi55;
assign w5427 = ~w5148 & ~w5426;
assign w5428 = pi14 & pi55;
assign w5429 = w5146 & w5428;
assign w5430 = ~w5427 & ~w5429;
assign w5431 = w5425 & ~w5430;
assign w5432 = ~w5425 & w5430;
assign w5433 = ~w5431 & ~w5432;
assign w5434 = w5424 & ~w5433;
assign w5435 = ~w5424 & w5433;
assign w5436 = ~w5434 & ~w5435;
assign w5437 = w5411 & w5436;
assign w5438 = ~w5411 & ~w5436;
assign w5439 = ~w5437 & ~w5438;
assign w5440 = w5373 & w5439;
assign w5441 = ~w5373 & ~w5439;
assign w5442 = ~w5440 & ~w5441;
assign w5443 = (~w5055 & w5052) | (~w5055 & w9052) | (w5052 & w9052);
assign w5444 = pi08 & pi60;
assign w5445 = pi09 & pi59;
assign w5446 = ~w5206 & ~w5445;
assign w5447 = pi10 & pi59;
assign w5448 = w5204 & w5447;
assign w5449 = ~w5446 & ~w5448;
assign w5450 = w5444 & w5449;
assign w5451 = ~w5444 & ~w5449;
assign w5452 = ~w5450 & ~w5451;
assign w5453 = w5215 & w5452;
assign w5454 = ~w5215 & ~w5452;
assign w5455 = ~w5453 & ~w5454;
assign w5456 = (w8970 & w5061) | (w8970 & w9053) | (w5061 & w9053);
assign w5457 = (w5455 & w8971) | (w5455 & w5067) | (w8971 & w5067);
assign w5458 = ~w5456 & ~w5457;
assign w5459 = w5443 & w5458;
assign w5460 = ~w5443 & ~w5458;
assign w5461 = ~w5459 & ~w5460;
assign w5462 = w5442 & ~w5461;
assign w5463 = ~w5442 & w5461;
assign w5464 = ~w5462 & ~w5463;
assign w5465 = w5307 & w5464;
assign w5466 = ~w5307 & ~w5464;
assign w5467 = ~w5465 & ~w5466;
assign w5468 = (w5467 & w5246) | (w5467 & w8972) | (w5246 & w8972);
assign w5469 = ~w5246 & w8973;
assign w5470 = ~w5468 & ~w5469;
assign w5471 = ~w5230 & ~w5233;
assign w5472 = ~w5224 & ~w5227;
assign w5473 = (~w5070 & ~w5072) | (~w5070 & w8974) | (~w5072 & w8974);
assign w5474 = w5472 & ~w5473;
assign w5475 = ~w5472 & w5473;
assign w5476 = ~w5474 & ~w5475;
assign w5477 = w5471 & w5476;
assign w5478 = ~w5471 & ~w5476;
assign w5479 = ~w5477 & ~w5478;
assign w5480 = w5470 & w5479;
assign w5481 = ~w5470 & ~w5479;
assign w5482 = ~w5480 & ~w5481;
assign w5483 = ~w5237 & ~w5248;
assign w5484 = ~w5482 & w5483;
assign w5485 = w5482 & ~w5483;
assign w5486 = ~w5484 & ~w5485;
assign w5487 = ~w5264 & w5486;
assign w5488 = w5264 & ~w5486;
assign w5489 = ~w5487 & ~w5488;
assign w5490 = (~w5484 & w5264) | (~w5484 & w9276) | (w5264 & w9276);
assign w5491 = ~w5462 & ~w5465;
assign w5492 = ~w5456 & ~w5459;
assign w5493 = (~w5302 & ~w5304) | (~w5302 & w8812) | (~w5304 & w8812);
assign w5494 = w5492 & ~w5493;
assign w5495 = ~w5492 & w5493;
assign w5496 = ~w5494 & ~w5495;
assign w5497 = ~w5491 & w5496;
assign w5498 = w5491 & ~w5496;
assign w5499 = ~w5497 & ~w5498;
assign w5500 = ~w5230 & ~w5474;
assign w5501 = ~w5233 & w5500;
assign w5502 = pi18 & pi51;
assign w5503 = pi22 & pi47;
assign w5504 = pi23 & pi46;
assign w5505 = ~w5312 & ~w5504;
assign w5506 = pi24 & pi46;
assign w5507 = w5310 & w5506;
assign w5508 = ~w5505 & ~w5507;
assign w5509 = w5503 & ~w5508;
assign w5510 = ~w5503 & w5508;
assign w5511 = ~w5509 & ~w5510;
assign w5512 = w5502 & ~w5511;
assign w5513 = ~w5502 & w5511;
assign w5514 = ~w5512 & ~w5513;
assign w5515 = pi19 & pi50;
assign w5516 = pi20 & pi49;
assign w5517 = ~w5324 & ~w5516;
assign w5518 = pi21 & pi49;
assign w5519 = w5322 & w5518;
assign w5520 = ~w5517 & ~w5519;
assign w5521 = w5515 & ~w5520;
assign w5522 = ~w5515 & w5520;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = w5514 & ~w5523;
assign w5525 = ~w5514 & w5523;
assign w5526 = ~w5524 & ~w5525;
assign w5527 = pi25 & pi44;
assign w5528 = pi29 & pi40;
assign w5529 = pi31 & pi38;
assign w5530 = pi30 & pi39;
assign w5531 = ~w5529 & w5530;
assign w5532 = w5529 & ~w5530;
assign w5533 = ~w5531 & ~w5532;
assign w5534 = w5528 & w5533;
assign w5535 = ~w5528 & ~w5533;
assign w5536 = ~w5534 & ~w5535;
assign w5537 = w5527 & w5536;
assign w5538 = ~w5527 & ~w5536;
assign w5539 = ~w5537 & ~w5538;
assign w5540 = pi26 & pi43;
assign w5541 = pi27 & pi42;
assign w5542 = ~w5359 & ~w5541;
assign w5543 = pi28 & pi42;
assign w5544 = w5357 & w5543;
assign w5545 = ~w5542 & ~w5544;
assign w5546 = w5540 & ~w5545;
assign w5547 = ~w5540 & w5545;
assign w5548 = ~w5546 & ~w5547;
assign w5549 = w5539 & ~w5548;
assign w5550 = ~w5539 & w5548;
assign w5551 = ~w5549 & ~w5550;
assign w5552 = w5448 & w5453;
assign w5553 = ~w5448 & ~w5453;
assign w5554 = ~w5552 & ~w5553;
assign w5555 = ~w5450 & ~w5554;
assign w5556 = w5551 & ~w5555;
assign w5557 = ~w5551 & w5555;
assign w5558 = ~w5556 & ~w5557;
assign w5559 = w5526 & w5558;
assign w5560 = ~w5526 & ~w5558;
assign w5561 = ~w5559 & ~w5560;
assign w5562 = (~w5422 & ~w5424) | (~w5422 & w8813) | (~w5424 & w8813);
assign w5563 = w5425 & ~w5427;
assign w5564 = ~w5429 & ~w5563;
assign w5565 = w5413 & ~w5415;
assign w5566 = ~w5417 & ~w5565;
assign w5567 = ~w5564 & ~w5566;
assign w5568 = w5564 & w5566;
assign w5569 = ~w5567 & ~w5568;
assign w5570 = ~w5562 & w5569;
assign w5571 = w5562 & ~w5569;
assign w5572 = ~w5570 & ~w5571;
assign w5573 = (~w5318 & ~w5320) | (~w5318 & w8634) | (~w5320 & w8634);
assign w5574 = w5321 & ~w5323;
assign w5575 = ~w5325 & ~w5574;
assign w5576 = w5309 & ~w5311;
assign w5577 = ~w5313 & ~w5576;
assign w5578 = ~w5575 & ~w5577;
assign w5579 = w5575 & w5577;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = ~w5573 & w5580;
assign w5582 = w5573 & ~w5580;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = (~w5353 & ~w5355) | (~w5353 & w8635) | (~w5355 & w8635);
assign w5585 = (~w5347 & ~w5349) | (~w5347 & w8814) | (~w5349 & w8814);
assign w5586 = w5356 & ~w5358;
assign w5587 = ~w5360 & ~w5586;
assign w5588 = ~w5585 & ~w5587;
assign w5589 = w5585 & w5587;
assign w5590 = ~w5588 & ~w5589;
assign w5591 = ~w5584 & w5590;
assign w5592 = w5584 & ~w5590;
assign w5593 = ~w5591 & ~w5592;
assign w5594 = w5583 & w5593;
assign w5595 = ~w5583 & ~w5593;
assign w5596 = ~w5594 & ~w5595;
assign w5597 = w5572 & w5596;
assign w5598 = ~w5572 & ~w5596;
assign w5599 = ~w5597 & ~w5598;
assign w5600 = pi11 & pi58;
assign w5601 = pi15 & pi54;
assign w5602 = pi16 & pi53;
assign w5603 = ~w5416 & ~w5602;
assign w5604 = pi17 & pi53;
assign w5605 = w5414 & w5604;
assign w5606 = ~w5603 & ~w5605;
assign w5607 = w5601 & ~w5606;
assign w5608 = ~w5601 & w5606;
assign w5609 = ~w5607 & ~w5608;
assign w5610 = w5600 & ~w5609;
assign w5611 = ~w5600 & w5609;
assign w5612 = ~w5610 & ~w5611;
assign w5613 = pi12 & pi57;
assign w5614 = pi13 & pi56;
assign w5615 = ~w5428 & ~w5614;
assign w5616 = pi14 & pi56;
assign w5617 = w5426 & w5616;
assign w5618 = ~w5615 & ~w5617;
assign w5619 = w5613 & ~w5618;
assign w5620 = ~w5613 & w5618;
assign w5621 = ~w5619 & ~w5620;
assign w5622 = w5612 & ~w5621;
assign w5623 = ~w5612 & w5621;
assign w5624 = ~w5622 & ~w5623;
assign w5625 = w5599 & w5624;
assign w5626 = ~w5599 & ~w5624;
assign w5627 = ~w5625 & ~w5626;
assign w5628 = w5561 & w5627;
assign w5629 = ~w5561 & ~w5627;
assign w5630 = ~w5628 & ~w5629;
assign w5631 = (~w5296 & ~w5293) | (~w5296 & w8815) | (~w5293 & w8815);
assign w5632 = pi08 & pi61;
assign w5633 = pi09 & pi60;
assign w5634 = ~w5447 & ~w5633;
assign w5635 = pi10 & pi60;
assign w5636 = w5445 & w5635;
assign w5637 = ~w5634 & ~w5636;
assign w5638 = w5632 & ~w5637;
assign w5639 = ~w5632 & w5637;
assign w5640 = ~w5638 & ~w5639;
assign w5641 = (~w5640 & w5290) | (~w5640 & w8975) | (w5290 & w8975);
assign w5642 = ~w5290 & w8976;
assign w5643 = ~w5641 & ~w5642;
assign w5644 = ~w5631 & w5643;
assign w5645 = w5631 & ~w5643;
assign w5646 = ~w5644 & ~w5645;
assign w5647 = w5630 & w5646;
assign w5648 = ~w5630 & ~w5646;
assign w5649 = ~w5647 & ~w5648;
assign w5650 = ~w5337 & ~w5340;
assign w5651 = pi06 & pi63;
assign w5652 = pi07 & pi62;
assign w5653 = w5651 & ~w5652;
assign w5654 = ~w5651 & w5652;
assign w5655 = ~w5653 & ~w5654;
assign w5656 = ~w5650 & ~w5655;
assign w5657 = w5650 & w5655;
assign w5658 = ~w5656 & ~w5657;
assign w5659 = (~w5379 & w5374) | (~w5379 & w8977) | (w5374 & w8977);
assign w5660 = (~w5400 & w5396) | (~w5400 & w8816) | (w5396 & w8816);
assign w5661 = (~w5390 & w5385) | (~w5390 & w8817) | (w5385 & w8817);
assign w5662 = ~w5660 & ~w5661;
assign w5663 = w5660 & w5661;
assign w5664 = ~w5662 & ~w5663;
assign w5665 = ~w5659 & w5664;
assign w5666 = w5659 & ~w5664;
assign w5667 = ~w5665 & ~w5666;
assign w5668 = w5658 & w5667;
assign w5669 = ~w5658 & ~w5667;
assign w5670 = ~w5668 & ~w5669;
assign w5671 = (~w5270 & ~w5281) | (~w5270 & w8978) | (~w5281 & w8978);
assign w5672 = (~w5276 & ~w5278) | (~w5276 & w8979) | (~w5278 & w8979);
assign w5673 = ~w5267 & ~w5672;
assign w5674 = w5267 & w5672;
assign w5675 = ~w5673 & ~w5674;
assign w5676 = ~w5671 & w5675;
assign w5677 = w5671 & ~w5675;
assign w5678 = ~w5676 & ~w5677;
assign w5679 = (~w5437 & ~w5439) | (~w5437 & w8752) | (~w5439 & w8752);
assign w5680 = ~w5368 & ~w5371;
assign w5681 = (~w5406 & ~w5408) | (~w5406 & w8980) | (~w5408 & w8980);
assign w5682 = ~w5680 & ~w5681;
assign w5683 = w5680 & w5681;
assign w5684 = ~w5682 & ~w5683;
assign w5685 = (w5439 & w9164) | (w5439 & w9165) | (w9164 & w9165);
assign w5686 = ~w5684 & w5679;
assign w5687 = ~w5685 & ~w5686;
assign w5688 = w5678 & w5687;
assign w5689 = ~w5678 & ~w5687;
assign w5690 = ~w5688 & ~w5689;
assign w5691 = w5670 & ~w5690;
assign w5692 = ~w5670 & w5690;
assign w5693 = ~w5691 & ~w5692;
assign w5694 = w5649 & ~w5693;
assign w5695 = ~w5649 & w5693;
assign w5696 = ~w5694 & ~w5695;
assign w5697 = ~w5501 & w8753;
assign w5698 = (~w5696 & w5501) | (~w5696 & w8754) | (w5501 & w8754);
assign w5699 = ~w5697 & ~w5698;
assign w5700 = w5499 & ~w5699;
assign w5701 = ~w5499 & w5699;
assign w5702 = ~w5700 & ~w5701;
assign w5703 = (~w5469 & ~w5470) | (~w5469 & w8755) | (~w5470 & w8755);
assign w5704 = w5702 & ~w5703;
assign w5705 = ~w5702 & w5703;
assign w5706 = ~w5704 & ~w5705;
assign w5707 = w5490 & ~w5706;
assign w5708 = (w5706 & w8756) | (w5706 & w5487) | (w8756 & w5487);
assign w5709 = ~w5707 & ~w5708;
assign w5710 = (~w5462 & w5493) | (~w5462 & w9054) | (w5493 & w9054);
assign w5711 = (~w5495 & w5465) | (~w5495 & w8757) | (w5465 & w8757);
assign w5712 = (~w5647 & w5693) | (~w5647 & w8818) | (w5693 & w8818);
assign w5713 = ~w5641 & ~w5644;
assign w5714 = (~w5689 & ~w5690) | (~w5689 & w8758) | (~w5690 & w8758);
assign w5715 = ~w5713 & w5714;
assign w5716 = w5713 & ~w5714;
assign w5717 = ~w5715 & ~w5716;
assign w5718 = ~w5712 & w5717;
assign w5719 = w5712 & ~w5717;
assign w5720 = ~w5718 & ~w5719;
assign w5721 = w5720 & w9277;
assign w5722 = ~w5567 & ~w5570;
assign w5723 = (~w5588 & w5584) | (~w5588 & w8759) | (w5584 & w8759);
assign w5724 = (~w5578 & w5573) | (~w5578 & w8760) | (w5573 & w8760);
assign w5725 = ~w5723 & ~w5724;
assign w5726 = w5723 & w5724;
assign w5727 = ~w5725 & ~w5726;
assign w5728 = ~w5722 & w5727;
assign w5729 = w5722 & ~w5727;
assign w5730 = ~w5728 & ~w5729;
assign w5731 = pi07 & pi63;
assign w5732 = pi08 & pi62;
assign w5733 = w5731 & ~w5732;
assign w5734 = ~w5731 & w5732;
assign w5735 = ~w5733 & ~w5734;
assign w5736 = w5552 & ~w5735;
assign w5737 = ~w5552 & w5735;
assign w5738 = ~w5736 & ~w5737;
assign w5739 = w5730 & w5738;
assign w5740 = ~w5730 & ~w5738;
assign w5741 = ~w5739 & ~w5740;
assign w5742 = (~w5656 & ~w5667) | (~w5656 & w8761) | (~w5667 & w8761);
assign w5743 = (~w5662 & ~w5664) | (~w5662 & w8762) | (~w5664 & w8762);
assign w5744 = ~w5653 & ~w5743;
assign w5745 = w5653 & w5743;
assign w5746 = ~w5744 & ~w5745;
assign w5747 = ~w5742 & w5746;
assign w5748 = w5742 & ~w5746;
assign w5749 = ~w5747 & ~w5748;
assign w5750 = (~w5625 & ~w5627) | (~w5625 & w8763) | (~w5627 & w8763);
assign w5751 = ~w5556 & ~w5559;
assign w5752 = (~w5594 & ~w5596) | (~w5594 & w8983) | (~w5596 & w8983);
assign w5753 = ~w5751 & ~w5752;
assign w5754 = w5751 & w5752;
assign w5755 = ~w5753 & ~w5754;
assign w5756 = (w5627 & w9166) | (w5627 & w9167) | (w9166 & w9167);
assign w5757 = ~w5755 & w5750;
assign w5758 = ~w5756 & ~w5757;
assign w5759 = w5749 & w5758;
assign w5760 = ~w5749 & ~w5758;
assign w5761 = ~w5759 & ~w5760;
assign w5762 = w5741 & w5761;
assign w5763 = ~w5741 & ~w5761;
assign w5764 = ~w5762 & ~w5763;
assign w5765 = pi25 & pi45;
assign w5766 = pi29 & pi41;
assign w5767 = pi31 & pi39;
assign w5768 = pi30 & pi40;
assign w5769 = ~w5767 & w5768;
assign w5770 = w5767 & ~w5768;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = w5766 & w5771;
assign w5773 = ~w5766 & ~w5771;
assign w5774 = ~w5772 & ~w5773;
assign w5775 = w5765 & w5774;
assign w5776 = ~w5765 & ~w5774;
assign w5777 = ~w5775 & ~w5776;
assign w5778 = pi26 & pi44;
assign w5779 = pi27 & pi43;
assign w5780 = ~w5543 & ~w5779;
assign w5781 = pi28 & pi43;
assign w5782 = w5541 & w5781;
assign w5783 = ~w5780 & ~w5782;
assign w5784 = w5778 & ~w5783;
assign w5785 = ~w5778 & w5783;
assign w5786 = ~w5784 & ~w5785;
assign w5787 = w5777 & ~w5786;
assign w5788 = ~w5777 & w5786;
assign w5789 = ~w5787 & ~w5788;
assign w5790 = w5632 & ~w5634;
assign w5791 = ~w5636 & ~w5790;
assign w5792 = w5789 & ~w5791;
assign w5793 = ~w5789 & w5791;
assign w5794 = ~w5792 & ~w5793;
assign w5795 = pi18 & pi52;
assign w5796 = pi22 & pi48;
assign w5797 = pi23 & pi47;
assign w5798 = ~w5506 & ~w5797;
assign w5799 = pi24 & pi47;
assign w5800 = w5504 & w5799;
assign w5801 = ~w5798 & ~w5800;
assign w5802 = w5796 & ~w5801;
assign w5803 = ~w5796 & w5801;
assign w5804 = ~w5802 & ~w5803;
assign w5805 = w5795 & ~w5804;
assign w5806 = ~w5795 & w5804;
assign w5807 = ~w5805 & ~w5806;
assign w5808 = pi19 & pi51;
assign w5809 = pi20 & pi50;
assign w5810 = ~w5518 & ~w5809;
assign w5811 = pi21 & pi50;
assign w5812 = w5516 & w5811;
assign w5813 = ~w5810 & ~w5812;
assign w5814 = w5808 & ~w5813;
assign w5815 = ~w5808 & w5813;
assign w5816 = ~w5814 & ~w5815;
assign w5817 = w5807 & ~w5816;
assign w5818 = ~w5807 & w5816;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = w5794 & w5819;
assign w5821 = ~w5794 & ~w5819;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = pi11 & pi59;
assign w5824 = pi15 & pi55;
assign w5825 = pi16 & pi54;
assign w5826 = ~w5604 & ~w5825;
assign w5827 = pi17 & pi54;
assign w5828 = w5602 & w5827;
assign w5829 = ~w5826 & ~w5828;
assign w5830 = w5824 & ~w5829;
assign w5831 = ~w5824 & w5829;
assign w5832 = ~w5830 & ~w5831;
assign w5833 = w5823 & ~w5832;
assign w5834 = ~w5823 & w5832;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = pi12 & pi58;
assign w5837 = pi13 & pi57;
assign w5838 = ~w5616 & ~w5837;
assign w5839 = pi14 & pi57;
assign w5840 = w5614 & w5839;
assign w5841 = ~w5838 & ~w5840;
assign w5842 = w5836 & ~w5841;
assign w5843 = ~w5836 & w5841;
assign w5844 = ~w5842 & ~w5843;
assign w5845 = w5835 & ~w5844;
assign w5846 = ~w5835 & w5844;
assign w5847 = ~w5845 & ~w5846;
assign w5848 = (~w5610 & ~w5612) | (~w5610 & w8636) | (~w5612 & w8636);
assign w5849 = w5613 & ~w5615;
assign w5850 = ~w5617 & ~w5849;
assign w5851 = w5601 & ~w5603;
assign w5852 = ~w5605 & ~w5851;
assign w5853 = ~w5850 & ~w5852;
assign w5854 = w5850 & w5852;
assign w5855 = ~w5853 & ~w5854;
assign w5856 = ~w5848 & w5855;
assign w5857 = w5848 & ~w5855;
assign w5858 = ~w5856 & ~w5857;
assign w5859 = (~w5512 & ~w5514) | (~w5512 & w8637) | (~w5514 & w8637);
assign w5860 = w5515 & ~w5517;
assign w5861 = ~w5519 & ~w5860;
assign w5862 = w5503 & ~w5505;
assign w5863 = ~w5507 & ~w5862;
assign w5864 = ~w5861 & ~w5863;
assign w5865 = w5861 & w5863;
assign w5866 = ~w5864 & ~w5865;
assign w5867 = ~w5859 & w5866;
assign w5868 = w5859 & ~w5866;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = (~w5537 & ~w5539) | (~w5537 & w8638) | (~w5539 & w8638);
assign w5871 = ~w5531 & ~w5534;
assign w5872 = w5540 & ~w5542;
assign w5873 = ~w5544 & ~w5872;
assign w5874 = ~w5871 & ~w5873;
assign w5875 = w5871 & w5873;
assign w5876 = ~w5874 & ~w5875;
assign w5877 = ~w5870 & w5876;
assign w5878 = w5870 & ~w5876;
assign w5879 = ~w5877 & ~w5878;
assign w5880 = w5869 & w5879;
assign w5881 = ~w5869 & ~w5879;
assign w5882 = ~w5880 & ~w5881;
assign w5883 = w5858 & w5882;
assign w5884 = ~w5858 & ~w5882;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = ~w5847 & ~w5885;
assign w5887 = w5847 & w5885;
assign w5888 = ~w5886 & ~w5887;
assign w5889 = ~w5822 & w5888;
assign w5890 = w5822 & ~w5888;
assign w5891 = ~w5889 & ~w5890;
assign w5892 = (~w5682 & w5679) | (~w5682 & w8819) | (w5679 & w8819);
assign w5893 = pi09 & pi61;
assign w5894 = ~w5635 & ~w5893;
assign w5895 = pi10 & pi61;
assign w5896 = w5633 & w5895;
assign w5897 = ~w5894 & ~w5896;
assign w5898 = ~w5676 & w8764;
assign w5899 = (w5897 & w5676) | (w5897 & w8765) | (w5676 & w8765);
assign w5900 = ~w5898 & ~w5899;
assign w5901 = w5892 & w5900;
assign w5902 = ~w5892 & ~w5900;
assign w5903 = ~w5901 & ~w5902;
assign w5904 = ~w5891 & ~w5903;
assign w5905 = w5891 & w5903;
assign w5906 = ~w5904 & ~w5905;
assign w5907 = w5764 & w5906;
assign w5908 = ~w5764 & ~w5906;
assign w5909 = ~w5907 & ~w5908;
assign w5910 = (w5909 & w5721) | (w5909 & w8766) | (w5721 & w8766);
assign w5911 = ~w5721 & w8767;
assign w5912 = ~w5910 & ~w5911;
assign w5913 = (~w5698 & ~w5699) | (~w5698 & w8984) | (~w5699 & w8984);
assign w5914 = w5912 & w5913;
assign w5915 = ~w5912 & ~w5913;
assign w5916 = ~w5914 & ~w5915;
assign w5917 = (w5264 & w9055) | (w5264 & w9056) | (w9055 & w9056);
assign w5918 = w5916 & ~w5917;
assign w5919 = ~w5916 & w5917;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = (w5264 & w9278) | (w5264 & w9279) | (w9278 & w9279);
assign w5922 = w5711 & w5720;
assign w5923 = ~w5922 & ~w5910;
assign w5924 = (~w5864 & w5859) | (~w5864 & w8820) | (w5859 & w8820);
assign w5925 = pi09 & pi62;
assign w5926 = pi11 & pi60;
assign w5927 = ~w5895 & ~w5926;
assign w5928 = pi11 & pi61;
assign w5929 = w5635 & w5928;
assign w5930 = ~w5927 & ~w5929;
assign w5931 = w5925 & ~w5930;
assign w5932 = ~w5925 & w5930;
assign w5933 = ~w5931 & ~w5932;
assign w5934 = ~w5924 & ~w5933;
assign w5935 = w5924 & w5933;
assign w5936 = ~w5934 & ~w5935;
assign w5937 = pi08 & pi63;
assign w5938 = (~w5874 & w5870) | (~w5874 & w8821) | (w5870 & w8821);
assign w5939 = w5937 & w5938;
assign w5940 = ~w5937 & ~w5938;
assign w5941 = ~w5939 & ~w5940;
assign w5942 = w5936 & ~w5941;
assign w5943 = ~w5936 & w5941;
assign w5944 = ~w5942 & ~w5943;
assign w5945 = (~w5736 & ~w5730) | (~w5736 & w8822) | (~w5730 & w8822);
assign w5946 = (~w5725 & ~w5727) | (~w5725 & w8823) | (~w5727 & w8823);
assign w5947 = ~w5733 & ~w5946;
assign w5948 = w5733 & w5946;
assign w5949 = ~w5947 & ~w5948;
assign w5950 = ~w5945 & w5949;
assign w5951 = w5945 & ~w5949;
assign w5952 = ~w5950 & ~w5951;
assign w5953 = (~w5886 & ~w5888) | (~w5886 & w8768) | (~w5888 & w8768);
assign w5954 = ~w5792 & ~w5820;
assign w5955 = (~w5880 & ~w5882) | (~w5880 & w8824) | (~w5882 & w8824);
assign w5956 = ~w5954 & ~w5955;
assign w5957 = w5954 & w5955;
assign w5958 = ~w5956 & ~w5957;
assign w5959 = w5958 & w5953;
assign w5960 = (w5888 & w9280) | (w5888 & w9281) | (w9280 & w9281);
assign w5961 = ~w5959 & ~w5960;
assign w5962 = w5952 & w5961;
assign w5963 = ~w5952 & ~w5961;
assign w5964 = ~w5962 & ~w5963;
assign w5965 = w5944 & w5964;
assign w5966 = ~w5944 & ~w5964;
assign w5967 = ~w5965 & ~w5966;
assign w5968 = pi25 & pi46;
assign w5969 = pi29 & pi42;
assign w5970 = pi31 & pi40;
assign w5971 = pi30 & pi41;
assign w5972 = ~w5970 & w5971;
assign w5973 = w5970 & ~w5971;
assign w5974 = ~w5972 & ~w5973;
assign w5975 = w5969 & w5974;
assign w5976 = ~w5969 & ~w5974;
assign w5977 = ~w5975 & ~w5976;
assign w5978 = w5968 & w5977;
assign w5979 = ~w5968 & ~w5977;
assign w5980 = ~w5978 & ~w5979;
assign w5981 = pi26 & pi45;
assign w5982 = pi27 & pi44;
assign w5983 = ~w5781 & ~w5982;
assign w5984 = pi28 & pi44;
assign w5985 = w5779 & w5984;
assign w5986 = ~w5983 & ~w5985;
assign w5987 = w5981 & ~w5986;
assign w5988 = ~w5981 & w5986;
assign w5989 = ~w5987 & ~w5988;
assign w5990 = w5980 & ~w5989;
assign w5991 = ~w5980 & w5989;
assign w5992 = ~w5990 & ~w5991;
assign w5993 = (~w5833 & ~w5835) | (~w5833 & w8639) | (~w5835 & w8639);
assign w5994 = w5836 & ~w5838;
assign w5995 = ~w5840 & ~w5994;
assign w5996 = w5824 & ~w5826;
assign w5997 = ~w5828 & ~w5996;
assign w5998 = ~w5995 & ~w5997;
assign w5999 = w5995 & w5997;
assign w6000 = ~w5998 & ~w5999;
assign w6001 = ~w5993 & w6000;
assign w6002 = w5993 & ~w6000;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = w5896 & w6003;
assign w6005 = ~w5896 & ~w6003;
assign w6006 = ~w6004 & ~w6005;
assign w6007 = w5992 & w6006;
assign w6008 = ~w5992 & ~w6006;
assign w6009 = ~w6007 & ~w6008;
assign w6010 = pi18 & pi53;
assign w6011 = pi22 & pi49;
assign w6012 = pi23 & pi48;
assign w6013 = ~w5799 & ~w6012;
assign w6014 = pi24 & pi48;
assign w6015 = w5797 & w6014;
assign w6016 = ~w6013 & ~w6015;
assign w6017 = w6011 & ~w6016;
assign w6018 = ~w6011 & w6016;
assign w6019 = ~w6017 & ~w6018;
assign w6020 = w6010 & ~w6019;
assign w6021 = ~w6010 & w6019;
assign w6022 = ~w6020 & ~w6021;
assign w6023 = pi19 & pi52;
assign w6024 = pi20 & pi51;
assign w6025 = ~w5811 & ~w6024;
assign w6026 = pi21 & pi51;
assign w6027 = w5809 & w6026;
assign w6028 = ~w6025 & ~w6027;
assign w6029 = w6023 & ~w6028;
assign w6030 = ~w6023 & w6028;
assign w6031 = ~w6029 & ~w6030;
assign w6032 = w6022 & ~w6031;
assign w6033 = ~w6022 & w6031;
assign w6034 = ~w6032 & ~w6033;
assign w6035 = (~w5805 & ~w5807) | (~w5805 & w8640) | (~w5807 & w8640);
assign w6036 = w5808 & ~w5810;
assign w6037 = ~w5812 & ~w6036;
assign w6038 = w5796 & ~w5798;
assign w6039 = ~w5800 & ~w6038;
assign w6040 = ~w6037 & ~w6039;
assign w6041 = w6037 & w6039;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = ~w6035 & w6042;
assign w6044 = w6035 & ~w6042;
assign w6045 = ~w6043 & ~w6044;
assign w6046 = (~w5853 & w5848) | (~w5853 & w8769) | (w5848 & w8769);
assign w6047 = (~w5775 & ~w5777) | (~w5775 & w8641) | (~w5777 & w8641);
assign w6048 = ~w5769 & ~w5772;
assign w6049 = w5778 & ~w5780;
assign w6050 = ~w5782 & ~w6049;
assign w6051 = ~w6048 & ~w6050;
assign w6052 = w6048 & w6050;
assign w6053 = ~w6051 & ~w6052;
assign w6054 = ~w6047 & w6053;
assign w6055 = w6047 & ~w6053;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = ~w6046 & w6056;
assign w6058 = w6046 & ~w6056;
assign w6059 = ~w6057 & ~w6058;
assign w6060 = w6045 & w6059;
assign w6061 = ~w6045 & ~w6059;
assign w6062 = ~w6060 & ~w6061;
assign w6063 = ~w6034 & ~w6062;
assign w6064 = w6034 & w6062;
assign w6065 = ~w6063 & ~w6064;
assign w6066 = ~w6009 & w6065;
assign w6067 = w6009 & ~w6065;
assign w6068 = ~w6066 & ~w6067;
assign w6069 = (~w5753 & w5750) | (~w5753 & w8825) | (w5750 & w8825);
assign w6070 = pi15 & pi56;
assign w6071 = pi16 & pi55;
assign w6072 = ~w5827 & ~w6071;
assign w6073 = pi17 & pi55;
assign w6074 = w5825 & w6073;
assign w6075 = ~w6072 & ~w6074;
assign w6076 = w6070 & ~w6075;
assign w6077 = ~w6070 & w6075;
assign w6078 = ~w6076 & ~w6077;
assign w6079 = pi12 & pi59;
assign w6080 = pi13 & pi58;
assign w6081 = ~w5839 & ~w6080;
assign w6082 = pi14 & pi58;
assign w6083 = w5837 & w6082;
assign w6084 = ~w6081 & ~w6083;
assign w6085 = w6079 & ~w6084;
assign w6086 = ~w6079 & w6084;
assign w6087 = ~w6085 & ~w6086;
assign w6088 = ~w6078 & ~w6087;
assign w6089 = w6078 & w6087;
assign w6090 = ~w6088 & ~w6089;
assign w6091 = ~w5747 & w8985;
assign w6092 = (w6090 & w5747) | (w6090 & w8986) | (w5747 & w8986);
assign w6093 = ~w6091 & ~w6092;
assign w6094 = w6069 & w6093;
assign w6095 = ~w6069 & ~w6093;
assign w6096 = ~w6094 & ~w6095;
assign w6097 = ~w6068 & ~w6096;
assign w6098 = w6068 & w6096;
assign w6099 = ~w6097 & ~w6098;
assign w6100 = w5967 & w6099;
assign w6101 = ~w5967 & ~w6099;
assign w6102 = ~w6100 & ~w6101;
assign w6103 = (~w5715 & w5712) | (~w5715 & w9170) | (w5712 & w9170);
assign w6104 = (~w5904 & ~w5764) | (~w5904 & w8826) | (~w5764 & w8826);
assign w6105 = ~w5898 & ~w5901;
assign w6106 = (~w5759 & ~w5761) | (~w5759 & w8827) | (~w5761 & w8827);
assign w6107 = w6105 & ~w6106;
assign w6108 = ~w6105 & w6106;
assign w6109 = ~w6107 & ~w6108;
assign w6110 = ~w6104 & w6109;
assign w6111 = w6104 & ~w6109;
assign w6112 = ~w6110 & ~w6111;
assign w6113 = ~w6103 & w6112;
assign w6114 = w6103 & ~w6112;
assign w6115 = ~w6113 & ~w6114;
assign w6116 = w6102 & w6115;
assign w6117 = ~w6102 & ~w6115;
assign w6118 = ~w6116 & ~w6117;
assign w6119 = w5923 & ~w6118;
assign w6120 = ~w5923 & w6118;
assign w6121 = ~w6119 & ~w6120;
assign w6122 = w5921 & ~w6121;
assign w6123 = ~w5921 & w6121;
assign w6124 = ~w6122 & ~w6123;
assign w6125 = ~w5915 & ~w6119;
assign w6126 = w5486 & w5706;
assign w6127 = w6125 & w6126;
assign w6128 = ~w5263 & w6127;
assign w6129 = w5484 & ~w5704;
assign w6130 = ~w5705 & ~w5914;
assign w6131 = ~w6120 & w9302;
assign w6132 = ~w6128 & w6131;
assign w6133 = ~w4262 & w5916;
assign w6134 = w6121 & w6133;
assign w6135 = w6126 & w6134;
assign w6136 = w5260 & w6135;
assign w6137 = ~w4520 & w6136;
assign w6138 = w6132 & ~w6137;
assign w6139 = (~w6113 & ~w6115) | (~w6113 & w8987) | (~w6115 & w8987);
assign w6140 = pi09 & pi63;
assign w6141 = pi10 & pi62;
assign w6142 = w6140 & ~w6141;
assign w6143 = ~w6140 & w6141;
assign w6144 = ~w6142 & ~w6143;
assign w6145 = (~w6051 & w6047) | (~w6051 & w8828) | (w6047 & w8828);
assign w6146 = pi13 & pi59;
assign w6147 = pi12 & pi60;
assign w6148 = ~w6146 & ~w6147;
assign w6149 = pi13 & pi60;
assign w6150 = w6079 & w6149;
assign w6151 = ~w6148 & ~w6150;
assign w6152 = w5928 & ~w6151;
assign w6153 = ~w5928 & w6151;
assign w6154 = ~w6152 & ~w6153;
assign w6155 = ~w6145 & ~w6154;
assign w6156 = w6145 & w6154;
assign w6157 = ~w6155 & ~w6156;
assign w6158 = ~w6144 & w6157;
assign w6159 = w6144 & ~w6157;
assign w6160 = ~w6158 & ~w6159;
assign w6161 = ~w5934 & ~w5942;
assign w6162 = w5925 & ~w5927;
assign w6163 = ~w5929 & ~w6162;
assign w6164 = ~w5939 & ~w6163;
assign w6165 = w5939 & w6163;
assign w6166 = ~w6164 & ~w6165;
assign w6167 = ~w6161 & w6166;
assign w6168 = w6161 & ~w6166;
assign w6169 = ~w6167 & ~w6168;
assign w6170 = (~w6063 & ~w6065) | (~w6063 & w8771) | (~w6065 & w8771);
assign w6171 = (~w6004 & ~w6006) | (~w6004 & w8829) | (~w6006 & w8829);
assign w6172 = (~w6057 & ~w6059) | (~w6057 & w8830) | (~w6059 & w8830);
assign w6173 = ~w6171 & ~w6172;
assign w6174 = w6171 & w6172;
assign w6175 = ~w6173 & ~w6174;
assign w6176 = w6170 & w6175;
assign w6177 = ~w6170 & ~w6175;
assign w6178 = ~w6176 & ~w6177;
assign w6179 = w6169 & w6178;
assign w6180 = ~w6169 & ~w6178;
assign w6181 = ~w6179 & ~w6180;
assign w6182 = w6160 & w6181;
assign w6183 = ~w6160 & ~w6181;
assign w6184 = ~w6182 & ~w6183;
assign w6185 = pi25 & pi47;
assign w6186 = pi29 & pi43;
assign w6187 = pi31 & pi41;
assign w6188 = pi30 & pi42;
assign w6189 = ~w6187 & w6188;
assign w6190 = w6187 & ~w6188;
assign w6191 = ~w6189 & ~w6190;
assign w6192 = w6186 & w6191;
assign w6193 = ~w6186 & ~w6191;
assign w6194 = ~w6192 & ~w6193;
assign w6195 = w6185 & w6194;
assign w6196 = ~w6185 & ~w6194;
assign w6197 = ~w6195 & ~w6196;
assign w6198 = pi26 & pi46;
assign w6199 = pi27 & pi45;
assign w6200 = ~w5984 & ~w6199;
assign w6201 = pi28 & pi45;
assign w6202 = w5982 & w6201;
assign w6203 = ~w6200 & ~w6202;
assign w6204 = w6198 & ~w6203;
assign w6205 = ~w6198 & w6203;
assign w6206 = ~w6204 & ~w6205;
assign w6207 = w6197 & ~w6206;
assign w6208 = ~w6197 & w6206;
assign w6209 = ~w6207 & ~w6208;
assign w6210 = w6079 & ~w6081;
assign w6211 = ~w6083 & ~w6210;
assign w6212 = w6070 & ~w6072;
assign w6213 = ~w6074 & ~w6212;
assign w6214 = ~w6211 & ~w6213;
assign w6215 = w6211 & w6213;
assign w6216 = ~w6214 & ~w6215;
assign w6217 = w6088 & w6216;
assign w6218 = ~w6088 & ~w6216;
assign w6219 = ~w6217 & ~w6218;
assign w6220 = (~w6020 & ~w6022) | (~w6020 & w8642) | (~w6022 & w8642);
assign w6221 = w6023 & ~w6025;
assign w6222 = ~w6027 & ~w6221;
assign w6223 = w6011 & ~w6013;
assign w6224 = ~w6015 & ~w6223;
assign w6225 = ~w6222 & ~w6224;
assign w6226 = w6222 & w6224;
assign w6227 = ~w6225 & ~w6226;
assign w6228 = ~w6220 & w6227;
assign w6229 = w6220 & ~w6227;
assign w6230 = ~w6228 & ~w6229;
assign w6231 = w6219 & w6230;
assign w6232 = ~w6219 & ~w6230;
assign w6233 = ~w6231 & ~w6232;
assign w6234 = w6209 & w6233;
assign w6235 = ~w6209 & ~w6233;
assign w6236 = ~w6234 & ~w6235;
assign w6237 = pi18 & pi54;
assign w6238 = pi22 & pi50;
assign w6239 = pi23 & pi49;
assign w6240 = ~w6014 & ~w6239;
assign w6241 = pi24 & pi49;
assign w6242 = w6012 & w6241;
assign w6243 = ~w6240 & ~w6242;
assign w6244 = w6238 & ~w6243;
assign w6245 = ~w6238 & w6243;
assign w6246 = ~w6244 & ~w6245;
assign w6247 = w6237 & ~w6246;
assign w6248 = ~w6237 & w6246;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = pi19 & pi53;
assign w6251 = pi20 & pi52;
assign w6252 = ~w6026 & ~w6251;
assign w6253 = pi21 & pi52;
assign w6254 = w6024 & w6253;
assign w6255 = ~w6252 & ~w6254;
assign w6256 = w6250 & ~w6255;
assign w6257 = ~w6250 & w6255;
assign w6258 = ~w6256 & ~w6257;
assign w6259 = w6249 & ~w6258;
assign w6260 = ~w6249 & w6258;
assign w6261 = ~w6259 & ~w6260;
assign w6262 = (~w5978 & ~w5980) | (~w5978 & w8772) | (~w5980 & w8772);
assign w6263 = (~w5972 & ~w5974) | (~w5972 & w8988) | (~w5974 & w8988);
assign w6264 = w5981 & ~w5983;
assign w6265 = ~w5985 & ~w6264;
assign w6266 = ~w6263 & ~w6265;
assign w6267 = w6263 & w6265;
assign w6268 = ~w6266 & ~w6267;
assign w6269 = ~w6262 & w6268;
assign w6270 = w6262 & ~w6268;
assign w6271 = ~w6269 & ~w6270;
assign w6272 = (~w6040 & w6035) | (~w6040 & w8643) | (w6035 & w8643);
assign w6273 = (~w5998 & w5993) | (~w5998 & w8644) | (w5993 & w8644);
assign w6274 = ~w6272 & ~w6273;
assign w6275 = w6272 & w6273;
assign w6276 = ~w6274 & ~w6275;
assign w6277 = w6271 & w6276;
assign w6278 = ~w6271 & ~w6276;
assign w6279 = ~w6277 & ~w6278;
assign w6280 = ~w6261 & ~w6279;
assign w6281 = w6261 & w6279;
assign w6282 = ~w6280 & ~w6281;
assign w6283 = ~w6236 & w6282;
assign w6284 = w6236 & ~w6282;
assign w6285 = ~w6283 & ~w6284;
assign w6286 = (~w5956 & ~w5953) | (~w5956 & w8645) | (~w5953 & w8645);
assign w6287 = pi15 & pi57;
assign w6288 = pi16 & pi56;
assign w6289 = ~w6073 & ~w6288;
assign w6290 = pi17 & pi56;
assign w6291 = w6071 & w6290;
assign w6292 = ~w6289 & ~w6291;
assign w6293 = w6287 & w6292;
assign w6294 = ~w6287 & ~w6292;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = w6082 & w6295;
assign w6297 = ~w6082 & ~w6295;
assign w6298 = ~w6296 & ~w6297;
assign w6299 = (w6298 & w5950) | (w6298 & w8646) | (w5950 & w8646);
assign w6300 = ~w5950 & w8647;
assign w6301 = ~w6299 & ~w6300;
assign w6302 = ~w6286 & w6301;
assign w6303 = w6286 & ~w6301;
assign w6304 = ~w6302 & ~w6303;
assign w6305 = ~w6285 & w6304;
assign w6306 = w6285 & ~w6304;
assign w6307 = ~w6305 & ~w6306;
assign w6308 = w6184 & w6307;
assign w6309 = ~w6184 & ~w6307;
assign w6310 = ~w6308 & ~w6309;
assign w6311 = (~w6107 & w6104) | (~w6107 & w9171) | (w6104 & w9171);
assign w6312 = (~w6097 & ~w5967) | (~w6097 & w8831) | (~w5967 & w8831);
assign w6313 = ~w6091 & ~w6094;
assign w6314 = (w5964 & w9172) | (w5964 & w9173) | (w9172 & w9173);
assign w6315 = ~w6313 & w9303;
assign w6316 = ~w6314 & ~w6315;
assign w6317 = ~w6312 & w6316;
assign w6318 = w6312 & ~w6316;
assign w6319 = ~w6317 & ~w6318;
assign w6320 = ~w6311 & w6319;
assign w6321 = w6311 & ~w6319;
assign w6322 = ~w6320 & ~w6321;
assign w6323 = w6310 & w6322;
assign w6324 = ~w6310 & ~w6322;
assign w6325 = ~w6323 & ~w6324;
assign w6326 = ~w6139 & w6325;
assign w6327 = w6139 & ~w6325;
assign w6328 = ~w6326 & ~w6327;
assign w6329 = (w6328 & w6137) | (w6328 & w8832) | (w6137 & w8832);
assign w6330 = w6138 & ~w6328;
assign w6331 = ~w6329 & ~w6330;
assign w6332 = (~w6137 & w8879) | (~w6137 & w8880) | (w8879 & w8880);
assign w6333 = (~w6320 & ~w6322) | (~w6320 & w8649) | (~w6322 & w8649);
assign w6334 = pi10 & pi63;
assign w6335 = pi11 & pi62;
assign w6336 = w6334 & ~w6335;
assign w6337 = ~w6334 & w6335;
assign w6338 = ~w6336 & ~w6337;
assign w6339 = pi12 & pi61;
assign w6340 = pi14 & pi59;
assign w6341 = ~w6149 & ~w6340;
assign w6342 = pi14 & pi60;
assign w6343 = w6146 & w6342;
assign w6344 = ~w6341 & ~w6343;
assign w6345 = w6339 & ~w6344;
assign w6346 = ~w6339 & w6344;
assign w6347 = ~w6345 & ~w6346;
assign w6348 = ~w6347 & w9304;
assign w6349 = (w6262 & w8989) | (w6262 & w8990) | (w8989 & w8990);
assign w6350 = ~w6348 & ~w6349;
assign w6351 = ~w6338 & w6350;
assign w6352 = w6338 & ~w6350;
assign w6353 = ~w6351 & ~w6352;
assign w6354 = (~w6155 & ~w6157) | (~w6155 & w8882) | (~w6157 & w8882);
assign w6355 = w5928 & ~w6148;
assign w6356 = ~w6150 & ~w6355;
assign w6357 = ~w6142 & ~w6356;
assign w6358 = w6142 & w6356;
assign w6359 = ~w6357 & ~w6358;
assign w6360 = ~w6354 & w6359;
assign w6361 = w6354 & ~w6359;
assign w6362 = ~w6360 & ~w6361;
assign w6363 = (~w6280 & ~w6282) | (~w6280 & w8773) | (~w6282 & w8773);
assign w6364 = (~w6231 & ~w6233) | (~w6231 & w8833) | (~w6233 & w8833);
assign w6365 = (~w6274 & ~w6276) | (~w6274 & w8883) | (~w6276 & w8883);
assign w6366 = ~w6364 & ~w6365;
assign w6367 = w6364 & w6365;
assign w6368 = ~w6366 & ~w6367;
assign w6369 = w6363 & w6368;
assign w6370 = ~w6363 & ~w6368;
assign w6371 = ~w6369 & ~w6370;
assign w6372 = w6362 & w6371;
assign w6373 = ~w6362 & ~w6371;
assign w6374 = ~w6372 & ~w6373;
assign w6375 = w6353 & w6374;
assign w6376 = ~w6353 & ~w6374;
assign w6377 = ~w6375 & ~w6376;
assign w6378 = (~w6173 & ~w6170) | (~w6173 & w8650) | (~w6170 & w8650);
assign w6379 = ~w6164 & ~w6167;
assign w6380 = pi15 & pi58;
assign w6381 = pi16 & pi57;
assign w6382 = ~w6290 & ~w6381;
assign w6383 = pi17 & pi57;
assign w6384 = w6288 & w6383;
assign w6385 = ~w6382 & ~w6384;
assign w6386 = w6380 & ~w6385;
assign w6387 = ~w6380 & w6385;
assign w6388 = ~w6386 & ~w6387;
assign w6389 = ~w6379 & ~w6388;
assign w6390 = w6379 & w6388;
assign w6391 = ~w6389 & ~w6390;
assign w6392 = ~w6378 & w6391;
assign w6393 = w6378 & ~w6391;
assign w6394 = ~w6392 & ~w6393;
assign w6395 = pi25 & pi48;
assign w6396 = pi29 & pi44;
assign w6397 = pi31 & pi42;
assign w6398 = pi30 & pi43;
assign w6399 = ~w6397 & w6398;
assign w6400 = w6397 & ~w6398;
assign w6401 = ~w6399 & ~w6400;
assign w6402 = w6396 & w6401;
assign w6403 = ~w6396 & ~w6401;
assign w6404 = ~w6402 & ~w6403;
assign w6405 = w6395 & w6404;
assign w6406 = ~w6395 & ~w6404;
assign w6407 = ~w6405 & ~w6406;
assign w6408 = pi26 & pi47;
assign w6409 = pi27 & pi46;
assign w6410 = ~w6201 & ~w6409;
assign w6411 = pi28 & pi46;
assign w6412 = w6199 & w6411;
assign w6413 = ~w6410 & ~w6412;
assign w6414 = w6408 & ~w6413;
assign w6415 = ~w6408 & w6413;
assign w6416 = ~w6414 & ~w6415;
assign w6417 = w6407 & ~w6416;
assign w6418 = ~w6407 & w6416;
assign w6419 = ~w6417 & ~w6418;
assign w6420 = (~w6247 & ~w6249) | (~w6247 & w8651) | (~w6249 & w8651);
assign w6421 = w6250 & ~w6252;
assign w6422 = ~w6254 & ~w6421;
assign w6423 = w6238 & ~w6240;
assign w6424 = ~w6242 & ~w6423;
assign w6425 = ~w6422 & ~w6424;
assign w6426 = w6422 & w6424;
assign w6427 = ~w6425 & ~w6426;
assign w6428 = ~w6420 & w6427;
assign w6429 = w6420 & ~w6427;
assign w6430 = ~w6428 & ~w6429;
assign w6431 = ~w6291 & ~w6296;
assign w6432 = w6295 & w8884;
assign w6433 = ~w6431 & ~w6432;
assign w6434 = ~w6293 & ~w6433;
assign w6435 = w6430 & ~w6434;
assign w6436 = ~w6430 & w6434;
assign w6437 = ~w6435 & ~w6436;
assign w6438 = w6419 & w6437;
assign w6439 = ~w6419 & ~w6437;
assign w6440 = ~w6438 & ~w6439;
assign w6441 = pi18 & pi55;
assign w6442 = pi22 & pi51;
assign w6443 = pi23 & pi50;
assign w6444 = ~w6241 & ~w6443;
assign w6445 = pi24 & pi50;
assign w6446 = w6239 & w6445;
assign w6447 = ~w6444 & ~w6446;
assign w6448 = w6442 & ~w6447;
assign w6449 = ~w6442 & w6447;
assign w6450 = ~w6448 & ~w6449;
assign w6451 = w6441 & ~w6450;
assign w6452 = ~w6441 & w6450;
assign w6453 = ~w6451 & ~w6452;
assign w6454 = pi19 & pi54;
assign w6455 = pi20 & pi53;
assign w6456 = ~w6253 & ~w6455;
assign w6457 = pi21 & pi53;
assign w6458 = w6251 & w6457;
assign w6459 = ~w6456 & ~w6458;
assign w6460 = w6454 & ~w6459;
assign w6461 = ~w6454 & w6459;
assign w6462 = ~w6460 & ~w6461;
assign w6463 = w6453 & ~w6462;
assign w6464 = ~w6453 & w6462;
assign w6465 = ~w6463 & ~w6464;
assign w6466 = (~w6195 & ~w6197) | (~w6195 & w8774) | (~w6197 & w8774);
assign w6467 = ~w6189 & ~w6192;
assign w6468 = w6198 & ~w6200;
assign w6469 = ~w6202 & ~w6468;
assign w6470 = ~w6467 & ~w6469;
assign w6471 = w6467 & w6469;
assign w6472 = ~w6470 & ~w6471;
assign w6473 = ~w6466 & w6472;
assign w6474 = w6466 & ~w6472;
assign w6475 = ~w6473 & ~w6474;
assign w6476 = (~w6225 & w6220) | (~w6225 & w8652) | (w6220 & w8652);
assign w6477 = ~w6214 & ~w6217;
assign w6478 = ~w6476 & ~w6477;
assign w6479 = w6476 & w6477;
assign w6480 = ~w6478 & ~w6479;
assign w6481 = w6475 & w6480;
assign w6482 = ~w6475 & ~w6480;
assign w6483 = ~w6481 & ~w6482;
assign w6484 = ~w6465 & ~w6483;
assign w6485 = w6465 & w6483;
assign w6486 = ~w6484 & ~w6485;
assign w6487 = ~w6440 & w6486;
assign w6488 = w6440 & ~w6486;
assign w6489 = ~w6487 & ~w6488;
assign w6490 = w6394 & ~w6489;
assign w6491 = ~w6394 & w6489;
assign w6492 = ~w6490 & ~w6491;
assign w6493 = w6377 & w6492;
assign w6494 = ~w6377 & ~w6492;
assign w6495 = ~w6493 & ~w6494;
assign w6496 = (~w6314 & w6312) | (~w6314 & w8653) | (w6312 & w8653);
assign w6497 = (~w6305 & ~w6184) | (~w6305 & w8654) | (~w6184 & w8654);
assign w6498 = ~w6299 & ~w6302;
assign w6499 = (w6181 & w9174) | (w6181 & w9175) | (w9174 & w9175);
assign w6500 = w6498 & w9305;
assign w6501 = ~w6499 & ~w6500;
assign w6502 = ~w6497 & w6501;
assign w6503 = w6497 & ~w6501;
assign w6504 = ~w6502 & ~w6503;
assign w6505 = ~w6496 & w6504;
assign w6506 = w6496 & ~w6504;
assign w6507 = ~w6505 & ~w6506;
assign w6508 = w6495 & w6507;
assign w6509 = ~w6495 & ~w6507;
assign w6510 = ~w6508 & ~w6509;
assign w6511 = w6333 & ~w6510;
assign w6512 = ~w6333 & w6510;
assign w6513 = ~w6511 & ~w6512;
assign w6514 = w6332 & ~w6513;
assign w6515 = ~w6332 & w6513;
assign w6516 = ~w6514 & ~w6515;
assign w6517 = (~w6505 & ~w6507) | (~w6505 & w8885) | (~w6507 & w8885);
assign w6518 = pi11 & pi63;
assign w6519 = pi12 & pi62;
assign w6520 = w6518 & ~w6519;
assign w6521 = ~w6518 & w6519;
assign w6522 = ~w6520 & ~w6521;
assign w6523 = (~w6470 & w6466) | (~w6470 & w8991) | (w6466 & w8991);
assign w6524 = pi13 & pi61;
assign w6525 = pi15 & pi59;
assign w6526 = ~w6342 & ~w6525;
assign w6527 = pi15 & pi60;
assign w6528 = w6340 & w6527;
assign w6529 = ~w6526 & ~w6528;
assign w6530 = w6524 & ~w6529;
assign w6531 = ~w6524 & w6529;
assign w6532 = ~w6530 & ~w6531;
assign w6533 = ~w6523 & ~w6532;
assign w6534 = w6523 & w6532;
assign w6535 = ~w6533 & ~w6534;
assign w6536 = ~w6522 & w6535;
assign w6537 = w6522 & ~w6535;
assign w6538 = ~w6536 & ~w6537;
assign w6539 = ~w6348 & ~w6351;
assign w6540 = w6339 & ~w6341;
assign w6541 = ~w6343 & ~w6540;
assign w6542 = ~w6336 & ~w6541;
assign w6543 = w6336 & w6541;
assign w6544 = ~w6542 & ~w6543;
assign w6545 = ~w6539 & w6544;
assign w6546 = w6539 & ~w6544;
assign w6547 = ~w6545 & ~w6546;
assign w6548 = (~w6484 & ~w6486) | (~w6484 & w8775) | (~w6486 & w8775);
assign w6549 = (~w6435 & ~w6437) | (~w6435 & w8834) | (~w6437 & w8834);
assign w6550 = (~w6478 & ~w6480) | (~w6478 & w8992) | (~w6480 & w8992);
assign w6551 = ~w6549 & ~w6550;
assign w6552 = w6549 & w6550;
assign w6553 = ~w6551 & ~w6552;
assign w6554 = w6548 & w6553;
assign w6555 = ~w6548 & ~w6553;
assign w6556 = ~w6554 & ~w6555;
assign w6557 = w6547 & w6556;
assign w6558 = ~w6547 & ~w6556;
assign w6559 = ~w6557 & ~w6558;
assign w6560 = w6538 & w6559;
assign w6561 = ~w6538 & ~w6559;
assign w6562 = ~w6560 & ~w6561;
assign w6563 = pi25 & pi49;
assign w6564 = pi29 & pi45;
assign w6565 = pi31 & pi43;
assign w6566 = pi30 & pi44;
assign w6567 = ~w6565 & w6566;
assign w6568 = w6565 & ~w6566;
assign w6569 = ~w6567 & ~w6568;
assign w6570 = w6564 & w6569;
assign w6571 = ~w6564 & ~w6569;
assign w6572 = ~w6570 & ~w6571;
assign w6573 = w6563 & w6572;
assign w6574 = ~w6563 & ~w6572;
assign w6575 = ~w6573 & ~w6574;
assign w6576 = pi26 & pi48;
assign w6577 = pi27 & pi47;
assign w6578 = ~w6411 & ~w6577;
assign w6579 = pi28 & pi47;
assign w6580 = w6409 & w6579;
assign w6581 = ~w6578 & ~w6580;
assign w6582 = w6576 & ~w6581;
assign w6583 = ~w6576 & w6581;
assign w6584 = ~w6582 & ~w6583;
assign w6585 = w6575 & ~w6584;
assign w6586 = ~w6575 & w6584;
assign w6587 = ~w6585 & ~w6586;
assign w6588 = (~w6451 & ~w6453) | (~w6451 & w8835) | (~w6453 & w8835);
assign w6589 = w6454 & ~w6456;
assign w6590 = ~w6458 & ~w6589;
assign w6591 = w6442 & ~w6444;
assign w6592 = ~w6446 & ~w6591;
assign w6593 = ~w6590 & ~w6592;
assign w6594 = w6590 & w6592;
assign w6595 = ~w6593 & ~w6594;
assign w6596 = ~w6588 & w6595;
assign w6597 = w6588 & ~w6595;
assign w6598 = ~w6596 & ~w6597;
assign w6599 = w6380 & ~w6382;
assign w6600 = ~w6384 & ~w6599;
assign w6601 = w6598 & ~w6600;
assign w6602 = ~w6598 & w6600;
assign w6603 = ~w6601 & ~w6602;
assign w6604 = w6587 & w6603;
assign w6605 = ~w6587 & ~w6603;
assign w6606 = ~w6604 & ~w6605;
assign w6607 = pi18 & pi56;
assign w6608 = pi22 & pi52;
assign w6609 = pi23 & pi51;
assign w6610 = ~w6445 & ~w6609;
assign w6611 = pi24 & pi51;
assign w6612 = w6443 & w6611;
assign w6613 = ~w6610 & ~w6612;
assign w6614 = w6608 & ~w6613;
assign w6615 = ~w6608 & w6613;
assign w6616 = ~w6614 & ~w6615;
assign w6617 = w6607 & ~w6616;
assign w6618 = ~w6607 & w6616;
assign w6619 = ~w6617 & ~w6618;
assign w6620 = pi19 & pi55;
assign w6621 = pi20 & pi54;
assign w6622 = ~w6457 & ~w6621;
assign w6623 = pi21 & pi54;
assign w6624 = w6455 & w6623;
assign w6625 = ~w6622 & ~w6624;
assign w6626 = w6620 & ~w6625;
assign w6627 = ~w6620 & w6625;
assign w6628 = ~w6626 & ~w6627;
assign w6629 = w6619 & ~w6628;
assign w6630 = ~w6619 & w6628;
assign w6631 = ~w6629 & ~w6630;
assign w6632 = (~w6405 & ~w6407) | (~w6405 & w8836) | (~w6407 & w8836);
assign w6633 = (~w6399 & ~w6401) | (~w6399 & w8993) | (~w6401 & w8993);
assign w6634 = w6408 & ~w6410;
assign w6635 = ~w6412 & ~w6634;
assign w6636 = ~w6633 & ~w6635;
assign w6637 = w6633 & w6635;
assign w6638 = ~w6636 & ~w6637;
assign w6639 = ~w6632 & w6638;
assign w6640 = w6632 & ~w6638;
assign w6641 = ~w6639 & ~w6640;
assign w6642 = (~w6420 & w8837) | (~w6420 & w8838) | (w8837 & w8838);
assign w6643 = (w6420 & w8839) | (w6420 & w8840) | (w8839 & w8840);
assign w6644 = ~w6642 & ~w6643;
assign w6645 = w6641 & w6644;
assign w6646 = ~w6641 & ~w6644;
assign w6647 = ~w6645 & ~w6646;
assign w6648 = w6631 & w6647;
assign w6649 = ~w6631 & ~w6647;
assign w6650 = ~w6648 & ~w6649;
assign w6651 = w6606 & w6650;
assign w6652 = ~w6606 & ~w6650;
assign w6653 = ~w6651 & ~w6652;
assign w6654 = (~w6366 & ~w6363) | (~w6366 & w8841) | (~w6363 & w8841);
assign w6655 = pi16 & pi58;
assign w6656 = ~w6383 & ~w6655;
assign w6657 = pi17 & pi58;
assign w6658 = w6381 & w6657;
assign w6659 = ~w6656 & ~w6658;
assign w6660 = ~w6357 & ~w6360;
assign w6661 = ~w6659 & w6660;
assign w6662 = w6659 & ~w6660;
assign w6663 = ~w6661 & ~w6662;
assign w6664 = w6654 & w6663;
assign w6665 = ~w6654 & ~w6663;
assign w6666 = ~w6664 & ~w6665;
assign w6667 = w6653 & ~w6666;
assign w6668 = ~w6653 & w6666;
assign w6669 = ~w6667 & ~w6668;
assign w6670 = w6562 & w6669;
assign w6671 = ~w6562 & ~w6669;
assign w6672 = ~w6670 & ~w6671;
assign w6673 = (~w6499 & w6497) | (~w6499 & w9176) | (w6497 & w9176);
assign w6674 = ~w6490 & ~w6493;
assign w6675 = ~w6389 & ~w6392;
assign w6676 = (~w6372 & ~w6374) | (~w6372 & w8842) | (~w6374 & w8842);
assign w6677 = ~w6675 & ~w6676;
assign w6678 = w6675 & w6676;
assign w6679 = ~w6677 & ~w6678;
assign w6680 = ~w6674 & w6679;
assign w6681 = w6674 & ~w6679;
assign w6682 = ~w6680 & ~w6681;
assign w6683 = ~w6673 & w6682;
assign w6684 = w6673 & ~w6682;
assign w6685 = ~w6683 & ~w6684;
assign w6686 = w6672 & w6685;
assign w6687 = ~w6672 & ~w6685;
assign w6688 = ~w6686 & ~w6687;
assign w6689 = ~w6517 & w6688;
assign w6690 = w6517 & ~w6688;
assign w6691 = ~w6689 & ~w6690;
assign w6692 = (w6137 & w8994) | (w6137 & w8995) | (w8994 & w8995);
assign w6693 = w6691 & w6692;
assign w6694 = ~w6691 & ~w6692;
assign w6695 = ~w6693 & ~w6694;
assign w6696 = (~w6137 & w9177) | (~w6137 & w9178) | (w9177 & w9178);
assign w6697 = (~w6683 & ~w6685) | (~w6683 & w8843) | (~w6685 & w8843);
assign w6698 = pi12 & pi63;
assign w6699 = pi16 & pi59;
assign w6700 = pi18 & pi57;
assign w6701 = ~w6657 & ~w6700;
assign w6702 = pi18 & pi58;
assign w6703 = w6383 & w6702;
assign w6704 = ~w6701 & ~w6703;
assign w6705 = w6699 & ~w6704;
assign w6706 = ~w6699 & w6704;
assign w6707 = ~w6705 & ~w6706;
assign w6708 = ~w6698 & ~w6707;
assign w6709 = w6698 & w6707;
assign w6710 = ~w6708 & ~w6709;
assign w6711 = pi13 & pi62;
assign w6712 = pi14 & pi61;
assign w6713 = ~w6527 & ~w6712;
assign w6714 = pi15 & pi61;
assign w6715 = w6342 & w6714;
assign w6716 = ~w6713 & ~w6715;
assign w6717 = w6711 & ~w6716;
assign w6718 = ~w6711 & w6716;
assign w6719 = ~w6717 & ~w6718;
assign w6720 = w6710 & ~w6719;
assign w6721 = ~w6710 & w6719;
assign w6722 = ~w6720 & ~w6721;
assign w6723 = ~w6533 & ~w6536;
assign w6724 = w6524 & ~w6526;
assign w6725 = ~w6528 & ~w6724;
assign w6726 = ~w6520 & ~w6725;
assign w6727 = w6520 & w6725;
assign w6728 = ~w6726 & ~w6727;
assign w6729 = ~w6723 & w6728;
assign w6730 = w6723 & ~w6728;
assign w6731 = ~w6729 & ~w6730;
assign w6732 = ~w6648 & ~w6651;
assign w6733 = (~w6601 & ~w6603) | (~w6601 & w8887) | (~w6603 & w8887);
assign w6734 = ~w6642 & ~w6645;
assign w6735 = ~w6733 & ~w6734;
assign w6736 = w6733 & w6734;
assign w6737 = ~w6735 & ~w6736;
assign w6738 = ~w6732 & w6737;
assign w6739 = w6732 & ~w6737;
assign w6740 = ~w6738 & ~w6739;
assign w6741 = w6731 & w6740;
assign w6742 = ~w6731 & ~w6740;
assign w6743 = ~w6741 & ~w6742;
assign w6744 = w6722 & w6743;
assign w6745 = ~w6722 & ~w6743;
assign w6746 = ~w6744 & ~w6745;
assign w6747 = pi25 & pi50;
assign w6748 = pi29 & pi46;
assign w6749 = pi31 & pi44;
assign w6750 = pi30 & pi45;
assign w6751 = ~w6749 & w6750;
assign w6752 = w6749 & ~w6750;
assign w6753 = ~w6751 & ~w6752;
assign w6754 = w6748 & w6753;
assign w6755 = ~w6748 & ~w6753;
assign w6756 = ~w6754 & ~w6755;
assign w6757 = w6747 & w6756;
assign w6758 = ~w6747 & ~w6756;
assign w6759 = ~w6757 & ~w6758;
assign w6760 = pi26 & pi49;
assign w6761 = pi27 & pi48;
assign w6762 = ~w6579 & ~w6761;
assign w6763 = pi28 & pi48;
assign w6764 = w6577 & w6763;
assign w6765 = ~w6762 & ~w6764;
assign w6766 = w6760 & ~w6765;
assign w6767 = ~w6760 & w6765;
assign w6768 = ~w6766 & ~w6767;
assign w6769 = w6759 & ~w6768;
assign w6770 = ~w6759 & w6768;
assign w6771 = ~w6769 & ~w6770;
assign w6772 = (~w6593 & w6588) | (~w6593 & w8888) | (w6588 & w8888);
assign w6773 = (~w6636 & w6632) | (~w6636 & w8889) | (w6632 & w8889);
assign w6774 = w6772 & w6773;
assign w6775 = ~w6772 & ~w6773;
assign w6776 = ~w6774 & ~w6775;
assign w6777 = w6771 & ~w6776;
assign w6778 = ~w6771 & w6776;
assign w6779 = ~w6777 & ~w6778;
assign w6780 = (~w6617 & ~w6619) | (~w6617 & w8844) | (~w6619 & w8844);
assign w6781 = w6620 & ~w6622;
assign w6782 = ~w6624 & ~w6781;
assign w6783 = w6608 & ~w6610;
assign w6784 = ~w6612 & ~w6783;
assign w6785 = ~w6782 & ~w6784;
assign w6786 = w6782 & w6784;
assign w6787 = ~w6785 & ~w6786;
assign w6788 = ~w6780 & w6787;
assign w6789 = w6780 & ~w6787;
assign w6790 = ~w6788 & ~w6789;
assign w6791 = (~w6573 & ~w6575) | (~w6573 & w8845) | (~w6575 & w8845);
assign w6792 = (~w6567 & ~w6569) | (~w6567 & w8996) | (~w6569 & w8996);
assign w6793 = w6576 & ~w6578;
assign w6794 = ~w6580 & ~w6793;
assign w6795 = ~w6792 & ~w6794;
assign w6796 = w6792 & w6794;
assign w6797 = ~w6795 & ~w6796;
assign w6798 = ~w6791 & w6797;
assign w6799 = w6791 & ~w6797;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = w6790 & w6800;
assign w6802 = ~w6790 & ~w6800;
assign w6803 = ~w6801 & ~w6802;
assign w6804 = w6658 & w6803;
assign w6805 = ~w6658 & ~w6803;
assign w6806 = ~w6804 & ~w6805;
assign w6807 = w6779 & w6806;
assign w6808 = ~w6779 & ~w6806;
assign w6809 = ~w6807 & ~w6808;
assign w6810 = (~w6551 & ~w6548) | (~w6551 & w8890) | (~w6548 & w8890);
assign w6811 = ~w6542 & ~w6545;
assign w6812 = pi19 & pi56;
assign w6813 = pi20 & pi55;
assign w6814 = ~w6623 & ~w6813;
assign w6815 = pi21 & pi55;
assign w6816 = w6621 & w6815;
assign w6817 = ~w6814 & ~w6816;
assign w6818 = w6812 & ~w6817;
assign w6819 = ~w6812 & w6817;
assign w6820 = ~w6818 & ~w6819;
assign w6821 = pi22 & pi53;
assign w6822 = pi23 & pi52;
assign w6823 = ~w6611 & ~w6822;
assign w6824 = pi24 & pi52;
assign w6825 = w6609 & w6824;
assign w6826 = ~w6823 & ~w6825;
assign w6827 = w6821 & ~w6826;
assign w6828 = ~w6821 & w6826;
assign w6829 = ~w6827 & ~w6828;
assign w6830 = ~w6820 & ~w6829;
assign w6831 = w6820 & w6829;
assign w6832 = ~w6830 & ~w6831;
assign w6833 = w6811 & ~w6832;
assign w6834 = ~w6811 & w6832;
assign w6835 = ~w6833 & ~w6834;
assign w6836 = w6810 & w6835;
assign w6837 = ~w6810 & ~w6835;
assign w6838 = ~w6836 & ~w6837;
assign w6839 = w6809 & ~w6838;
assign w6840 = ~w6809 & w6838;
assign w6841 = ~w6839 & ~w6840;
assign w6842 = w6746 & w6841;
assign w6843 = ~w6746 & ~w6841;
assign w6844 = ~w6842 & ~w6843;
assign w6845 = (~w6677 & w6674) | (~w6677 & w8846) | (w6674 & w8846);
assign w6846 = (~w6667 & ~w6562) | (~w6667 & w8847) | (~w6562 & w8847);
assign w6847 = ~w6661 & ~w6664;
assign w6848 = (w6559 & w9179) | (w6559 & w9180) | (w9179 & w9180);
assign w6849 = ~w6847 & w9306;
assign w6850 = ~w6848 & ~w6849;
assign w6851 = ~w6846 & w6850;
assign w6852 = w6846 & ~w6850;
assign w6853 = ~w6851 & ~w6852;
assign w6854 = ~w6845 & w6853;
assign w6855 = w6845 & ~w6853;
assign w6856 = ~w6854 & ~w6855;
assign w6857 = w6844 & w6856;
assign w6858 = ~w6844 & ~w6856;
assign w6859 = ~w6857 & ~w6858;
assign w6860 = ~w6697 & w6859;
assign w6861 = w6697 & ~w6859;
assign w6862 = ~w6860 & ~w6861;
assign w6863 = w6696 & ~w6862;
assign w6864 = ~w6696 & w6862;
assign w6865 = ~w6863 & ~w6864;
assign w6866 = w6326 & ~w6511;
assign w6867 = ~w6512 & ~w6689;
assign w6868 = ~w6866 & w6867;
assign w6869 = ~w6690 & w6862;
assign w6870 = (~w6860 & w6868) | (~w6860 & w8656) | (w6868 & w8656);
assign w6871 = w6328 & ~w6511;
assign w6872 = w6871 & w8891;
assign w6873 = (~w4520 & w9181) | (~w4520 & w9182) | (w9181 & w9182);
assign w6874 = (~w6854 & ~w6856) | (~w6854 & w8997) | (~w6856 & w8997);
assign w6875 = pi14 & pi62;
assign w6876 = pi20 & pi56;
assign w6877 = pi19 & pi57;
assign w6878 = ~w6876 & ~w6877;
assign w6879 = pi20 & pi57;
assign w6880 = w6812 & w6879;
assign w6881 = ~w6878 & ~w6880;
assign w6882 = w6702 & ~w6881;
assign w6883 = ~w6702 & w6881;
assign w6884 = ~w6882 & ~w6883;
assign w6885 = w6875 & ~w6884;
assign w6886 = ~w6875 & w6884;
assign w6887 = ~w6885 & ~w6886;
assign w6888 = pi17 & pi59;
assign w6889 = pi16 & pi60;
assign w6890 = ~w6888 & ~w6889;
assign w6891 = pi17 & pi60;
assign w6892 = w6699 & w6891;
assign w6893 = ~w6890 & ~w6892;
assign w6894 = w6714 & ~w6893;
assign w6895 = ~w6714 & w6893;
assign w6896 = ~w6894 & ~w6895;
assign w6897 = w6887 & ~w6896;
assign w6898 = ~w6887 & w6896;
assign w6899 = ~w6897 & ~w6898;
assign w6900 = ~w6708 & ~w6720;
assign w6901 = w6711 & ~w6713;
assign w6902 = ~w6715 & ~w6901;
assign w6903 = w6699 & ~w6701;
assign w6904 = ~w6703 & ~w6903;
assign w6905 = ~w6902 & ~w6904;
assign w6906 = w6902 & w6904;
assign w6907 = ~w6905 & ~w6906;
assign w6908 = ~w6900 & w6907;
assign w6909 = w6900 & ~w6907;
assign w6910 = ~w6908 & ~w6909;
assign w6911 = (~w6777 & ~w6806) | (~w6777 & w8892) | (~w6806 & w8892);
assign w6912 = (~w6801 & ~w6803) | (~w6801 & w8850) | (~w6803 & w8850);
assign w6913 = ~w6774 & ~w6912;
assign w6914 = w6774 & w6912;
assign w6915 = ~w6913 & ~w6914;
assign w6916 = ~w6911 & w6915;
assign w6917 = w6911 & ~w6915;
assign w6918 = ~w6916 & ~w6917;
assign w6919 = w6910 & w6918;
assign w6920 = ~w6910 & ~w6918;
assign w6921 = ~w6919 & ~w6920;
assign w6922 = w6899 & w6921;
assign w6923 = ~w6899 & ~w6921;
assign w6924 = ~w6922 & ~w6923;
assign w6925 = w6812 & ~w6814;
assign w6926 = ~w6816 & ~w6925;
assign w6927 = w6821 & ~w6823;
assign w6928 = ~w6825 & ~w6927;
assign w6929 = ~w6926 & ~w6928;
assign w6930 = w6926 & w6928;
assign w6931 = ~w6929 & ~w6930;
assign w6932 = w6830 & w6931;
assign w6933 = ~w6830 & ~w6931;
assign w6934 = ~w6932 & ~w6933;
assign w6935 = (~w6785 & w6780) | (~w6785 & w8893) | (w6780 & w8893);
assign w6936 = (~w6757 & ~w6759) | (~w6757 & w8851) | (~w6759 & w8851);
assign w6937 = (~w6751 & ~w6753) | (~w6751 & w8998) | (~w6753 & w8998);
assign w6938 = w6760 & ~w6762;
assign w6939 = ~w6764 & ~w6938;
assign w6940 = ~w6937 & ~w6939;
assign w6941 = w6937 & w6939;
assign w6942 = ~w6940 & ~w6941;
assign w6943 = ~w6936 & w6942;
assign w6944 = w6936 & ~w6942;
assign w6945 = ~w6943 & ~w6944;
assign w6946 = ~w6935 & w6945;
assign w6947 = w6935 & ~w6945;
assign w6948 = ~w6946 & ~w6947;
assign w6949 = w6934 & w6948;
assign w6950 = ~w6934 & ~w6948;
assign w6951 = ~w6949 & ~w6950;
assign w6952 = pi25 & pi51;
assign w6953 = pi29 & pi47;
assign w6954 = pi31 & pi45;
assign w6955 = pi30 & pi46;
assign w6956 = ~w6954 & w6955;
assign w6957 = w6954 & ~w6955;
assign w6958 = ~w6956 & ~w6957;
assign w6959 = w6953 & w6958;
assign w6960 = ~w6953 & ~w6958;
assign w6961 = ~w6959 & ~w6960;
assign w6962 = w6952 & w6961;
assign w6963 = ~w6952 & ~w6961;
assign w6964 = ~w6962 & ~w6963;
assign w6965 = pi26 & pi50;
assign w6966 = pi27 & pi49;
assign w6967 = ~w6763 & ~w6966;
assign w6968 = pi28 & pi49;
assign w6969 = w6761 & w6968;
assign w6970 = ~w6967 & ~w6969;
assign w6971 = w6965 & ~w6970;
assign w6972 = ~w6965 & w6970;
assign w6973 = ~w6971 & ~w6972;
assign w6974 = w6964 & ~w6973;
assign w6975 = ~w6964 & w6973;
assign w6976 = ~w6974 & ~w6975;
assign w6977 = pi13 & pi63;
assign w6978 = (w6791 & w8999) | (w6791 & w9000) | (w8999 & w9000);
assign w6979 = ~w6977 & w9307;
assign w6980 = ~w6978 & ~w6979;
assign w6981 = w6976 & ~w6980;
assign w6982 = ~w6976 & w6980;
assign w6983 = ~w6981 & ~w6982;
assign w6984 = w6951 & w6983;
assign w6985 = ~w6951 & ~w6983;
assign w6986 = ~w6984 & ~w6985;
assign w6987 = (~w6735 & w6732) | (~w6735 & w8895) | (w6732 & w8895);
assign w6988 = (~w6726 & w6723) | (~w6726 & w8852) | (w6723 & w8852);
assign w6989 = pi22 & pi54;
assign w6990 = pi23 & pi53;
assign w6991 = ~w6824 & ~w6990;
assign w6992 = pi24 & pi53;
assign w6993 = w6822 & w6992;
assign w6994 = ~w6991 & ~w6993;
assign w6995 = w6989 & w6994;
assign w6996 = ~w6989 & ~w6994;
assign w6997 = ~w6995 & ~w6996;
assign w6998 = w6815 & w6997;
assign w6999 = ~w6815 & ~w6997;
assign w7000 = ~w6998 & ~w6999;
assign w7001 = ~w6988 & w7000;
assign w7002 = w6988 & ~w7000;
assign w7003 = ~w7001 & ~w7002;
assign w7004 = ~w6987 & w7003;
assign w7005 = w6987 & ~w7003;
assign w7006 = ~w7004 & ~w7005;
assign w7007 = w6986 & w7006;
assign w7008 = ~w6986 & ~w7006;
assign w7009 = ~w7007 & ~w7008;
assign w7010 = w6924 & w7009;
assign w7011 = ~w6924 & ~w7009;
assign w7012 = ~w7010 & ~w7011;
assign w7013 = (~w6848 & w6846) | (~w6848 & w9183) | (w6846 & w9183);
assign w7014 = (~w6839 & ~w6746) | (~w6839 & w8896) | (~w6746 & w8896);
assign w7015 = ~w6833 & ~w6836;
assign w7016 = (w6743 & w9184) | (w6743 & w9185) | (w9184 & w9185);
assign w7017 = ~w7015 & w9308;
assign w7018 = ~w7016 & ~w7017;
assign w7019 = ~w7014 & w7018;
assign w7020 = w7014 & ~w7018;
assign w7021 = ~w7019 & ~w7020;
assign w7022 = ~w7013 & w7021;
assign w7023 = w7013 & ~w7021;
assign w7024 = ~w7022 & ~w7023;
assign w7025 = w7012 & w7024;
assign w7026 = ~w7012 & ~w7024;
assign w7027 = ~w7025 & ~w7026;
assign w7028 = ~w6874 & w7027;
assign w7029 = w6874 & ~w7027;
assign w7030 = ~w7028 & ~w7029;
assign w7031 = (w7030 & w6873) | (w7030 & w8854) | (w6873 & w8854);
assign w7032 = ~w6873 & w9282;
assign w7033 = ~w7031 & ~w7032;
assign w7034 = (~w6137 & w9001) | (~w6137 & w9002) | (w9001 & w9002);
assign w7035 = (~w7022 & ~w7024) | (~w7022 & w8855) | (~w7024 & w8855);
assign w7036 = pi15 & pi62;
assign w7037 = pi19 & pi58;
assign w7038 = pi21 & pi56;
assign w7039 = ~w6879 & ~w7038;
assign w7040 = pi21 & pi57;
assign w7041 = w6876 & w7040;
assign w7042 = ~w7039 & ~w7041;
assign w7043 = w7037 & ~w7042;
assign w7044 = ~w7037 & w7042;
assign w7045 = ~w7043 & ~w7044;
assign w7046 = w7036 & ~w7045;
assign w7047 = ~w7036 & w7045;
assign w7048 = ~w7046 & ~w7047;
assign w7049 = pi16 & pi61;
assign w7050 = pi18 & pi59;
assign w7051 = ~w6891 & ~w7050;
assign w7052 = pi18 & pi60;
assign w7053 = w6888 & w7052;
assign w7054 = ~w7051 & ~w7053;
assign w7055 = w7049 & ~w7054;
assign w7056 = ~w7049 & w7054;
assign w7057 = ~w7055 & ~w7056;
assign w7058 = w7048 & ~w7057;
assign w7059 = ~w7048 & w7057;
assign w7060 = ~w7058 & ~w7059;
assign w7061 = (~w6981 & ~w6951) | (~w6981 & w8899) | (~w6951 & w8899);
assign w7062 = (~w6946 & ~w6948) | (~w6946 & w8900) | (~w6948 & w8900);
assign w7063 = ~w6978 & ~w7062;
assign w7064 = w6978 & w7062;
assign w7065 = ~w7063 & ~w7064;
assign w7066 = ~w7061 & w7065;
assign w7067 = w7061 & ~w7065;
assign w7068 = ~w7066 & ~w7067;
assign w7069 = ~w6885 & ~w6897;
assign w7070 = w6714 & ~w6890;
assign w7071 = ~w6892 & ~w7070;
assign w7072 = w6702 & ~w6878;
assign w7073 = ~w6880 & ~w7072;
assign w7074 = ~w7071 & ~w7073;
assign w7075 = w7071 & w7073;
assign w7076 = ~w7074 & ~w7075;
assign w7077 = ~w7069 & w7076;
assign w7078 = w7069 & ~w7076;
assign w7079 = ~w7077 & ~w7078;
assign w7080 = w7068 & w7079;
assign w7081 = ~w7068 & ~w7079;
assign w7082 = ~w7080 & ~w7081;
assign w7083 = w7060 & w7082;
assign w7084 = ~w7060 & ~w7082;
assign w7085 = ~w7083 & ~w7084;
assign w7086 = ~w6929 & ~w6932;
assign w7087 = (~w6962 & ~w6964) | (~w6962 & w8856) | (~w6964 & w8856);
assign w7088 = (~w6956 & ~w6958) | (~w6956 & w9003) | (~w6958 & w9003);
assign w7089 = w6965 & ~w6967;
assign w7090 = ~w6969 & ~w7089;
assign w7091 = ~w7088 & ~w7090;
assign w7092 = w7088 & w7090;
assign w7093 = ~w7091 & ~w7092;
assign w7094 = ~w7087 & w7093;
assign w7095 = w7087 & ~w7093;
assign w7096 = ~w7094 & ~w7095;
assign w7097 = ~w7086 & w7096;
assign w7098 = w7086 & ~w7096;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = ~w6993 & ~w6998;
assign w7101 = w6993 & w6998;
assign w7102 = ~w7100 & ~w7101;
assign w7103 = ~w6995 & ~w7102;
assign w7104 = w7099 & ~w7103;
assign w7105 = ~w7099 & w7103;
assign w7106 = ~w7104 & ~w7105;
assign w7107 = pi25 & pi52;
assign w7108 = pi29 & pi48;
assign w7109 = pi31 & pi46;
assign w7110 = pi30 & pi47;
assign w7111 = ~w7109 & w7110;
assign w7112 = w7109 & ~w7110;
assign w7113 = ~w7111 & ~w7112;
assign w7114 = w7108 & w7113;
assign w7115 = ~w7108 & ~w7113;
assign w7116 = ~w7114 & ~w7115;
assign w7117 = w7107 & w7116;
assign w7118 = ~w7107 & ~w7116;
assign w7119 = ~w7117 & ~w7118;
assign w7120 = pi26 & pi51;
assign w7121 = pi27 & pi50;
assign w7122 = ~w6968 & ~w7121;
assign w7123 = pi28 & pi50;
assign w7124 = w6966 & w7123;
assign w7125 = ~w7122 & ~w7124;
assign w7126 = w7120 & ~w7125;
assign w7127 = ~w7120 & w7125;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = w7119 & ~w7128;
assign w7130 = ~w7119 & w7128;
assign w7131 = ~w7129 & ~w7130;
assign w7132 = pi14 & pi63;
assign w7133 = (w6936 & w9004) | (w6936 & w9005) | (w9004 & w9005);
assign w7134 = ~w7132 & w9309;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = w7131 & ~w7135;
assign w7137 = ~w7131 & w7135;
assign w7138 = ~w7136 & ~w7137;
assign w7139 = w7106 & w7138;
assign w7140 = ~w7106 & ~w7138;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = ~w6905 & ~w6908;
assign w7143 = pi22 & pi55;
assign w7144 = pi23 & pi54;
assign w7145 = ~w6992 & ~w7144;
assign w7146 = pi24 & pi54;
assign w7147 = w6990 & w7146;
assign w7148 = ~w7145 & ~w7147;
assign w7149 = w7143 & ~w7148;
assign w7150 = ~w7143 & w7148;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = ~w7142 & ~w7151;
assign w7153 = w7142 & w7151;
assign w7154 = ~w7152 & ~w7153;
assign w7155 = (w7154 & w6916) | (w7154 & w9006) | (w6916 & w9006);
assign w7156 = ~w6916 & w9007;
assign w7157 = ~w7155 & ~w7156;
assign w7158 = w7141 & w7157;
assign w7159 = ~w7141 & ~w7157;
assign w7160 = ~w7158 & ~w7159;
assign w7161 = w7085 & w7160;
assign w7162 = ~w7085 & ~w7160;
assign w7163 = ~w7161 & ~w7162;
assign w7164 = (~w7016 & w7014) | (~w7016 & w8857) | (w7014 & w8857);
assign w7165 = ~w7007 & ~w7010;
assign w7166 = (~w6919 & ~w6921) | (~w6919 & w8858) | (~w6921 & w8858);
assign w7167 = ~w7001 & ~w7004;
assign w7168 = ~w7166 & ~w7167;
assign w7169 = w7166 & w7167;
assign w7170 = ~w7168 & ~w7169;
assign w7171 = ~w7165 & w7170;
assign w7172 = w7165 & ~w7170;
assign w7173 = ~w7171 & ~w7172;
assign w7174 = ~w7164 & w7173;
assign w7175 = w7164 & ~w7173;
assign w7176 = ~w7174 & ~w7175;
assign w7177 = w7163 & w7176;
assign w7178 = ~w7163 & ~w7176;
assign w7179 = ~w7177 & ~w7178;
assign w7180 = w7035 & ~w7179;
assign w7181 = ~w7035 & w7179;
assign w7182 = ~w7180 & ~w7181;
assign w7183 = w7034 & w7182;
assign w7184 = ~w7034 & ~w7182;
assign w7185 = ~w7183 & ~w7184;
assign w7186 = (~w7174 & ~w7176) | (~w7174 & w9008) | (~w7176 & w9008);
assign w7187 = w7143 & ~w7145;
assign w7188 = ~w7147 & ~w7187;
assign w7189 = (~w7117 & ~w7119) | (~w7117 & w8859) | (~w7119 & w8859);
assign w7190 = ~w7111 & ~w7114;
assign w7191 = w7120 & ~w7122;
assign w7192 = ~w7124 & ~w7191;
assign w7193 = ~w7190 & ~w7192;
assign w7194 = w7190 & w7192;
assign w7195 = ~w7193 & ~w7194;
assign w7196 = ~w7189 & w7195;
assign w7197 = w7189 & ~w7195;
assign w7198 = ~w7196 & ~w7197;
assign w7199 = w7101 & ~w7198;
assign w7200 = ~w7101 & w7198;
assign w7201 = ~w7199 & ~w7200;
assign w7202 = ~w7188 & ~w7201;
assign w7203 = w7188 & w7201;
assign w7204 = ~w7202 & ~w7203;
assign w7205 = pi25 & pi53;
assign w7206 = pi29 & pi49;
assign w7207 = pi31 & pi47;
assign w7208 = pi30 & pi48;
assign w7209 = ~w7207 & w7208;
assign w7210 = w7207 & ~w7208;
assign w7211 = ~w7209 & ~w7210;
assign w7212 = w7206 & w7211;
assign w7213 = ~w7206 & ~w7211;
assign w7214 = ~w7212 & ~w7213;
assign w7215 = w7205 & w7214;
assign w7216 = ~w7205 & ~w7214;
assign w7217 = ~w7215 & ~w7216;
assign w7218 = pi26 & pi52;
assign w7219 = pi27 & pi51;
assign w7220 = ~w7123 & ~w7219;
assign w7221 = pi28 & pi51;
assign w7222 = w7121 & w7221;
assign w7223 = ~w7220 & ~w7222;
assign w7224 = w7218 & ~w7223;
assign w7225 = ~w7218 & w7223;
assign w7226 = ~w7224 & ~w7225;
assign w7227 = w7217 & ~w7226;
assign w7228 = ~w7217 & w7226;
assign w7229 = ~w7227 & ~w7228;
assign w7230 = pi15 & pi63;
assign w7231 = (w7087 & w9009) | (w7087 & w9010) | (w9009 & w9010);
assign w7232 = ~w7230 & w9310;
assign w7233 = ~w7231 & ~w7232;
assign w7234 = w7229 & ~w7233;
assign w7235 = ~w7229 & w7233;
assign w7236 = ~w7234 & ~w7235;
assign w7237 = w7204 & w7236;
assign w7238 = ~w7204 & ~w7236;
assign w7239 = ~w7237 & ~w7238;
assign w7240 = pi23 & pi55;
assign w7241 = ~w7146 & ~w7240;
assign w7242 = pi24 & pi55;
assign w7243 = w7144 & w7242;
assign w7244 = ~w7241 & ~w7243;
assign w7245 = ~w7074 & ~w7077;
assign w7246 = w7244 & ~w7245;
assign w7247 = ~w7244 & w7245;
assign w7248 = ~w7246 & ~w7247;
assign w7249 = (w7248 & w7066) | (w7248 & w9011) | (w7066 & w9011);
assign w7250 = ~w7066 & w9012;
assign w7251 = ~w7249 & ~w7250;
assign w7252 = w7239 & w7251;
assign w7253 = ~w7239 & ~w7251;
assign w7254 = ~w7252 & ~w7253;
assign w7255 = pi16 & pi62;
assign w7256 = pi20 & pi58;
assign w7257 = pi22 & pi56;
assign w7258 = ~w7040 & ~w7257;
assign w7259 = pi22 & pi57;
assign w7260 = w7038 & w7259;
assign w7261 = ~w7258 & ~w7260;
assign w7262 = w7256 & ~w7261;
assign w7263 = ~w7256 & w7261;
assign w7264 = ~w7262 & ~w7263;
assign w7265 = w7255 & ~w7264;
assign w7266 = ~w7255 & w7264;
assign w7267 = ~w7265 & ~w7266;
assign w7268 = pi17 & pi61;
assign w7269 = pi19 & pi59;
assign w7270 = ~w7052 & ~w7269;
assign w7271 = pi19 & pi60;
assign w7272 = w7050 & w7271;
assign w7273 = ~w7270 & ~w7272;
assign w7274 = w7268 & ~w7273;
assign w7275 = ~w7268 & w7273;
assign w7276 = ~w7274 & ~w7275;
assign w7277 = w7267 & ~w7276;
assign w7278 = ~w7267 & w7276;
assign w7279 = ~w7277 & ~w7278;
assign w7280 = (~w7136 & ~w7106) | (~w7136 & w8903) | (~w7106 & w8903);
assign w7281 = (~w7097 & ~w7099) | (~w7097 & w8904) | (~w7099 & w8904);
assign w7282 = ~w7133 & ~w7281;
assign w7283 = w7133 & w7281;
assign w7284 = ~w7282 & ~w7283;
assign w7285 = ~w7280 & w7284;
assign w7286 = w7280 & ~w7284;
assign w7287 = ~w7285 & ~w7286;
assign w7288 = ~w7046 & ~w7058;
assign w7289 = w7049 & ~w7051;
assign w7290 = ~w7053 & ~w7289;
assign w7291 = w7037 & ~w7039;
assign w7292 = ~w7041 & ~w7291;
assign w7293 = ~w7290 & ~w7292;
assign w7294 = w7290 & w7292;
assign w7295 = ~w7293 & ~w7294;
assign w7296 = ~w7288 & w7295;
assign w7297 = w7288 & ~w7295;
assign w7298 = ~w7296 & ~w7297;
assign w7299 = w7287 & w7298;
assign w7300 = ~w7287 & ~w7298;
assign w7301 = ~w7299 & ~w7300;
assign w7302 = w7279 & w7301;
assign w7303 = ~w7279 & ~w7301;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = w7254 & w7304;
assign w7306 = ~w7254 & ~w7304;
assign w7307 = ~w7305 & ~w7306;
assign w7308 = (~w7168 & w7165) | (~w7168 & w9013) | (w7165 & w9013);
assign w7309 = (~w7158 & ~w7085) | (~w7158 & w9014) | (~w7085 & w9014);
assign w7310 = ~w7152 & ~w7155;
assign w7311 = (~w7080 & ~w7082) | (~w7080 & w9015) | (~w7082 & w9015);
assign w7312 = ~w7310 & ~w7311;
assign w7313 = w7310 & w7311;
assign w7314 = ~w7312 & ~w7313;
assign w7315 = ~w7309 & w7314;
assign w7316 = w7309 & ~w7314;
assign w7317 = ~w7315 & ~w7316;
assign w7318 = ~w7308 & w7317;
assign w7319 = w7308 & ~w7317;
assign w7320 = ~w7318 & ~w7319;
assign w7321 = w7307 & w7320;
assign w7322 = ~w7307 & ~w7320;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = ~w7186 & w7323;
assign w7325 = w7186 & ~w7323;
assign w7326 = ~w7324 & ~w7325;
assign w7327 = (w6137 & w9186) | (w6137 & w9187) | (w9186 & w9187);
assign w7328 = w7326 & ~w7327;
assign w7329 = ~w7326 & w7327;
assign w7330 = ~w7328 & ~w7329;
assign w7331 = ~w7318 & ~w7321;
assign w7332 = pi16 & pi63;
assign w7333 = pi17 & pi62;
assign w7334 = pi18 & pi61;
assign w7335 = ~w7333 & ~w7334;
assign w7336 = pi18 & pi62;
assign w7337 = w7268 & w7336;
assign w7338 = ~w7335 & ~w7337;
assign w7339 = w7332 & ~w7338;
assign w7340 = ~w7332 & w7338;
assign w7341 = ~w7339 & ~w7340;
assign w7342 = w7243 & w7341;
assign w7343 = ~w7243 & ~w7341;
assign w7344 = ~w7342 & ~w7343;
assign w7345 = (~w7193 & w7189) | (~w7193 & w9059) | (w7189 & w9059);
assign w7346 = (~w7215 & ~w7217) | (~w7215 & w9016) | (~w7217 & w9016);
assign w7347 = ~w7209 & ~w7212;
assign w7348 = w7218 & ~w7220;
assign w7349 = ~w7222 & ~w7348;
assign w7350 = ~w7347 & ~w7349;
assign w7351 = w7347 & w7349;
assign w7352 = ~w7350 & ~w7351;
assign w7353 = ~w7346 & w7352;
assign w7354 = w7346 & ~w7352;
assign w7355 = ~w7353 & ~w7354;
assign w7356 = w7345 & ~w7355;
assign w7357 = ~w7345 & w7355;
assign w7358 = ~w7356 & ~w7357;
assign w7359 = w7344 & ~w7358;
assign w7360 = ~w7344 & w7358;
assign w7361 = ~w7359 & ~w7360;
assign w7362 = ~w7293 & ~w7296;
assign w7363 = pi29 & pi50;
assign w7364 = pi31 & pi48;
assign w7365 = pi30 & pi49;
assign w7366 = ~w7364 & w7365;
assign w7367 = w7364 & ~w7365;
assign w7368 = ~w7366 & ~w7367;
assign w7369 = w7363 & w7368;
assign w7370 = ~w7363 & ~w7368;
assign w7371 = ~w7369 & ~w7370;
assign w7372 = pi26 & pi53;
assign w7373 = pi27 & pi52;
assign w7374 = ~w7221 & ~w7373;
assign w7375 = pi28 & pi52;
assign w7376 = w7219 & w7375;
assign w7377 = ~w7374 & ~w7376;
assign w7378 = w7372 & ~w7377;
assign w7379 = ~w7372 & w7377;
assign w7380 = ~w7378 & ~w7379;
assign w7381 = w7371 & ~w7380;
assign w7382 = ~w7371 & w7380;
assign w7383 = ~w7381 & ~w7382;
assign w7384 = ~w7362 & w7383;
assign w7385 = w7362 & ~w7383;
assign w7386 = ~w7384 & ~w7385;
assign w7387 = (w7386 & w7285) | (w7386 & w9017) | (w7285 & w9017);
assign w7388 = ~w7285 & w9018;
assign w7389 = ~w7387 & ~w7388;
assign w7390 = w7361 & w7389;
assign w7391 = ~w7361 & ~w7389;
assign w7392 = ~w7390 & ~w7391;
assign w7393 = pi23 & pi56;
assign w7394 = pi25 & pi54;
assign w7395 = ~w7242 & ~w7394;
assign w7396 = pi25 & pi55;
assign w7397 = w7146 & w7396;
assign w7398 = ~w7395 & ~w7397;
assign w7399 = w7393 & ~w7398;
assign w7400 = ~w7393 & w7398;
assign w7401 = ~w7399 & ~w7400;
assign w7402 = w7271 & ~w7401;
assign w7403 = ~w7271 & w7401;
assign w7404 = ~w7402 & ~w7403;
assign w7405 = pi20 & pi59;
assign w7406 = pi21 & pi58;
assign w7407 = ~w7259 & ~w7406;
assign w7408 = pi22 & pi58;
assign w7409 = w7040 & w7408;
assign w7410 = ~w7407 & ~w7409;
assign w7411 = w7405 & ~w7410;
assign w7412 = ~w7405 & w7410;
assign w7413 = ~w7411 & ~w7412;
assign w7414 = w7404 & ~w7413;
assign w7415 = ~w7404 & w7413;
assign w7416 = ~w7414 & ~w7415;
assign w7417 = ~w7265 & ~w7277;
assign w7418 = w7268 & ~w7270;
assign w7419 = ~w7272 & ~w7418;
assign w7420 = w7256 & ~w7258;
assign w7421 = ~w7260 & ~w7420;
assign w7422 = ~w7419 & ~w7421;
assign w7423 = w7419 & w7421;
assign w7424 = ~w7422 & ~w7423;
assign w7425 = ~w7417 & w7424;
assign w7426 = w7417 & ~w7424;
assign w7427 = ~w7425 & ~w7426;
assign w7428 = (~w7234 & ~w7204) | (~w7234 & w8905) | (~w7204 & w8905);
assign w7429 = ~w7231 & w9311;
assign w7430 = (w7201 & w9019) | (w7201 & w9020) | (w9019 & w9020);
assign w7431 = ~w7429 & ~w7430;
assign w7432 = ~w7428 & w7431;
assign w7433 = w7428 & ~w7431;
assign w7434 = ~w7432 & ~w7433;
assign w7435 = w7427 & w7434;
assign w7436 = ~w7427 & ~w7434;
assign w7437 = ~w7435 & ~w7436;
assign w7438 = w7416 & w7437;
assign w7439 = ~w7416 & ~w7437;
assign w7440 = ~w7438 & ~w7439;
assign w7441 = w7392 & w7440;
assign w7442 = ~w7392 & ~w7440;
assign w7443 = ~w7441 & ~w7442;
assign w7444 = ~w7312 & ~w7315;
assign w7445 = (~w7252 & ~w7304) | (~w7252 & w9021) | (~w7304 & w9021);
assign w7446 = ~w7246 & ~w7249;
assign w7447 = (~w7299 & ~w7301) | (~w7299 & w9022) | (~w7301 & w9022);
assign w7448 = ~w7446 & ~w7447;
assign w7449 = w7446 & w7447;
assign w7450 = ~w7448 & ~w7449;
assign w7451 = ~w7445 & w7450;
assign w7452 = w7445 & ~w7450;
assign w7453 = ~w7451 & ~w7452;
assign w7454 = ~w7444 & w7453;
assign w7455 = w7444 & ~w7453;
assign w7456 = ~w7454 & ~w7455;
assign w7457 = w7443 & w7456;
assign w7458 = ~w7443 & ~w7456;
assign w7459 = ~w7457 & ~w7458;
assign w7460 = ~w7331 & w7459;
assign w7461 = w7331 & ~w7459;
assign w7462 = ~w7460 & ~w7461;
assign w7463 = w7030 & w7182;
assign w7464 = ~w7325 & w7463;
assign w7465 = w7028 & ~w7180;
assign w7466 = ~w7181 & ~w7324;
assign w7467 = ~w7465 & w7466;
assign w7468 = ~w7325 & ~w7467;
assign w7469 = (~w7468 & w6870) | (~w7468 & w8907) | (w6870 & w8907);
assign w7470 = w6132 & w7469;
assign w7471 = ~w6137 & w7470;
assign w7472 = w7326 & w7463;
assign w7473 = w6872 & w7472;
assign w7474 = w7469 & ~w7473;
assign w7475 = ~w7474 & w9312;
assign w7476 = w7462 & w9313;
assign w7477 = ~w7475 & ~w7476;
assign w7478 = (~w7454 & ~w7456) | (~w7454 & w9060) | (~w7456 & w9060);
assign w7479 = pi21 & pi59;
assign w7480 = pi27 & pi53;
assign w7481 = pi26 & pi54;
assign w7482 = ~w7480 & ~w7481;
assign w7483 = pi27 & pi54;
assign w7484 = w7372 & w7483;
assign w7485 = ~w7482 & ~w7484;
assign w7486 = w7396 & ~w7485;
assign w7487 = ~w7396 & w7485;
assign w7488 = ~w7486 & ~w7487;
assign w7489 = w7479 & ~w7488;
assign w7490 = ~w7479 & w7488;
assign w7491 = ~w7489 & ~w7490;
assign w7492 = pi24 & pi56;
assign w7493 = pi23 & pi57;
assign w7494 = ~w7492 & ~w7493;
assign w7495 = pi24 & pi57;
assign w7496 = w7393 & w7495;
assign w7497 = ~w7494 & ~w7496;
assign w7498 = w7408 & ~w7497;
assign w7499 = ~w7408 & w7497;
assign w7500 = ~w7498 & ~w7499;
assign w7501 = w7491 & ~w7500;
assign w7502 = ~w7491 & w7500;
assign w7503 = ~w7501 & ~w7502;
assign w7504 = ~w7402 & ~w7414;
assign w7505 = w7405 & ~w7407;
assign w7506 = ~w7409 & ~w7505;
assign w7507 = w7393 & ~w7395;
assign w7508 = ~w7397 & ~w7507;
assign w7509 = ~w7506 & ~w7508;
assign w7510 = w7506 & w7508;
assign w7511 = ~w7509 & ~w7510;
assign w7512 = ~w7504 & w7511;
assign w7513 = w7504 & ~w7511;
assign w7514 = ~w7512 & ~w7513;
assign w7515 = (~w7342 & w7358) | (~w7342 & w9061) | (w7358 & w9061);
assign w7516 = ~w7337 & ~w7340;
assign w7517 = ~w7356 & ~w7516;
assign w7518 = w7356 & w7516;
assign w7519 = ~w7517 & ~w7518;
assign w7520 = ~w7515 & w7519;
assign w7521 = w7515 & ~w7519;
assign w7522 = ~w7520 & ~w7521;
assign w7523 = w7514 & w7522;
assign w7524 = ~w7514 & ~w7522;
assign w7525 = ~w7523 & ~w7524;
assign w7526 = w7503 & w7525;
assign w7527 = ~w7503 & ~w7525;
assign w7528 = ~w7526 & ~w7527;
assign w7529 = ~w7366 & ~w7369;
assign w7530 = w7372 & ~w7374;
assign w7531 = ~w7376 & ~w7530;
assign w7532 = ~w7529 & ~w7531;
assign w7533 = w7529 & w7531;
assign w7534 = ~w7532 & ~w7533;
assign w7535 = w7381 & w7534;
assign w7536 = ~w7381 & ~w7534;
assign w7537 = ~w7535 & ~w7536;
assign w7538 = pi20 & pi60;
assign w7539 = pi19 & pi61;
assign w7540 = ~w7538 & ~w7539;
assign w7541 = pi20 & pi61;
assign w7542 = w7271 & w7541;
assign w7543 = ~w7540 & ~w7542;
assign w7544 = w7336 & ~w7543;
assign w7545 = ~w7336 & w7543;
assign w7546 = ~w7544 & ~w7545;
assign w7547 = w7537 & ~w7546;
assign w7548 = ~w7537 & w7546;
assign w7549 = ~w7547 & ~w7548;
assign w7550 = pi17 & pi63;
assign w7551 = (~w7350 & w7346) | (~w7350 & w9062) | (w7346 & w9062);
assign w7552 = w7550 & w7551;
assign w7553 = ~w7550 & ~w7551;
assign w7554 = ~w7552 & ~w7553;
assign w7555 = w7549 & ~w7554;
assign w7556 = ~w7549 & w7554;
assign w7557 = ~w7555 & ~w7556;
assign w7558 = (~w7429 & w7428) | (~w7429 & w9023) | (w7428 & w9023);
assign w7559 = ~w7422 & ~w7425;
assign w7560 = pi29 & pi51;
assign w7561 = pi31 & pi49;
assign w7562 = pi30 & pi50;
assign w7563 = ~w7561 & w7562;
assign w7564 = w7561 & ~w7562;
assign w7565 = ~w7563 & ~w7564;
assign w7566 = w7560 & w7565;
assign w7567 = ~w7560 & ~w7565;
assign w7568 = ~w7566 & ~w7567;
assign w7569 = w7375 & w7568;
assign w7570 = ~w7375 & ~w7568;
assign w7571 = ~w7569 & ~w7570;
assign w7572 = ~w7559 & w7571;
assign w7573 = w7559 & ~w7571;
assign w7574 = ~w7572 & ~w7573;
assign w7575 = ~w7558 & w7574;
assign w7576 = w7558 & ~w7574;
assign w7577 = ~w7575 & ~w7576;
assign w7578 = w7557 & w7577;
assign w7579 = ~w7557 & ~w7577;
assign w7580 = ~w7578 & ~w7579;
assign w7581 = w7528 & w7580;
assign w7582 = ~w7528 & ~w7580;
assign w7583 = ~w7581 & ~w7582;
assign w7584 = ~w7448 & ~w7451;
assign w7585 = (~w7390 & ~w7440) | (~w7390 & w9024) | (~w7440 & w9024);
assign w7586 = ~w7384 & ~w7387;
assign w7587 = (~w7435 & ~w7437) | (~w7435 & w9025) | (~w7437 & w9025);
assign w7588 = ~w7586 & ~w7587;
assign w7589 = w7586 & w7587;
assign w7590 = ~w7588 & ~w7589;
assign w7591 = ~w7585 & w7590;
assign w7592 = w7585 & ~w7590;
assign w7593 = ~w7591 & ~w7592;
assign w7594 = ~w7584 & w7593;
assign w7595 = w7584 & ~w7593;
assign w7596 = ~w7594 & ~w7595;
assign w7597 = w7583 & w7596;
assign w7598 = ~w7583 & ~w7596;
assign w7599 = ~w7597 & ~w7598;
assign w7600 = ~w7478 & w7599;
assign w7601 = w7478 & ~w7599;
assign w7602 = ~w7600 & ~w7601;
assign w7603 = (w9064 & w9284) | (w9064 & w9285) | (w9284 & w9285);
assign w7604 = ~w7461 & w7602;
assign w7605 = (w6137 & w9190) | (w6137 & w9191) | (w9190 & w9191);
assign w7606 = ~w7603 & ~w7605;
assign w7607 = (~w7594 & ~w7596) | (~w7594 & w9067) | (~w7596 & w9067);
assign w7608 = pi22 & pi59;
assign w7609 = pi26 & pi55;
assign w7610 = pi28 & pi53;
assign w7611 = ~w7483 & ~w7610;
assign w7612 = pi28 & pi54;
assign w7613 = w7480 & w7612;
assign w7614 = ~w7611 & ~w7613;
assign w7615 = w7609 & ~w7614;
assign w7616 = ~w7609 & w7614;
assign w7617 = ~w7615 & ~w7616;
assign w7618 = w7608 & ~w7617;
assign w7619 = ~w7608 & w7617;
assign w7620 = ~w7618 & ~w7619;
assign w7621 = pi23 & pi58;
assign w7622 = pi25 & pi56;
assign w7623 = ~w7495 & ~w7622;
assign w7624 = pi25 & pi57;
assign w7625 = w7492 & w7624;
assign w7626 = ~w7623 & ~w7625;
assign w7627 = w7621 & ~w7626;
assign w7628 = ~w7621 & w7626;
assign w7629 = ~w7627 & ~w7628;
assign w7630 = w7620 & ~w7629;
assign w7631 = ~w7620 & w7629;
assign w7632 = ~w7630 & ~w7631;
assign w7633 = ~w7489 & ~w7501;
assign w7634 = w7408 & ~w7494;
assign w7635 = ~w7496 & ~w7634;
assign w7636 = w7396 & ~w7482;
assign w7637 = ~w7484 & ~w7636;
assign w7638 = ~w7635 & ~w7637;
assign w7639 = w7635 & w7637;
assign w7640 = ~w7638 & ~w7639;
assign w7641 = ~w7633 & w7640;
assign w7642 = w7633 & ~w7640;
assign w7643 = ~w7641 & ~w7642;
assign w7644 = ~w7547 & ~w7555;
assign w7645 = w7336 & ~w7540;
assign w7646 = ~w7542 & ~w7645;
assign w7647 = ~w7552 & ~w7646;
assign w7648 = w7552 & w7646;
assign w7649 = ~w7647 & ~w7648;
assign w7650 = ~w7644 & w7649;
assign w7651 = w7644 & ~w7649;
assign w7652 = ~w7650 & ~w7651;
assign w7653 = w7643 & w7652;
assign w7654 = ~w7643 & ~w7652;
assign w7655 = ~w7653 & ~w7654;
assign w7656 = w7632 & w7655;
assign w7657 = ~w7632 & ~w7655;
assign w7658 = ~w7656 & ~w7657;
assign w7659 = w7563 & w7569;
assign w7660 = ~w7563 & ~w7569;
assign w7661 = ~w7659 & ~w7660;
assign w7662 = ~w7566 & ~w7661;
assign w7663 = pi19 & pi62;
assign w7664 = pi21 & pi60;
assign w7665 = ~w7541 & ~w7664;
assign w7666 = pi21 & pi61;
assign w7667 = w7538 & w7666;
assign w7668 = ~w7665 & ~w7667;
assign w7669 = w7663 & ~w7668;
assign w7670 = ~w7663 & w7668;
assign w7671 = ~w7669 & ~w7670;
assign w7672 = ~w7662 & ~w7671;
assign w7673 = w7662 & w7671;
assign w7674 = ~w7672 & ~w7673;
assign w7675 = pi18 & pi63;
assign w7676 = ~w7532 & ~w7535;
assign w7677 = w7675 & w7676;
assign w7678 = ~w7675 & ~w7676;
assign w7679 = ~w7677 & ~w7678;
assign w7680 = w7674 & ~w7679;
assign w7681 = ~w7674 & w7679;
assign w7682 = ~w7680 & ~w7681;
assign w7683 = ~w7517 & ~w7520;
assign w7684 = ~w7509 & ~w7512;
assign w7685 = pi29 & pi52;
assign w7686 = pi31 & pi50;
assign w7687 = pi30 & pi51;
assign w7688 = ~w7686 & w7687;
assign w7689 = w7686 & ~w7687;
assign w7690 = ~w7688 & ~w7689;
assign w7691 = w7685 & w7690;
assign w7692 = ~w7685 & ~w7690;
assign w7693 = ~w7691 & ~w7692;
assign w7694 = ~w7684 & w7693;
assign w7695 = w7684 & ~w7693;
assign w7696 = ~w7694 & ~w7695;
assign w7697 = ~w7683 & w7696;
assign w7698 = w7683 & ~w7696;
assign w7699 = ~w7697 & ~w7698;
assign w7700 = w7682 & w7699;
assign w7701 = ~w7682 & ~w7699;
assign w7702 = ~w7700 & ~w7701;
assign w7703 = w7658 & w7702;
assign w7704 = ~w7658 & ~w7702;
assign w7705 = ~w7703 & ~w7704;
assign w7706 = ~w7588 & ~w7591;
assign w7707 = (~w7578 & ~w7580) | (~w7578 & w9068) | (~w7580 & w9068);
assign w7708 = ~w7523 & ~w7526;
assign w7709 = ~w7572 & ~w7575;
assign w7710 = ~w7708 & ~w7709;
assign w7711 = w7708 & w7709;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = ~w7707 & w7712;
assign w7714 = w7707 & ~w7712;
assign w7715 = ~w7713 & ~w7714;
assign w7716 = ~w7706 & w7715;
assign w7717 = w7706 & ~w7715;
assign w7718 = ~w7716 & ~w7717;
assign w7719 = w7705 & w7718;
assign w7720 = ~w7705 & ~w7718;
assign w7721 = ~w7719 & ~w7720;
assign w7722 = w7607 & ~w7721;
assign w7723 = ~w7607 & w7721;
assign w7724 = ~w7722 & ~w7723;
assign w7725 = w8779 & ~w7605;
assign w7726 = ~w7724 & w9314;
assign w7727 = ~w7725 & ~w7726;
assign w7728 = (~w7716 & ~w7718) | (~w7716 & w9069) | (~w7718 & w9069);
assign w7729 = pi23 & pi59;
assign w7730 = pi27 & pi55;
assign w7731 = pi29 & pi53;
assign w7732 = ~w7612 & ~w7731;
assign w7733 = pi29 & pi54;
assign w7734 = w7610 & w7733;
assign w7735 = ~w7732 & ~w7734;
assign w7736 = w7730 & ~w7735;
assign w7737 = ~w7730 & w7735;
assign w7738 = ~w7736 & ~w7737;
assign w7739 = w7729 & ~w7738;
assign w7740 = ~w7729 & w7738;
assign w7741 = ~w7739 & ~w7740;
assign w7742 = pi24 & pi58;
assign w7743 = pi26 & pi56;
assign w7744 = ~w7624 & ~w7743;
assign w7745 = pi26 & pi57;
assign w7746 = w7622 & w7745;
assign w7747 = ~w7744 & ~w7746;
assign w7748 = w7742 & ~w7747;
assign w7749 = ~w7742 & w7747;
assign w7750 = ~w7748 & ~w7749;
assign w7751 = w7741 & ~w7750;
assign w7752 = ~w7741 & w7750;
assign w7753 = ~w7751 & ~w7752;
assign w7754 = ~w7618 & ~w7630;
assign w7755 = w7621 & ~w7623;
assign w7756 = ~w7625 & ~w7755;
assign w7757 = w7609 & ~w7611;
assign w7758 = ~w7613 & ~w7757;
assign w7759 = ~w7756 & ~w7758;
assign w7760 = w7756 & w7758;
assign w7761 = ~w7759 & ~w7760;
assign w7762 = ~w7754 & w7761;
assign w7763 = w7754 & ~w7761;
assign w7764 = ~w7762 & ~w7763;
assign w7765 = ~w7672 & ~w7680;
assign w7766 = w7663 & ~w7665;
assign w7767 = ~w7667 & ~w7766;
assign w7768 = ~w7677 & ~w7767;
assign w7769 = w7677 & w7767;
assign w7770 = ~w7768 & ~w7769;
assign w7771 = ~w7765 & w7770;
assign w7772 = w7765 & ~w7770;
assign w7773 = ~w7771 & ~w7772;
assign w7774 = w7764 & w7773;
assign w7775 = ~w7764 & ~w7773;
assign w7776 = ~w7774 & ~w7775;
assign w7777 = w7753 & w7776;
assign w7778 = ~w7753 & ~w7776;
assign w7779 = ~w7777 & ~w7778;
assign w7780 = pi19 & pi63;
assign w7781 = ~w7659 & w7780;
assign w7782 = w7659 & ~w7780;
assign w7783 = ~w7781 & ~w7782;
assign w7784 = ~w7688 & ~w7691;
assign w7785 = pi20 & pi62;
assign w7786 = pi22 & pi60;
assign w7787 = ~w7666 & ~w7786;
assign w7788 = pi22 & pi61;
assign w7789 = w7664 & w7788;
assign w7790 = ~w7787 & ~w7789;
assign w7791 = w7785 & ~w7790;
assign w7792 = ~w7785 & w7790;
assign w7793 = ~w7791 & ~w7792;
assign w7794 = ~w7784 & ~w7793;
assign w7795 = w7784 & w7793;
assign w7796 = ~w7794 & ~w7795;
assign w7797 = ~w7783 & w7796;
assign w7798 = w7783 & ~w7796;
assign w7799 = ~w7797 & ~w7798;
assign w7800 = ~w7647 & ~w7650;
assign w7801 = ~w7638 & ~w7641;
assign w7802 = pi31 & pi51;
assign w7803 = pi30 & pi52;
assign w7804 = ~w7802 & w7803;
assign w7805 = w7802 & ~w7803;
assign w7806 = ~w7804 & ~w7805;
assign w7807 = ~w7801 & w7806;
assign w7808 = w7801 & ~w7806;
assign w7809 = ~w7807 & ~w7808;
assign w7810 = ~w7800 & w7809;
assign w7811 = w7800 & ~w7809;
assign w7812 = ~w7810 & ~w7811;
assign w7813 = w7799 & w7812;
assign w7814 = ~w7799 & ~w7812;
assign w7815 = ~w7813 & ~w7814;
assign w7816 = w7779 & w7815;
assign w7817 = ~w7779 & ~w7815;
assign w7818 = ~w7816 & ~w7817;
assign w7819 = ~w7710 & ~w7713;
assign w7820 = ~w7700 & ~w7703;
assign w7821 = ~w7653 & ~w7656;
assign w7822 = ~w7694 & ~w7697;
assign w7823 = ~w7821 & ~w7822;
assign w7824 = w7821 & w7822;
assign w7825 = ~w7823 & ~w7824;
assign w7826 = ~w7820 & w7825;
assign w7827 = w7820 & ~w7825;
assign w7828 = ~w7826 & ~w7827;
assign w7829 = ~w7819 & w7828;
assign w7830 = w7819 & ~w7828;
assign w7831 = ~w7829 & ~w7830;
assign w7832 = w7818 & w7831;
assign w7833 = ~w7818 & ~w7831;
assign w7834 = ~w7832 & ~w7833;
assign w7835 = ~w7728 & w7834;
assign w7836 = w7728 & ~w7834;
assign w7837 = ~w7835 & ~w7836;
assign w7838 = w7837 & w9315;
assign w7839 = (w7471 & w9192) | (w7471 & w9193) | (w9192 & w9193);
assign w7840 = ~w7838 & ~w7839;
assign w7841 = ~w7829 & ~w7832;
assign w7842 = pi25 & pi58;
assign w7843 = pi31 & pi52;
assign w7844 = pi30 & pi53;
assign w7845 = ~w7843 & w7844;
assign w7846 = w7843 & ~w7844;
assign w7847 = ~w7845 & ~w7846;
assign w7848 = w7733 & w7847;
assign w7849 = ~w7733 & ~w7847;
assign w7850 = ~w7848 & ~w7849;
assign w7851 = w7842 & w7850;
assign w7852 = ~w7842 & ~w7850;
assign w7853 = ~w7851 & ~w7852;
assign w7854 = pi27 & pi56;
assign w7855 = pi28 & pi55;
assign w7856 = ~w7854 & ~w7855;
assign w7857 = pi28 & pi56;
assign w7858 = w7730 & w7857;
assign w7859 = ~w7856 & ~w7858;
assign w7860 = w7745 & ~w7859;
assign w7861 = ~w7745 & w7859;
assign w7862 = ~w7860 & ~w7861;
assign w7863 = w7853 & ~w7862;
assign w7864 = ~w7853 & w7862;
assign w7865 = ~w7863 & ~w7864;
assign w7866 = ~w7794 & ~w7797;
assign w7867 = w7785 & ~w7787;
assign w7868 = ~w7789 & ~w7867;
assign w7869 = ~w7781 & ~w7868;
assign w7870 = w7781 & w7868;
assign w7871 = ~w7869 & ~w7870;
assign w7872 = ~w7866 & w7871;
assign w7873 = w7866 & ~w7871;
assign w7874 = ~w7872 & ~w7873;
assign w7875 = ~w7739 & ~w7751;
assign w7876 = w7742 & ~w7744;
assign w7877 = ~w7746 & ~w7876;
assign w7878 = w7730 & ~w7732;
assign w7879 = ~w7734 & ~w7878;
assign w7880 = ~w7877 & ~w7879;
assign w7881 = w7877 & w7879;
assign w7882 = ~w7880 & ~w7881;
assign w7883 = ~w7875 & w7882;
assign w7884 = w7875 & ~w7882;
assign w7885 = ~w7883 & ~w7884;
assign w7886 = w7874 & w7885;
assign w7887 = ~w7874 & ~w7885;
assign w7888 = ~w7886 & ~w7887;
assign w7889 = w7865 & w7888;
assign w7890 = ~w7865 & ~w7888;
assign w7891 = ~w7889 & ~w7890;
assign w7892 = pi20 & pi63;
assign w7893 = pi21 & pi62;
assign w7894 = w7892 & ~w7893;
assign w7895 = ~w7892 & w7893;
assign w7896 = ~w7894 & ~w7895;
assign w7897 = pi23 & pi60;
assign w7898 = pi24 & pi59;
assign w7899 = ~w7897 & ~w7898;
assign w7900 = pi24 & pi60;
assign w7901 = w7729 & w7900;
assign w7902 = ~w7899 & ~w7901;
assign w7903 = w7788 & ~w7902;
assign w7904 = ~w7788 & w7902;
assign w7905 = ~w7903 & ~w7904;
assign w7906 = ~w7896 & ~w7905;
assign w7907 = w7896 & w7905;
assign w7908 = ~w7906 & ~w7907;
assign w7909 = ~w7768 & ~w7771;
assign w7910 = ~w7759 & ~w7762;
assign w7911 = w7804 & ~w7910;
assign w7912 = ~w7804 & w7910;
assign w7913 = ~w7911 & ~w7912;
assign w7914 = ~w7909 & w7913;
assign w7915 = w7909 & ~w7913;
assign w7916 = ~w7914 & ~w7915;
assign w7917 = w7908 & w7916;
assign w7918 = ~w7908 & ~w7916;
assign w7919 = ~w7917 & ~w7918;
assign w7920 = w7891 & w7919;
assign w7921 = ~w7891 & ~w7919;
assign w7922 = ~w7920 & ~w7921;
assign w7923 = ~w7823 & ~w7826;
assign w7924 = ~w7813 & ~w7816;
assign w7925 = ~w7774 & ~w7777;
assign w7926 = ~w7807 & ~w7810;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = w7925 & w7926;
assign w7929 = ~w7927 & ~w7928;
assign w7930 = ~w7924 & w7929;
assign w7931 = w7924 & ~w7929;
assign w7932 = ~w7930 & ~w7931;
assign w7933 = ~w7923 & w7932;
assign w7934 = w7923 & ~w7932;
assign w7935 = ~w7933 & ~w7934;
assign w7936 = w7922 & w7935;
assign w7937 = ~w7922 & ~w7935;
assign w7938 = ~w7936 & ~w7937;
assign w7939 = ~w7841 & w7938;
assign w7940 = w7841 & ~w7938;
assign w7941 = ~w7939 & ~w7940;
assign w7942 = (w7471 & w9194) | (w7471 & w9195) | (w9194 & w9195);
assign w7943 = (w9072 & w9073) | (w9072 & w9315) | (w9073 & w9315);
assign w7944 = ~w7942 & ~w7943;
assign w7945 = ~w7600 & ~w7723;
assign w7946 = ~w7722 & ~w7836;
assign w7947 = ~w7945 & w7946;
assign w7948 = ~w7835 & ~w7939;
assign w7949 = (~w7940 & w7947) | (~w7940 & w9074) | (w7947 & w9074);
assign w7950 = w7724 & w7837;
assign w7951 = w7941 & w7950;
assign w7952 = w7604 & w7951;
assign w7953 = (w6137 & w9196) | (w6137 & w9197) | (w9196 & w9197);
assign w7954 = ~w7933 & ~w7936;
assign w7955 = pi25 & pi59;
assign w7956 = pi29 & pi55;
assign w7957 = pi31 & pi53;
assign w7958 = pi30 & pi54;
assign w7959 = ~w7957 & w7958;
assign w7960 = w7957 & ~w7958;
assign w7961 = ~w7959 & ~w7960;
assign w7962 = w7956 & w7961;
assign w7963 = ~w7956 & ~w7961;
assign w7964 = ~w7962 & ~w7963;
assign w7965 = w7955 & w7964;
assign w7966 = ~w7955 & ~w7964;
assign w7967 = ~w7965 & ~w7966;
assign w7968 = pi26 & pi58;
assign w7969 = pi27 & pi57;
assign w7970 = ~w7857 & ~w7969;
assign w7971 = pi28 & pi57;
assign w7972 = w7854 & w7971;
assign w7973 = ~w7970 & ~w7972;
assign w7974 = w7968 & ~w7973;
assign w7975 = ~w7968 & w7973;
assign w7976 = ~w7974 & ~w7975;
assign w7977 = w7967 & ~w7976;
assign w7978 = ~w7967 & w7976;
assign w7979 = ~w7977 & ~w7978;
assign w7980 = w7788 & ~w7899;
assign w7981 = ~w7901 & ~w7980;
assign w7982 = ~w7894 & ~w7981;
assign w7983 = w7894 & w7981;
assign w7984 = ~w7982 & ~w7983;
assign w7985 = w7906 & w7984;
assign w7986 = ~w7906 & ~w7984;
assign w7987 = ~w7985 & ~w7986;
assign w7988 = ~w7851 & ~w7863;
assign w7989 = ~w7845 & ~w7848;
assign w7990 = w7745 & ~w7856;
assign w7991 = ~w7858 & ~w7990;
assign w7992 = ~w7989 & ~w7991;
assign w7993 = w7989 & w7991;
assign w7994 = ~w7992 & ~w7993;
assign w7995 = ~w7988 & w7994;
assign w7996 = w7988 & ~w7994;
assign w7997 = ~w7995 & ~w7996;
assign w7998 = w7987 & w7997;
assign w7999 = ~w7987 & ~w7997;
assign w8000 = ~w7998 & ~w7999;
assign w8001 = w7979 & w8000;
assign w8002 = ~w7979 & ~w8000;
assign w8003 = ~w8001 & ~w8002;
assign w8004 = pi21 & pi63;
assign w8005 = pi22 & pi62;
assign w8006 = pi23 & pi61;
assign w8007 = ~w7900 & ~w8006;
assign w8008 = pi24 & pi61;
assign w8009 = w7897 & w8008;
assign w8010 = ~w8007 & ~w8009;
assign w8011 = w8005 & w8010;
assign w8012 = ~w8005 & ~w8010;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = w8004 & ~w8013;
assign w8015 = ~w8004 & w8013;
assign w8016 = ~w8014 & ~w8015;
assign w8017 = ~w7869 & ~w7872;
assign w8018 = ~w7880 & ~w7883;
assign w8019 = w8017 & w8018;
assign w8020 = ~w8017 & ~w8018;
assign w8021 = ~w8019 & ~w8020;
assign w8022 = w8016 & ~w8021;
assign w8023 = ~w8016 & w8021;
assign w8024 = ~w8022 & ~w8023;
assign w8025 = w8003 & w8024;
assign w8026 = ~w8003 & ~w8024;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = ~w7927 & ~w7930;
assign w8029 = ~w7917 & ~w7920;
assign w8030 = ~w7886 & ~w7889;
assign w8031 = ~w7911 & ~w7914;
assign w8032 = ~w8030 & ~w8031;
assign w8033 = w8030 & w8031;
assign w8034 = ~w8032 & ~w8033;
assign w8035 = ~w8029 & w8034;
assign w8036 = w8029 & ~w8034;
assign w8037 = ~w8035 & ~w8036;
assign w8038 = ~w8028 & w8037;
assign w8039 = w8028 & ~w8037;
assign w8040 = ~w8038 & ~w8039;
assign w8041 = w8027 & w8040;
assign w8042 = ~w8027 & ~w8040;
assign w8043 = ~w8041 & ~w8042;
assign w8044 = ~w7954 & w8043;
assign w8045 = w7954 & ~w8043;
assign w8046 = ~w8044 & ~w8045;
assign w8047 = w8046 & w9316;
assign w8048 = (w7471 & w9198) | (w7471 & w9199) | (w9198 & w9199);
assign w8049 = ~w8047 & ~w8048;
assign w8050 = ~w8038 & ~w8041;
assign w8051 = pi22 & pi63;
assign w8052 = pi23 & pi62;
assign w8053 = ~w8008 & ~w8052;
assign w8054 = pi24 & pi62;
assign w8055 = w8006 & w8054;
assign w8056 = ~w8053 & ~w8055;
assign w8057 = w8051 & ~w8056;
assign w8058 = ~w8051 & w8056;
assign w8059 = ~w8057 & ~w8058;
assign w8060 = ~w7982 & ~w7985;
assign w8061 = ~w7992 & ~w7995;
assign w8062 = w8060 & w8061;
assign w8063 = ~w8060 & ~w8061;
assign w8064 = ~w8062 & ~w8063;
assign w8065 = ~w8059 & w8064;
assign w8066 = w8059 & ~w8064;
assign w8067 = ~w8065 & ~w8066;
assign w8068 = pi25 & pi60;
assign w8069 = pi29 & pi56;
assign w8070 = pi31 & pi54;
assign w8071 = pi30 & pi55;
assign w8072 = ~w8070 & w8071;
assign w8073 = w8070 & ~w8071;
assign w8074 = ~w8072 & ~w8073;
assign w8075 = w8069 & w8074;
assign w8076 = ~w8069 & ~w8074;
assign w8077 = ~w8075 & ~w8076;
assign w8078 = w8068 & w8077;
assign w8079 = ~w8068 & ~w8077;
assign w8080 = ~w8078 & ~w8079;
assign w8081 = pi26 & pi59;
assign w8082 = pi27 & pi58;
assign w8083 = ~w7971 & ~w8082;
assign w8084 = pi28 & pi58;
assign w8085 = w7969 & w8084;
assign w8086 = ~w8083 & ~w8085;
assign w8087 = w8081 & ~w8086;
assign w8088 = ~w8081 & w8086;
assign w8089 = ~w8087 & ~w8088;
assign w8090 = w8080 & ~w8089;
assign w8091 = ~w8080 & w8089;
assign w8092 = ~w8090 & ~w8091;
assign w8093 = ~w7965 & ~w7977;
assign w8094 = ~w7959 & ~w7962;
assign w8095 = w7968 & ~w7970;
assign w8096 = ~w7972 & ~w8095;
assign w8097 = ~w8094 & ~w8096;
assign w8098 = w8094 & w8096;
assign w8099 = ~w8097 & ~w8098;
assign w8100 = ~w8093 & w8099;
assign w8101 = w8093 & ~w8099;
assign w8102 = ~w8100 & ~w8101;
assign w8103 = w8009 & w8015;
assign w8104 = ~w8009 & ~w8015;
assign w8105 = ~w8103 & ~w8104;
assign w8106 = ~w8011 & ~w8105;
assign w8107 = w8102 & ~w8106;
assign w8108 = ~w8102 & w8106;
assign w8109 = ~w8107 & ~w8108;
assign w8110 = w8092 & w8109;
assign w8111 = ~w8092 & ~w8109;
assign w8112 = ~w8110 & ~w8111;
assign w8113 = w8067 & ~w8112;
assign w8114 = ~w8067 & w8112;
assign w8115 = ~w8113 & ~w8114;
assign w8116 = ~w8032 & ~w8035;
assign w8117 = ~w8022 & ~w8025;
assign w8118 = ~w7998 & ~w8001;
assign w8119 = ~w8019 & ~w8118;
assign w8120 = w8019 & w8118;
assign w8121 = ~w8119 & ~w8120;
assign w8122 = ~w8117 & w8121;
assign w8123 = w8117 & ~w8121;
assign w8124 = ~w8122 & ~w8123;
assign w8125 = ~w8116 & w8124;
assign w8126 = w8116 & ~w8124;
assign w8127 = ~w8125 & ~w8126;
assign w8128 = ~w8115 & w8127;
assign w8129 = w8115 & ~w8127;
assign w8130 = ~w8128 & ~w8129;
assign w8131 = w8050 & ~w8130;
assign w8132 = ~w8050 & w8130;
assign w8133 = ~w8131 & ~w8132;
assign w8134 = (w7471 & w9200) | (w7471 & w9201) | (w9200 & w9201);
assign w8135 = (w9075 & w9076) | (w9075 & w9316) | (w9076 & w9316);
assign w8136 = ~w8134 & ~w8135;
assign w8137 = w8044 & ~w8131;
assign w8138 = ~w8132 & ~w8137;
assign w8139 = ~w8045 & ~w8131;
assign w8140 = ~w8132 & ~w8139;
assign w8141 = ~w8125 & ~w8128;
assign w8142 = pi25 & pi61;
assign w8143 = pi29 & pi57;
assign w8144 = pi31 & pi55;
assign w8145 = pi30 & pi56;
assign w8146 = ~w8144 & w8145;
assign w8147 = w8144 & ~w8145;
assign w8148 = ~w8146 & ~w8147;
assign w8149 = w8143 & w8148;
assign w8150 = ~w8143 & ~w8148;
assign w8151 = ~w8149 & ~w8150;
assign w8152 = w8142 & w8151;
assign w8153 = ~w8142 & ~w8151;
assign w8154 = ~w8152 & ~w8153;
assign w8155 = pi26 & pi60;
assign w8156 = pi27 & pi59;
assign w8157 = ~w8084 & ~w8156;
assign w8158 = pi28 & pi59;
assign w8159 = w8082 & w8158;
assign w8160 = ~w8157 & ~w8159;
assign w8161 = w8155 & ~w8160;
assign w8162 = ~w8155 & w8160;
assign w8163 = ~w8161 & ~w8162;
assign w8164 = w8154 & ~w8163;
assign w8165 = ~w8154 & w8163;
assign w8166 = ~w8164 & ~w8165;
assign w8167 = ~w8078 & ~w8090;
assign w8168 = ~w8072 & ~w8075;
assign w8169 = w8081 & ~w8083;
assign w8170 = ~w8085 & ~w8169;
assign w8171 = ~w8168 & ~w8170;
assign w8172 = w8168 & w8170;
assign w8173 = ~w8171 & ~w8172;
assign w8174 = ~w8167 & w8173;
assign w8175 = w8167 & ~w8173;
assign w8176 = ~w8174 & ~w8175;
assign w8177 = ~w8055 & ~w8058;
assign w8178 = w8176 & ~w8177;
assign w8179 = ~w8176 & w8177;
assign w8180 = ~w8178 & ~w8179;
assign w8181 = w8166 & w8180;
assign w8182 = ~w8166 & ~w8180;
assign w8183 = ~w8181 & ~w8182;
assign w8184 = pi23 & pi63;
assign w8185 = w8054 & ~w8184;
assign w8186 = ~w8054 & w8184;
assign w8187 = ~w8185 & ~w8186;
assign w8188 = ~w8097 & ~w8100;
assign w8189 = ~w8103 & w8188;
assign w8190 = w8103 & ~w8188;
assign w8191 = ~w8189 & ~w8190;
assign w8192 = w8187 & ~w8191;
assign w8193 = ~w8187 & w8191;
assign w8194 = ~w8192 & ~w8193;
assign w8195 = w8183 & w8194;
assign w8196 = ~w8183 & ~w8194;
assign w8197 = ~w8195 & ~w8196;
assign w8198 = ~w8119 & ~w8122;
assign w8199 = ~w8065 & ~w8113;
assign w8200 = ~w8107 & ~w8110;
assign w8201 = ~w8062 & ~w8200;
assign w8202 = w8062 & w8200;
assign w8203 = ~w8201 & ~w8202;
assign w8204 = w8199 & w8203;
assign w8205 = ~w8199 & ~w8203;
assign w8206 = ~w8204 & ~w8205;
assign w8207 = ~w8198 & w8206;
assign w8208 = w8198 & ~w8206;
assign w8209 = ~w8207 & ~w8208;
assign w8210 = w8197 & w8209;
assign w8211 = ~w8197 & ~w8209;
assign w8212 = ~w8210 & ~w8211;
assign w8213 = ~w8141 & w8212;
assign w8214 = w8141 & ~w8212;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = (w7471 & w9202) | (w7471 & w9203) | (w9202 & w9203);
assign w8217 = ~w8215 & w9317;
assign w8218 = ~w8216 & ~w8217;
assign w8219 = ~w8207 & ~w8210;
assign w8220 = pi29 & pi58;
assign w8221 = pi31 & pi56;
assign w8222 = pi30 & pi57;
assign w8223 = ~w8221 & w8222;
assign w8224 = w8221 & ~w8222;
assign w8225 = ~w8223 & ~w8224;
assign w8226 = w8220 & w8225;
assign w8227 = ~w8220 & ~w8225;
assign w8228 = ~w8226 & ~w8227;
assign w8229 = pi26 & pi61;
assign w8230 = pi27 & pi60;
assign w8231 = ~w8158 & ~w8230;
assign w8232 = pi28 & pi60;
assign w8233 = w8156 & w8232;
assign w8234 = ~w8231 & ~w8233;
assign w8235 = w8229 & ~w8234;
assign w8236 = ~w8229 & w8234;
assign w8237 = ~w8235 & ~w8236;
assign w8238 = w8228 & ~w8237;
assign w8239 = ~w8228 & w8237;
assign w8240 = ~w8238 & ~w8239;
assign w8241 = pi24 & pi63;
assign w8242 = pi25 & pi62;
assign w8243 = w8241 & ~w8242;
assign w8244 = ~w8241 & w8242;
assign w8245 = ~w8243 & ~w8244;
assign w8246 = w8240 & ~w8245;
assign w8247 = ~w8240 & w8245;
assign w8248 = ~w8246 & ~w8247;
assign w8249 = ~w8171 & ~w8174;
assign w8250 = ~w8152 & ~w8164;
assign w8251 = ~w8146 & ~w8149;
assign w8252 = w8155 & ~w8157;
assign w8253 = ~w8159 & ~w8252;
assign w8254 = ~w8251 & ~w8253;
assign w8255 = w8251 & w8253;
assign w8256 = ~w8254 & ~w8255;
assign w8257 = ~w8250 & w8256;
assign w8258 = w8250 & ~w8256;
assign w8259 = ~w8257 & ~w8258;
assign w8260 = ~w8249 & w8259;
assign w8261 = w8249 & ~w8259;
assign w8262 = ~w8260 & ~w8261;
assign w8263 = w8185 & w8262;
assign w8264 = ~w8185 & ~w8262;
assign w8265 = ~w8263 & ~w8264;
assign w8266 = w8248 & w8265;
assign w8267 = ~w8248 & ~w8265;
assign w8268 = ~w8266 & ~w8267;
assign w8269 = ~w8201 & ~w8204;
assign w8270 = ~w8192 & ~w8195;
assign w8271 = ~w8178 & ~w8181;
assign w8272 = ~w8189 & ~w8271;
assign w8273 = w8189 & w8271;
assign w8274 = ~w8272 & ~w8273;
assign w8275 = ~w8270 & w8274;
assign w8276 = w8270 & ~w8274;
assign w8277 = ~w8275 & ~w8276;
assign w8278 = ~w8269 & w8277;
assign w8279 = w8269 & ~w8277;
assign w8280 = ~w8278 & ~w8279;
assign w8281 = w8268 & w8280;
assign w8282 = ~w8268 & ~w8280;
assign w8283 = ~w8281 & ~w8282;
assign w8284 = ~w8219 & w8283;
assign w8285 = w8219 & ~w8283;
assign w8286 = ~w8284 & ~w8285;
assign w8287 = (w7471 & w9204) | (w7471 & w9205) | (w9204 & w9205);
assign w8288 = ~w8214 & w8286;
assign w8289 = (w9197 & w9286) | (w9197 & w9287) | (w9286 & w9287);
assign w8290 = ~w8287 & ~w8289;
assign w8291 = ~w8278 & ~w8281;
assign w8292 = ~w8272 & ~w8275;
assign w8293 = ~w8246 & ~w8266;
assign w8294 = ~w8260 & ~w8263;
assign w8295 = ~w8243 & ~w8294;
assign w8296 = w8243 & w8294;
assign w8297 = ~w8295 & ~w8296;
assign w8298 = ~w8293 & w8297;
assign w8299 = w8293 & ~w8297;
assign w8300 = ~w8298 & ~w8299;
assign w8301 = ~w8292 & w8300;
assign w8302 = w8292 & ~w8300;
assign w8303 = ~w8301 & ~w8302;
assign w8304 = pi29 & pi59;
assign w8305 = pi31 & pi57;
assign w8306 = pi30 & pi58;
assign w8307 = ~w8305 & w8306;
assign w8308 = w8305 & ~w8306;
assign w8309 = ~w8307 & ~w8308;
assign w8310 = w8304 & w8309;
assign w8311 = ~w8304 & ~w8309;
assign w8312 = ~w8310 & ~w8311;
assign w8313 = w8232 & w8312;
assign w8314 = ~w8232 & ~w8312;
assign w8315 = ~w8313 & ~w8314;
assign w8316 = pi25 & pi63;
assign w8317 = pi27 & pi61;
assign w8318 = pi26 & pi62;
assign w8319 = ~w8317 & ~w8318;
assign w8320 = pi27 & pi62;
assign w8321 = w8229 & w8320;
assign w8322 = ~w8319 & ~w8321;
assign w8323 = w8316 & ~w8322;
assign w8324 = ~w8316 & w8322;
assign w8325 = ~w8323 & ~w8324;
assign w8326 = w8315 & w8325;
assign w8327 = ~w8315 & ~w8325;
assign w8328 = ~w8326 & ~w8327;
assign w8329 = ~w8254 & ~w8257;
assign w8330 = ~w8223 & ~w8226;
assign w8331 = w8229 & ~w8231;
assign w8332 = ~w8233 & ~w8331;
assign w8333 = ~w8330 & ~w8332;
assign w8334 = w8330 & w8332;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = w8238 & w8335;
assign w8337 = ~w8238 & ~w8335;
assign w8338 = ~w8336 & ~w8337;
assign w8339 = w8329 & ~w8338;
assign w8340 = ~w8329 & w8338;
assign w8341 = ~w8339 & ~w8340;
assign w8342 = w8328 & ~w8341;
assign w8343 = ~w8328 & w8341;
assign w8344 = ~w8342 & ~w8343;
assign w8345 = w8303 & w8344;
assign w8346 = ~w8303 & ~w8344;
assign w8347 = ~w8345 & ~w8346;
assign w8348 = ~w8291 & w8347;
assign w8349 = w8291 & ~w8347;
assign w8350 = ~w8348 & ~w8349;
assign w8351 = (w9197 & w9288) | (w9197 & w9289) | (w9288 & w9289);
assign w8352 = (w7471 & w9206) | (w7471 & w9207) | (w9206 & w9207);
assign w8353 = ~w8351 & ~w8352;
assign w8354 = ~w8301 & ~w8345;
assign w8355 = pi29 & pi60;
assign w8356 = pi31 & pi58;
assign w8357 = pi30 & pi59;
assign w8358 = ~w8356 & w8357;
assign w8359 = w8356 & ~w8357;
assign w8360 = ~w8358 & ~w8359;
assign w8361 = w8355 & w8360;
assign w8362 = ~w8355 & ~w8360;
assign w8363 = ~w8361 & ~w8362;
assign w8364 = pi26 & pi63;
assign w8365 = pi28 & pi61;
assign w8366 = ~w8320 & ~w8365;
assign w8367 = pi28 & pi62;
assign w8368 = w8317 & w8367;
assign w8369 = ~w8366 & ~w8368;
assign w8370 = w8364 & ~w8369;
assign w8371 = ~w8364 & w8369;
assign w8372 = ~w8370 & ~w8371;
assign w8373 = w8363 & w8372;
assign w8374 = ~w8363 & ~w8372;
assign w8375 = ~w8373 & ~w8374;
assign w8376 = w8307 & w8313;
assign w8377 = ~w8307 & ~w8313;
assign w8378 = ~w8376 & ~w8377;
assign w8379 = ~w8310 & ~w8378;
assign w8380 = ~w8333 & ~w8336;
assign w8381 = w8379 & w8380;
assign w8382 = ~w8379 & ~w8380;
assign w8383 = ~w8381 & ~w8382;
assign w8384 = w8375 & ~w8383;
assign w8385 = ~w8375 & w8383;
assign w8386 = ~w8384 & ~w8385;
assign w8387 = ~w8295 & ~w8298;
assign w8388 = ~w8326 & ~w8342;
assign w8389 = ~w8321 & ~w8324;
assign w8390 = ~w8339 & ~w8389;
assign w8391 = w8339 & w8389;
assign w8392 = ~w8390 & ~w8391;
assign w8393 = ~w8388 & w8392;
assign w8394 = w8388 & ~w8392;
assign w8395 = ~w8393 & ~w8394;
assign w8396 = ~w8387 & w8395;
assign w8397 = w8387 & ~w8395;
assign w8398 = ~w8396 & ~w8397;
assign w8399 = w8386 & w8398;
assign w8400 = ~w8386 & ~w8398;
assign w8401 = ~w8399 & ~w8400;
assign w8402 = w8354 & ~w8401;
assign w8403 = ~w8354 & w8401;
assign w8404 = ~w8402 & ~w8403;
assign w8405 = (~w7953 & w9080) | (~w7953 & w9081) | (w9080 & w9081);
assign w8406 = (w7953 & w9082) | (w7953 & w9083) | (w9082 & w9083);
assign w8407 = ~w8405 & ~w8406;
assign w8408 = w8350 & w8404;
assign w8409 = ~w8348 & ~w8403;
assign w8410 = ~w8402 & ~w8409;
assign w8411 = ~w8408 & ~w8410;
assign w8412 = ~w8284 & ~w8410;
assign w8413 = ~w8396 & ~w8399;
assign w8414 = ~w8358 & ~w8361;
assign w8415 = ~w8376 & ~w8414;
assign w8416 = pi31 & pi59;
assign w8417 = pi30 & pi60;
assign w8418 = ~w8416 & w8417;
assign w8419 = w8416 & ~w8417;
assign w8420 = ~w8418 & ~w8419;
assign w8421 = pi27 & pi63;
assign w8422 = pi29 & pi61;
assign w8423 = ~w8367 & ~w8422;
assign w8424 = pi29 & pi62;
assign w8425 = w8365 & w8424;
assign w8426 = ~w8423 & ~w8425;
assign w8427 = w8421 & ~w8426;
assign w8428 = ~w8421 & w8426;
assign w8429 = ~w8427 & ~w8428;
assign w8430 = w8420 & w8429;
assign w8431 = ~w8420 & ~w8429;
assign w8432 = ~w8430 & ~w8431;
assign w8433 = ~w8415 & w8432;
assign w8434 = w8415 & ~w8432;
assign w8435 = ~w8433 & ~w8434;
assign w8436 = ~w8390 & ~w8393;
assign w8437 = ~w8373 & ~w8384;
assign w8438 = ~w8368 & ~w8371;
assign w8439 = ~w8381 & ~w8438;
assign w8440 = w8381 & w8438;
assign w8441 = ~w8439 & ~w8440;
assign w8442 = ~w8437 & w8441;
assign w8443 = w8437 & ~w8441;
assign w8444 = ~w8442 & ~w8443;
assign w8445 = ~w8436 & w8444;
assign w8446 = w8436 & ~w8444;
assign w8447 = ~w8445 & ~w8446;
assign w8448 = w8435 & w8447;
assign w8449 = ~w8435 & ~w8447;
assign w8450 = ~w8448 & ~w8449;
assign w8451 = ~w8413 & w8450;
assign w8452 = w8413 & ~w8450;
assign w8453 = ~w8451 & ~w8452;
assign w8454 = (~w7471 & w9208) | (~w7471 & w9209) | (w9208 & w9209);
assign w8455 = ~w8410 & w8453;
assign w8456 = (w7471 & w9210) | (w7471 & w9211) | (w9210 & w9211);
assign w8457 = ~w8454 & ~w8456;
assign w8458 = ~w8445 & ~w8448;
assign w8459 = pi28 & pi63;
assign w8460 = ~w8418 & w8459;
assign w8461 = w8418 & ~w8459;
assign w8462 = ~w8460 & ~w8461;
assign w8463 = pi31 & pi60;
assign w8464 = pi30 & pi61;
assign w8465 = ~w8463 & w8464;
assign w8466 = w8463 & ~w8464;
assign w8467 = ~w8465 & ~w8466;
assign w8468 = w8424 & w8467;
assign w8469 = ~w8424 & ~w8467;
assign w8470 = ~w8468 & ~w8469;
assign w8471 = ~w8462 & w8470;
assign w8472 = w8462 & ~w8470;
assign w8473 = ~w8471 & ~w8472;
assign w8474 = ~w8439 & ~w8442;
assign w8475 = ~w8430 & ~w8433;
assign w8476 = ~w8425 & ~w8428;
assign w8477 = ~w8414 & ~w8476;
assign w8478 = w8414 & w8476;
assign w8479 = ~w8477 & ~w8478;
assign w8480 = ~w8475 & w8479;
assign w8481 = w8475 & ~w8479;
assign w8482 = ~w8480 & ~w8481;
assign w8483 = ~w8474 & w8482;
assign w8484 = w8474 & ~w8482;
assign w8485 = ~w8483 & ~w8484;
assign w8486 = w8473 & w8485;
assign w8487 = ~w8473 & ~w8485;
assign w8488 = ~w8486 & ~w8487;
assign w8489 = ~w8458 & w8488;
assign w8490 = w8458 & ~w8488;
assign w8491 = ~w8489 & ~w8490;
assign w8492 = (w7953 & w9086) | (w7953 & w9087) | (w9086 & w9087);
assign w8493 = ~w8451 & ~w8491;
assign w8494 = w8451 & w8491;
assign w8495 = ~w8493 & ~w8494;
assign w8496 = (~w7953 & w9088) | (~w7953 & w9089) | (w9088 & w9089);
assign w8497 = ~w8492 & ~w8496;
assign w8498 = ~w8483 & ~w8486;
assign w8499 = ~w8465 & ~w8468;
assign w8500 = ~w8460 & ~w8499;
assign w8501 = w8460 & w8499;
assign w8502 = ~w8500 & ~w8501;
assign w8503 = w8471 & w8502;
assign w8504 = ~w8471 & ~w8502;
assign w8505 = ~w8503 & ~w8504;
assign w8506 = ~w8477 & ~w8480;
assign w8507 = w8505 & ~w8506;
assign w8508 = ~w8505 & w8506;
assign w8509 = ~w8507 & ~w8508;
assign w8510 = pi29 & pi63;
assign w8511 = pi31 & pi61;
assign w8512 = pi30 & pi62;
assign w8513 = w8511 & ~w8512;
assign w8514 = ~w8511 & w8512;
assign w8515 = ~w8513 & ~w8514;
assign w8516 = w8510 & ~w8515;
assign w8517 = ~w8510 & w8515;
assign w8518 = ~w8516 & ~w8517;
assign w8519 = w8509 & ~w8518;
assign w8520 = ~w8509 & w8518;
assign w8521 = ~w8519 & ~w8520;
assign w8522 = ~w8498 & w8521;
assign w8523 = w8498 & ~w8521;
assign w8524 = ~w8522 & ~w8523;
assign w8525 = ~w8452 & ~w8490;
assign w8526 = ~w8455 & w8525;
assign w8527 = ~w8489 & ~w8526;
assign w8528 = ~w8284 & w8527;
assign w8529 = w8408 & w8525;
assign w8530 = w8527 & ~w8529;
assign w8531 = (w9197 & w9290) | (w9197 & w9291) | (w9290 & w9291);
assign w8532 = (w7471 & w9212) | (w7471 & w9213) | (w9212 & w9213);
assign w8533 = ~w8531 & ~w8532;
assign w8534 = ~w8507 & ~w8519;
assign w8535 = ~w8500 & ~w8503;
assign w8536 = ~w8510 & w8514;
assign w8537 = pi31 & pi63;
assign w8538 = ~w8512 & w8537;
assign w8539 = w8422 & w8538;
assign w8540 = ~w8536 & ~w8539;
assign w8541 = ~w8535 & w8540;
assign w8542 = w8535 & ~w8540;
assign w8543 = ~w8541 & ~w8542;
assign w8544 = pi31 & pi62;
assign w8545 = pi30 & pi63;
assign w8546 = w8544 & ~w8545;
assign w8547 = ~w8544 & w8545;
assign w8548 = ~w8546 & ~w8547;
assign w8549 = w8543 & w8548;
assign w8550 = ~w8543 & ~w8548;
assign w8551 = ~w8549 & ~w8550;
assign w8552 = w8534 & ~w8551;
assign w8553 = ~w8534 & w8551;
assign w8554 = ~w8552 & ~w8553;
assign w8555 = w8522 & ~w8554;
assign w8556 = ~w8522 & w8554;
assign w8557 = ~w8555 & ~w8556;
assign w8558 = (~w7953 & w9091) | (~w7953 & w9092) | (w9091 & w9092);
assign w8559 = w8524 & w8554;
assign w8560 = (w9197 & w9292) | (w9197 & w9293) | (w9292 & w9293);
assign w8561 = ~w8558 & ~w8560;
assign w8562 = ~w8541 & ~w8549;
assign w8563 = ~w8536 & ~w8538;
assign w8564 = w8562 & w8563;
assign w8565 = ~w8562 & ~w8563;
assign w8566 = ~w8564 & ~w8565;
assign w8567 = ~w8552 & ~w8556;
assign w8568 = ~w8566 & ~w8567;
assign w8569 = w8566 & w8567;
assign w8570 = ~w8568 & ~w8569;
assign w8571 = (~w7953 & w9093) | (~w7953 & w9094) | (w9093 & w9094);
assign w8572 = (w7953 & w9095) | (w7953 & w9096) | (w9095 & w9096);
assign w8573 = ~w8571 & ~w8572;
assign w8574 = ~w8565 & ~w8567;
assign w8575 = (~w7953 & w9097) | (~w7953 & w9098) | (w9097 & w9098);
assign w8576 = ~w8564 & ~w8575;
assign w8577 = ~w1 & ~w9;
assign w8578 = w15 & ~w29;
assign w8579 = w35 & ~w56;
assign w8580 = ~w268 & ~w262;
assign w8581 = ~w275 & ~w274;
assign w8582 = w310 & ~w295;
assign w8583 = ~w349 & ~w382;
assign w8584 = ~w478 & ~w476;
assign w8585 = ~w448 & ~w446;
assign w8586 = (~w472 & ~w483) | (~w472 & w8662) | (~w483 & w8662);
assign w8587 = w440 & ~w558;
assign w8588 = w768 & ~w757;
assign w8589 = ~w1068 & ~w1067;
assign w8590 = ~w1410 & ~w1408;
assign w8591 = w1520 & ~w1509;
assign w8592 = ~w1543 & ~w1541;
assign w8593 = ~w1443 & ~w1564;
assign w8594 = w1443 & w1564;
assign w8595 = w1734 & ~w1723;
assign w8596 = ~w1715 & ~w1717;
assign w8597 = (~w1889 & w1723) | (~w1889 & w8663) | (w1723 & w8663);
assign w8598 = ~w1888 & w2026;
assign w8599 = ~w2029 & ~w2030;
assign w8600 = w1924 & ~w1913;
assign w8601 = w1862 & ~w1851;
assign w8602 = w2060 & ~w2049;
assign w8603 = w2087 & ~w2076;
assign w8604 = w2292 & ~w2281;
assign w8605 = w2250 & ~w2239;
assign w8606 = (~w2465 & w2281) | (~w2465 & w8664) | (w2281 & w8664);
assign w8607 = ~w2413 & ~w2412;
assign w8608 = w2758 & ~w2747;
assign w8609 = w2961 & ~w2950;
assign w8610 = w2985 & ~w2974;
assign w8611 = w3093 & ~w3082;
assign w8612 = w3065 & ~w3054;
assign w8613 = w3349 & ~w3338;
assign w8614 = w3373 & ~w3362;
assign w8615 = w3723 & ~w3712;
assign w8616 = w3691 & ~w3680;
assign w8617 = w3592 & ~w3581;
assign w8618 = w3616 & ~w3605;
assign w8619 = w3899 & ~w3888;
assign w8620 = w3780 & ~w3769;
assign w8621 = w4114 & ~w4103;
assign w8622 = w4034 & ~w4023;
assign w8623 = w4083 & ~w4072;
assign w8624 = w4059 & ~w4048;
assign w8625 = w4289 & ~w4278;
assign w8626 = w4548 & ~w4536;
assign w8627 = w4597 & ~w4585;
assign w8628 = w4573 & ~w4561;
assign w8629 = w4847 & ~w4836;
assign w8630 = w4797 & ~w4786;
assign w8631 = w4822 & ~w4811;
assign w8632 = w5125 & ~w5114;
assign w8633 = w5097 & ~w5086;
assign w8634 = w5329 & ~w5318;
assign w8635 = w5364 & ~w5353;
assign w8636 = w5621 & ~w5610;
assign w8637 = w5523 & ~w5512;
assign w8638 = w5548 & ~w5537;
assign w8639 = w5844 & ~w5833;
assign w8640 = w5816 & ~w5805;
assign w8641 = w5786 & ~w5775;
assign w8642 = w6031 & ~w6020;
assign w8643 = ~w6042 & ~w6040;
assign w8644 = ~w6000 & ~w5998;
assign w8645 = ~w5958 & ~w5956;
assign w8646 = w5947 & w6298;
assign w8647 = ~w5947 & ~w6298;
assign w8648 = (~w5944 & ~w5961) | (~w5944 & w9099) | (~w5961 & w9099);
assign w8649 = ~w6310 & ~w6320;
assign w8650 = ~w6175 & ~w6173;
assign w8651 = w6258 & ~w6247;
assign w8652 = ~w6227 & ~w6225;
assign w8653 = ~w6316 & ~w6314;
assign w8654 = ~w6307 & ~w6305;
assign w8655 = (~w6160 & ~w6178) | (~w6160 & w9100) | (~w6178 & w9100);
assign w8656 = ~w6869 & ~w6860;
assign w8657 = w7952 & w7460;
assign w8658 = (w7952 & ~w7474) | (w7952 & w8657) | (~w7474 & w8657);
assign w8659 = (~w8140 & w7949) | (~w8140 & w9101) | (w7949 & w9101);
assign w8660 = ~w8213 & w8140;
assign w8661 = ~w8213 & ~w8659;
assign w8662 = ~w344 & ~w472;
assign w8663 = w1888 & ~w1889;
assign w8664 = w2464 & ~w2465;
assign w8665 = w193 & ~w162;
assign w8666 = ~w190 & ~w178;
assign w8667 = ~w158 & ~w156;
assign w8668 = w252 & ~w242;
assign w8669 = ~w341 & ~w339;
assign w8670 = ~w359 & ~w361;
assign w8671 = ~w367 & w478;
assign w8672 = w367 & ~w478;
assign w8673 = w469 & ~w458;
assign w8674 = ~w450 & ~w452;
assign w8675 = w550 & w476;
assign w8676 = w550 & ~w8584;
assign w8677 = ~w594 & ~w589;
assign w8678 = w525 & ~w514;
assign w8679 = ~w506 & ~w508;
assign w8680 = w617 & ~w606;
assign w8681 = w722 & ~w711;
assign w8682 = ~w932 & ~w927;
assign w8683 = w843 & w984;
assign w8684 = ~w845 & w986;
assign w8685 = w888 & ~w876;
assign w8686 = ~w1038 & ~w1036;
assign w8687 = w969 & ~w957;
assign w8688 = w1017 & ~w1005;
assign w8689 = w1140 & ~w1129;
assign w8690 = (~w1067 & w1286) | (~w1067 & w9214) | (w1286 & w9214);
assign w8691 = ~w1287 & w8589;
assign w8692 = ~w1286 & w9215;
assign w8693 = w1287 & ~w8589;
assign w8694 = ~w1403 & ~w1401;
assign w8695 = ~w1419 & w1624;
assign w8696 = ~w1536 & ~w1534;
assign w8697 = ~w1548 & ~w1550;
assign w8698 = ~w1756 & ~w1754;
assign w8699 = ~w1694 & ~w1693;
assign w8700 = ~w1749 & ~w1747;
assign w8701 = ~w1765 & ~w1975;
assign w8702 = w1765 & w1975;
assign w8703 = ~w2026 & ~w1889;
assign w8704 = ~w2026 & w8597;
assign w8705 = ~w1877 & ~w1875;
assign w8706 = (w1883 & w1893) | (w1883 & w9216) | (w1893 & w9216);
assign w8707 = ~w2098 & ~w2097;
assign w8708 = ~w2108 & ~w2106;
assign w8709 = w2090 & ~w2112;
assign w8710 = ~w2330 & w2429;
assign w8711 = ~w2064 & ~w2328;
assign w8712 = ~w2261 & ~w2259;
assign w8713 = ~w2307 & ~w2305;
assign w8714 = ~w2511 & ~w2509;
assign w8715 = ~w2471 & ~w2465;
assign w8716 = ~w2471 & w8606;
assign w8717 = w2455 & ~w2444;
assign w8718 = w2713 & ~w2702;
assign w8719 = ~w2739 & ~w2741;
assign w8720 = w2685 & ~w2674;
assign w8721 = ~w3017 & ~w3030;
assign w8722 = ~w2826 & ~w2824;
assign w8723 = w2926 & ~w2925;
assign w8724 = ~w3026 & ~w3024;
assign w8725 = (~w3264 & w3036) | (~w3264 & w8782) | (w3036 & w8782);
assign w8726 = (~w3099 & ~w3137) | (~w3099 & w8867) | (~w3137 & w8867);
assign w8727 = (~w3386 & ~w3424) | (~w3386 & w8868) | (~w3424 & w8868);
assign w8728 = ~w3415 & ~w3413;
assign w8729 = ~w3405 & ~w3403;
assign w8730 = ~w3650 & ~w3648;
assign w8731 = (w3631 & ~w3669) | (w3631 & w8869) | (~w3669 & w8869);
assign w8732 = ~w3753 & w4009;
assign w8733 = w3829 & ~w3818;
assign w8734 = ~w3857 & ~w3855;
assign w8735 = ~w3846 & ~w3844;
assign w8736 = w3805 & ~w3794;
assign w8737 = ~w3868 & ~w3866;
assign w8738 = ~w3931 & ~w3929;
assign w8739 = (~w3838 & ~w3877) | (~w3838 & w8870) | (~w3877 & w8870);
assign w8740 = (w4092 & ~w4145) | (w4092 & w8871) | (~w4145 & w8871);
assign w8741 = w4366 & ~w4355;
assign w8742 = w4338 & ~w4327;
assign w8743 = ~w4439 & ~w4437;
assign w8744 = ~w4458 & ~w4456;
assign w8745 = (~w4344 & ~w4403) | (~w4344 & w8872) | (~w4403 & w8872);
assign w8746 = w4628 & ~w4616;
assign w8747 = ~w4708 & ~w4706;
assign w8748 = ~w4952 & ~w4950;
assign w8749 = ~w4875 & ~w4873;
assign w8750 = ~w4934 & ~w4932;
assign w8751 = (w5131 & w5195) | (w5131 & w9102) | (w5195 & w9102);
assign w8752 = (~w5373 & ~w5411) | (~w5373 & w9103) | (~w5411 & w9103);
assign w8753 = ~w5475 & w5696;
assign w8754 = w5475 & ~w5696;
assign w8755 = ~w5479 & ~w5469;
assign w8756 = w5484 & w5706;
assign w8757 = ~w5710 & ~w5495;
assign w8758 = (w5670 & w5687) | (w5670 & w9104) | (w5687 & w9104);
assign w8759 = ~w5590 & ~w5588;
assign w8760 = ~w5580 & ~w5578;
assign w8761 = ~w5658 & ~w5656;
assign w8762 = w5659 & ~w5662;
assign w8763 = (~w5561 & ~w5599) | (~w5561 & w9105) | (~w5599 & w9105);
assign w8764 = ~w5673 & ~w5897;
assign w8765 = w5673 & w5897;
assign w8766 = ~w5720 & w9106;
assign w8767 = (~w5909 & w5720) | (~w5909 & w9107) | (w5720 & w9107);
assign w8768 = (w5822 & w5885) | (w5822 & w9217) | (w5885 & w9217);
assign w8769 = ~w5855 & ~w5853;
assign w8770 = ~w6130 & w6125;
assign w8771 = w6009 & ~w6063;
assign w8772 = w5989 & ~w5978;
assign w8773 = w6236 & ~w6280;
assign w8774 = w6206 & ~w6195;
assign w8775 = w6440 & ~w6484;
assign w8776 = ~w6427 & ~w6425;
assign w8777 = w7604 & w7460;
assign w8778 = (w7604 & ~w7474) | (w7604 & w8777) | (~w7474 & w8777);
assign w8779 = ~w7600 & w7724;
assign w8780 = w8288 & ~w8660;
assign w8781 = w8288 & ~w8661;
assign w8782 = w3263 & ~w3264;
assign w8783 = w4004 & ~w4261;
assign w8784 = ~w4262 & w4261;
assign w8785 = ~w4262 & ~w8783;
assign w8786 = w4499 & ~w4510;
assign w8787 = w4475 & ~w4674;
assign w8788 = ~w4475 & w4674;
assign w8789 = ~w4487 & ~w4485;
assign w8790 = ~w4442 & ~w4445;
assign w8791 = (w4472 & w4490) | (w4472 & w8873) | (w4490 & w8873);
assign w8792 = ~w4752 & ~w4763;
assign w8793 = ~w4731 & ~w4729;
assign w8794 = ~w4305 & ~w4579;
assign w8795 = ~w4690 & ~w4688;
assign w8796 = ~w4700 & ~w4721;
assign w8797 = (w4606 & w4663) | (w4606 & w9108) | (w4663 & w9108);
assign w8798 = ~w4759 & ~w4757;
assign w8799 = ~w4684 & ~w4682;
assign w8800 = (w4726 & w4743) | (w4726 & w8874) | (w4743 & w8874);
assign w8801 = w5042 & ~w4932;
assign w8802 = w5042 & w8750;
assign w8803 = (~w4856 & ~w4884) | (~w4856 & w9109) | (~w4884 & w9109);
assign w8804 = ~w4944 & ~w4965;
assign w8805 = w5258 & w5257;
assign w8806 = (~w5251 & ~w5253) | (~w5251 & w8875) | (~w5253 & w8875);
assign w8807 = ~w5038 & ~w5036;
assign w8808 = ~w5186 & ~w5184;
assign w8809 = ~w5048 & ~w5046;
assign w8810 = w5023 & ~w5026;
assign w8811 = w5153 & ~w5142;
assign w8812 = ~w5284 & ~w5302;
assign w8813 = w5433 & ~w5422;
assign w8814 = ~w5344 & ~w5347;
assign w8815 = ~w5298 & ~w5296;
assign w8816 = ~w5402 & ~w5400;
assign w8817 = ~w5392 & ~w5390;
assign w8818 = ~w5649 & ~w5647;
assign w8819 = ~w5684 & ~w5682;
assign w8820 = ~w5866 & ~w5864;
assign w8821 = ~w5876 & ~w5874;
assign w8822 = ~w5738 & ~w5736;
assign w8823 = w5722 & ~w5725;
assign w8824 = ~w5858 & ~w5880;
assign w8825 = ~w5755 & ~w5753;
assign w8826 = ~w5906 & ~w5904;
assign w8827 = (~w5741 & ~w5758) | (~w5741 & w9110) | (~w5758 & w9110);
assign w8828 = ~w6053 & ~w6051;
assign w8829 = ~w5992 & ~w6004;
assign w8830 = ~w6045 & ~w6057;
assign w8831 = ~w6099 & ~w6097;
assign w8832 = (w6328 & w6128) | (w6328 & w8876) | (w6128 & w8876);
assign w8833 = (~w6209 & ~w6230) | (~w6209 & w9111) | (~w6230 & w9111);
assign w8834 = (~w6419 & ~w6430) | (~w6419 & w9112) | (~w6430 & w9112);
assign w8835 = w6462 & ~w6451;
assign w8836 = w6416 & ~w6405;
assign w8837 = w6432 & w6425;
assign w8838 = w6432 & ~w8776;
assign w8839 = ~w6432 & ~w6425;
assign w8840 = ~w6432 & w8776;
assign w8841 = ~w6368 & ~w6366;
assign w8842 = (~w6353 & ~w6371) | (~w6353 & w9113) | (~w6371 & w9113);
assign w8843 = (~w6672 & ~w6682) | (~w6672 & w9218) | (~w6682 & w9218);
assign w8844 = w6628 & ~w6617;
assign w8845 = w6584 & ~w6573;
assign w8846 = ~w6679 & ~w6677;
assign w8847 = ~w6669 & ~w6667;
assign w8848 = (~w6538 & ~w6556) | (~w6538 & w9114) | (~w6556 & w9114);
assign w8849 = (w6872 & w6128) | (w6872 & w9115) | (w6128 & w9115);
assign w8850 = ~w6658 & ~w6801;
assign w8851 = w6768 & ~w6757;
assign w8852 = ~w6728 & ~w6726;
assign w8853 = (~w6722 & ~w6740) | (~w6722 & w9116) | (~w6740 & w9116);
assign w8854 = ~w6870 & w7030;
assign w8855 = ~w7012 & ~w7022;
assign w8856 = w6973 & ~w6962;
assign w8857 = ~w7018 & ~w7016;
assign w8858 = ~w6899 & ~w6919;
assign w8859 = w7128 & ~w7117;
assign w8860 = ~w8779 & ~w7722;
assign w8861 = ~w8284 & ~w8780;
assign w8862 = ~w8284 & ~w8781;
assign w8863 = w8412 & ~w8780;
assign w8864 = w8412 & ~w8781;
assign w8865 = w8528 & ~w8780;
assign w8866 = w8528 & ~w8781;
assign w8867 = ~w3162 & ~w3099;
assign w8868 = ~w3449 & ~w3386;
assign w8869 = ~w3694 & w3631;
assign w8870 = ~w3902 & ~w3838;
assign w8871 = w4117 & w4092;
assign w8872 = ~w4369 & ~w4344;
assign w8873 = w4480 & w4472;
assign w8874 = w4734 & w4726;
assign w8875 = w5014 & ~w5251;
assign w8876 = ~w6131 & w6328;
assign w8877 = w5260 & w8784;
assign w8878 = w5260 & w8785;
assign w8879 = ~w6326 & ~w6328;
assign w8880 = ~w6326 & ~w8832;
assign w8881 = ~w6268 & ~w6266;
assign w8882 = w6144 & ~w6155;
assign w8883 = ~w6271 & ~w6274;
assign w8884 = w6082 & w6291;
assign w8885 = ~w6495 & ~w6505;
assign w8886 = w6512 & ~w6511;
assign w8887 = (~w6587 & ~w6598) | (~w6587 & w9117) | (~w6598 & w9117);
assign w8888 = ~w6595 & ~w6593;
assign w8889 = ~w6638 & ~w6636;
assign w8890 = ~w6553 & ~w6551;
assign w8891 = w6867 & w6869;
assign w8892 = ~w6779 & ~w6777;
assign w8893 = ~w6787 & ~w6785;
assign w8894 = ~w6797 & ~w6795;
assign w8895 = ~w6737 & ~w6735;
assign w8896 = ~w6841 & ~w6839;
assign w8897 = ~w7028 & ~w7030;
assign w8898 = (~w7028 & w6870) | (~w7028 & w8897) | (w6870 & w8897);
assign w8899 = ~w6983 & ~w6981;
assign w8900 = ~w6934 & ~w6946;
assign w8901 = ~w6942 & ~w6940;
assign w8902 = ~w7093 & ~w7091;
assign w8903 = ~w7138 & ~w7136;
assign w8904 = w7103 & ~w7097;
assign w8905 = ~w7236 & ~w7234;
assign w8906 = w7188 & ~w7101;
assign w8907 = ~w7464 & ~w7468;
assign w8908 = (~w7722 & w8860) | (~w7722 & w8777) | (w8860 & w8777);
assign w8909 = (~w7722 & w8860) | (~w7722 & w8778) | (w8860 & w8778);
assign w8910 = ~w7949 & ~w8657;
assign w8911 = (w7474 & w9219) | (w7474 & w8910) | (w9219 & w8910);
assign w8912 = w8350 & ~w8861;
assign w8913 = w8350 & ~w8862;
assign w8914 = ~w8411 & ~w8863;
assign w8915 = ~w8411 & ~w8864;
assign w8916 = ~w8530 & ~w8865;
assign w8917 = ~w8530 & ~w8866;
assign w8918 = w2906 & ~w2895;
assign w8919 = ~w2966 & ~w2968;
assign w8920 = ~w3216 & ~w2925;
assign w8921 = ~w3216 & w8723;
assign w8922 = w3293 & w3126;
assign w8923 = (w3293 & w3128) | (w3293 & w8922) | (w3128 & w8922);
assign w8924 = ~w3293 & ~w3126;
assign w8925 = ~w3128 & w8924;
assign w8926 = w3159 & ~w3148;
assign w8927 = ~w3046 & ~w3048;
assign w8928 = w3446 & ~w3435;
assign w8929 = ~w3354 & ~w3356;
assign w8930 = ~w3318 & ~w3316;
assign w8931 = ~w3536 & ~w3534;
assign w8932 = ~w3597 & ~w3599;
assign w8933 = w3940 & w3658;
assign w8934 = (w3940 & w3660) | (w3940 & w8933) | (w3660 & w8933);
assign w8935 = ~w3940 & ~w3658;
assign w8936 = ~w3660 & w8935;
assign w8937 = ~w3555 & ~w3553;
assign w8938 = w3556 & ~w3559;
assign w8939 = ~w3735 & ~w3733;
assign w8940 = (~w3567 & ~w3539) | (~w3567 & w9118) | (~w3539 & w9118);
assign w8941 = ~w3973 & ~w3972;
assign w8942 = ~w3946 & ~w3944;
assign w8943 = ~w3947 & ~w3950;
assign w8944 = ~w3924 & ~w3922;
assign w8945 = (w3957 & ~w3976) | (w3957 & w9119) | (~w3976 & w9119);
assign w8946 = ~w4232 & ~w4230;
assign w8947 = ~w4064 & ~w4066;
assign w8948 = ~w4187 & ~w4190;
assign w8949 = w4487 & w8740;
assign w8950 = w4487 & ~w4146;
assign w8951 = ~w4487 & ~w8740;
assign w8952 = ~w4487 & w4146;
assign w8953 = ~w4177 & ~w4175;
assign w8954 = (w4217 & w4235) | (w4217 & w9120) | (w4235 & w9120);
assign w8955 = w4519 & w8784;
assign w8956 = ~w8783 & w9121;
assign w8957 = ~w4477 & w8788;
assign w8958 = ~w4377 & ~w4375;
assign w8959 = w5000 & ~w8800;
assign w8960 = w5000 & w4745;
assign w8961 = (~w4997 & ~w5006) | (~w4997 & w9122) | (~w5006 & w9122);
assign w8962 = ~w5003 & ~w5001;
assign w8963 = ~w4976 & ~w4974;
assign w8964 = w5263 & ~w8878;
assign w8965 = w5263 & ~w8877;
assign w8966 = w5162 & ~w5269;
assign w8967 = ~w5162 & w5269;
assign w8968 = ~w5167 & ~w5190;
assign w8969 = ~w5077 & ~w5080;
assign w8970 = ~w5064 & ~w5455;
assign w8971 = w5064 & w5455;
assign w8972 = w5242 & w5467;
assign w8973 = ~w5242 & ~w5467;
assign w8974 = ~w5051 & ~w5070;
assign w8975 = w5287 & ~w5640;
assign w8976 = ~w5287 & w5640;
assign w8977 = ~w5381 & ~w5379;
assign w8978 = ~w5272 & ~w5270;
assign w8979 = w5273 & ~w5276;
assign w8980 = ~w5384 & ~w5406;
assign w8981 = w8756 & w5706;
assign w8982 = (w5706 & w8756) | (w5706 & w5486) | (w8756 & w5486);
assign w8983 = ~w5572 & ~w5594;
assign w8984 = w5499 & ~w5698;
assign w8985 = ~w5744 & ~w6090;
assign w8986 = w5744 & w6090;
assign w8987 = ~w6102 & ~w6113;
assign w8988 = ~w5969 & ~w5972;
assign w8989 = w6347 & ~w6266;
assign w8990 = w6347 & w8881;
assign w8991 = ~w6472 & ~w6470;
assign w8992 = ~w6475 & ~w6478;
assign w8993 = ~w6396 & ~w6399;
assign w8994 = (~w6511 & w8886) | (~w6511 & ~w8879) | (w8886 & ~w8879);
assign w8995 = (w8832 & w9123) | (w8832 & w9124) | (w9123 & w9124);
assign w8996 = ~w6564 & ~w6567;
assign w8997 = ~w6844 & ~w6854;
assign w8998 = ~w6748 & ~w6751;
assign w8999 = w6977 & ~w6795;
assign w9000 = w6977 & w8894;
assign w9001 = (w8897 & w8898) | (w8897 & ~w6872) | (w8898 & ~w6872);
assign w9002 = (w8897 & w8898) | (w8897 & ~w8849) | (w8898 & ~w8849);
assign w9003 = ~w6953 & ~w6956;
assign w9004 = w7132 & ~w6940;
assign w9005 = w7132 & w8901;
assign w9006 = w6913 & w7154;
assign w9007 = ~w6913 & ~w7154;
assign w9008 = ~w7163 & ~w7174;
assign w9009 = w7230 & ~w7091;
assign w9010 = w7230 & w8902;
assign w9011 = w7063 & w7248;
assign w9012 = ~w7063 & ~w7248;
assign w9013 = ~w7170 & ~w7168;
assign w9014 = ~w7160 & ~w7158;
assign w9015 = ~w7060 & ~w7080;
assign w9016 = w7226 & ~w7215;
assign w9017 = w7282 & w7386;
assign w9018 = ~w7282 & ~w7386;
assign w9019 = w7231 & ~w7101;
assign w9020 = w7231 & w8906;
assign w9021 = ~w7254 & ~w7252;
assign w9022 = ~w7279 & ~w7299;
assign w9023 = ~w7431 & ~w7429;
assign w9024 = ~w7392 & ~w7390;
assign w9025 = ~w7416 & ~w7435;
assign w9026 = ~w7837 & ~w7835;
assign w9027 = ~w8046 & ~w8044;
assign w9028 = ~w8213 & ~w9077;
assign w9029 = (w7474 & w9220) | (w7474 & w9028) | (w9220 & w9028);
assign w9030 = (w8861 & w8862) | (w8861 & ~w8657) | (w8862 & ~w8657);
assign w9031 = (w7474 & w9221) | (w7474 & w9030) | (w9221 & w9030);
assign w9032 = ~w8348 & ~w8912;
assign w9033 = ~w8348 & ~w8913;
assign w9034 = w8453 & w8914;
assign w9035 = w8453 & w8915;
assign w9036 = w8524 & w8916;
assign w9037 = w8524 & w8917;
assign w9038 = w8559 & w8916;
assign w9039 = w8559 & w8917;
assign w9040 = ~w4517 & ~w8955;
assign w9041 = (~w4517 & ~w9121) | (~w4517 & w9222) | (~w9121 & w9222);
assign w9042 = ~w4740 & ~w4738;
assign w9043 = ~w4643 & ~w4641;
assign w9044 = ~w4693 & ~w4695;
assign w9045 = w4712 & ~w4715;
assign w9046 = ~w4677 & ~w4675;
assign w9047 = w4770 & ~w4769;
assign w9048 = ~w4985 & ~w4983;
assign w9049 = ~w5223 & ~w4974;
assign w9050 = ~w5223 & w8963;
assign w9051 = ~w4970 & ~w4990;
assign w9052 = ~w5057 & ~w5055;
assign w9053 = ~w5066 & w8970;
assign w9054 = ~w5492 & ~w5462;
assign w9055 = ~w5705 & ~w8982;
assign w9056 = ~w5705 & ~w8981;
assign w9057 = ~w6691 & ~w6689;
assign w9058 = w7181 & ~w7180;
assign w9059 = ~w7195 & ~w7193;
assign w9060 = ~w7443 & ~w7454;
assign w9061 = ~w7344 & ~w7342;
assign w9062 = ~w7352 & ~w7350;
assign w9063 = w7474 & ~w7460;
assign w9064 = (~w7460 & w9063) | (~w7460 & w7470) | (w9063 & w7470);
assign w9065 = ~w7600 & ~w8777;
assign w9066 = (w7474 & w9223) | (w7474 & w9065) | (w9223 & w9065);
assign w9067 = ~w7583 & ~w7594;
assign w9068 = ~w7528 & ~w7578;
assign w9069 = ~w7705 & ~w7716;
assign w9070 = ~w7941 & ~w7835;
assign w9071 = ~w7941 & w9026;
assign w9072 = w7941 & w7835;
assign w9073 = w7941 & ~w9026;
assign w9074 = ~w7948 & ~w7940;
assign w9075 = w8133 & w8044;
assign w9076 = w8133 & ~w9027;
assign w9077 = (~w8140 & w8659) | (~w8140 & w8657) | (w8659 & w8657);
assign w9078 = (~w8140 & w8659) | (~w8140 & w8658) | (w8659 & w8658);
assign w9079 = w8214 & ~w8286;
assign w9080 = w8404 & w9032;
assign w9081 = w8404 & w9033;
assign w9082 = ~w8404 & ~w9032;
assign w9083 = ~w8404 & ~w9033;
assign w9084 = (w8914 & w8915) | (w8914 & w8657) | (w8915 & w8657);
assign w9085 = ~w8408 & w8455;
assign w9086 = ~w8491 & w9034;
assign w9087 = ~w8491 & w9035;
assign w9088 = w8495 & ~w9034;
assign w9089 = w8495 & ~w9035;
assign w9090 = (w8916 & w8917) | (w8916 & w8657) | (w8917 & w8657);
assign w9091 = w8557 & ~w9036;
assign w9092 = w8557 & ~w9037;
assign w9093 = ~w8570 & ~w9038;
assign w9094 = ~w8570 & ~w9039;
assign w9095 = w8566 & w9038;
assign w9096 = w8566 & w9039;
assign w9097 = w8574 & ~w9038;
assign w9098 = w8574 & ~w9039;
assign w9099 = ~w5952 & ~w5944;
assign w9100 = ~w6169 & ~w6160;
assign w9101 = ~w8138 & ~w8140;
assign w9102 = w5156 & w5131;
assign w9103 = ~w5436 & ~w5373;
assign w9104 = w5678 & w5670;
assign w9105 = ~w5624 & ~w5561;
assign w9106 = w5711 & w5909;
assign w9107 = ~w5711 & ~w5909;
assign w9108 = w4631 & w4606;
assign w9109 = ~w4909 & ~w4856;
assign w9110 = ~w5749 & ~w5741;
assign w9111 = ~w6219 & ~w6209;
assign w9112 = w6434 & ~w6419;
assign w9113 = ~w6362 & ~w6353;
assign w9114 = ~w6547 & ~w6538;
assign w9115 = ~w6131 & w6872;
assign w9116 = ~w6731 & ~w6722;
assign w9117 = w6600 & ~w6587;
assign w9118 = ~w3530 & ~w3567;
assign w9119 = w3967 & w3957;
assign w9120 = w4226 & w4217;
assign w9121 = ~w4262 & w4519;
assign w9122 = w4998 & ~w4997;
assign w9123 = w8886 | ~w6511;
assign w9124 = (~w6511 & w8886) | (~w6511 & w6326) | (w8886 & w6326);
assign w9125 = w2501 & ~w2490;
assign w9126 = ~w2996 & ~w2994;
assign w9127 = ~w2917 & ~w2915;
assign w9128 = ~w3107 & ~w3105;
assign w9129 = ~w3118 & ~w3116;
assign w9130 = ~w3214 & ~w3212;
assign w9131 = w3215 & ~w3217;
assign w9132 = ~w3110 & ~w3132;
assign w9133 = w3318 & ~w8726;
assign w9134 = w3318 & w3163;
assign w9135 = ~w3291 & ~w3289;
assign w9136 = w3292 & ~w3294;
assign w9137 = ~w3397 & ~w3419;
assign w9138 = w3536 & ~w8727;
assign w9139 = w3536 & w3450;
assign w9140 = ~w3394 & ~w3392;
assign w9141 = ~w3639 & ~w3637;
assign w9142 = ~w3642 & ~w3664;
assign w9143 = ~w3973 & ~w8731;
assign w9144 = ~w3973 & w3695;
assign w9145 = w3962 & w4167;
assign w9146 = ~w3962 & ~w4167;
assign w9147 = ~w3849 & ~w3872;
assign w9148 = w4232 & ~w8739;
assign w9149 = w4232 & w3903;
assign w9150 = ~w3992 & ~w3990;
assign w9151 = w4221 & w4422;
assign w9152 = ~w4221 & ~w4422;
assign w9153 = ~w4136 & ~w4134;
assign w9154 = ~w4125 & ~w4123;
assign w9155 = ~w4203 & ~w4201;
assign w9156 = ~w4184 & ~w4182;
assign w9157 = ~w4037 & ~w4087;
assign w9158 = ~w4251 & ~w4249;
assign w9159 = ~w4244 & ~w4255;
assign w9160 = ~w4505 & ~w4503;
assign w9161 = (~w4769 & w9047) | (~w4769 & ~w9040) | (w9047 & ~w9040);
assign w9162 = (~w4769 & w9047) | (~w4769 & ~w9041) | (w9047 & ~w9041);
assign w9163 = ~w4927 & ~w4925;
assign w9164 = w5684 & ~w8752;
assign w9165 = w5684 & w5437;
assign w9166 = w5755 & ~w8763;
assign w9167 = w5755 & w5625;
assign w9168 = w5916 & ~w9056;
assign w9169 = w5916 & ~w9055;
assign w9170 = ~w5717 & ~w5715;
assign w9171 = ~w6109 & ~w6107;
assign w9172 = w6313 & ~w8648;
assign w9173 = w6313 & w5962;
assign w9174 = ~w6498 & ~w8655;
assign w9175 = ~w6498 & w6179;
assign w9176 = ~w6501 & ~w6499;
assign w9177 = (~w6689 & w9057) | (~w6689 & ~w8994) | (w9057 & ~w8994);
assign w9178 = (~w8832 & w9224) | (~w8832 & w9225) | (w9224 & w9225);
assign w9179 = w6847 & ~w8848;
assign w9180 = w6847 & w6557;
assign w9181 = w8849 & w6872;
assign w9182 = (w6872 & w8849) | (w6872 & w6136) | (w8849 & w6136);
assign w9183 = ~w6850 & ~w6848;
assign w9184 = w7015 & ~w8853;
assign w9185 = w7015 & w6741;
assign w9186 = (w8849 & w9226) | (w8849 & w9227) | (w9226 & w9227);
assign w9187 = (~w7180 & w9058) | (~w7180 & ~w9001) | (w9058 & ~w9001);
assign w9188 = ~w7470 & ~w7474;
assign w9189 = w7461 & ~w7602;
assign w9190 = (w8777 & ~w7474) | (w8777 & w9228) | (~w7474 & w9228);
assign w9191 = (w8777 & w8778) | (w8777 & ~w7470) | (w8778 & ~w7470);
assign w9192 = ~w7837 & ~w8908;
assign w9193 = ~w7837 & ~w8909;
assign w9194 = ~w7941 & w9318;
assign w9195 = (w9070 & w9071) | (w9070 & ~w8909) | (w9071 & ~w8909);
assign w9196 = (w8657 & ~w7474) | (w8657 & w9229) | (~w7474 & w9229);
assign w9197 = (w8657 & w8658) | (w8657 & ~w7470) | (w8658 & ~w7470);
assign w9198 = ~w8046 & w8910;
assign w9199 = ~w8046 & w8911;
assign w9200 = ~w8133 & w9319;
assign w9201 = ~w8133 & w9320;
assign w9202 = w8215 & ~w9077;
assign w9203 = w8215 & ~w9078;
assign w9204 = (~w8286 & w9079) | (~w8286 & w9028) | (w9079 & w9028);
assign w9205 = (~w8286 & w9079) | (~w8286 & w9029) | (w9079 & w9029);
assign w9206 = ~w8350 & w9030;
assign w9207 = ~w8350 & w9031;
assign w9208 = (w8658 & w9230) | (w8658 & w9231) | (w9230 & w9231);
assign w9209 = ~w8453 & w9084;
assign w9210 = (w8455 & w9085) | (w8455 & w9030) | (w9085 & w9030);
assign w9211 = (w8455 & w9085) | (w8455 & w9031) | (w9085 & w9031);
assign w9212 = (~w8658 & w9232) | (~w8658 & w9233) | (w9232 & w9233);
assign w9213 = ~w8524 & ~w9090;
assign w9214 = w1072 & ~w1067;
assign w9215 = ~w1072 & w1067;
assign w9216 = w1762 & w1883;
assign w9217 = w5847 & w5822;
assign w9218 = w6673 & ~w6672;
assign w9219 = ~w7949 & ~w7952;
assign w9220 = ~w8213 & w9321;
assign w9221 = (w8861 & w8862) | (w8861 & ~w7952) | (w8862 & ~w7952);
assign w9222 = w8783 & ~w4517;
assign w9223 = ~w7600 & ~w7604;
assign w9224 = (~w6689 & w9057) | (~w6689 & ~w9124) | (w9057 & ~w9124);
assign w9225 = (~w6689 & w9057) | (~w6689 & ~w9123) | (w9057 & ~w9123);
assign w9226 = (~w7180 & w9058) | (~w7180 & ~w8897) | (w9058 & ~w8897);
assign w9227 = (~w7180 & w9058) | (~w7180 & ~w8898) | (w9058 & ~w8898);
assign w9228 = w8777 | w7604;
assign w9229 = w8657 | w7952;
assign w9230 = ~w8453 & w8914;
assign w9231 = ~w8453 & w8915;
assign w9232 = ~w8524 & ~w8916;
assign w9233 = ~w8524 & ~w8917;
assign w9234 = w631 & ~w630;
assign w9235 = ~w654 & ~w653;
assign w9236 = ~w749 & ~w751;
assign w9237 = ~w744 & ~w742;
assign w9238 = ~w905 & ~w903;
assign w9239 = ~w838 & ~w860;
assign w9240 = ~w856 & ~w854;
assign w9241 = ~w1028 & ~w1026;
assign w9242 = w1020 & ~w1045;
assign w9243 = ~w1161 & ~w1159;
assign w9244 = ~w1182 & ~w1180;
assign w9245 = w1143 & ~w1166;
assign w9246 = w1174 & ~w1186;
assign w9247 = ~w1233 & ~w1231;
assign w9248 = w1223 & ~w1211;
assign w9249 = ~w1312 & ~w1301;
assign w9250 = ~w1331 & ~w1330;
assign w9251 = w1416 & ~w1623;
assign w9252 = w1623 & ~w1417;
assign w9253 = ~w1501 & ~w1503;
assign w9254 = ~w1871 & ~w1754;
assign w9255 = ~w1871 & w8698;
assign w9256 = w1781 & w1930;
assign w9257 = ~w1781 & ~w1930;
assign w9258 = ~w1825 & ~w1823;
assign w9259 = ~w1990 & ~w2002;
assign w9260 = ~w1936 & ~w1934;
assign w9261 = w1961 & ~w1983;
assign w9262 = ~w1996 & ~w1994;
assign w9263 = w1976 & w2129;
assign w9264 = ~w1976 & ~w2129;
assign w9265 = w2137 & ~w8706;
assign w9266 = w2137 & w1895;
assign w9267 = ~w2008 & ~w1836;
assign w9268 = ~w2202 & w2403;
assign w9269 = w3752 & w2405;
assign w9270 = w8783 & ~w4261;
assign w9271 = (~w4261 & w8783) | (~w4261 & ~w3754) | (w8783 & ~w3754);
assign w9272 = w5015 & w9162;
assign w9273 = w5015 & w9161;
assign w9274 = ~w5298 & ~w8751;
assign w9275 = ~w5298 & w5196;
assign w9276 = ~w5486 & ~w5484;
assign w9277 = ~w5494 & ~w5497;
assign w9278 = ~w5914 & ~w9169;
assign w9279 = ~w5914 & ~w9168;
assign w9280 = ~w5958 & ~w8768;
assign w9281 = ~w5958 & w5886;
assign w9282 = w6870 & ~w7030;
assign w9283 = ~w7462 & w6137;
assign w9284 = (~w7602 & w9189) | (~w7602 & ~w6137) | (w9189 & ~w6137);
assign w9285 = (~w7602 & w9189) | (~w7602 & w9063) | (w9189 & w9063);
assign w9286 = w8288 & w9322;
assign w9287 = w8288 & w9323;
assign w9288 = w8350 & w9324;
assign w9289 = w8350 & w9325;
assign w9290 = (w9036 & w9037) | (w9036 & w6137) | (w9037 & w6137);
assign w9291 = (w9036 & w9037) | (w9036 & w9196) | (w9037 & w9196);
assign w9292 = (w9038 & w9039) | (w9038 & w6137) | (w9039 & w6137);
assign w9293 = (w9038 & w9039) | (w9038 & w9196) | (w9039 & w9196);
assign w9294 = (~w476 & w8584) | (~w476 & ~w480) | (w8584 & ~w480);
assign w9295 = (w1754 & ~w8698) | (w1754 & ~w1750) | (~w8698 & ~w1750);
assign w9296 = (w8706 & ~w1895) | (w8706 & ~w1896) | (~w1895 & ~w1896);
assign w9297 = (w2925 & ~w8723) | (w2925 & ~w2921) | (~w8723 & ~w2921);
assign w9298 = (w4261 & ~w8783) | (w4261 & ~w4010) | (~w8783 & ~w4010);
assign w9299 = (w8800 & ~w4745) | (w8800 & ~w4746) | (~w4745 & ~w4746);
assign w9300 = (w4932 & ~w8750) | (w4932 & ~w4928) | (~w8750 & ~w4928);
assign w9301 = (w4974 & ~w8963) | (w4974 & ~w4971) | (~w8963 & ~w4971);
assign w9302 = (~w6125 & ~w6129) | (~w6125 & ~w8770) | (~w6129 & ~w8770);
assign w9303 = (w8648 & ~w5962) | (w8648 & ~w5964) | (~w5962 & ~w5964);
assign w9304 = (w6266 & ~w8881) | (w6266 & ~w6262) | (~w8881 & ~w6262);
assign w9305 = (w8655 & ~w6179) | (w8655 & ~w6181) | (~w6179 & ~w6181);
assign w9306 = (w8848 & ~w6557) | (w8848 & ~w6559) | (~w6557 & ~w6559);
assign w9307 = (w6795 & ~w8894) | (w6795 & ~w6791) | (~w8894 & ~w6791);
assign w9308 = (w8853 & ~w6741) | (w8853 & ~w6743) | (~w6741 & ~w6743);
assign w9309 = (w6940 & ~w8901) | (w6940 & ~w6936) | (~w8901 & ~w6936);
assign w9310 = (w7091 & ~w8902) | (w7091 & ~w7087) | (~w8902 & ~w7087);
assign w9311 = (w7101 & ~w8906) | (w7101 & ~w7201) | (~w8906 & ~w7201);
assign w9312 = (~w7470 & ~w7462) | (~w7470 & w9283) | (~w7462 & w9283);
assign w9313 = (w7474 & ~w6137) | (w7474 & ~w9188) | (~w6137 & ~w9188);
assign w9314 = (~w9065 & ~w9066) | (~w9065 & ~w7471) | (~w9066 & ~w7471);
assign w9315 = (w8908 & w8909) | (w8908 & ~w7471) | (w8909 & ~w7471);
assign w9316 = (~w8910 & ~w8911) | (~w8910 & ~w7471) | (~w8911 & ~w7471);
assign w9317 = (w9077 & w9078) | (w9077 & ~w7471) | (w9078 & ~w7471);
assign w9318 = (~w7835 & w9026) | (~w7835 & ~w8908) | (w9026 & ~w8908);
assign w9319 = (~w8044 & w9027) | (~w8044 & w8910) | (w9027 & w8910);
assign w9320 = (~w8044 & w9027) | (~w8044 & w8911) | (w9027 & w8911);
assign w9321 = (w8140 & ~w8659) | (w8140 & ~w7952) | (~w8659 & ~w7952);
assign w9322 = (~w8660 & ~w8661) | (~w8660 & w6137) | (~w8661 & w6137);
assign w9323 = (~w8660 & ~w8661) | (~w8660 & w9196) | (~w8661 & w9196);
assign w9324 = (~w8861 & ~w8862) | (~w8861 & w6137) | (~w8862 & w6137);
assign w9325 = (~w8861 & ~w8862) | (~w8861 & w9196) | (~w8862 & w9196);
assign one = 1;
assign po00 = w3;// level 3
assign po01 = w14;// level 7
assign po02 = w34;// level 9
assign po03 = w61;// level 11
assign po04 = w97;// level 13
assign po05 = ~w150;// level 16
assign po06 = ~w205;// level 17
assign po07 = w267;// level 19
assign po08 = w337;// level 19
assign po09 = ~w412;// level 21
assign po10 = w501;// level 22
assign po11 = ~w593;// level 24
assign po12 = ~w698;// level 25
assign po13 = w812;// level 27
assign po14 = w931;// level 28
assign po15 = ~w1061;// level 28
assign po16 = w1200;// level 30
assign po17 = ~w1344;// level 32
assign po18 = w1498;// level 34
assign po19 = w1661;// level 36
assign po20 = w1840;// level 31
assign po21 = ~w2014;// level 33
assign po22 = w2206;// level 35
assign po23 = ~w2402;// level 34
assign po24 = w2608;// level 34
assign po25 = w2819;// level 36
assign po26 = w3042;// level 38
assign po27 = ~w3268;// level 40
assign po28 = w3509;// level 37
assign po29 = w3751;// level 39
assign po30 = w4008;// level 38
assign po31 = ~w4267;// level 39
assign po32 = w4524;// level 40
assign po33 = w4774;// level 39
assign po34 = w5019;// level 40
assign po35 = w5256;// level 41
assign po36 = w5489;// level 40
assign po37 = w5709;// level 41
assign po38 = w5920;// level 41
assign po39 = w6124;// level 41
assign po40 = w6331;// level 40
assign po41 = w6516;// level 41
assign po42 = w6695;// level 41
assign po43 = w6865;// level 41
assign po44 = w7033;// level 41
assign po45 = ~w7185;// level 41
assign po46 = ~w7330;// level 41
assign po47 = ~w7477;// level 41
assign po48 = w7606;// level 40
assign po49 = ~w7727;// level 41
assign po50 = w7840;// level 41
assign po51 = w7944;// level 41
assign po52 = w8049;// level 41
assign po53 = w8136;// level 41
assign po54 = ~w8218;// level 41
assign po55 = w8290;// level 41
assign po56 = w8353;// level 41
assign po57 = ~w8407;// level 41
assign po58 = ~w8457;// level 41
assign po59 = ~w8497;// level 41
assign po60 = w8533;// level 41
assign po61 = w8561;// level 41
assign po62 = w8573;// level 41
assign po63 = ~w8576;// level 41
assign po64 = ~w8576;// level 41
endmodule
