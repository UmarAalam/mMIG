// Benchmark "usb_funct" written by ABC on Wed Apr 29 13:54:56 2015

module usb_funct ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457,
    pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466,
    pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475,
    pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484,
    pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493,
    pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502,
    pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511,
    pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520,
    pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529,
    pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538,
    pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547,
    pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556,
    pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565,
    pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574,
    pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583,
    pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592,
    pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601,
    pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610,
    pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619,
    pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628,
    pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637,
    pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646,
    pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655,
    pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664,
    pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673,
    pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682,
    pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691,
    pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700,
    pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709,
    pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718,
    pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727,
    pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736,
    pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745,
    pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754,
    pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763,
    pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772,
    pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781,
    pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790,
    pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799,
    pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808,
    pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817,
    pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826,
    pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835,
    pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844,
    pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853,
    pi1854, pi1855, pi1856, pi1857, pi1858, pi1859,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511,
    po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520,
    po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529,
    po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538,
    po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547,
    po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556,
    po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565,
    po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574,
    po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583,
    po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592,
    po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601,
    po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610,
    po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619,
    po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628,
    po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637,
    po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646,
    po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655,
    po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664,
    po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673,
    po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682,
    po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691,
    po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700,
    po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709,
    po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718,
    po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727,
    po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736,
    po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745,
    po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754,
    po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763,
    po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772,
    po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781,
    po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790,
    po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799,
    po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808,
    po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817,
    po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826,
    po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835,
    po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844,
    po1845  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456,
    pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465,
    pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474,
    pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483,
    pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492,
    pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501,
    pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510,
    pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519,
    pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528,
    pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537,
    pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546,
    pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555,
    pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564,
    pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573,
    pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582,
    pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591,
    pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600,
    pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609,
    pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618,
    pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627,
    pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636,
    pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645,
    pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654,
    pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663,
    pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672,
    pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681,
    pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690,
    pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699,
    pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708,
    pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717,
    pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726,
    pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735,
    pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744,
    pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753,
    pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762,
    pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771,
    pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780,
    pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789,
    pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798,
    pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807,
    pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816,
    pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825,
    pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834,
    pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843,
    pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852,
    pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519,
    po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528,
    po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537,
    po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546,
    po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555,
    po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564,
    po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573,
    po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582,
    po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591,
    po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600,
    po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609,
    po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618,
    po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627,
    po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636,
    po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645,
    po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654,
    po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663,
    po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672,
    po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681,
    po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690,
    po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699,
    po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708,
    po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717,
    po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726,
    po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735,
    po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744,
    po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753,
    po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762,
    po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771,
    po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780,
    po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789,
    po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798,
    po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807,
    po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816,
    po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825,
    po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834,
    po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843,
    po1844, po1845;
  wire n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
    n3728, n3729, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3758, n3759,
    n3761, n3762, n3764, n3765, n3767, n3768, n3770, n3771, n3773, n3774,
    n3776, n3777, n3779, n3780, n3782, n3783, n3785, n3786, n3788, n3789,
    n3791, n3792, n3794, n3795, n3797, n3798, n3800, n3801, n3803, n3804,
    n3806, n3807, n3809, n3810, n3812, n3813, n3815, n3816, n3818, n3819,
    n3821, n3822, n3824, n3825, n3827, n3828, n3830, n3831, n3833, n3834,
    n3836, n3837, n3839, n3840, n3842, n3843, n3845, n3846, n3848, n3849,
    n3851, n3852, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3866, n3867, n3869, n3870, n3872, n3873, n3875,
    n3876, n3878, n3879, n3881, n3882, n3884, n3885, n3887, n3888, n3890,
    n3891, n3893, n3894, n3896, n3897, n3899, n3900, n3902, n3903, n3905,
    n3906, n3908, n3909, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4114, n4115, n4117, n4118, n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4161, n4162, n4163, n4164, n4165, n4166,
    n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4332, n4333, n4334, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
    n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
    n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4536, n4537, n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4663, n4664, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
    n4673, n4674, n4675, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4686, n4687, n4688, n4689, n4690, n4691, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
    n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
    n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
    n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4787, n4788,
    n4789, n4790, n4791, n4792, n4794, n4795, n4796, n4797, n4798, n4799,
    n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4813, n4814, n4815, n4816, n4817, n4818, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
    n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5006, n5007, n5008, n5010, n5011, n5012, n5014, n5015,
    n5016, n5018, n5019, n5020, n5022, n5023, n5024, n5026, n5027, n5028,
    n5030, n5031, n5032, n5034, n5035, n5036, n5038, n5039, n5040, n5042,
    n5043, n5044, n5046, n5047, n5048, n5050, n5051, n5052, n5054, n5055,
    n5056, n5058, n5059, n5060, n5062, n5063, n5064, n5065, n5066, n5067,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5077, n5078, n5079,
    n5080, n5082, n5083, n5084, n5085, n5086, n5087, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5101, n5102,
    n5103, n5104, n5105, n5106, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5118, n5119, n5120, n5121, n5122, n5123, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5145, n5146, n5147,
    n5148, n5149, n5150, n5151, n5152, n5153, n5155, n5156, n5157, n5158,
    n5159, n5160, n5161, n5162, n5163, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
    n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5202,
    n5203, n5204, n5205, n5206, n5207, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5221, n5222, n5224, n5225, n5226,
    n5227, n5229, n5231, n5232, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
    n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
    n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
    n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
    n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
    n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
    n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5453,
    n5454, n5455, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
    n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
    n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
    n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
    n5609, n5610, n5611, n5612, n5613, n5614, n5616, n5617, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
    n5643, n5644, n5646, n5647, n5648, n5649, n5650, n5651, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
    n5666, n5667, n5668, n5669, n5672, n5673, n5674, n5675, n5676, n5677,
    n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5699,
    n5700, n5702, n5703, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5714, n5715, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5726, n5727, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
    n5736, n5738, n5739, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
    n5748, n5749, n5751, n5752, n5754, n5755, n5756, n5757, n5758, n5759,
    n5760, n5761, n5762, n5764, n5765, n5767, n5768, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5777, n5778, n5780, n5781, n5782, n5783,
    n5784, n5785, n5786, n5787, n5788, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
    n5816, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
    n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882, n5884, n5885, n5886, n5887,
    n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
    n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
    n6044, n6045, n6046, n6047, n6048, n6049, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6083, n6085, n6086, n6087,
    n6089, n6090, n6092, n6093, n6095, n6096, n6098, n6099, n6100, n6102,
    n6103, n6104, n6106, n6107, n6108, n6110, n6111, n6112, n6114, n6115,
    n6116, n6118, n6119, n6120, n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6144, n6145, n6146, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6157, n6158, n6159, n6160, n6161,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6183,
    n6184, n6185, n6187, n6188, n6189, n6191, n6192, n6193, n6195, n6196,
    n6197, n6199, n6200, n6201, n6203, n6204, n6205, n6207, n6208, n6209,
    n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6228, n6230, n6231, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6263, n6264, n6265,
    n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
    n6287, n6288, n6289, n6290, n6291, n6293, n6294, n6296, n6297, n6298,
    n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6309,
    n6311, n6313, n6314, n6316, n6317, n6319, n6320, n6322, n6323, n6325,
    n6326, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6414, n6415, n6416, n6417, n6418,
    n6420, n6421, n6422, n6424, n6425, n6427, n6428, n6429, n6430, n6431,
    n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
    n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
    n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6583,
    n6584, n6586, n6587, n6589, n6590, n6592, n6593, n6595, n6596, n6597,
    n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6608, n6609,
    n6611, n6612, n6614, n6615, n6617, n6618, n6620, n6621, n6623, n6624,
    n6626, n6627, n6629, n6630, n6632, n6633, n6635, n6636, n6638, n6639,
    n6641, n6642, n6644, n6645, n6647, n6648, n6650, n6651, n6653, n6654,
    n6656, n6657, n6659, n6660, n6662, n6663, n6665, n6666, n6668, n6669,
    n6671, n6672, n6674, n6675, n6677, n6678, n6680, n6681, n6683, n6684,
    n6686, n6687, n6689, n6690, n6692, n6693, n6695, n6696, n6697, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
    n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
    n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6789, n6790, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
    n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
    n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6876, n6877, n6878, n6880, n6881, n6884, n6885, n6886,
    n6887, n6888, n6889, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
    n6911, n6912, n6913, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
    n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7010, n7011,
    n7012, n7013, n7014, n7015, n7016, n7017, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
    n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7055, n7056,
    n7057, n7059, n7060, n7061, n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7132, n7133,
    n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
    n7145, n7146, n7147, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
    n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7231, n7232, n7233, n7234,
    n7235, n7236, n7237, n7238, n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7262, n7263, n7264, n7265, n7266, n7267,
    n7269, n7270, n7271, n7272, n7273, n7275, n7276, n7277, n7278, n7279,
    n7281, n7282, n7283, n7284, n7285, n7287, n7288, n7289, n7290, n7291,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7383, n7384, n7385,
    n7386, n7387, n7388, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
    n7470, n7471, n7472, n7474, n7475, n7476, n7478, n7479, n7480, n7482,
    n7483, n7484, n7486, n7487, n7488, n7490, n7491, n7493, n7494, n7495,
    n7497, n7499, n7500, n7501, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7514, n7515, n7516, n7518, n7519, n7520,
    n7522, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7532, n7533,
    n7534, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
    n7646, n7647, n7648, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7707,
    n7708, n7710, n7711, n7712, n7713, n7714, n7716, n7717, n7718, n7720,
    n7721, n7722, n7724, n7725, n7726, n7728, n7729, n7730, n7732, n7733,
    n7734, n7736, n7737, n7738, n7739, n7741, n7742, n7743, n7744, n7746,
    n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7755, n7756, n7758,
    n7759, n7760, n7761, n7763, n7764, n7765, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7787, n7788, n7789, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7813, n7814,
    n7815, n7816, n7818, n7819, n7821, n7822, n7823, n7825, n7826, n7827,
    n7828, n7829, n7830, n7832, n7833, n7834, n7835, n7836, n7837, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7875, n7876, n7877, n7878, n7880, n7881, n7882, n7883, n7885, n7886,
    n7887, n7888, n7889, n7891, n7892, n7893, n7894, n7895, n7897, n7898,
    n7900, n7901, n7902, n7904, n7905, n7906, n7907, n7908, n7909, n7911,
    n7912, n7913, n7914, n7916, n7917, n7918, n7919, n7920, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940, n7942, n7943, n7944, n7945,
    n7946, n7947, n7949, n7950, n7952, n7953, n7954, n7955, n7956, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994, n7996, n7997, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8020, n8021,
    n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038, n8040, n8041, n8042, n8043,
    n8044, n8045, n8046, n8047, n8048, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
    n8088, n8089, n8090, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
    n8110, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8122, n8123, n8124, n8125, n8126, n8127, n8129, n8130, n8131, n8132,
    n8133, n8134, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8146, n8147, n8148, n8149, n8150, n8151, n8153, n8154, n8155,
    n8156, n8157, n8158, n8160, n8161, n8162, n8163, n8164, n8165, n8167,
    n8168, n8169, n8170, n8171, n8172, n8174, n8175, n8176, n8177, n8178,
    n8179, n8181, n8182, n8183, n8184, n8185, n8186, n8188, n8190, n8191,
    n8193, n8194, n8195, n8197, n8198, n8199, n8200, n8201, n8202, n8204,
    n8205, n8206, n8207, n8208, n8209, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8233, n8234, n8235, n8236, n8237,
    n8238, n8239, n8240, n8241, n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
    n8260, n8261, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
    n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8379, n8380, n8381,
    n8382, n8383, n8385, n8386, n8387, n8388, n8389, n8390, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8413, n8414, n8415,
    n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8551, n8552, n8553, n8554, n8555, n8556, n8558,
    n8559, n8560, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
    n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8602, n8603,
    n8604, n8605, n8606, n8607, n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
    n8626, n8627, n8629, n8630, n8631, n8632, n8633, n8634, n8636, n8637,
    n8638, n8639, n8640, n8641, n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8653, n8654, n8655, n8656, n8657, n8658, n8660,
    n8661, n8662, n8663, n8664, n8665, n8667, n8668, n8669, n8670, n8671,
    n8672, n8674, n8675, n8676, n8677, n8678, n8679, n8681, n8682, n8683,
    n8684, n8685, n8686, n8688, n8689, n8690, n8691, n8692, n8693, n8695,
    n8696, n8697, n8698, n8699, n8700, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
    n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
    n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
    n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
    n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
    n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
    n9012, n9013, n9014, n9015, n9016, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9097, n9098, n9099, n9100, n9101, n9102, n9104, n9105, n9106, n9107,
    n9108, n9109, n9111, n9112, n9113, n9114, n9115, n9116, n9118, n9119,
    n9120, n9121, n9122, n9123, n9125, n9126, n9127, n9128, n9129, n9130,
    n9132, n9133, n9134, n9135, n9136, n9137, n9139, n9140, n9141, n9142,
    n9143, n9144, n9146, n9147, n9148, n9149, n9150, n9151, n9153, n9154,
    n9155, n9156, n9157, n9158, n9160, n9161, n9162, n9163, n9164, n9165,
    n9167, n9168, n9169, n9170, n9171, n9172, n9174, n9175, n9176, n9177,
    n9178, n9179, n9181, n9182, n9183, n9184, n9185, n9186, n9188, n9189,
    n9190, n9191, n9192, n9193, n9195, n9196, n9197, n9198, n9199, n9200,
    n9202, n9203, n9204, n9205, n9206, n9207, n9209, n9210, n9211, n9212,
    n9213, n9214, n9216, n9217, n9218, n9219, n9220, n9221, n9223, n9224,
    n9225, n9226, n9227, n9228, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
    n9280, n9281, n9282, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9407, n9408, n9409, n9410, n9411, n9412,
    n9413, n9414, n9415, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
    n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9490, n9491, n9492, n9493, n9494, n9495, n9497, n9498,
    n9499, n9500, n9501, n9502, n9504, n9505, n9506, n9507, n9508, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9528, n9529, n9530, n9531, n9532,
    n9533, n9534, n9535, n9536, n9538, n9539, n9540, n9541, n9542, n9543,
    n9544, n9545, n9546, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9581, n9582, n9583, n9584, n9585, n9586, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
    n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9614, n9615, n9616, n9617, n9618, n9619,
    n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9628, n9629, n9630,
    n9631, n9632, n9633, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9645, n9646, n9647, n9648, n9649, n9650, n9652, n9653,
    n9654, n9655, n9656, n9657, n9659, n9660, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
    n9676, n9677, n9678, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
    n9698, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
    n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9751, n9752, n9753,
    n9754, n9755, n9756, n9758, n9759, n9760, n9761, n9762, n9763, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9785, n9786, n9787,
    n9788, n9789, n9790, n9792, n9793, n9794, n9795, n9796, n9797, n9799,
    n9800, n9801, n9802, n9803, n9804, n9806, n9807, n9808, n9809, n9810,
    n9811, n9813, n9814, n9815, n9816, n9817, n9818, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
    n9833, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9860, n9861, n9862, n9863, n9864,
    n9865, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
    n9896, n9897, n9898, n9899, n9901, n9902, n9903, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9928,
    n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
    n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
    n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
    n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10026, n10027,
    n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10036, n10037,
    n10038, n10039, n10040, n10041, n10043, n10044, n10045, n10046, n10047,
    n10048, n10050, n10051, n10052, n10053, n10054, n10055, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
    n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10127, n10128, n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
    n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
    n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
    n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10230,
    n10231, n10232, n10233, n10234, n10235, n10237, n10238, n10239, n10240,
    n10241, n10242, n10244, n10245, n10246, n10247, n10248, n10249, n10251,
    n10252, n10253, n10254, n10255, n10256, n10258, n10259, n10260, n10261,
    n10262, n10263, n10265, n10266, n10267, n10268, n10269, n10270, n10272,
    n10273, n10274, n10275, n10276, n10277, n10279, n10280, n10281, n10282,
    n10283, n10284, n10286, n10287, n10288, n10289, n10290, n10291, n10293,
    n10294, n10295, n10296, n10297, n10298, n10300, n10301, n10302, n10303,
    n10304, n10305, n10307, n10308, n10309, n10310, n10311, n10312, n10314,
    n10315, n10316, n10317, n10318, n10319, n10321, n10322, n10323, n10324,
    n10325, n10326, n10328, n10329, n10330, n10331, n10332, n10333, n10335,
    n10336, n10337, n10338, n10339, n10340, n10342, n10343, n10344, n10345,
    n10346, n10347, n10349, n10350, n10351, n10352, n10353, n10354, n10356,
    n10357, n10358, n10359, n10360, n10361, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10386,
    n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
    n10396, n10397, n10398, n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10414, n10415,
    n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
    n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10498, n10499, n10500, n10501, n10502, n10503,
    n10504, n10505, n10506, n10508, n10509, n10510, n10511, n10512, n10513,
    n10514, n10515, n10516, n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10528, n10529, n10530, n10531, n10532, n10533,
    n10534, n10535, n10536, n10538, n10539, n10540, n10541, n10542, n10543,
    n10544, n10545, n10546, n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10618, n10619, n10620, n10621, n10622, n10623,
    n10624, n10625, n10626, n10628, n10629, n10630, n10631, n10632, n10633,
    n10634, n10635, n10636, n10638, n10639, n10640, n10641, n10642, n10643,
    n10644, n10645, n10646, n10648, n10649, n10650, n10651, n10652, n10653,
    n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
    n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10710, n10711, n10712,
    n10713, n10714, n10715, n10717, n10718, n10719, n10720, n10721, n10722,
    n10724, n10725, n10726, n10727, n10728, n10729, n10731, n10732, n10733,
    n10734, n10735, n10736, n10738, n10739, n10740, n10741, n10742, n10743,
    n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
    n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
    n10764, n10765, n10766, n10767, n10768, n10769, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779, n10781, n10782, n10783,
    n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
    n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
    n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
    n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849, n10851, n10852, n10853,
    n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
    n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
    n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
    n10908, n10909, n10910, n10912, n10913, n10914, n10915, n10916, n10917,
    n10918, n10919, n10920, n10922, n10923, n10924, n10925, n10926, n10927,
    n10928, n10929, n10930, n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10942, n10943, n10944, n10945, n10946, n10947,
    n10948, n10949, n10950, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10972, n10973, n10974, n10975, n10976, n10977,
    n10978, n10979, n10980, n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11006,
    n11007, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
    n11026, n11027, n11028, n11029, n11030, n11032, n11033, n11034, n11035,
    n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
    n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
    n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
    n11063, n11064, n11065, n11066, n11067, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
    n11148, n11149, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11206, n11207, n11208, n11209, n11210, n11211, n11213, n11214,
    n11215, n11216, n11217, n11218, n11220, n11221, n11222, n11223, n11224,
    n11225, n11227, n11228, n11229, n11230, n11231, n11232, n11234, n11235,
    n11236, n11237, n11238, n11239, n11241, n11242, n11243, n11244, n11245,
    n11246, n11248, n11249, n11250, n11251, n11252, n11253, n11255, n11256,
    n11257, n11258, n11259, n11260, n11262, n11263, n11264, n11265, n11266,
    n11267, n11269, n11270, n11271, n11272, n11273, n11274, n11276, n11277,
    n11278, n11279, n11280, n11281, n11283, n11284, n11285, n11286, n11287,
    n11288, n11290, n11291, n11292, n11293, n11294, n11295, n11297, n11298,
    n11299, n11300, n11301, n11302, n11304, n11305, n11306, n11307, n11308,
    n11309, n11311, n11312, n11313, n11314, n11315, n11316, n11318, n11319,
    n11320, n11321, n11322, n11323, n11324, n11325, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
    n11378, n11379, n11380, n11382, n11383, n11384, n11385, n11386, n11387,
    n11388, n11389, n11390, n11391, n11392, n11393, n11395, n11396, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11418,
    n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11508,
    n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11568,
    n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11598,
    n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11618,
    n11619, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11631, n11632, n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11648, n11649,
    n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11661, n11662, n11663, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
    n11698, n11699, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
    n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11746,
    n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
    n11766, n11767, n11768, n11769, n11770, n11772, n11773, n11774, n11775,
    n11776, n11777, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
    n11786, n11787, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11801, n11802, n11803, n11804, n11805,
    n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
    n11815, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11827, n11828, n11829, n11830, n11831, n11832, n11834, n11835,
    n11836, n11837, n11838, n11840, n11841, n11842, n11843, n11844, n11845,
    n11847, n11848, n11849, n11850, n11851, n11852, n11854, n11855, n11856,
    n11857, n11858, n11859, n11861, n11862, n11863, n11864, n11865, n11866,
    n11868, n11869, n11870, n11871, n11872, n11873, n11875, n11876, n11877,
    n11878, n11879, n11880, n11881, n11882, n11883, n11885, n11886, n11887,
    n11888, n11889, n11890, n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11916,
    n11917, n11919, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
    n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942, n11944, n11945, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
    n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11982, n11983, n11984, n11985,
    n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
    n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
    n12004, n12005, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
    n12014, n12015, n12016, n12017, n12018, n12019, n12021, n12022, n12023,
    n12024, n12025, n12026, n12028, n12029, n12030, n12031, n12032, n12033,
    n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12049, n12050, n12051, n12052, n12053,
    n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12063,
    n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
    n12073, n12074, n12075, n12076, n12078, n12079, n12080, n12081, n12082,
    n12083, n12084, n12085, n12086, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12098, n12099, n12100, n12101, n12102,
    n12103, n12104, n12105, n12106, n12108, n12109, n12110, n12111, n12112,
    n12113, n12114, n12115, n12116, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12128, n12129, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
    n12143, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12206, n12207,
    n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
    n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
    n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
    n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
    n12244, n12245, n12246, n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12278, n12279, n12281, n12282,
    n12283, n12284, n12285, n12286, n12288, n12289, n12290, n12291, n12292,
    n12293, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12314, n12315, n12316, n12317, n12318, n12319, n12321, n12322,
    n12323, n12324, n12325, n12326, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12396,
    n12397, n12398, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
    n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
    n12425, n12426, n12427, n12428, n12429, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
    n12444, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
    n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
    n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
    n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
    n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
    n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
    n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
    n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
    n12526, n12527, n12528, n12529, n12530, n12531, n12533, n12534, n12535,
    n12536, n12537, n12538, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12554, n12555,
    n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
    n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
    n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12583,
    n12584, n12585, n12586, n12587, n12588, n12590, n12591, n12592, n12593,
    n12594, n12595, n12597, n12598, n12599, n12600, n12601, n12602, n12604,
    n12605, n12606, n12607, n12608, n12609, n12611, n12612, n12613, n12614,
    n12615, n12616, n12618, n12619, n12620, n12621, n12622, n12623, n12625,
    n12626, n12627, n12628, n12629, n12630, n12632, n12633, n12634, n12635,
    n12636, n12637, n12639, n12640, n12641, n12642, n12643, n12644, n12646,
    n12647, n12648, n12649, n12650, n12651, n12653, n12654, n12655, n12656,
    n12657, n12658, n12660, n12661, n12662, n12663, n12664, n12665, n12667,
    n12668, n12669, n12670, n12671, n12672, n12674, n12675, n12676, n12677,
    n12678, n12679, n12681, n12682, n12683, n12684, n12685, n12686, n12688,
    n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
    n12698, n12699, n12700, n12701, n12702, n12704, n12705, n12706, n12707,
    n12708, n12709, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
    n12757, n12758, n12759, n12760, n12762, n12763, n12764, n12765, n12766,
    n12767, n12768, n12769, n12770, n12772, n12773, n12775, n12776, n12777,
    n12778, n12779, n12780, n12781, n12782, n12784, n12785, n12786, n12787,
    n12788, n12789, n12791, n12792, n12793, n12794, n12795, n12796, n12798,
    n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
    n12808, n12809, n12810, n12811, n12813, n12814, n12815, n12816, n12817,
    n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12827,
    n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
    n12846, n12847, n12848, n12849, n12850, n12851, n12853, n12854, n12855,
    n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
    n12865, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
    n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
    n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
    n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
    n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
    n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
    n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
    n12947, n12948, n12949, n12950, n12951, n12952, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
    n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
    n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
    n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
    n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
    n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
    n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
    n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
    n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
    n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
    n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
    n13057, n13058, n13059, n13060, n13061, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110, n13112, n13113, n13114,
    n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
    n13124, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
    n13134, n13135, n13136, n13137, n13138, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
    n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
    n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
    n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
    n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
    n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
    n13254, n13255, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
    n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
    n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
    n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
    n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
    n13300, n13301, n13302, n13304, n13305, n13306, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
    n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
    n13330, n13331, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
    n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
    n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
    n13394, n13395, n13396, n13397, n13398, n13400, n13401, n13402, n13404,
    n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
    n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
    n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
    n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
    n13441, n13442, n13443, n13444, n13445, n13447, n13448, n13449, n13450,
    n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
    n13470, n13471, n13472, n13473, n13474, n13475, n13477, n13478, n13479,
    n13481, n13482, n13483, n13485, n13486, n13487, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497, n13499, n13500, n13501,
    n13502, n13503, n13504, n13506, n13507, n13508, n13509, n13510, n13511,
    n13512, n13513, n13514, n13516, n13517, n13518, n13519, n13520, n13521,
    n13522, n13523, n13524, n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13546, n13547, n13548, n13549, n13550, n13551,
    n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
    n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
    n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
    n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
    n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602, n13604, n13605, n13606,
    n13608, n13609, n13610, n13611, n13612, n13613, n13615, n13616, n13617,
    n13618, n13619, n13620, n13622, n13623, n13624, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13635, n13636, n13637, n13638,
    n13639, n13640, n13641, n13642, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
    n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
    n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13757, n13758, n13759, n13760, n13761, n13762,
    n13763, n13764, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13793,
    n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
    n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
    n13813, n13814, n13815, n13816, n13819, n13820, n13821, n13822, n13823,
    n13824, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
    n13835, n13836, n13837, n13838, n13839, n13840, n13842, n13843, n13844,
    n13846, n13847, n13848, n13850, n13851, n13852, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13872, n13873, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13884, n13885, n13886, n13887,
    n13888, n13889, n13890, n13891, n13893, n13894, n13895, n13896, n13897,
    n13898, n13899, n13900, n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
    n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
    n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
    n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
    n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
    n13981, n13982, n13983, n13984, n13986, n13987, n13988, n13990, n13991,
    n13992, n13994, n13995, n13996, n13998, n13999, n14000, n14001, n14002,
    n14003, n14004, n14005, n14007, n14008, n14010, n14011, n14013, n14014,
    n14015, n14017, n14018, n14020, n14021, n14022, n14023, n14024, n14025,
    n14026, n14028, n14029, n14030, n14031, n14032, n14034, n14035, n14036,
    n14038, n14039, n14040, n14042, n14043, n14044, n14046, n14047, n14048,
    n14051, n14052, n14053, n14055, n14056, n14057, n14059, n14060, n14062,
    n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
    n14123, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
    n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14143,
    n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14152, n14153,
    n14154, n14155, n14156, n14157, n14158, n14159, n14161, n14162, n14163,
    n14164, n14165, n14166, n14167, n14168, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14188, n14189, n14190, n14191, n14192, n14193,
    n14194, n14195, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
    n14204, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
    n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14224,
    n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
    n14285, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
    n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14305,
    n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14314, n14315,
    n14316, n14317, n14318, n14319, n14320, n14321, n14323, n14324, n14325,
    n14326, n14327, n14328, n14329, n14330, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14341, n14342, n14343, n14344, n14345,
    n14346, n14347, n14348, n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
    n14366, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
    n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14386,
    n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
    n14447, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
    n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14476, n14477,
    n14478, n14479, n14480, n14481, n14482, n14483, n14485, n14486, n14487,
    n14488, n14489, n14490, n14491, n14492, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14503, n14504, n14505, n14506, n14507,
    n14508, n14509, n14510, n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
    n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14548,
    n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14575, n14576, n14577, n14578,
    n14579, n14580, n14581, n14582, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
    n14609, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
    n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14638, n14639,
    n14640, n14641, n14642, n14643, n14644, n14645, n14647, n14648, n14649,
    n14650, n14651, n14652, n14653, n14654, n14656, n14657, n14658, n14659,
    n14661, n14662, n14663, n14665, n14666, n14667, n14668, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677, n14679, n14680, n14681,
    n14682, n14683, n14684, n14685, n14686, n14688, n14689, n14690, n14691,
    n14692, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
    n14703, n14704, n14705, n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14716, n14717, n14718, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14729, n14730, n14731, n14732, n14733,
    n14734, n14735, n14736, n14738, n14739, n14741, n14742, n14744, n14745,
    n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
    n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
    n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
    n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
    n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
    n14791, n14792, n14794, n14795, n14797, n14798, n14799, n14800, n14801,
    n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
    n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14847,
    n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
    n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
    n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
    n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
    n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
    n14893, n14894, n14895, n14897, n14898, n14900, n14901, n14903, n14904,
    n14906, n14907, n14909, n14910, n14911, n14912, n14913, n14915, n14916,
    n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
    n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
    n14963, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
    n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
    n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15014, n15015, n15016, n15017, n15018,
    n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
    n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
    n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15063, n15064,
    n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
    n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
    n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15161, n15162, n15163, n15164, n15165,
    n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
    n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
    n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
    n15211, n15212, n15213, n15214, n15215, n15217, n15218, n15219, n15220,
    n15222, n15223, n15225, n15226, n15228, n15229, n15231, n15232, n15234,
    n15235, n15237, n15238, n15240, n15241, n15243, n15244, n15246, n15247,
    n15249, n15250, n15252, n15253, n15255, n15256, n15258, n15259, n15261,
    n15262, n15263, n15264, n15265, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
    n15281, n15282, n15283, n15284, n15285, n15286, n15288, n15289, n15291,
    n15292, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15308, n15309, n15311, n15312,
    n15313, n15314, n15315, n15316, n15317, n15319, n15320, n15322, n15323,
    n15325, n15326, n15328, n15329, n15331, n15332, n15334, n15335, n15337,
    n15338, n15340, n15341, n15343, n15344, n15346, n15347, n15349, n15350,
    n15352, n15353, n15355, n15356, n15358, n15359, n15361, n15362, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15374,
    n15375, n15376, n15377, n15379, n15380, n15381, n15382, n15384, n15385,
    n15386, n15388, n15389, n15390, n15392, n15393, n15395, n15396, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
    n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
    n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15542, n15543, n15544, n15545,
    n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
    n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
    n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15590, n15591,
    n15593, n15594, n15596, n15597, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
    n15613, n15614, n15615, n15617, n15618, n15620, n15621, n15623, n15624,
    n15625, n15626, n15627, n15629, n15630, n15632, n15633, n15636, n15637,
    n15639, n15640, n15642, n15643, n15644, n15646, n15647, n15649, n15651,
    n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
    n15661, n15662, n15663, n15664, n15666, n15667, n15668, n15669, n15671,
    n15672, n15673, n15675, n15676, n15677, n15678, n15680, n15681, n15683,
    n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15697, n15698, n15700, n15701, n15702, n15705,
    n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
    n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
    n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
    n15733, n15734, n15735, n15736, n15737, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15761,
    n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
    n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
    n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
    n15790, n15791, n15792, n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823, n15825, n15826, n15827,
    n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
    n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
    n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
    n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
    n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
    n15883, n15884, n15885, n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
    n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15930,
    n15931, n15932, n15933, n15934, n15936, n15938, n15940, n15942, n15943,
    n15945, n15946, n15948, n15950, n15951, n15953, n15954, n15955, n15956,
    n15958, n15959, n15960, n15962, n15963, n15964, n15965, n15967, n15968,
    n15969, n15970, n15971, n15974, n15975, n15977, n15978, n15980, n15981,
    n15983, n15984, n15986, n15987, n15989, n15990, n15992, n15993, n15995,
    n15996, n15998, n15999, n16001, n16002, n16004, n16005, n16007, n16008,
    n16010, n16011, n16013, n16014, n16016, n16017, n16019, n16020, n16022,
    n16023, n16025, n16026, n16027, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
    n16043, n16044, n16045, n16046, n16047, n16048, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
    n16063, n16064, n16065, n16067, n16068, n16069, n16070, n16071, n16072,
    n16073, n16074, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
    n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
    n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
    n16112, n16113, n16115, n16116, n16117, n16118, n16120, n16121, n16122,
    n16124, n16125, n16126, n16128, n16129, n16130, n16132, n16133, n16134,
    n16136, n16137, n16138, n16139, n16141, n16142, n16143, n16145, n16146,
    n16147, n16149, n16150, n16151, n16153, n16154, n16155, n16156, n16158,
    n16159, n16160, n16162, n16163, n16164, n16166, n16167, n16168, n16170,
    n16171, n16173, n16174, n16176, n16177, n16179, n16180, n16181, n16182,
    n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
    n16193, n16194, n16195, n16196, n16198, n16199, n16201, n16202, n16204,
    n16205, n16207, n16208, n16210, n16211, n16213, n16214, n16216, n16217,
    n16218, n16219, n16220, n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16232, n16234, n16235, n16237, n16238, n16239, n16241,
    n16242, n16243, n16244, n16246, n16247, n16248, n16250, n16251, n16253,
    n16254, n16255, n16257, n16258, n16260, n16261, n16263, n16264, n16266,
    n16267, n16268, n16269, n16270, n16272, n16273, n16274, n16275, n16276,
    n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
    n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
    n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
    n16304, n16305, n16306, n16308, n16309, n16310, n16311, n16312, n16313,
    n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
    n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
    n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
    n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16380, n16381, n16383, n16384, n16386, n16387, n16389, n16390,
    n16392, n16393, n16395, n16396, n16398, n16399, n16400, n16401, n16402,
    n16403, n16404, n16406, n16407, n16408, n16410, n16411, n16412, n16414,
    n16415, n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
    n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16451, n16452,
    n16454, n16455, n16456, n16458, n16459, n16461, n16462, n16463, n16465,
    n16466, n16468, n16469, n16470, n16472, n16473, n16474, n16476, n16477,
    n16478, n16480, n16481, n16482, n16484, n16485, n16487, n16488, n16489,
    n16491, n16492, n16493, n16495, n16496, n16498, n16499, n16501, n16502,
    n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
    n16513, n16515, n16516, n16519, n16520, n16521, n16522, n16523, n16525,
    n16526, n16527, n16528, n16529, n16531, n16532, n16533, n16535, n16536,
    n16538, n16539, n16540, n16542, n16543, n16544, n16546, n16547, n16548,
    n16550, n16551, n16552, n16554, n16555, n16556, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
    n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
    n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
    n16588, n16589, n16590, n16591, n16592, n16593, n16595, n16596, n16597,
    n16599, n16600, n16601, n16603, n16604, n16605, n16607, n16608, n16609,
    n16611, n16612, n16613, n16615, n16616, n16617, n16619, n16620, n16621,
    n16623, n16624, n16625, n16627, n16628, n16629, n16631, n16632, n16633,
    n16635, n16636, n16637, n16639, n16640, n16641, n16643, n16644, n16645,
    n16647, n16648, n16649, n16651, n16652, n16653, n16655, n16656, n16657,
    n16659, n16660, n16661, n16663, n16664, n16665, n16667, n16668, n16669,
    n16671, n16672, n16673, n16675, n16676, n16677, n16679, n16680, n16681,
    n16683, n16684, n16685, n16687, n16688, n16689, n16691, n16692, n16693,
    n16695, n16696, n16697, n16699, n16700, n16701, n16703, n16704, n16705,
    n16707, n16708, n16709, n16711, n16712, n16713, n16715, n16716, n16717,
    n16719, n16720, n16721, n16723, n16724, n16725, n16727, n16728, n16729,
    n16731, n16732, n16733, n16735, n16736, n16737, n16739, n16740, n16741,
    n16743, n16744, n16745, n16747, n16748, n16749, n16751, n16752, n16753,
    n16755, n16756, n16757, n16759, n16760, n16761, n16763, n16764, n16765,
    n16767, n16768, n16769, n16771, n16772, n16773, n16775, n16776, n16777,
    n16779, n16780, n16781, n16783, n16784, n16785, n16787, n16788, n16790,
    n16791, n16793, n16794, n16796, n16797, n16799, n16800, n16802, n16803,
    n16805, n16806, n16808, n16809, n16811, n16812, n16814, n16815, n16817,
    n16818, n16820, n16821, n16823, n16824, n16826, n16827, n16829, n16830,
    n16832, n16833, n16834, n16835, n16836, n16837, n16839, n16840, n16842,
    n16843, n16845, n16846, n16848, n16849, n16851, n16852, n16854, n16855,
    n16857, n16858, n16860, n16861, n16863, n16864, n16866, n16867, n16869,
    n16870, n16872, n16873, n16875, n16876, n16878, n16879, n16881, n16882,
    n16884, n16885, n16887, n16888, n16890, n16891, n16893, n16894, n16896,
    n16897, n16898, n16899, n16900, n16902, n16903, n16905, n16906, n16908,
    n16909, n16911, n16912, n16914, n16915, n16917, n16918, n16920, n16921,
    n16923, n16924, n16926, n16927, n16929, n16930, n16932, n16933, n16935,
    n16936, n16938, n16939, n16941, n16942, n16944, n16945, n16947, n16948,
    n16950, n16951, n16953, n16954, n16956, n16957, n16959, n16960, n16962,
    n16963, n16965, n16966, n16967, n16968, n16969, n16971, n16972, n16974,
    n16975, n16977, n16978, n16980, n16981, n16983, n16984, n16986, n16987,
    n16989, n16990, n16992, n16993, n16995, n16996, n16998, n16999, n17001,
    n17002, n17004, n17005, n17007, n17008, n17010, n17011, n17013, n17014,
    n17016, n17017, n17019, n17020, n17022, n17023, n17025, n17026, n17027,
    n17028, n17029, n17031, n17032, n17034, n17035, n17036, n17038, n17039,
    n17040, n17042, n17043, n17044, n17046, n17047, n17048, n17050, n17051,
    n17052, n17054, n17055, n17058, n17059, n17060, n17062, n17063, n17064,
    n17066, n17067, n17068, n17070, n17071, n17073, n17074, n17076, n17077,
    n17079, n17080, n17082, n17083, n17084, n17086, n17087, n17088, n17090,
    n17091, n17093, n17094, n17096, n17097, n17099, n17100, n17102, n17103,
    n17105, n17106, n17109, n17110, n17111, n17113, n17114, n17115, n17117,
    n17118, n17120, n17121, n17122, n17124, n17125, n17126, n17128, n17129,
    n17130, n17132, n17133, n17134, n17136, n17137, n17138, n17140, n17141,
    n17142, n17144, n17145, n17146, n17148, n17149, n17150, n17152, n17153,
    n17155, n17156, n17158, n17159, n17160, n17162, n17163, n17165, n17166,
    n17167, n17169, n17170, n17171, n17173, n17174, n17176, n17177, n17178,
    n17180, n17181, n17182, n17184, n17185, n17186, n17188, n17189, n17190,
    n17192, n17193, n17194, n17196, n17197, n17199, n17200, n17202, n17203,
    n17204, n17206, n17207, n17209, n17210, n17212, n17213, n17214, n17216,
    n17217, n17219, n17220, n17222, n17223, n17225, n17226, n17228, n17229,
    n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
    n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
    n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
    n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
    n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
    n17276, n17277, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
    n17286, n17287, n17288, n17290, n17291, n17292, n17294, n17295, n17296,
    n17298, n17299, n17300, n17302, n17303, n17304, n17306, n17307, n17309,
    n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
    n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
    n17346, n17347, n17348, n17349, n17350, n17351, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
    n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
    n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
    n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
    n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
    n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
    n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17479, n17480, n17481, n17482, n17483, n17484,
    n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
    n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
    n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17521,
    n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
    n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
    n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
    n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
    n17558, n17559, n17560, n17561, n17562, n17563, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
    n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
    n17604, n17605, n17606, n17607, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
    n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
    n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
    n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
    n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
    n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
    n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
    n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
    n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
    n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
    n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
    n17779, n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
    n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
    n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17827, n17828, n17830, n17831, n17832, n17833, n17835, n17836,
    n17837, n17838, n17840, n17841, n17842, n17843, n17845, n17846, n17847,
    n17848, n17850, n17851, n17852, n17854, n17855, n17857, n17858, n17860,
    n17861, n17863, n17865, n17866, n17868, n17869, n17871, n17872, n17874,
    n17875, n17876, n17878, n17879, n17880, n17882, n17883, n17884, n17886,
    n17887, n17888, n17890, n17891, n17892, n17894, n17895, n17896, n17898,
    n17899, n17900, n17902, n17903, n17904, n17906, n17907, n17908, n17910,
    n17911, n17912, n17914, n17915, n17916, n17918, n17919, n17920, n17922,
    n17923, n17925, n17926, n17928, n17929, n17931, n17932, n17934, n17935,
    n17937, n17938, n17940, n17941, n17943, n17944, n17945, n17947, n17948,
    n17949, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
    n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
    n17996, n17997, n17998, n17999, n18001, n18002, n18003, n18005, n18006,
    n18008, n18009, n18011, n18012, n18014, n18015, n18016, n18018, n18019,
    n18021, n18022, n18023, n18024, n18026, n18027, n18028, n18030, n18031,
    n18032, n18033, n18035, n18036, n18037, n18039, n18040, n18041, n18043,
    n18044, n18045, n18047, n18048, n18049, n18051, n18052, n18053, n18055,
    n18056, n18057, n18059, n18060, n18061, n18063, n18064, n18065, n18067,
    n18069, n18070, n18071, n18073, n18074, n18075, n18076, n18078, n18079,
    n18080, n18082, n18083, n18084, n18086, n18087, n18088, n18090, n18091,
    n18092, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
    n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
    n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
    n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
    n18222, n18223, n18224, n18225, n18226, n18227, n18229, n18230, n18231,
    n18233, n18234, n18235, n18236, n18237, n18238, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18270,
    n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
    n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
    n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
    n18298, n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18330, n18331, n18332, n18333, n18335, n18336,
    n18337, n18339, n18340, n18341, n18343, n18344, n18345, n18347, n18348,
    n18349, n18351, n18352, n18353, n18355, n18356, n18357, n18359, n18360,
    n18361, n18363, n18364, n18365, n18367, n18368, n18369, n18370, n18372,
    n18373, n18374, n18376, n18377, n18378, n18380, n18381, n18382, n18384,
    n18385, n18386, n18388, n18389, n18390, n18392, n18393, n18394, n18396,
    n18397, n18398, n18400, n18401, n18402, n18404, n18405, n18406, n18407,
    n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
    n18426, n18427, n18428, n18429, n18431, n18432, n18433, n18435, n18436,
    n18437, n18439, n18440, n18441, n18443, n18444, n18445, n18447, n18448,
    n18449, n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18476, n18477,
    n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
    n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495,
    n18496, n18497, n18498, n18499, n18501, n18502, n18503, n18505, n18506,
    n18507, n18508, n18510, n18511, n18512, n18514, n18515, n18516, n18518,
    n18519, n18520, n18522, n18523, n18524, n18526, n18527, n18528, n18530,
    n18531, n18532, n18534, n18535, n18536, n18538, n18539, n18540, n18542,
    n18543, n18544, n18546, n18547, n18548, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
    n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18604, n18605, n18606, n18607, n18608, n18609,
    n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
    n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634, n18636, n18637, n18638,
    n18640, n18641, n18642, n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18655, n18656, n18657, n18658, n18659,
    n18660, n18662, n18663, n18665, n18666, n18667, n18669, n18670, n18672,
    n18673, n18675, n18676, n18678, n18679, n18680, n18682, n18683, n18684,
    n18686, n18687, n18688, n18690, n18691, n18692, n18694, n18695, n18696,
    n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18705, n18706,
    n18707, n18708, n18709, n18710, n18711, n18712, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722, n18724, n18726, n18727,
    n18728, n18729, n18730, n18731, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18743, n18744, n18745, n18747, n18748, n18749, n18751,
    n18752, n18753, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18774, n18775, n18776, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18798, n18799, n18800, n18801,
    n18803, n18804, n18805, n18806, n18808, n18809, n18810, n18811, n18813,
    n18814, n18815, n18816, n18818, n18819, n18821, n18822, n18823, n18824,
    n18825, n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18835,
    n18836, n18837, n18838, n18840, n18841, n18843, n18844, n18845, n18846,
    n18847, n18848, n18850, n18851, n18853, n18854, n18855, n18856, n18858,
    n18859, n18860, n18861, n18862, n18863, n18864, n18866, n18867, n18869,
    n18870, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
    n18882, n18883, n18884, n18885, n18886, n18887, n18889, n18890, n18891,
    n18892, n18893, n18894, n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
    n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
    n18922, n18923, n18924, n18925, n18926, n18927, n18930, n18931, n18933,
    n18935, n18936, n18938, n18939, n18941, n18942, n18943, n18944, n18945,
    n18946, n18948, n18949, n18950, n18951, n18953, n18954, n18955, n18956,
    n18957, n18959, n18960, n18961, n18962, n18964, n18965, n18967, n18969,
    n18970, n18972, n18973, n18975, n18976, n18977, n18978, n18980, n18981,
    n18982, n18983, n18986, n18987, n18989, n18991, n18992, n18994, n18995,
    n18996, n18997, n18999, n19000, n19001, n19002, n19004, n19005, n19007,
    n19008, n19009, n19011, n19013, n19014, n19015, n19017, n19018, n19019,
    n19021, n19022, n19023, n19025, n19026, n19027, n19029, n19030, n19031,
    n19032, n19033, n19034, n19039, n19040, n19042, n19043, n19045, n19046,
    n19048, n19050, n19051, n19052, n19054, n19055, n19056, n19058, n19059,
    n19061, n19062, n19063, n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19074, n19075, n19077, n19078, n19079, n19080, n19081, n19082,
    n19084, n19085, n19086, n19087, n19089, n19090, n19091, n19092, n19093,
    n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
    n19114, n19115, n19116, n19118, n19120, n19123, n19124, n19125, n19126,
    n19127, n19129, n19130, n19131, n19133, n19134, n19135, n19137, n19138,
    n19139, n19141, n19142, n19143, n19145, n19146, n19147, n19149, n19150,
    n19152, n19153, n19154, n19155, n19156, n19157, n19159, n19160, n19162,
    n19164, n19165, n19166, n19168, n19170, n19172, n19174, n19176, n19177,
    n19178, n19179, n19180, n19182, n19184, n19185, n19186, n19187, n19188,
    n19190, n19191, n19193, n19194, n19196, n19197, n19198, n19200, n19201,
    n19202, n19204, n19205, n19206, n19208, n19209, n19210, n19212, n19213,
    n19215, n19216, n19217, n19219, n19220, n19221, n19223, n19224, n19225,
    n19227, n19228, n19229, n19231, n19232, n19234, n19235, n19237, n19238,
    n19239, n19241, n19242, n19244, n19245, n19247, n19248, n19250, n19251,
    n19253, n19257, n19258, n19260, n19261, n19263, n19264, n19266, n19267,
    n19269, n19270, n19272, n19274, n19275, n19277, n19278, n19280, n19281,
    n19283, n19284, n19286, n19287, n19289, n19290, n19292, n19293, n19295,
    n19296, n19298, n19299, n19301, n19302, n19304, n19305, n19308, n19309,
    n19311, n19312, n19314, n19315, n19317, n19318, n19320, n19321, n19323,
    n19324, n19326, n19327, n19329, n19330, n19332, n19333, n19335, n19336,
    n19338, n19339, n19341, n19342, n19344, n19345, n19347, n19348, n19350,
    n19351, n19353, n19354, n19356, n19357, n19358, n19359, n19360, n19361,
    n19362, n19363, n19364, n19365, n19366, n19367, n19369, n19370, n19371,
    n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
    n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
    n19391, n19392, n19393, n19395, n19396, n19398, n19399, n19401, n19402,
    n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
    n19422, n19423, n19424, n19425, n19427, n19428, n19429, n19430, n19431,
    n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
    n19451, n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19466, n19467, n19468, n19469, n19470,
    n19471, n19473, n19475, n19477, n19482, n19484, n19485, n19487, n19488,
    n19489, n19491, n19492, n19494, n19495, n19497, n19498, n19500, n19501,
    n19503, n19504, n19506, n19507, n19509, n19510, n19512, n19513, n19515,
    n19516, n19518, n19519, n19521, n19522, n19524, n19525, n19527, n19528,
    n19530, n19531, n19533, n19534, n19536, n19537, n19539, n19540, n19542,
    n19543, n19545, n19546, n19548, n19549, n19551, n19552, n19554, n19555,
    n19557, n19558, n19560, n19561, n19563, n19564, n19566, n19567, n19569,
    n19570, n19572, n19573, n19575, n19576, n19578, n19579, n19581, n19582,
    n19584, n19585, n19587, n19591, n19593, n19594, n19595, n19598, n19599;
  assign n3708 = ~pi1091 & ~pi1370;
  assign n3709 = ~pi0409 & ~pi1088;
  assign n3710 = n3708 & n3709;
  assign n3711 = ~pi0660 & n3710;
  assign n3712 = ~pi0336 & n3711;
  assign n3713 = ~pi0309 & n3712;
  assign n3714 = pi1090 & n3713;
  assign n3715 = ~pi0309 & ~pi1090;
  assign n3716 = ~pi0336 & ~pi0660;
  assign n3717 = n3715 & n3716;
  assign n3718 = n3709 & n3717;
  assign n3719 = pi1091 & n3718;
  assign n3720 = ~pi1370 & n3719;
  assign n3721 = ~pi1091 & n3717;
  assign n3722 = ~pi0409 & n3721;
  assign n3723 = ~pi1370 & n3722;
  assign n3724 = pi1088 & n3723;
  assign n3725 = ~n3720 & ~n3724;
  assign n3726 = ~n3714 & ~n3725;
  assign n3727 = ~pi0138 & n3714;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~pi1101 & ~n3728;
  assign po1210 = pi0196 | n3729;
  assign n3731 = pi0646 & ~po1210;
  assign n3732 = ~pi0634 & ~pi0677;
  assign n3733 = ~pi1401 & n3732;
  assign n3734 = ~pi0619 & ~pi0702;
  assign n3735 = n3733 & n3734;
  assign n3736 = pi0716 & n3735;
  assign n3737 = ~n3731 & n3736;
  assign n3738 = pi1688 & pi1748;
  assign n3739 = pi1773 & n3738;
  assign n3740 = pi1688 & ~pi1748;
  assign n3741 = pi1773 & n3740;
  assign n3742 = ~n3739 & ~n3741;
  assign n3743 = ~pi0716 & ~pi1401;
  assign n3744 = n3732 & n3743;
  assign n3745 = ~pi0702 & n3744;
  assign n3746 = pi0619 & n3745;
  assign n3747 = ~n3742 & n3746;
  assign n3748 = ~n3737 & ~n3747;
  assign n3749 = pi0702 & n3744;
  assign n3750 = ~pi0619 & n3749;
  assign n3751 = ~n3731 & n3750;
  assign n3752 = n3748 & ~n3751;
  assign n3753 = ~n3731 & n3752;
  assign n3754 = ~po1210 & ~n3753;
  assign n3755 = pi0156 & ~n3754;
  assign n3756 = pi1774 & n3754;
  assign po0032 = n3755 | n3756;
  assign n3758 = pi0146 & ~n3754;
  assign n3759 = pi1775 & n3754;
  assign po0033 = n3758 | n3759;
  assign n3761 = pi0175 & ~n3754;
  assign n3762 = pi1776 & n3754;
  assign po0034 = n3761 | n3762;
  assign n3764 = pi0177 & ~n3754;
  assign n3765 = pi1777 & n3754;
  assign po0035 = n3764 | n3765;
  assign n3767 = pi0178 & ~n3754;
  assign n3768 = pi1778 & n3754;
  assign po0036 = n3767 | n3768;
  assign n3770 = pi0144 & ~n3754;
  assign n3771 = pi1779 & n3754;
  assign po0037 = n3770 | n3771;
  assign n3773 = pi0179 & ~n3754;
  assign n3774 = pi1780 & n3754;
  assign po0038 = n3773 | n3774;
  assign n3776 = pi0180 & ~n3754;
  assign n3777 = pi1781 & n3754;
  assign po0039 = n3776 | n3777;
  assign n3779 = pi0181 & ~n3754;
  assign n3780 = pi1782 & n3754;
  assign po0040 = n3779 | n3780;
  assign n3782 = pi0182 & ~n3754;
  assign n3783 = pi1783 & n3754;
  assign po0041 = n3782 | n3783;
  assign n3785 = pi0157 & ~n3754;
  assign n3786 = pi1784 & n3754;
  assign po0042 = n3785 | n3786;
  assign n3788 = pi0159 & ~n3754;
  assign n3789 = pi1785 & n3754;
  assign po0043 = n3788 | n3789;
  assign n3791 = pi0158 & ~n3754;
  assign n3792 = pi1786 & n3754;
  assign po0044 = n3791 | n3792;
  assign n3794 = pi0160 & ~n3754;
  assign n3795 = pi1787 & n3754;
  assign po0045 = n3794 | n3795;
  assign n3797 = pi0161 & ~n3754;
  assign n3798 = pi1788 & n3754;
  assign po0046 = n3797 | n3798;
  assign n3800 = pi0162 & ~n3754;
  assign n3801 = pi1789 & n3754;
  assign po0047 = n3800 | n3801;
  assign n3803 = pi0147 & ~n3754;
  assign n3804 = pi1790 & n3754;
  assign po0048 = n3803 | n3804;
  assign n3806 = pi0163 & ~n3754;
  assign n3807 = pi1791 & n3754;
  assign po0049 = n3806 | n3807;
  assign n3809 = pi0164 & ~n3754;
  assign n3810 = pi1792 & n3754;
  assign po0050 = n3809 | n3810;
  assign n3812 = pi0165 & ~n3754;
  assign n3813 = pi1793 & n3754;
  assign po0051 = n3812 | n3813;
  assign n3815 = pi0166 & ~n3754;
  assign n3816 = pi1794 & n3754;
  assign po0052 = n3815 | n3816;
  assign n3818 = pi0167 & ~n3754;
  assign n3819 = pi1795 & n3754;
  assign po0053 = n3818 | n3819;
  assign n3821 = pi0168 & ~n3754;
  assign n3822 = pi1796 & n3754;
  assign po0054 = n3821 | n3822;
  assign n3824 = pi0169 & ~n3754;
  assign n3825 = pi1797 & n3754;
  assign po0055 = n3824 | n3825;
  assign n3827 = pi0170 & ~n3754;
  assign n3828 = pi1798 & n3754;
  assign po0056 = n3827 | n3828;
  assign n3830 = pi0171 & ~n3754;
  assign n3831 = pi1799 & n3754;
  assign po0057 = n3830 | n3831;
  assign n3833 = pi0172 & ~n3754;
  assign n3834 = pi1800 & n3754;
  assign po0058 = n3833 | n3834;
  assign n3836 = pi0145 & ~n3754;
  assign n3837 = pi1801 & n3754;
  assign po0059 = n3836 | n3837;
  assign n3839 = pi0173 & ~n3754;
  assign n3840 = pi1802 & n3754;
  assign po0060 = n3839 | n3840;
  assign n3842 = pi0174 & ~n3754;
  assign n3843 = pi1803 & n3754;
  assign po0061 = n3842 | n3843;
  assign n3845 = pi0141 & ~n3754;
  assign n3846 = pi1804 & n3754;
  assign po0062 = n3845 | n3846;
  assign n3848 = pi0176 & ~n3754;
  assign n3849 = pi1805 & n3754;
  assign po0063 = n3848 | n3849;
  assign n3851 = ~pi1858 & pi1859;
  assign n3852 = pi1038 & pi1683;
  assign po0072 = n3851 | n3852;
  assign n3854 = ~pi0702 & ~pi0716;
  assign n3855 = n3733 & n3854;
  assign n3856 = ~n3731 & ~n3855;
  assign n3857 = pi0702 & n3856;
  assign n3858 = ~pi0702 & n3739;
  assign n3859 = n3855 & n3858;
  assign n3860 = ~n3857 & ~n3859;
  assign n3861 = ~n3752 & ~n3860;
  assign n3862 = n3754 & n3861;
  assign n3863 = ~pi1669 & ~n3754;
  assign n3864 = po1210 & n3863;
  assign po0075 = n3862 | n3864;
  assign n3866 = pi0038 & ~n3754;
  assign n3867 = pi1758 & n3754;
  assign po0094 = n3866 | n3867;
  assign n3869 = pi0044 & ~n3754;
  assign n3870 = pi1759 & n3754;
  assign po0095 = n3869 | n3870;
  assign n3872 = pi0040 & ~n3754;
  assign n3873 = pi1760 & n3754;
  assign po0096 = n3872 | n3873;
  assign n3875 = pi0039 & ~n3754;
  assign n3876 = pi1761 & n3754;
  assign po0097 = n3875 | n3876;
  assign n3878 = pi0041 & ~n3754;
  assign n3879 = pi1762 & n3754;
  assign po0098 = n3878 | n3879;
  assign n3881 = pi0034 & ~n3754;
  assign n3882 = pi1763 & n3754;
  assign po0099 = n3881 | n3882;
  assign n3884 = pi0035 & ~n3754;
  assign n3885 = pi1764 & n3754;
  assign po0100 = n3884 | n3885;
  assign n3887 = pi0036 & ~n3754;
  assign n3888 = pi1765 & n3754;
  assign po0101 = n3887 | n3888;
  assign n3890 = pi0037 & ~n3754;
  assign n3891 = pi1766 & n3754;
  assign po0102 = n3890 | n3891;
  assign n3893 = pi0045 & ~n3754;
  assign n3894 = pi1767 & n3754;
  assign po0103 = n3893 | n3894;
  assign n3896 = pi0042 & ~n3754;
  assign n3897 = pi1768 & n3754;
  assign po0104 = n3896 | n3897;
  assign n3899 = pi0031 & ~n3754;
  assign n3900 = pi1769 & n3754;
  assign po0105 = n3899 | n3900;
  assign n3902 = pi0043 & ~n3754;
  assign n3903 = pi1770 & n3754;
  assign po0106 = n3902 | n3903;
  assign n3905 = pi0032 & ~n3754;
  assign n3906 = pi1771 & n3754;
  assign po0107 = n3905 | n3906;
  assign n3908 = pi0033 & ~n3754;
  assign n3909 = pi1772 & n3754;
  assign po0108 = n3908 | n3909;
  assign po1733 = pi0096 | pi1018;
  assign po0179 = ~pi0093 | po1733;
  assign n3913 = pi0068 & po0179;
  assign n3914 = ~pi1753 & ~n3913;
  assign n3915 = pi1667 & n3914;
  assign n3916 = pi0000 & n3915;
  assign n3917 = ~pi0004 & ~pi0005;
  assign n3918 = pi0004 & pi0005;
  assign n3919 = ~n3917 & ~n3918;
  assign n3920 = ~pi0065 & pi0093;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = ~pi0055 & ~pi0059;
  assign n3923 = ~pi1429 & n3922;
  assign n3924 = ~pi1422 & n3923;
  assign n3925 = pi0061 & n3924;
  assign n3926 = ~pi0061 & ~pi1422;
  assign n3927 = ~pi0059 & n3926;
  assign n3928 = pi0055 & n3927;
  assign n3929 = ~pi1429 & n3928;
  assign n3930 = pi0058 & pi1692;
  assign n3931 = ~po1733 & n3930;
  assign n3932 = n3929 & n3931;
  assign n3933 = ~n3925 & ~n3932;
  assign n3934 = pi1422 & n3923;
  assign n3935 = ~pi0061 & n3934;
  assign n3936 = pi0059 & n3926;
  assign n3937 = ~pi0055 & n3936;
  assign n3938 = ~pi1429 & n3937;
  assign n3939 = po1733 & n3938;
  assign n3940 = ~pi0094 & po1733;
  assign n3941 = n3938 & n3940;
  assign n3942 = ~n3939 & ~n3941;
  assign n3943 = n3922 & n3926;
  assign n3944 = pi1429 & n3943;
  assign n3945 = n3942 & ~n3944;
  assign n3946 = ~n3935 & n3945;
  assign n3947 = n3933 & n3946;
  assign n3948 = pi0055 & pi1692;
  assign n3949 = pi0058 & n3948;
  assign n3950 = ~pi0874 & ~n3949;
  assign n3951 = ~pi0152 & n3950;
  assign n3952 = pi0152 & ~n3950;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~pi0193 & ~pi0874;
  assign n3955 = pi0055 & n3930;
  assign n3956 = n3954 & ~n3955;
  assign n3957 = ~pi0874 & ~n3955;
  assign n3958 = pi0152 & pi0199;
  assign n3959 = ~pi0193 & n3958;
  assign n3960 = pi0193 & ~n3958;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~n3957 & n3961;
  assign n3963 = ~n3956 & ~n3962;
  assign n3964 = ~pi0199 & n3950;
  assign n3965 = ~pi0152 & pi0199;
  assign n3966 = ~n3950 & ~n3965;
  assign n3967 = pi0152 & ~pi0199;
  assign n3968 = n3966 & ~n3967;
  assign n3969 = ~n3964 & ~n3968;
  assign n3970 = ~n3963 & n3969;
  assign n3971 = n3953 & n3970;
  assign n3972 = pi1644 & n3971;
  assign n3973 = ~pi0193 & n3957;
  assign n3974 = ~n3962 & ~n3973;
  assign n3975 = ~n3965 & ~n3967;
  assign n3976 = ~n3950 & n3975;
  assign n3977 = ~n3964 & ~n3976;
  assign n3978 = ~n3974 & ~n3977;
  assign n3979 = n3953 & n3978;
  assign n3980 = pi1664 & n3979;
  assign n3981 = ~n3972 & ~n3980;
  assign n3982 = ~n3953 & n3970;
  assign n3983 = pi1638 & n3982;
  assign n3984 = ~n3953 & n3978;
  assign n3985 = pi1645 & n3984;
  assign n3986 = ~n3983 & ~n3985;
  assign n3987 = n3981 & n3986;
  assign n3988 = n3963 & n3969;
  assign n3989 = n3953 & n3988;
  assign n3990 = pi1585 & n3989;
  assign n3991 = n3963 & ~n3977;
  assign n3992 = n3953 & n3991;
  assign n3993 = pi1614 & n3992;
  assign n3994 = ~n3990 & ~n3993;
  assign n3995 = ~n3953 & n3988;
  assign n3996 = pi1563 & n3995;
  assign n3997 = ~n3953 & n3991;
  assign n3998 = pi1586 & n3997;
  assign n3999 = ~n3996 & ~n3998;
  assign n4000 = n3994 & n3999;
  assign n4001 = n3987 & n4000;
  assign n4002 = n3947 & ~n4001;
  assign n4003 = ~pi1692 & n3935;
  assign n4004 = ~n3925 & ~n4003;
  assign n4005 = ~n3932 & n4004;
  assign n4006 = pi1422 & pi1692;
  assign n4007 = ~n3944 & ~n4006;
  assign n4008 = n4005 & n4007;
  assign n4009 = pi0982 & n4008;
  assign n4010 = pi0052 & n4005;
  assign n4011 = ~pi0779 & ~n4005;
  assign n4012 = ~n4010 & ~n4011;
  assign n4013 = ~n4008 & ~n4012;
  assign n4014 = ~n4009 & ~n4013;
  assign n4015 = ~n3947 & ~n4014;
  assign n4016 = ~n4002 & ~n4015;
  assign n4017 = n3920 & n4016;
  assign n4018 = ~n3921 & ~n4017;
  assign n4019 = ~n3914 & n4018;
  assign po0110 = n3916 | n4019;
  assign n4021 = pi0001 & n3915;
  assign n4022 = pi0004 & ~pi0005;
  assign n4023 = ~pi0004 & pi0005;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = ~n3920 & ~n4024;
  assign n4026 = pi1658 & n3984;
  assign n4027 = pi1633 & n3971;
  assign n4028 = ~n4026 & ~n4027;
  assign n4029 = pi1663 & n3979;
  assign n4030 = pi1636 & n3982;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = pi1575 & n3997;
  assign n4033 = pi1600 & n3992;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = pi1601 & n3995;
  assign n4036 = pi1573 & n3989;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = n4034 & n4037;
  assign n4039 = n4031 & n4038;
  assign n4040 = n4028 & n4039;
  assign n4041 = n3947 & ~n4040;
  assign n4042 = pi0025 & ~n4005;
  assign n4043 = pi0013 & n4005;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = ~n4008 & ~n4044;
  assign n4046 = ~pi0982 & n4008;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = ~n3947 & ~n4047;
  assign n4049 = ~n4041 & ~n4048;
  assign n4050 = n3920 & n4049;
  assign n4051 = ~n4025 & ~n4050;
  assign n4052 = ~n3914 & n4051;
  assign po0111 = n4021 | n4052;
  assign n4054 = pi0002 & n3915;
  assign n4055 = pi0005 & ~n3920;
  assign n4056 = pi1584 & n3989;
  assign n4057 = pi1632 & n3984;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = pi1641 & n3979;
  assign n4060 = pi1648 & n3971;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = pi1610 & n3992;
  assign n4063 = pi1589 & n3997;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n4061 & n4064;
  assign n4066 = pi1591 & n3995;
  assign n4067 = pi1640 & n3982;
  assign n4068 = ~n4066 & ~n4067;
  assign n4069 = n4065 & n4068;
  assign n4070 = n4058 & n4069;
  assign n4071 = n3947 & ~n4070;
  assign n4072 = pi1016 & n4008;
  assign n4073 = pi0060 & n4005;
  assign n4074 = ~pi0778 & ~n4005;
  assign n4075 = ~n4073 & ~n4074;
  assign n4076 = ~n4008 & ~n4075;
  assign n4077 = ~n4072 & ~n4076;
  assign n4078 = ~n3947 & ~n4077;
  assign n4079 = ~n4071 & ~n4078;
  assign n4080 = n3920 & n4079;
  assign n4081 = ~n4055 & ~n4080;
  assign n4082 = ~n3914 & n4081;
  assign po0112 = n4054 | n4082;
  assign n4084 = pi0003 & n3915;
  assign n4085 = pi1659 & n3982;
  assign n4086 = pi1643 & n3971;
  assign n4087 = pi1635 & n3984;
  assign n4088 = ~n4086 & ~n4087;
  assign n4089 = pi1595 & n3997;
  assign n4090 = pi1593 & n3992;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = pi1649 & n3979;
  assign n4093 = n4091 & ~n4092;
  assign n4094 = pi1599 & n3995;
  assign n4095 = pi1574 & n3989;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = n4093 & n4096;
  assign n4098 = n4088 & n4097;
  assign n4099 = ~n4085 & n4098;
  assign n4100 = n3947 & ~n4099;
  assign n4101 = ~pi0054 & ~n4005;
  assign n4102 = pi0010 & n4005;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~n4008 & ~n4103;
  assign n4105 = ~pi1016 & n4008;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = ~n3947 & ~n4106;
  assign n4108 = ~n4100 & ~n4107;
  assign n4109 = n3920 & n4108;
  assign n4110 = ~pi0005 & ~n3920;
  assign n4111 = ~n4109 & ~n4110;
  assign n4112 = ~n3914 & n4111;
  assign po0113 = n4084 | n4112;
  assign n4114 = ~pi1229 & ~pi1236;
  assign n4115 = pi1227 & ~pi1228;
  assign po1676 = n4114 & n4115;
  assign n4117 = pi1470 & po1676;
  assign n4118 = ~pi1229 & pi1236;
  assign po1678 = n4115 & n4118;
  assign n4120 = pi1471 & po1678;
  assign n4121 = ~n4117 & ~n4120;
  assign n4122 = ~pi0771 & ~pi0801;
  assign n4123 = ~n4121 & n4122;
  assign n4124 = pi1470 & pi1471;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = ~pi0771 & pi0801;
  assign n4127 = ~pi0385 & n4126;
  assign n4128 = pi0771 & ~pi0801;
  assign n4129 = ~pi0125 & n4128;
  assign n4130 = ~n4127 & ~n4129;
  assign n4131 = pi0796 & ~n4122;
  assign n4132 = ~n4130 & n4131;
  assign n4133 = n4125 & ~n4132;
  assign n4134 = pi1229 & ~pi1236;
  assign n4135 = n4115 & n4134;
  assign n4136 = pi0352 & ~n4135;
  assign n4137 = ~pi0780 & pi0798;
  assign n4138 = n4136 & ~n4137;
  assign n4139 = ~n4133 & n4138;
  assign n4140 = ~pi0088 & ~pi0092;
  assign n4141 = ~pi0110 & ~pi0111;
  assign n4142 = ~pi0095 & ~pi0112;
  assign n4143 = n4141 & n4142;
  assign n4144 = ~pi0089 & ~pi0108;
  assign n4145 = n4143 & n4144;
  assign n4146 = ~pi0109 & n4145;
  assign n4147 = n4140 & n4146;
  assign n4148 = ~pi0110 & n4147;
  assign n4149 = pi0780 & ~pi0798;
  assign n4150 = n4148 & ~n4149;
  assign n4151 = n4139 & n4150;
  assign n4152 = ~pi0725 & ~pi0743;
  assign n4153 = pi0006 & pi0008;
  assign n4154 = pi1479 & n4153;
  assign n4155 = ~pi0625 & n4154;
  assign n4156 = n4152 & ~n4155;
  assign n4157 = pi0110 & ~n4147;
  assign n4158 = ~n4156 & n4157;
  assign n4159 = ~pi0138 & n4158;
  assign po0114 = n4151 | n4159;
  assign n4161 = n4138 & n4148;
  assign n4162 = n4149 & n4161;
  assign n4163 = n4154 & n4157;
  assign n4164 = ~pi0138 & ~pi0625;
  assign n4165 = n4152 & n4164;
  assign n4166 = n4163 & n4165;
  assign po0115 = n4162 | n4166;
  assign n4168 = pi1458 & n4122;
  assign n4169 = ~pi0796 & ~pi1471;
  assign n4170 = ~pi0767 & ~pi1470;
  assign n4171 = n4169 & ~n4170;
  assign n4172 = ~n4122 & n4171;
  assign n4173 = ~n4168 & ~n4172;
  assign n4174 = ~pi0776 & ~n4173;
  assign n4175 = pi0024 & n4173;
  assign n4176 = ~n4131 & n4175;
  assign n4177 = ~pi1470 & ~n4132;
  assign n4178 = ~n4176 & n4177;
  assign po0116 = n4174 | ~n4178;
  assign n4180 = pi1493 & n4122;
  assign n4181 = ~n4128 & ~n4180;
  assign n4182 = n4131 & ~n4181;
  assign n4183 = ~n4126 & ~n4168;
  assign n4184 = pi0192 & ~n4183;
  assign n4185 = ~n4182 & n4184;
  assign n4186 = ~pi0740 & ~n4185;
  assign n4187 = ~pi1099 & ~n4186;
  assign n4188 = pi0740 & n4185;
  assign n4189 = pi0877 & n4182;
  assign n4190 = pi0236 & n4183;
  assign n4191 = pi0189 & ~n4183;
  assign n4192 = ~n4190 & ~n4191;
  assign n4193 = ~n4182 & ~n4192;
  assign n4194 = ~n4189 & ~n4193;
  assign n4195 = ~pi0739 & n4194;
  assign n4196 = pi0759 & n4182;
  assign n4197 = pi0135 & ~n4183;
  assign n4198 = ~n4182 & n4197;
  assign n4199 = ~n4182 & n4183;
  assign n4200 = pi0243 & n4199;
  assign n4201 = ~n4198 & ~n4200;
  assign n4202 = ~pi0875 & n4201;
  assign n4203 = ~n4196 & n4202;
  assign n4204 = ~n4195 & ~n4203;
  assign n4205 = pi0190 & ~n4183;
  assign n4206 = ~n4182 & n4205;
  assign n4207 = ~pi0864 & ~n4206;
  assign n4208 = pi0191 & ~n4182;
  assign n4209 = ~n4183 & n4208;
  assign n4210 = pi0774 & ~n4209;
  assign n4211 = ~n4207 & ~n4210;
  assign n4212 = pi0242 & n4199;
  assign n4213 = pi0809 & n4182;
  assign n4214 = pi0132 & ~n4182;
  assign n4215 = ~n4183 & n4214;
  assign n4216 = ~n4213 & ~n4215;
  assign n4217 = ~n4212 & n4216;
  assign n4218 = ~pi0868 & n4217;
  assign n4219 = pi0224 & n4199;
  assign n4220 = pi0810 & n4182;
  assign n4221 = pi0134 & ~n4182;
  assign n4222 = ~n4183 & n4221;
  assign n4223 = ~n4220 & ~n4222;
  assign n4224 = ~n4219 & n4223;
  assign n4225 = ~pi0869 & n4224;
  assign n4226 = ~n4218 & ~n4225;
  assign n4227 = pi0241 & n4199;
  assign n4228 = pi0808 & n4182;
  assign n4229 = pi0133 & ~n4182;
  assign n4230 = ~n4183 & n4229;
  assign n4231 = ~n4228 & ~n4230;
  assign n4232 = ~n4227 & n4231;
  assign n4233 = ~pi0867 & n4232;
  assign n4234 = pi0755 & n4182;
  assign n4235 = pi0221 & n4183;
  assign n4236 = pi0151 & ~n4183;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~n4182 & ~n4237;
  assign n4239 = ~n4234 & ~n4238;
  assign n4240 = ~pi0945 & n4239;
  assign n4241 = ~n4233 & ~n4240;
  assign n4242 = n4226 & n4241;
  assign n4243 = n4211 & n4242;
  assign n4244 = pi0804 & n4182;
  assign n4245 = pi0238 & n4183;
  assign n4246 = pi0150 & ~n4183;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = ~n4182 & ~n4247;
  assign n4249 = ~n4244 & ~n4248;
  assign n4250 = ~pi0940 & n4249;
  assign n4251 = pi0240 & n4183;
  assign n4252 = pi0188 & ~n4183;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4182 & ~n4253;
  assign n4255 = pi0807 & n4182;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = ~pi0742 & n4256;
  assign n4258 = pi0239 & n4183;
  assign n4259 = pi0149 & ~n4183;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4182 & ~n4260;
  assign n4262 = pi0806 & n4182;
  assign n4263 = ~pi0741 & ~n4262;
  assign n4264 = ~n4261 & n4263;
  assign n4265 = ~n4257 & ~n4264;
  assign n4266 = pi0859 & n4182;
  assign n4267 = pi0187 & ~n4183;
  assign n4268 = pi0257 & n4183;
  assign n4269 = ~n4267 & ~n4268;
  assign n4270 = ~n4182 & ~n4269;
  assign n4271 = ~n4266 & ~n4270;
  assign n4272 = ~pi0895 & ~n4271;
  assign n4273 = pi0750 & n4182;
  assign n4274 = pi0237 & n4183;
  assign n4275 = pi0148 & ~n4183;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n4182 & ~n4276;
  assign n4278 = ~n4273 & ~n4277;
  assign n4279 = ~pi0946 & n4278;
  assign n4280 = n4272 & ~n4279;
  assign n4281 = n4265 & n4280;
  assign n4282 = ~n4250 & n4281;
  assign n4283 = pi0742 & ~n4256;
  assign n4284 = ~n4261 & ~n4262;
  assign n4285 = pi0741 & ~n4284;
  assign n4286 = ~n4257 & n4285;
  assign n4287 = ~n4283 & ~n4286;
  assign n4288 = pi0946 & ~n4278;
  assign n4289 = ~n4250 & n4288;
  assign n4290 = pi0940 & ~n4249;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = n4265 & ~n4291;
  assign n4293 = n4287 & ~n4292;
  assign n4294 = ~n4282 & n4293;
  assign n4295 = n4243 & ~n4294;
  assign n4296 = n4204 & n4295;
  assign n4297 = pi0869 & ~n4224;
  assign n4298 = pi0868 & ~n4217;
  assign n4299 = ~n4225 & n4298;
  assign n4300 = ~n4297 & ~n4299;
  assign n4301 = pi0867 & ~n4232;
  assign n4302 = pi0945 & ~n4239;
  assign n4303 = ~n4233 & n4302;
  assign n4304 = ~n4301 & ~n4303;
  assign n4305 = n4226 & ~n4304;
  assign n4306 = n4300 & ~n4305;
  assign n4307 = n4204 & ~n4306;
  assign n4308 = pi0739 & ~n4194;
  assign n4309 = ~n4196 & ~n4198;
  assign n4310 = ~n4200 & n4309;
  assign n4311 = pi0875 & ~n4310;
  assign n4312 = ~n4195 & n4311;
  assign n4313 = ~n4308 & ~n4312;
  assign n4314 = ~n4307 & n4313;
  assign n4315 = n4211 & ~n4314;
  assign n4316 = pi0864 & n4206;
  assign n4317 = ~n4210 & n4316;
  assign n4318 = ~pi0774 & n4209;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = ~n4315 & n4319;
  assign n4321 = ~n4296 & n4320;
  assign n4322 = ~n4188 & n4321;
  assign n4323 = n4187 & n4322;
  assign n4324 = ~n4296 & ~n4315;
  assign n4325 = n4319 & n4324;
  assign n4326 = ~n4186 & ~n4188;
  assign n4327 = ~pi1099 & ~n4326;
  assign n4328 = ~n4325 & n4327;
  assign n4329 = ~pi0815 & pi1099;
  assign n4330 = ~n4328 & ~n4329;
  assign po0117 = n4323 | ~n4330;
  assign n4332 = pi0024 & ~n4173;
  assign n4333 = pi0672 & n4173;
  assign n4334 = ~n4332 & ~n4333;
  assign po0118 = pi1471 | ~n4334;
  assign n4336 = ~pi0066 & ~pi1625;
  assign n4337 = pi1542 & n4336;
  assign n4338 = n3955 & n4005;
  assign n4339 = ~n4337 & ~n4338;
  assign n4340 = pi0009 & n4339;
  assign n4341 = n4040 & n4099;
  assign n4342 = ~n4040 & ~n4099;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = pi0025 & pi0053;
  assign n4345 = ~pi0025 & ~pi0053;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = n4343 & n4346;
  assign n4348 = ~n4343 & ~n4346;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = n3987 & ~n4070;
  assign n4351 = n4000 & n4350;
  assign n4352 = ~n4057 & ~n4066;
  assign n4353 = ~n4063 & ~n4067;
  assign n4354 = n4352 & n4353;
  assign n4355 = ~n4056 & ~n4062;
  assign n4356 = n4061 & n4355;
  assign n4357 = n4354 & n4356;
  assign n4358 = ~n4001 & n4357;
  assign n4359 = ~n4351 & ~n4358;
  assign n4360 = pi1642 & n3984;
  assign n4361 = pi1662 & n3979;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = pi1598 & n3995;
  assign n4364 = pi1592 & n3989;
  assign n4365 = ~n4363 & ~n4364;
  assign n4366 = n4362 & n4365;
  assign n4367 = pi1655 & n3982;
  assign n4368 = pi1634 & n3971;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = pi1606 & n3997;
  assign n4371 = pi1588 & n3992;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = n4369 & n4372;
  assign n4374 = n4366 & n4373;
  assign n4375 = pi1596 & n3997;
  assign n4376 = pi1615 & n3992;
  assign n4377 = ~n4375 & ~n4376;
  assign n4378 = pi1577 & n3995;
  assign n4379 = pi1609 & n3989;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = n4377 & n4380;
  assign n4382 = pi1652 & n3971;
  assign n4383 = pi1654 & n3982;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = pi1660 & n3979;
  assign n4386 = pi1646 & n3984;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = n4384 & n4387;
  assign n4389 = n4381 & n4388;
  assign n4390 = n4374 & n4389;
  assign n4391 = ~n4374 & ~n4389;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = n4359 & n4392;
  assign n4394 = ~n4359 & ~n4392;
  assign n4395 = ~n4393 & ~n4394;
  assign n4396 = n4349 & n4395;
  assign n4397 = ~n4349 & ~n4395;
  assign n4398 = ~n4396 & ~n4397;
  assign n4399 = pi0779 & ~pi0878;
  assign n4400 = ~pi0779 & pi0878;
  assign n4401 = ~n4399 & ~n4400;
  assign n4402 = ~pi0054 & pi0777;
  assign n4403 = pi0054 & ~pi0777;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4401 & n4404;
  assign n4406 = n4401 & ~n4404;
  assign n4407 = ~n4405 & ~n4406;
  assign n4408 = pi0747 & pi0778;
  assign n4409 = ~pi0747 & ~pi0778;
  assign n4410 = ~n4408 & ~n4409;
  assign n4411 = pi1650 & n3984;
  assign n4412 = pi1605 & n3995;
  assign n4413 = ~n4411 & ~n4412;
  assign n4414 = pi1647 & n3979;
  assign n4415 = pi1576 & n3989;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = n4413 & n4416;
  assign n4418 = pi1656 & n3982;
  assign n4419 = pi1590 & n3992;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = pi1587 & n3997;
  assign n4422 = pi1639 & n3971;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = n4420 & n4423;
  assign n4425 = n4417 & n4424;
  assign n4426 = pi1653 & n3979;
  assign n4427 = pi1661 & n3971;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = pi1657 & n3982;
  assign n4430 = pi1651 & n3984;
  assign n4431 = ~n4429 & ~n4430;
  assign n4432 = n4428 & n4431;
  assign n4433 = pi1602 & n3989;
  assign n4434 = pi1597 & n3992;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = pi1603 & n3995;
  assign n4437 = pi1564 & n3997;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = n4435 & n4438;
  assign n4440 = n4432 & n4439;
  assign n4441 = ~n4425 & n4440;
  assign n4442 = n4417 & ~n4440;
  assign n4443 = n4424 & n4442;
  assign n4444 = ~n4441 & ~n4443;
  assign n4445 = pi0009 & n4444;
  assign n4446 = ~pi0009 & ~n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = n4410 & n4447;
  assign n4449 = ~n4410 & ~n4447;
  assign n4450 = ~n4448 & ~n4449;
  assign n4451 = n4407 & n4450;
  assign n4452 = ~n4407 & ~n4450;
  assign n4453 = ~n4451 & ~n4452;
  assign n4454 = ~n4398 & n4453;
  assign n4455 = n4398 & ~n4453;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~n4339 & ~n4456;
  assign n4458 = pi1625 & po1733;
  assign n4459 = ~n4457 & ~n4458;
  assign po0119 = n4340 | ~n4459;
  assign n4461 = ~pi0010 & n4339;
  assign n4462 = ~pi0777 & pi0878;
  assign n4463 = pi0777 & ~pi0878;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = pi0054 & n4464;
  assign n4466 = ~pi0054 & ~n4464;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = n4099 & n4392;
  assign n4469 = ~n4099 & ~n4392;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = ~n4467 & n4470;
  assign n4472 = n4467 & ~n4470;
  assign n4473 = ~n4471 & ~n4472;
  assign n4474 = ~pi0778 & pi0779;
  assign n4475 = pi0778 & ~pi0779;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = pi0009 & ~pi0747;
  assign n4478 = ~pi0009 & pi0747;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = ~n4359 & n4444;
  assign n4481 = n4359 & ~n4444;
  assign n4482 = ~n4480 & ~n4481;
  assign n4483 = n4479 & n4482;
  assign n4484 = ~n4479 & ~n4482;
  assign n4485 = ~n4483 & ~n4484;
  assign n4486 = n4476 & n4485;
  assign n4487 = ~n4476 & ~n4485;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = ~n4473 & n4488;
  assign n4490 = n4473 & ~n4488;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = ~n4339 & ~n4491;
  assign n4493 = ~n4458 & ~n4492;
  assign po0120 = n4461 | ~n4493;
  assign n4495 = ~n4186 & n4318;
  assign n4496 = ~n4188 & ~n4495;
  assign n4497 = ~n4186 & ~n4210;
  assign n4498 = ~n4207 & n4308;
  assign n4499 = ~n4316 & ~n4498;
  assign n4500 = ~n4195 & ~n4207;
  assign n4501 = n4225 & ~n4297;
  assign n4502 = ~n4203 & ~n4501;
  assign n4503 = ~n4218 & n4301;
  assign n4504 = ~n4298 & ~n4503;
  assign n4505 = ~n4297 & n4504;
  assign n4506 = n4502 & ~n4505;
  assign n4507 = ~n4311 & ~n4506;
  assign n4508 = n4500 & ~n4507;
  assign n4509 = n4499 & ~n4508;
  assign n4510 = n4497 & ~n4509;
  assign n4511 = n4496 & ~n4510;
  assign n4512 = ~n4250 & ~n4264;
  assign n4513 = ~n4280 & ~n4288;
  assign n4514 = n4512 & ~n4513;
  assign n4515 = ~n4264 & n4290;
  assign n4516 = ~n4285 & ~n4515;
  assign n4517 = ~n4514 & n4516;
  assign n4518 = ~n4240 & ~n4257;
  assign n4519 = ~n4517 & n4518;
  assign n4520 = ~n4240 & n4283;
  assign n4521 = ~n4302 & ~n4520;
  assign n4522 = ~n4519 & n4521;
  assign n4523 = ~n4203 & ~n4225;
  assign n4524 = ~n4218 & ~n4233;
  assign n4525 = n4523 & n4524;
  assign n4526 = ~n4522 & n4525;
  assign n4527 = n4497 & n4500;
  assign n4528 = n4526 & n4527;
  assign n4529 = n4511 & ~n4528;
  assign n4530 = pi0865 & n4529;
  assign n4531 = ~pi0865 & ~n4529;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~pi1099 & ~n4532;
  assign n4534 = ~pi0870 & pi1099;
  assign po0121 = n4533 | n4534;
  assign n4536 = pi0024 & n4183;
  assign n4537 = pi0029 & ~n4183;
  assign po0122 = n4536 | n4537;
  assign n4539 = ~pi0013 & n4339;
  assign n4540 = ~n4476 & n4479;
  assign n4541 = n4476 & ~n4479;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = pi0025 & pi0054;
  assign n4544 = ~pi0025 & ~pi0054;
  assign n4545 = ~n4543 & ~n4544;
  assign n4546 = n4464 & ~n4545;
  assign n4547 = ~n4464 & n4545;
  assign n4548 = ~n4546 & ~n4547;
  assign n4549 = ~n4542 & n4548;
  assign n4550 = n4542 & ~n4548;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = n4343 & ~n4392;
  assign n4553 = ~n4343 & n4392;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = ~n4482 & n4554;
  assign n4556 = n4482 & ~n4554;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~n4551 & n4557;
  assign n4559 = n4551 & ~n4557;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~n4339 & ~n4560;
  assign n4562 = ~n4458 & ~n4561;
  assign po0123 = n4539 | ~n4562;
  assign n4564 = ~n4210 & ~n4318;
  assign n4565 = ~n4521 & n4524;
  assign n4566 = n4504 & ~n4565;
  assign n4567 = n4518 & n4524;
  assign n4568 = ~n4517 & n4567;
  assign n4569 = n4566 & ~n4568;
  assign n4570 = n4500 & n4523;
  assign n4571 = ~n4569 & n4570;
  assign n4572 = ~n4203 & n4297;
  assign n4573 = ~n4311 & ~n4572;
  assign n4574 = n4500 & ~n4573;
  assign n4575 = n4499 & ~n4574;
  assign n4576 = ~n4571 & n4575;
  assign n4577 = n4564 & n4576;
  assign n4578 = ~n4564 & ~n4576;
  assign n4579 = ~n4577 & ~n4578;
  assign n4580 = ~pi1099 & ~n4579;
  assign n4581 = ~pi0814 & pi1099;
  assign po0124 = n4580 | n4581;
  assign n4583 = pi0865 & pi0866;
  assign n4584 = ~n4496 & n4583;
  assign n4585 = n4497 & n4583;
  assign n4586 = ~n4575 & n4585;
  assign n4587 = ~n4584 & ~n4586;
  assign n4588 = n4570 & n4585;
  assign n4589 = ~n4569 & n4588;
  assign n4590 = n4587 & ~n4589;
  assign n4591 = pi0775 & ~n4590;
  assign n4592 = ~pi0775 & n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~pi1099 & ~n4593;
  assign n4595 = ~pi0817 & pi1099;
  assign po0125 = n4594 | n4595;
  assign n4597 = ~n4195 & ~n4308;
  assign n4598 = n4507 & ~n4526;
  assign n4599 = n4597 & n4598;
  assign n4600 = ~n4597 & ~n4598;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~pi1099 & ~n4601;
  assign n4603 = ~pi0812 & pi1099;
  assign po0126 = n4602 | n4603;
  assign n4605 = pi0017 & n3915;
  assign n4606 = pi0878 & ~n4005;
  assign n4607 = ~pi0051 & n4005;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = ~n3947 & ~n4008;
  assign n4610 = n4608 & n4609;
  assign n4611 = n3947 & ~n4374;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = ~n3914 & ~n4612;
  assign n4614 = ~n3914 & ~n3920;
  assign n4615 = ~n4613 & ~n4614;
  assign po0127 = n4605 | ~n4615;
  assign n4617 = ~pi0816 & pi1099;
  assign n4618 = pi0865 & n4188;
  assign n4619 = pi0865 & ~n4186;
  assign n4620 = ~n4319 & n4619;
  assign n4621 = ~n4618 & ~n4620;
  assign n4622 = n4211 & n4619;
  assign n4623 = n4204 & ~n4300;
  assign n4624 = n4313 & ~n4623;
  assign n4625 = n4622 & ~n4624;
  assign n4626 = n4621 & ~n4625;
  assign n4627 = n4204 & n4226;
  assign n4628 = n4622 & n4627;
  assign n4629 = ~n4250 & ~n4279;
  assign n4630 = n4272 & n4629;
  assign n4631 = ~n4289 & ~n4630;
  assign n4632 = ~n4290 & n4631;
  assign n4633 = n4265 & ~n4632;
  assign n4634 = n4241 & n4633;
  assign n4635 = n4241 & ~n4287;
  assign n4636 = n4304 & ~n4635;
  assign n4637 = ~n4634 & n4636;
  assign n4638 = n4628 & ~n4637;
  assign n4639 = n4626 & ~n4638;
  assign n4640 = pi0866 & ~n4639;
  assign n4641 = ~pi0866 & n4639;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = ~pi1099 & n4642;
  assign po0128 = n4617 | n4643;
  assign n4645 = ~n4207 & ~n4316;
  assign n4646 = n4627 & ~n4637;
  assign n4647 = n4624 & ~n4646;
  assign n4648 = n4645 & n4647;
  assign n4649 = ~n4645 & ~n4647;
  assign n4650 = ~n4648 & ~n4649;
  assign n4651 = ~pi1099 & ~n4650;
  assign n4652 = ~pi0813 & pi1099;
  assign po0129 = n4651 | n4652;
  assign n4654 = pi0020 & n3915;
  assign n4655 = n3947 & ~n4440;
  assign n4656 = pi0048 & n4005;
  assign n4657 = ~pi0747 & ~n4005;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n3947 & ~n4658;
  assign n4660 = ~n4655 & ~n4659;
  assign n4661 = ~n3947 & n4008;
  assign n4662 = n4660 & ~n4661;
  assign n4663 = ~n3914 & ~n4662;
  assign n4664 = ~n4614 & ~n4663;
  assign po0130 = n4654 | ~n4664;
  assign n4666 = pi0021 & n3915;
  assign n4667 = ~n3914 & n3920;
  assign n4668 = n3947 & n4425;
  assign n4669 = pi0009 & ~n4005;
  assign n4670 = pi0053 & n4005;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = ~n3947 & ~n4671;
  assign n4673 = ~n4668 & ~n4672;
  assign n4674 = ~n4661 & ~n4673;
  assign n4675 = n4667 & ~n4674;
  assign po0131 = n4666 | n4675;
  assign n4677 = ~n4203 & ~n4311;
  assign n4678 = n4242 & ~n4294;
  assign n4679 = n4306 & ~n4678;
  assign n4680 = n4677 & n4679;
  assign n4681 = ~n4677 & ~n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = ~pi1099 & ~n4682;
  assign n4684 = ~pi0834 & pi1099;
  assign po0132 = n4683 | n4684;
  assign n4686 = ~n4233 & ~n4301;
  assign n4687 = ~n4522 & ~n4686;
  assign n4688 = n4522 & n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~pi1099 & ~n4689;
  assign n4691 = ~pi0832 & pi1099;
  assign po0133 = n4690 | n4691;
  assign n4693 = pi0086 & pi0281;
  assign n4694 = pi0200 & n4693;
  assign n4695 = ~pi0218 & ~pi0877;
  assign n4696 = ~pi0355 & ~pi0809;
  assign n4697 = ~pi0280 & ~pi0810;
  assign n4698 = ~pi0353 & ~pi0759;
  assign n4699 = ~pi0759 & ~pi0810;
  assign n4700 = ~pi0280 & ~pi0353;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~n4698 & n4701;
  assign n4703 = ~n4697 & n4702;
  assign n4704 = n4696 & ~n4703;
  assign n4705 = ~pi0355 & ~pi0431;
  assign n4706 = ~pi0808 & n4705;
  assign n4707 = ~pi0808 & ~pi0809;
  assign n4708 = ~pi0431 & n4707;
  assign n4709 = ~n4706 & ~n4708;
  assign n4710 = ~n4703 & ~n4709;
  assign n4711 = ~n4704 & ~n4710;
  assign n4712 = ~pi0810 & n4700;
  assign n4713 = ~pi0353 & n4699;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = ~pi0280 & ~pi0759;
  assign n4716 = n4714 & ~n4715;
  assign n4717 = n4711 & n4716;
  assign n4718 = pi0218 & pi0877;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = ~n4695 & ~n4719;
  assign n4721 = n4694 & n4720;
  assign n4722 = ~pi0355 & ~pi0808;
  assign n4723 = ~pi0431 & ~pi0809;
  assign n4724 = ~n4705 & ~n4707;
  assign n4725 = ~n4723 & n4724;
  assign n4726 = ~n4722 & n4725;
  assign n4727 = ~n4718 & ~n4726;
  assign n4728 = ~n4703 & n4727;
  assign n4729 = n4721 & ~n4728;
  assign n4730 = pi0333 & ~pi0807;
  assign n4731 = pi0620 & ~pi0755;
  assign n4732 = pi0333 & pi0620;
  assign n4733 = ~pi0755 & ~pi0807;
  assign n4734 = ~n4732 & ~n4733;
  assign n4735 = ~n4731 & n4734;
  assign n4736 = ~n4730 & n4735;
  assign n4737 = ~pi0804 & ~pi0806;
  assign n4738 = ~pi0673 & n4737;
  assign n4739 = ~pi0545 & ~pi0673;
  assign n4740 = ~pi0804 & n4739;
  assign n4741 = ~n4738 & ~n4740;
  assign n4742 = ~pi0545 & ~pi0806;
  assign n4743 = n4741 & ~n4742;
  assign n4744 = ~n4736 & ~n4743;
  assign n4745 = ~pi0807 & n4732;
  assign n4746 = pi0620 & n4733;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = pi0333 & ~pi0755;
  assign n4749 = n4721 & ~n4748;
  assign n4750 = n4747 & n4749;
  assign n4751 = ~n4744 & n4750;
  assign n4752 = pi0726 & pi0750;
  assign n4753 = pi1358 & ~n4752;
  assign n4754 = pi0750 & pi0859;
  assign n4755 = ~pi0726 & ~n4754;
  assign n4756 = ~n4753 & ~n4755;
  assign n4757 = ~pi0750 & ~pi0859;
  assign n4758 = n4756 & ~n4757;
  assign n4759 = ~n4736 & ~n4758;
  assign n4760 = ~pi0545 & ~pi0804;
  assign n4761 = ~pi0673 & ~pi0806;
  assign n4762 = ~n4737 & ~n4739;
  assign n4763 = ~n4761 & n4762;
  assign n4764 = ~n4760 & n4763;
  assign n4765 = n4759 & ~n4764;
  assign n4766 = n4751 & ~n4765;
  assign po0134 = n4729 | n4766;
  assign n4768 = ~pi0025 & n4339;
  assign n4769 = ~pi0013 & ~pi0747;
  assign n4770 = pi0013 & pi0747;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = n4447 & ~n4771;
  assign n4773 = ~n4447 & n4771;
  assign n4774 = ~n4772 & ~n4773;
  assign n4775 = ~n4339 & ~n4774;
  assign n4776 = ~n4768 & ~n4775;
  assign po0135 = n4458 | ~n4776;
  assign n4778 = pi0026 & n3915;
  assign n4779 = pi0777 & ~n4005;
  assign n4780 = ~pi0050 & n4005;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = n4609 & n4781;
  assign n4783 = n3947 & ~n4389;
  assign n4784 = ~n4782 & ~n4783;
  assign n4785 = n4667 & ~n4784;
  assign po0136 = n4778 | n4785;
  assign n4787 = ~n4225 & ~n4297;
  assign n4788 = n4569 & n4787;
  assign n4789 = ~n4569 & ~n4787;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = ~pi1099 & ~n4790;
  assign n4792 = ~pi0833 & pi1099;
  assign po0137 = n4791 | n4792;
  assign n4794 = ~n4240 & ~n4302;
  assign n4795 = n4294 & n4794;
  assign n4796 = ~n4294 & ~n4794;
  assign n4797 = ~n4795 & ~n4796;
  assign n4798 = ~pi1099 & ~n4797;
  assign n4799 = ~pi0831 & pi1099;
  assign po0138 = n4798 | n4799;
  assign n4801 = pi0355 & pi0431;
  assign n4802 = pi0280 & n4801;
  assign n4803 = pi0353 & n4802;
  assign n4804 = n4693 & n4803;
  assign n4805 = pi0200 & n4804;
  assign n4806 = pi0218 & n4805;
  assign n4807 = ~pi1358 & n4806;
  assign n4808 = pi0545 & n4807;
  assign n4809 = pi0673 & n4808;
  assign n4810 = pi0726 & n4809;
  assign n4811 = ~pi0333 & ~pi0620;
  assign po0139 = n4810 & n4811;
  assign n4813 = ~n4218 & ~n4298;
  assign n4814 = n4637 & n4813;
  assign n4815 = ~n4637 & ~n4813;
  assign n4816 = ~n4814 & ~n4815;
  assign n4817 = ~pi1099 & ~n4816;
  assign n4818 = ~pi0757 & pi1099;
  assign po0140 = n4817 | n4818;
  assign n4820 = ~pi0097 & ~pi0121;
  assign n4821 = pi1101 & pi1579;
  assign n4822 = pi0031 & ~n4821;
  assign n4823 = pi0036 & pi0037;
  assign n4824 = pi0038 & pi0040;
  assign n4825 = pi0044 & n4824;
  assign n4826 = pi0039 & n4825;
  assign n4827 = pi0034 & pi0035;
  assign n4828 = pi0041 & n4827;
  assign n4829 = n4826 & n4828;
  assign n4830 = n4823 & n4829;
  assign n4831 = pi0042 & n4830;
  assign n4832 = pi0045 & n4831;
  assign n4833 = pi0031 & n4832;
  assign n4834 = ~pi0031 & ~n4832;
  assign n4835 = ~n4833 & ~n4834;
  assign n4836 = n4821 & n4835;
  assign n4837 = ~n4822 & ~n4836;
  assign n4838 = pi0042 & ~n4821;
  assign n4839 = pi0037 & pi0045;
  assign n4840 = pi0035 & pi0036;
  assign n4841 = pi0034 & pi0041;
  assign n4842 = n4826 & n4841;
  assign n4843 = n4840 & n4842;
  assign n4844 = n4839 & n4843;
  assign n4845 = pi0042 & n4844;
  assign n4846 = ~pi0042 & ~n4844;
  assign n4847 = ~n4845 & ~n4846;
  assign n4848 = n4821 & n4847;
  assign n4849 = ~n4838 & ~n4848;
  assign n4850 = pi0102 & n4849;
  assign n4851 = ~pi0102 & ~n4849;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = n4823 & n4827;
  assign n4854 = pi0038 & pi0044;
  assign n4855 = pi0040 & n4854;
  assign n4856 = pi0041 & n4855;
  assign n4857 = pi0039 & n4856;
  assign n4858 = n4853 & n4857;
  assign n4859 = pi0045 & ~n4858;
  assign n4860 = ~pi0045 & n4858;
  assign n4861 = ~n4859 & ~n4860;
  assign n4862 = n4821 & ~n4861;
  assign n4863 = pi0045 & ~n4821;
  assign n4864 = ~n4862 & ~n4863;
  assign n4865 = pi0120 & n4864;
  assign n4866 = ~pi0120 & ~n4864;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4852 & ~n4867;
  assign n4869 = pi0031 & pi0042;
  assign n4870 = n4839 & n4869;
  assign n4871 = pi0041 & n4826;
  assign n4872 = pi0034 & n4871;
  assign n4873 = n4840 & n4872;
  assign n4874 = n4870 & n4873;
  assign n4875 = pi0043 & ~n4874;
  assign n4876 = ~pi0043 & n4874;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = n4821 & ~n4877;
  assign n4879 = pi0043 & ~n4821;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = ~pi0113 & n4880;
  assign n4882 = pi0113 & ~n4880;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = n4868 & ~n4883;
  assign n4885 = pi0036 & ~n4821;
  assign n4886 = pi0036 & n4829;
  assign n4887 = ~pi0036 & ~n4829;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = n4821 & n4888;
  assign n4890 = ~n4885 & ~n4889;
  assign n4891 = pi0245 & n4890;
  assign n4892 = ~pi0245 & ~n4890;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = pi0035 & ~n4821;
  assign n4895 = pi0035 & n4842;
  assign n4896 = ~pi0035 & ~n4842;
  assign n4897 = ~n4895 & ~n4896;
  assign n4898 = n4821 & n4897;
  assign n4899 = ~n4894 & ~n4898;
  assign n4900 = pi0140 & n4899;
  assign n4901 = ~pi0140 & ~n4899;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = pi0041 & ~n4821;
  assign n4904 = ~pi0041 & ~n4826;
  assign n4905 = ~n4871 & ~n4904;
  assign n4906 = n4821 & n4905;
  assign n4907 = ~n4903 & ~n4906;
  assign n4908 = pi0215 & n4907;
  assign n4909 = ~pi0215 & ~n4907;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = ~n4902 & ~n4910;
  assign n4912 = ~n4893 & n4911;
  assign n4913 = pi0037 & ~n4821;
  assign n4914 = pi0037 & n4873;
  assign n4915 = ~pi0037 & ~n4873;
  assign n4916 = ~n4914 & ~n4915;
  assign n4917 = n4821 & n4916;
  assign n4918 = ~n4913 & ~n4917;
  assign n4919 = pi0139 & n4918;
  assign n4920 = ~pi0139 & ~n4918;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = pi0034 & ~n4821;
  assign n4923 = pi0034 & n4857;
  assign n4924 = ~pi0034 & ~n4857;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = n4821 & n4925;
  assign n4927 = ~n4922 & ~n4926;
  assign n4928 = pi0216 & n4927;
  assign n4929 = ~pi0216 & ~n4927;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = ~n4921 & ~n4930;
  assign n4932 = n4912 & n4931;
  assign n4933 = n4884 & n4932;
  assign n4934 = ~pi0038 & pi0044;
  assign n4935 = pi0038 & ~pi0044;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = n4821 & ~n4936;
  assign n4938 = pi0044 & ~n4821;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = pi0361 & n4939;
  assign n4941 = ~pi0361 & ~n4939;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = pi0038 & ~n4821;
  assign n4944 = ~pi0038 & n4821;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = pi0701 & n4945;
  assign n4947 = ~pi0701 & ~n4945;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = pi0039 & ~n4821;
  assign n4950 = ~pi0039 & ~n4825;
  assign n4951 = ~n4826 & ~n4950;
  assign n4952 = n4821 & n4951;
  assign n4953 = ~n4949 & ~n4952;
  assign n4954 = pi0282 & n4953;
  assign n4955 = ~pi0282 & ~n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = pi0040 & ~n4821;
  assign n4958 = ~pi0040 & ~n4854;
  assign n4959 = ~n4855 & ~n4958;
  assign n4960 = n4821 & n4959;
  assign n4961 = ~n4957 & ~n4960;
  assign n4962 = pi0260 & n4961;
  assign n4963 = ~pi0260 & ~n4961;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n4956 & ~n4964;
  assign n4966 = ~n4948 & n4965;
  assign n4967 = ~n4942 & n4966;
  assign n4968 = pi0033 & ~n4821;
  assign n4969 = n4844 & n4869;
  assign n4970 = pi0032 & n4969;
  assign n4971 = pi0043 & n4970;
  assign n4972 = ~pi0033 & n4971;
  assign n4973 = pi0033 & ~n4971;
  assign n4974 = ~n4972 & ~n4973;
  assign n4975 = n4821 & ~n4974;
  assign n4976 = ~n4968 & ~n4975;
  assign n4977 = pi0091 & ~n4976;
  assign n4978 = ~pi0091 & n4976;
  assign n4979 = ~n4977 & ~n4978;
  assign n4980 = n4967 & ~n4979;
  assign n4981 = pi0032 & ~n4821;
  assign n4982 = pi0045 & n4853;
  assign n4983 = n4857 & n4982;
  assign n4984 = pi0042 & n4983;
  assign n4985 = pi0043 & n4984;
  assign n4986 = pi0031 & n4985;
  assign n4987 = pi0032 & n4986;
  assign n4988 = ~pi0032 & ~n4986;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = n4821 & n4989;
  assign n4991 = ~n4981 & ~n4990;
  assign n4992 = pi0090 & n4991;
  assign n4993 = ~pi0090 & ~n4991;
  assign n4994 = ~n4992 & ~n4993;
  assign n4995 = pi0122 & n4837;
  assign n4996 = ~pi0122 & ~n4837;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = n4994 & ~n4997;
  assign n4999 = n4131 & n4998;
  assign n5000 = n4980 & n4999;
  assign n5001 = n4933 & n5000;
  assign n5002 = ~n4837 & ~n5001;
  assign n5003 = n4820 & n5002;
  assign n5004 = pi1001 & ~n4820;
  assign po0141 = n5003 | n5004;
  assign n5006 = ~n4991 & ~n5001;
  assign n5007 = n4820 & n5006;
  assign n5008 = ~pi1003 & ~n4820;
  assign po0142 = n5007 | n5008;
  assign n5010 = ~n4976 & ~n5001;
  assign n5011 = n4820 & n5010;
  assign n5012 = ~pi1004 & ~n4820;
  assign po0143 = n5011 | n5012;
  assign n5014 = ~n4927 & ~n5001;
  assign n5015 = n4820 & n5014;
  assign n5016 = ~pi1009 & ~n4820;
  assign po0145 = n5015 | n5016;
  assign n5018 = ~n4899 & ~n5001;
  assign n5019 = n4820 & n5018;
  assign n5020 = ~pi1010 & ~n4820;
  assign po0146 = n5019 | n5020;
  assign n5022 = ~n4890 & ~n5001;
  assign n5023 = n4820 & n5022;
  assign n5024 = ~pi1011 & ~n4820;
  assign po0147 = n5023 | n5024;
  assign n5026 = ~n4918 & ~n5001;
  assign n5027 = n4820 & n5026;
  assign n5028 = pi1012 & ~n4820;
  assign po0148 = n5027 | n5028;
  assign n5030 = ~n4945 & ~n5001;
  assign n5031 = n4820 & n5030;
  assign n5032 = pi0999 & ~n4820;
  assign po0149 = n5031 | n5032;
  assign n5034 = ~n4953 & ~n5001;
  assign n5035 = n4820 & n5034;
  assign n5036 = pi1007 & ~n4820;
  assign po0150 = n5035 | n5036;
  assign n5038 = ~n4961 & ~n5001;
  assign n5039 = n4820 & n5038;
  assign n5040 = pi1006 & ~n4820;
  assign po0151 = n5039 | n5040;
  assign n5042 = ~n4907 & ~n5001;
  assign n5043 = n4820 & n5042;
  assign n5044 = ~pi1008 & ~n4820;
  assign po0152 = n5043 | n5044;
  assign n5046 = ~n4849 & ~n5001;
  assign n5047 = n4820 & n5046;
  assign n5048 = ~pi1000 & ~n4820;
  assign po0153 = n5047 | n5048;
  assign n5050 = ~n4880 & ~n5001;
  assign n5051 = n4820 & n5050;
  assign n5052 = ~pi1002 & ~n4820;
  assign po0154 = n5051 | n5052;
  assign n5054 = ~n4939 & ~n5001;
  assign n5055 = n4820 & n5054;
  assign n5056 = pi1005 & ~n4820;
  assign po0155 = n5055 | n5056;
  assign n5058 = ~n4864 & ~n5001;
  assign n5059 = n4820 & n5058;
  assign n5060 = ~pi1013 & ~n4820;
  assign po0156 = n5059 | n5060;
  assign n5062 = ~n4257 & ~n4283;
  assign n5063 = ~n4517 & ~n5062;
  assign n5064 = n4517 & n5062;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = ~pi1099 & ~n5065;
  assign n5067 = ~pi0830 & pi1099;
  assign po0157 = n5066 | n5067;
  assign n5069 = pi1549 & ~pi1753;
  assign n5070 = pi0047 & n5069;
  assign n5071 = ~pi1692 & n3944;
  assign n5072 = pi1692 & n3935;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = ~n3929 & n3942;
  assign n5075 = ~n3925 & n5074;
  assign po0173 = n3935 | ~n5075;
  assign n5077 = pi1667 & ~po0173;
  assign n5078 = pi0093 & n5077;
  assign n5079 = n5073 & n5078;
  assign n5080 = ~n5070 & n5079;
  assign po0158 = pi1747 & ~n5080;
  assign n5082 = ~pi0048 & n4339;
  assign n5083 = n4359 & ~n4476;
  assign n5084 = ~n4359 & n4476;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = ~n4339 & ~n5085;
  assign n5087 = ~n5082 & ~n5086;
  assign po0159 = n4458 | ~n5087;
  assign n5089 = ~n4264 & ~n4285;
  assign n5090 = ~n4632 & ~n5089;
  assign n5091 = n4632 & n5089;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = pi0012 & n4131;
  assign n5094 = pi0095 & ~n5093;
  assign n5095 = ~n5092 & n5094;
  assign n5096 = pi0983 & ~pi1099;
  assign n5097 = ~pi0756 & pi1099;
  assign n5098 = ~n5096 & ~n5097;
  assign n5099 = ~n5094 & ~n5098;
  assign po0160 = n5095 | n5099;
  assign n5101 = ~pi0050 & n4339;
  assign n5102 = ~n4343 & ~n4545;
  assign n5103 = n4343 & n4545;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = ~n4339 & ~n5104;
  assign n5106 = ~n5101 & ~n5105;
  assign po0161 = n4458 | ~n5106;
  assign n5108 = ~pi0051 & n4339;
  assign n5109 = n4099 & ~n4389;
  assign n5110 = ~n4099 & n4389;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = ~n4404 & n5111;
  assign n5113 = n4404 & ~n5111;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = ~n4339 & ~n5114;
  assign n5116 = ~n5108 & ~n5115;
  assign po0162 = n4458 | ~n5116;
  assign n5118 = ~pi0052 & n4339;
  assign n5119 = ~n4392 & ~n4464;
  assign n5120 = n4392 & n4464;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = ~n4339 & ~n5121;
  assign n5123 = ~n5118 & ~n5122;
  assign po0163 = n4458 | ~n5123;
  assign n5125 = pi0053 & n4339;
  assign n5126 = ~n4070 & n4440;
  assign n5127 = n4070 & ~n4440;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = n4410 & n5128;
  assign n5130 = ~n4410 & ~n5128;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = ~n4339 & ~n5131;
  assign n5133 = ~n5125 & ~n5132;
  assign po0164 = n4458 | ~n5133;
  assign n5135 = pi0054 & n4339;
  assign n5136 = ~pi0010 & n4425;
  assign n5137 = pi0010 & ~n4425;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = pi0009 & n5138;
  assign n5140 = ~pi0009 & ~n5138;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = ~n4339 & ~n5141;
  assign n5143 = ~n5135 & ~n5142;
  assign po0165 = n4458 | ~n5143;
  assign n5145 = n3929 & ~n3931;
  assign n5146 = pi0055 & n5145;
  assign n5147 = pi0055 & ~pi1692;
  assign n5148 = n3944 & n5147;
  assign n5149 = ~pi0055 & ~po1733;
  assign n5150 = n3938 & ~n3940;
  assign n5151 = ~n5149 & n5150;
  assign n5152 = ~n5148 & ~n5151;
  assign n5153 = ~n5146 & n5152;
  assign po0166 = pi1747 & ~n5153;
  assign n5155 = ~n4250 & ~n4290;
  assign n5156 = ~n4513 & ~n5155;
  assign n5157 = n4513 & n5155;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = n5094 & ~n5158;
  assign n5160 = pi0894 & ~pi1099;
  assign n5161 = ~pi0828 & pi1099;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~n5094 & ~n5162;
  assign po0167 = n5159 | n5163;
  assign n5165 = ~n4279 & ~n4288;
  assign n5166 = n4272 & n5165;
  assign n5167 = ~n4272 & ~n5165;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = n5094 & n5168;
  assign n5170 = ~pi1099 & ~n4131;
  assign n5171 = ~pi0012 & ~pi0805;
  assign n5172 = pi0767 & pi0805;
  assign n5173 = ~pi0767 & ~pi0805;
  assign n5174 = ~n5172 & ~n5173;
  assign n5175 = pi0012 & ~n5174;
  assign n5176 = ~n5171 & ~n5175;
  assign n5177 = ~n5094 & ~n5176;
  assign n5178 = n5170 & n5177;
  assign n5179 = pi1099 & ~n5094;
  assign n5180 = ~pi0820 & n5179;
  assign n5181 = ~n5178 & ~n5180;
  assign po0168 = n5169 | ~n5181;
  assign n5183 = ~pi0059 & ~pi1692;
  assign n5184 = n3944 & ~n5183;
  assign n5185 = pi0059 & n3935;
  assign n5186 = ~pi1692 & n5185;
  assign n5187 = pi0059 & n5150;
  assign n5188 = ~po1733 & n5187;
  assign n5189 = pi1747 & ~n5188;
  assign n5190 = ~n5186 & n5189;
  assign po0170 = n5184 | ~n5190;
  assign n5192 = ~pi0060 & n4339;
  assign n5193 = n4001 & ~n4374;
  assign n5194 = ~n4001 & n4374;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = ~n4401 & n5195;
  assign n5197 = n4401 & ~n5195;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~n4339 & ~n5198;
  assign n5200 = ~n5192 & ~n5199;
  assign po0171 = n4458 | ~n5200;
  assign n5202 = pi0061 & n3944;
  assign n5203 = ~pi1692 & n5202;
  assign n5204 = pi0061 & ~po1733;
  assign n5205 = n3938 & n5204;
  assign n5206 = ~n3941 & ~n5205;
  assign n5207 = ~n5203 & n5206;
  assign po0172 = pi1747 & ~n5207;
  assign po0174 = ~pi0086 & ~pi1099;
  assign n5210 = ~pi0012 & pi0767;
  assign n5211 = pi0012 & ~pi0767;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = n5170 & ~n5212;
  assign n5214 = ~pi0811 & pi1099;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = ~n5094 & ~n5215;
  assign n5217 = pi0895 & n4271;
  assign n5218 = ~n4272 & ~n5217;
  assign n5219 = n5094 & n5218;
  assign po0175 = n5216 | n5219;
  assign n5221 = pi0065 & ~pi1692;
  assign n5222 = pi0093 & ~n5221;
  assign po0176 = pi1747 & ~n5222;
  assign n5224 = pi1747 & n5073;
  assign n5225 = pi0066 & ~n4458;
  assign n5226 = ~pi0094 & n4458;
  assign n5227 = ~n5225 & ~n5226;
  assign po0177 = n5224 & ~n5227;
  assign n5229 = ~pi1227 & ~pi1228;
  assign po1690 = n4134 & n5229;
  assign n5231 = pi1479 & po1690;
  assign n5232 = pi1229 & pi1236;
  assign po1688 = n4115 & n5232;
  assign n5234 = ~po1676 & ~po1688;
  assign n5235 = n4122 & ~n5234;
  assign n5236 = ~n4128 & ~n5235;
  assign n5237 = po1678 & n4122;
  assign n5238 = ~n4126 & ~n5237;
  assign n5239 = n5236 & n5238;
  assign n5240 = pi0067 & n5239;
  assign n5241 = ~n5231 & n5240;
  assign n5242 = n4133 & n4138;
  assign n5243 = n5241 & n5242;
  assign n5244 = ~pi0111 & ~pi0112;
  assign n5245 = ~pi0110 & n5244;
  assign n5246 = ~pi0095 & n5245;
  assign n5247 = ~pi0108 & ~pi0109;
  assign n5248 = ~pi0089 & ~pi0092;
  assign n5249 = n5247 & n5248;
  assign n5250 = n5246 & n5249;
  assign n5251 = pi0067 & ~pi0088;
  assign n5252 = n5250 & n5251;
  assign n5253 = ~n4149 & n5252;
  assign n5254 = n5243 & n5253;
  assign n5255 = pi0067 & n5252;
  assign n5256 = ~n4138 & n5255;
  assign n5257 = ~n5254 & ~n5256;
  assign n5258 = ~pi1227 & pi1228;
  assign n5259 = n4114 & n5258;
  assign n5260 = pi1233 & n5259;
  assign n5261 = pi0067 & ~n5260;
  assign n5262 = ~pi1417 & ~n5261;
  assign n5263 = n5246 & n5248;
  assign n5264 = ~pi0067 & ~pi0088;
  assign n5265 = pi0108 & n5264;
  assign n5266 = ~pi0109 & n5265;
  assign n5267 = n5263 & n5266;
  assign n5268 = ~n5262 & n5267;
  assign n5269 = n5257 & ~n5268;
  assign n5270 = ~pi0095 & n5264;
  assign n5271 = n5244 & n5249;
  assign n5272 = n5270 & n5271;
  assign n5273 = pi0110 & n5272;
  assign n5274 = ~n4165 & n5273;
  assign n5275 = n5269 & ~n5274;
  assign n5276 = ~pi0110 & n5270;
  assign n5277 = n5249 & n5276;
  assign n5278 = ~pi0111 & pi0112;
  assign n5279 = n5277 & n5278;
  assign n5280 = ~pi0108 & n5264;
  assign n5281 = pi0109 & n5280;
  assign n5282 = n5263 & n5281;
  assign n5283 = pi0138 & n5282;
  assign n5284 = ~n5279 & ~n5283;
  assign n5285 = pi1043 & pi1068;
  assign n5286 = ~pi1043 & ~pi1068;
  assign n5287 = ~n5285 & ~n5286;
  assign n5288 = ~pi1049 & pi1096;
  assign n5289 = pi1049 & ~pi1096;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~pi1041 & pi1069;
  assign n5292 = pi1041 & ~pi1069;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = n5290 & n5293;
  assign n5295 = ~pi1039 & pi1094;
  assign n5296 = pi1039 & ~pi1094;
  assign n5297 = ~n5295 & ~n5296;
  assign n5298 = ~pi1040 & pi1095;
  assign n5299 = pi1040 & ~pi1095;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = n5297 & n5300;
  assign n5302 = n5294 & n5301;
  assign n5303 = ~n5287 & n5302;
  assign n5304 = pi1233 & n5303;
  assign n5305 = ~pi1479 & po1690;
  assign n5306 = n4118 & n5229;
  assign n5307 = ~n5305 & ~n5306;
  assign n5308 = pi1234 & n5307;
  assign n5309 = n5304 & n5308;
  assign n5310 = ~pi1313 & pi1318;
  assign n5311 = pi1313 & ~pi1318;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = pi1042 & ~pi1044;
  assign n5314 = ~pi1042 & pi1044;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~pi1039 & pi1040;
  assign n5317 = pi1039 & ~pi1040;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = pi1041 & ~pi1049;
  assign n5320 = ~pi1041 & pi1049;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = n5318 & n5321;
  assign n5323 = ~n5318 & ~n5321;
  assign n5324 = ~n5322 & ~n5323;
  assign n5325 = n5315 & n5324;
  assign n5326 = ~n5315 & ~n5324;
  assign n5327 = ~n5325 & ~n5326;
  assign n5328 = n5312 & n5327;
  assign n5329 = ~n5312 & ~n5327;
  assign n5330 = ~n5328 & ~n5329;
  assign n5331 = pi1336 & n5330;
  assign n5332 = ~pi1336 & ~n5330;
  assign n5333 = ~n5331 & ~n5332;
  assign n5334 = ~pi1044 & ~pi1317;
  assign n5335 = pi1044 & pi1317;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = pi1017 & n5321;
  assign n5338 = ~pi1017 & ~n5321;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = ~n5318 & n5339;
  assign n5341 = n5318 & ~n5339;
  assign n5342 = ~n5340 & ~n5341;
  assign n5343 = n5336 & n5342;
  assign n5344 = ~n5336 & ~n5342;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = pi1335 & n5345;
  assign n5347 = ~pi1335 & ~n5345;
  assign n5348 = ~n5346 & ~n5347;
  assign n5349 = pi1044 & ~pi1318;
  assign n5350 = ~pi1044 & pi1318;
  assign n5351 = ~n5349 & ~n5350;
  assign n5352 = ~pi1042 & pi1043;
  assign n5353 = pi1042 & ~pi1043;
  assign n5354 = ~n5352 & ~n5353;
  assign n5355 = ~n5351 & n5354;
  assign n5356 = n5351 & ~n5354;
  assign n5357 = ~n5355 & ~n5356;
  assign n5358 = ~n5318 & ~n5357;
  assign n5359 = n5318 & n5357;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = pi1337 & n5360;
  assign n5362 = ~pi1337 & ~n5360;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = pi1043 & ~pi1049;
  assign n5365 = ~pi1043 & pi1049;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = pi1017 & ~pi1313;
  assign n5368 = ~pi1017 & pi1313;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = ~n5366 & n5369;
  assign n5371 = n5366 & ~n5369;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = ~n5318 & n5372;
  assign n5374 = n5318 & ~n5372;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = pi1334 & n5375;
  assign n5377 = ~pi1334 & ~n5375;
  assign n5378 = ~n5376 & ~n5377;
  assign n5379 = ~pi1039 & pi1041;
  assign n5380 = pi1039 & ~pi1041;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = pi1017 & ~pi1042;
  assign n5383 = ~pi1017 & pi1042;
  assign n5384 = ~n5382 & ~n5383;
  assign n5385 = ~n5381 & n5384;
  assign n5386 = n5381 & ~n5384;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = pi1317 & n5387;
  assign n5389 = ~pi1317 & ~n5387;
  assign n5390 = ~n5388 & ~n5389;
  assign n5391 = pi1285 & n5390;
  assign n5392 = ~pi1285 & ~n5390;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394 = n5378 & n5393;
  assign n5395 = ~n5363 & n5394;
  assign n5396 = ~n5348 & n5395;
  assign n5397 = ~n5333 & n5396;
  assign po1002 = pi1233 & ~n5397;
  assign n5399 = ~pi1017 & pi1098;
  assign n5400 = pi1017 & ~pi1098;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = n4134 & n5258;
  assign n5403 = n5229 & n5232;
  assign n5404 = ~n5402 & ~n5403;
  assign n5405 = ~n4118 & ~n5232;
  assign n5406 = n5258 & ~n5405;
  assign n5407 = ~n5259 & ~n5406;
  assign n5408 = n5404 & n5407;
  assign n5409 = ~pi1042 & pi1097;
  assign n5410 = pi1042 & ~pi1097;
  assign n5411 = ~n5409 & ~n5410;
  assign n5412 = n5408 & n5411;
  assign n5413 = n5401 & n5412;
  assign n5414 = ~po1002 & n5413;
  assign po0462 = n5309 & n5414;
  assign n5416 = pi1747 & ~po0462;
  assign n5417 = ~pi0067 & pi0088;
  assign n5418 = n5250 & n5417;
  assign n5419 = n5416 & ~n5418;
  assign n5420 = ~pi0382 & ~pi0695;
  assign n5421 = ~pi0696 & n5420;
  assign n5422 = pi0647 & n5421;
  assign n5423 = ~pi1626 & ~pi1627;
  assign po1526 = n5422 & ~n5423;
  assign n5425 = pi0727 & ~pi0731;
  assign n5426 = ~pi0732 & ~pi0744;
  assign n5427 = ~pi0730 & ~pi0737;
  assign n5428 = ~pi0723 & ~pi0738;
  assign n5429 = n5427 & n5428;
  assign n5430 = n5426 & n5429;
  assign n5431 = n5425 & n5430;
  assign n5432 = ~pi0722 & pi0729;
  assign n5433 = pi0733 & n5432;
  assign n5434 = pi0746 & n5433;
  assign n5435 = ~pi0736 & ~pi0745;
  assign n5436 = n5434 & n5435;
  assign n5437 = ~pi0734 & n5436;
  assign n5438 = ~pi0735 & n5437;
  assign n5439 = n5431 & n5438;
  assign n5440 = po1526 & ~n5439;
  assign n5441 = pi1416 & ~n5440;
  assign n5442 = ~pi0138 & n5441;
  assign n5443 = pi0067 & ~po1526;
  assign n5444 = n5442 & ~n5443;
  assign n5445 = ~pi0109 & n5280;
  assign n5446 = n5246 & n5445;
  assign n5447 = pi0089 & n5446;
  assign n5448 = ~pi0092 & n5447;
  assign n5449 = ~n5444 & n5448;
  assign n5450 = n5419 & ~n5449;
  assign n5451 = n5284 & n5450;
  assign po0178 = ~n5275 | ~n5451;
  assign n5453 = n4147 & ~n5238;
  assign n5454 = ~n4149 & ~n5231;
  assign n5455 = n5453 & n5454;
  assign po0232 = n5242 & n5455;
  assign n5457 = ~pi0121 & ~po0232;
  assign n5458 = pi0826 & n4173;
  assign n5459 = pi0849 & ~n4173;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = pi0827 & n4173;
  assign n5462 = pi0850 & ~n4173;
  assign n5463 = ~n5461 & ~n5462;
  assign n5464 = n5460 & n5463;
  assign n5465 = pi0877 & n5463;
  assign n5466 = ~n5464 & ~n5465;
  assign n5467 = pi0762 & n4173;
  assign n5468 = pi0749 & ~n4173;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = ~pi0852 & ~n4173;
  assign n5471 = ~pi0768 & n4173;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = n5469 & ~n5472;
  assign n5474 = ~n5466 & n5473;
  assign n5475 = pi0877 & n5460;
  assign n5476 = pi0772 & n4173;
  assign n5477 = pi0810 & ~n5476;
  assign n5478 = pi0748 & ~n4173;
  assign n5479 = n5477 & ~n5478;
  assign n5480 = pi0848 & ~n4173;
  assign n5481 = pi0825 & n4173;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = pi0759 & n5482;
  assign n5484 = ~n5479 & ~n5483;
  assign n5485 = ~n5475 & n5484;
  assign n5486 = pi0845 & ~n4173;
  assign n5487 = pi0822 & n4173;
  assign n5488 = ~n5486 & ~n5487;
  assign n5489 = pi0770 & n4173;
  assign n5490 = pi0751 & ~n4173;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = ~n5488 & ~n5491;
  assign n5493 = ~pi0807 & n5492;
  assign n5494 = ~pi0755 & ~n5488;
  assign n5495 = n4733 & ~n5491;
  assign n5496 = ~n5494 & ~n5495;
  assign n5497 = pi0755 & n5488;
  assign n5498 = pi0807 & ~n5489;
  assign n5499 = ~n5490 & n5498;
  assign n5500 = ~n5497 & ~n5499;
  assign n5501 = pi0844 & ~n4173;
  assign n5502 = pi0821 & n4173;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = ~pi0806 & ~n5503;
  assign n5505 = n5500 & n5504;
  assign n5506 = n5496 & ~n5505;
  assign n5507 = ~n5493 & n5506;
  assign n5508 = pi0806 & n5503;
  assign n5509 = n5500 & ~n5508;
  assign n5510 = pi0819 & n4173;
  assign n5511 = pi0842 & ~n4173;
  assign n5512 = ~n5510 & ~n5511;
  assign n5513 = ~pi0804 & ~n5512;
  assign n5514 = n5509 & n5513;
  assign n5515 = n5507 & ~n5514;
  assign n5516 = ~pi0806 & ~n5512;
  assign n5517 = ~pi0804 & ~n5503;
  assign n5518 = ~n5503 & ~n5512;
  assign n5519 = ~n4737 & ~n5518;
  assign n5520 = ~n5517 & n5519;
  assign n5521 = ~n5516 & n5520;
  assign n5522 = ~pi0841 & ~n4173;
  assign n5523 = ~pi0818 & n4173;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = n4754 & ~n5524;
  assign n5526 = pi0871 & n4173;
  assign n5527 = pi0754 & ~n4173;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = ~pi0750 & ~n5523;
  assign n5530 = ~n5522 & n5529;
  assign n5531 = n5528 & ~n5530;
  assign n5532 = ~n5525 & ~n5531;
  assign n5533 = ~n4757 & ~n5532;
  assign n5534 = ~n5521 & ~n5533;
  assign n5535 = n5500 & n5534;
  assign n5536 = n5515 & ~n5535;
  assign n5537 = pi0823 & n4173;
  assign n5538 = pi0846 & ~n4173;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = pi0824 & n4173;
  assign n5541 = pi0809 & ~n5540;
  assign n5542 = pi0847 & ~n4173;
  assign n5543 = n5541 & ~n5542;
  assign n5544 = ~n5539 & ~n5543;
  assign n5545 = ~n5540 & ~n5542;
  assign n5546 = ~pi0808 & ~n5545;
  assign n5547 = ~n4707 & ~n5546;
  assign n5548 = ~n5544 & n5547;
  assign n5549 = ~n5536 & ~n5548;
  assign n5550 = n5485 & n5549;
  assign n5551 = ~n5476 & ~n5478;
  assign n5552 = ~n5482 & ~n5551;
  assign n5553 = ~pi0810 & n5552;
  assign n5554 = ~pi0759 & ~n5482;
  assign n5555 = n4699 & ~n5551;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = ~n5553 & n5556;
  assign n5558 = ~pi0809 & ~n5545;
  assign n5559 = n5484 & n5558;
  assign n5560 = n5557 & ~n5559;
  assign n5561 = pi0809 & n5545;
  assign n5562 = n5484 & ~n5561;
  assign n5563 = ~pi0808 & ~n5539;
  assign n5564 = n5562 & n5563;
  assign n5565 = n5560 & ~n5564;
  assign n5566 = ~n5475 & ~n5565;
  assign n5567 = ~n5550 & ~n5566;
  assign n5568 = n5474 & n5567;
  assign n5569 = ~n5460 & n5568;
  assign n5570 = pi0877 & ~n5568;
  assign po0300 = n5569 | n5570;
  assign n5572 = ~n5457 & po0300;
  assign n5573 = ~pi0077 & ~pi0078;
  assign n5574 = ~pi0071 & ~pi0079;
  assign n5575 = n5573 & n5574;
  assign n5576 = ~pi0073 & ~pi0076;
  assign n5577 = n5575 & n5576;
  assign n5578 = ~pi0080 & ~pi0081;
  assign n5579 = ~pi0082 & ~pi0083;
  assign n5580 = n5578 & n5579;
  assign n5581 = n5577 & n5580;
  assign n5582 = pi0069 & ~n5581;
  assign n5583 = ~pi0069 & n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = pi1091 & pi1101;
  assign n5586 = ~pi0070 & ~pi0075;
  assign n5587 = ~pi0069 & ~pi0074;
  assign n5588 = n5586 & n5587;
  assign n5589 = n5580 & n5588;
  assign po1655 = n5577 & n5589;
  assign n5591 = n3955 & ~po1655;
  assign n5592 = ~n5585 & ~n5591;
  assign n5593 = ~n5584 & ~n5592;
  assign n5594 = pi0069 & n5592;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = n5457 & ~n5595;
  assign n5597 = ~n5572 & ~n5596;
  assign po0180 = ~pi1747 | ~n5597;
  assign po0302 = ~n5469 & n5568;
  assign n5600 = ~n5457 & po0302;
  assign n5601 = n5579 & n5587;
  assign n5602 = ~pi0077 & n5576;
  assign n5603 = ~pi0078 & n5602;
  assign n5604 = n5578 & n5603;
  assign n5605 = n5574 & n5604;
  assign n5606 = n5601 & n5605;
  assign n5607 = pi0070 & ~n5606;
  assign n5608 = ~pi0070 & n5606;
  assign n5609 = ~n5607 & ~n5608;
  assign n5610 = ~n5592 & ~n5609;
  assign n5611 = pi0070 & n5592;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = n5457 & ~n5612;
  assign n5614 = ~n5600 & ~n5613;
  assign po0181 = ~pi1747 | ~n5614;
  assign n5616 = ~n5491 & n5568;
  assign n5617 = pi0807 & ~n5568;
  assign po0299 = n5616 | n5617;
  assign n5619 = ~n5457 & po0299;
  assign n5620 = pi0071 & ~n5603;
  assign n5621 = ~pi0071 & n5603;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~n5592 & ~n5622;
  assign n5624 = pi0071 & n5592;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = n5457 & ~n5625;
  assign n5627 = ~n5619 & ~n5626;
  assign po0182 = ~pi1747 | ~n5627;
  assign n5629 = pi0072 & pi1747;
  assign n5630 = ~pi1839 & n5629;
  assign n5631 = ~pi1080 & pi1132;
  assign n5632 = pi1541 & n5631;
  assign n5633 = pi0072 & n5632;
  assign n5634 = pi0137 & pi1492;
  assign n5635 = pi0072 & n5634;
  assign n5636 = ~n5631 & n5635;
  assign n5637 = ~n5633 & ~n5636;
  assign n5638 = pi1747 & ~n5637;
  assign n5639 = ~n5630 & ~n5638;
  assign n5640 = ~pi0711 & pi1747;
  assign n5641 = ~pi1608 & n5640;
  assign po0184 = ~n5639 | n5641;
  assign n5643 = n5524 & n5568;
  assign n5644 = pi0859 & ~n5568;
  assign po0298 = n5643 | n5644;
  assign n5646 = ~n5457 & ~po0298;
  assign n5647 = pi0073 & ~n5592;
  assign n5648 = ~pi0073 & n5592;
  assign n5649 = ~n5647 & ~n5648;
  assign n5650 = n5457 & ~n5649;
  assign n5651 = ~n5646 & ~n5650;
  assign po0185 = ~pi1747 | n5651;
  assign po0301 = ~n5463 & n5568;
  assign n5654 = ~n5457 & ~po0301;
  assign n5655 = ~pi0069 & ~pi0083;
  assign n5656 = ~pi0081 & ~pi0082;
  assign n5657 = ~pi0078 & ~pi0080;
  assign n5658 = n5602 & n5657;
  assign n5659 = n5574 & n5658;
  assign n5660 = n5656 & n5659;
  assign n5661 = n5655 & n5660;
  assign n5662 = pi0074 & n5661;
  assign n5663 = ~pi0074 & ~n5661;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = ~n5592 & n5664;
  assign n5666 = pi0074 & n5592;
  assign n5667 = ~n5665 & ~n5666;
  assign n5668 = n5457 & n5667;
  assign n5669 = ~n5654 & ~n5668;
  assign po0186 = ~pi1747 | n5669;
  assign po0303 = n5472 & n5568;
  assign n5672 = ~n5457 & ~po0303;
  assign n5673 = ~pi0070 & ~pi0074;
  assign n5674 = ~pi0071 & ~pi0078;
  assign n5675 = n5602 & n5674;
  assign n5676 = ~pi0079 & n5675;
  assign n5677 = ~pi0082 & n5578;
  assign n5678 = n5676 & n5677;
  assign n5679 = n5673 & n5678;
  assign n5680 = n5655 & n5679;
  assign n5681 = pi0075 & n5680;
  assign n5682 = ~pi0075 & ~n5680;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = ~n5592 & n5683;
  assign n5685 = pi0075 & n5592;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = n5457 & n5686;
  assign n5688 = ~n5672 & ~n5687;
  assign po0187 = ~pi1747 | n5688;
  assign n5690 = pi0073 & pi0076;
  assign n5691 = ~n5576 & ~n5690;
  assign n5692 = ~n5592 & ~n5691;
  assign n5693 = pi0076 & n5592;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = n5457 & ~n5694;
  assign n5696 = ~n5528 & n5568;
  assign n5697 = pi0750 & ~n5568;
  assign po0259 = n5696 | n5697;
  assign n5699 = ~n5457 & po0259;
  assign n5700 = ~n5695 & ~n5699;
  assign po0188 = ~pi1747 | ~n5700;
  assign n5702 = n5512 & n5568;
  assign n5703 = ~pi0804 & ~n5568;
  assign po0261 = ~n5702 & ~n5703;
  assign n5705 = ~n5457 & ~po0261;
  assign n5706 = pi0077 & ~n5576;
  assign n5707 = ~n5602 & ~n5706;
  assign n5708 = ~n5592 & ~n5707;
  assign n5709 = pi0077 & n5592;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = n5457 & n5710;
  assign n5712 = ~n5705 & ~n5711;
  assign po0189 = ~pi1747 | n5712;
  assign n5714 = ~n5503 & n5568;
  assign n5715 = pi0806 & ~n5568;
  assign po0260 = n5714 | n5715;
  assign n5717 = ~n5457 & ~po0260;
  assign n5718 = pi0078 & ~n5602;
  assign n5719 = ~n5603 & ~n5718;
  assign n5720 = ~n5592 & ~n5719;
  assign n5721 = pi0078 & n5592;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = n5457 & n5722;
  assign n5724 = ~n5717 & ~n5723;
  assign po0190 = ~pi1747 | n5724;
  assign n5726 = ~n5488 & n5568;
  assign n5727 = pi0755 & ~n5568;
  assign po0262 = n5726 | n5727;
  assign n5729 = ~n5457 & ~po0262;
  assign n5730 = pi0079 & ~n5675;
  assign n5731 = ~n5676 & ~n5730;
  assign n5732 = ~n5592 & ~n5731;
  assign n5733 = pi0079 & n5592;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = n5457 & n5734;
  assign n5736 = ~n5729 & ~n5735;
  assign po0191 = ~pi1747 | n5736;
  assign n5738 = ~n5539 & n5568;
  assign n5739 = pi0808 & ~n5568;
  assign po0244 = n5738 | n5739;
  assign n5741 = ~n5457 & ~po0244;
  assign n5742 = pi0080 & n5577;
  assign n5743 = ~pi0080 & ~n5577;
  assign n5744 = ~n5742 & ~n5743;
  assign n5745 = ~n5592 & n5744;
  assign n5746 = pi0080 & n5592;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = n5457 & n5747;
  assign n5749 = ~n5741 & ~n5748;
  assign po0192 = ~pi1747 | n5749;
  assign n5751 = ~n5545 & n5568;
  assign n5752 = pi0809 & ~n5568;
  assign po0243 = n5751 | n5752;
  assign n5754 = ~n5457 & ~po0243;
  assign n5755 = pi0081 & n5659;
  assign n5756 = ~pi0081 & ~n5659;
  assign n5757 = ~n5755 & ~n5756;
  assign n5758 = ~n5592 & n5757;
  assign n5759 = pi0081 & n5592;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = n5457 & n5760;
  assign n5762 = ~n5754 & ~n5761;
  assign po0193 = ~pi1747 | n5762;
  assign n5764 = ~n5551 & n5568;
  assign n5765 = pi0810 & ~n5568;
  assign po0245 = n5764 | n5765;
  assign n5767 = ~n5457 & ~po0245;
  assign n5768 = pi0082 & n5605;
  assign n5769 = ~pi0082 & ~n5605;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~n5592 & n5770;
  assign n5772 = pi0082 & n5592;
  assign n5773 = ~n5771 & ~n5772;
  assign n5774 = n5457 & n5773;
  assign n5775 = ~n5767 & ~n5774;
  assign po0194 = ~pi1747 | n5775;
  assign n5777 = ~n5482 & n5568;
  assign n5778 = pi0759 & ~n5568;
  assign po0246 = n5777 | n5778;
  assign n5780 = ~n5457 & ~po0246;
  assign n5781 = pi0083 & n5678;
  assign n5782 = ~pi0083 & ~n5678;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = ~n5592 & n5783;
  assign n5785 = pi0083 & n5592;
  assign n5786 = ~n5784 & ~n5785;
  assign n5787 = n5457 & n5786;
  assign n5788 = ~n5780 & ~n5787;
  assign po0195 = ~pi1747 | n5788;
  assign n5790 = pi0084 & pi1747;
  assign n5791 = ~pi1840 & n5790;
  assign n5792 = ~pi1144 & pi1259;
  assign n5793 = pi1538 & n5792;
  assign n5794 = pi0084 & n5793;
  assign n5795 = pi0142 & pi1491;
  assign n5796 = pi0084 & n5795;
  assign n5797 = ~n5792 & n5796;
  assign n5798 = ~n5794 & ~n5797;
  assign n5799 = pi1747 & ~n5798;
  assign n5800 = ~n5791 & ~n5799;
  assign n5801 = ~pi0713 & pi1747;
  assign n5802 = ~pi1583 & n5801;
  assign po0196 = ~n5800 | n5802;
  assign n5804 = pi0085 & pi1747;
  assign n5805 = ~pi1838 & n5804;
  assign n5806 = ~pi1256 & pi1257;
  assign n5807 = pi1540 & n5806;
  assign n5808 = pi0085 & n5807;
  assign n5809 = pi0143 & pi1477;
  assign n5810 = pi0085 & n5809;
  assign n5811 = ~n5806 & n5810;
  assign n5812 = ~n5808 & ~n5811;
  assign n5813 = pi1747 & ~n5812;
  assign n5814 = ~n5805 & ~n5813;
  assign n5815 = ~pi0676 & pi1747;
  assign n5816 = ~pi1607 & n5815;
  assign po0197 = ~n5814 | n5816;
  assign n5818 = pi0123 & ~n5472;
  assign n5819 = ~pi0123 & n5472;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = ~pi0126 & n5463;
  assign n5822 = ~pi0127 & n5469;
  assign n5823 = ~n5821 & ~n5822;
  assign n5824 = ~pi0119 & n5460;
  assign n5825 = pi0101 & ~n5482;
  assign n5826 = ~n5824 & n5825;
  assign n5827 = pi0119 & ~n5460;
  assign n5828 = ~n5826 & ~n5827;
  assign n5829 = n5823 & ~n5828;
  assign n5830 = pi0126 & ~n5463;
  assign n5831 = ~pi0127 & ~n5830;
  assign n5832 = n5469 & ~n5830;
  assign n5833 = pi0127 & ~n5469;
  assign n5834 = n5822 & ~n5833;
  assign n5835 = ~n5832 & ~n5834;
  assign n5836 = ~n5831 & n5835;
  assign n5837 = ~n5829 & ~n5836;
  assign n5838 = ~pi0101 & n5482;
  assign n5839 = ~n5824 & ~n5838;
  assign n5840 = n5823 & n5839;
  assign n5841 = pi0100 & ~n5551;
  assign n5842 = ~pi0100 & n5551;
  assign n5843 = pi0099 & ~n5545;
  assign n5844 = ~n5842 & n5843;
  assign n5845 = ~n5841 & ~n5844;
  assign n5846 = ~pi0099 & n5545;
  assign n5847 = ~n5842 & ~n5846;
  assign n5848 = pi0098 & ~n5539;
  assign n5849 = ~pi0098 & n5539;
  assign n5850 = pi0107 & ~n5488;
  assign n5851 = ~n5849 & n5850;
  assign n5852 = ~n5848 & ~n5851;
  assign n5853 = n5847 & ~n5852;
  assign n5854 = n5845 & ~n5853;
  assign n5855 = ~pi0106 & n5503;
  assign n5856 = ~pi0117 & n5491;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = ~pi0103 & ~n5524;
  assign n5859 = ~pi0104 & n5528;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~pi0105 & n5512;
  assign n5862 = n5860 & ~n5861;
  assign n5863 = pi0105 & ~n5512;
  assign n5864 = pi0104 & ~n5528;
  assign n5865 = ~n5861 & n5864;
  assign n5866 = ~n5863 & ~n5865;
  assign n5867 = ~n5862 & n5866;
  assign n5868 = n5857 & ~n5867;
  assign n5869 = pi0117 & ~n5491;
  assign n5870 = pi0106 & ~n5503;
  assign n5871 = ~n5856 & n5870;
  assign n5872 = ~n5869 & ~n5871;
  assign n5873 = ~n5868 & n5872;
  assign n5874 = ~pi0107 & n5488;
  assign n5875 = ~n5849 & ~n5874;
  assign n5876 = n5847 & n5875;
  assign n5877 = ~n5873 & n5876;
  assign n5878 = n5854 & ~n5877;
  assign n5879 = n5840 & ~n5878;
  assign n5880 = n5837 & ~n5879;
  assign n5881 = ~n5820 & n5880;
  assign n5882 = n5820 & ~n5880;
  assign po0198 = n5881 | n5882;
  assign n5884 = pi0087 & pi1747;
  assign n5885 = ~pi1841 & n5884;
  assign n5886 = ~pi1112 & pi1113;
  assign n5887 = pi1539 & n5886;
  assign n5888 = pi0087 & n5887;
  assign n5889 = pi0184 & pi1520;
  assign n5890 = pi0087 & n5889;
  assign n5891 = ~n5886 & n5890;
  assign n5892 = ~n5888 & ~n5891;
  assign n5893 = pi1747 & ~n5892;
  assign n5894 = ~n5885 & ~n5893;
  assign n5895 = ~pi0721 & pi1747;
  assign n5896 = ~pi1604 & n5895;
  assign po0199 = ~n5894 | n5896;
  assign n5898 = ~pi0089 & pi0092;
  assign n5899 = n5446 & n5898;
  assign n5900 = pi1251 & n5899;
  assign n5901 = pi0088 & n5900;
  assign n5902 = pi0088 & n5239;
  assign n5903 = ~n4149 & ~n5902;
  assign n5904 = ~n5231 & n5903;
  assign n5905 = n4138 & ~n5904;
  assign n5906 = ~n4139 & ~n5905;
  assign n5907 = n5252 & ~n5906;
  assign n5908 = pi0088 & n5252;
  assign n5909 = ~n4138 & n5908;
  assign n5910 = ~n5907 & ~n5909;
  assign n5911 = ~n5901 & n5910;
  assign po0200 = n5416 & ~n5911;
  assign n5913 = n5442 & n5448;
  assign n5914 = pi0089 & n5913;
  assign n5915 = ~po1526 & n5914;
  assign n5916 = pi0089 & pi1251;
  assign n5917 = n5899 & n5916;
  assign n5918 = ~pi0089 & ~n4138;
  assign n5919 = ~pi0089 & n5236;
  assign n5920 = n5238 & n5454;
  assign n5921 = n4133 & n5920;
  assign n5922 = ~n5919 & n5921;
  assign n5923 = n4138 & ~n5922;
  assign n5924 = ~n5918 & ~n5923;
  assign n5925 = n5252 & n5924;
  assign n5926 = ~n5917 & ~n5925;
  assign n5927 = ~n5915 & n5926;
  assign po0201 = n5416 & ~n5927;
  assign n5929 = pi1001 & n5472;
  assign n5930 = ~pi1001 & ~n5472;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = pi1000 & n5469;
  assign n5933 = pi1013 & n5463;
  assign n5934 = pi1010 & n5551;
  assign n5935 = pi1009 & n5545;
  assign n5936 = pi1008 & n5539;
  assign n5937 = ~pi1007 & n5488;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = ~n5935 & n5938;
  assign n5940 = ~n5934 & n5939;
  assign n5941 = pi1006 & ~n5491;
  assign n5942 = ~pi1006 & n5491;
  assign n5943 = pi1005 & ~n5503;
  assign n5944 = ~n5942 & n5943;
  assign n5945 = ~n5941 & ~n5944;
  assign n5946 = pi0999 & ~n5512;
  assign n5947 = ~pi0999 & n5512;
  assign n5948 = pi0998 & ~n5528;
  assign n5949 = ~n5947 & n5948;
  assign n5950 = ~n5946 & ~n5949;
  assign n5951 = ~pi1005 & n5503;
  assign n5952 = ~n5942 & ~n5951;
  assign n5953 = ~n5950 & n5952;
  assign n5954 = pi0997 & n5524;
  assign n5955 = ~pi0998 & n5528;
  assign n5956 = n5954 & ~n5955;
  assign n5957 = n5952 & n5956;
  assign n5958 = ~n5947 & n5957;
  assign n5959 = ~n5953 & ~n5958;
  assign n5960 = n5945 & n5959;
  assign n5961 = n5940 & ~n5960;
  assign n5962 = ~pi1010 & ~n5551;
  assign n5963 = ~pi1009 & ~n5545;
  assign n5964 = ~n5934 & n5963;
  assign n5965 = ~n5962 & ~n5964;
  assign n5966 = ~pi1008 & ~n5539;
  assign n5967 = pi1007 & ~n5488;
  assign n5968 = ~n5936 & n5967;
  assign n5969 = ~n5966 & ~n5968;
  assign n5970 = ~n5934 & ~n5935;
  assign n5971 = ~n5969 & n5970;
  assign n5972 = n5965 & ~n5971;
  assign n5973 = ~n5961 & n5972;
  assign n5974 = ~pi1012 & n5460;
  assign n5975 = pi1011 & n5482;
  assign n5976 = ~n5974 & ~n5975;
  assign n5977 = ~n5973 & n5976;
  assign n5978 = ~n5933 & n5977;
  assign n5979 = ~n5932 & n5978;
  assign n5980 = ~pi1000 & ~n5469;
  assign n5981 = pi1012 & ~n5460;
  assign n5982 = ~pi1011 & ~n5482;
  assign n5983 = ~n5974 & n5982;
  assign n5984 = ~n5981 & ~n5983;
  assign n5985 = ~n5933 & ~n5984;
  assign n5986 = ~pi1013 & ~n5463;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = ~n5932 & ~n5987;
  assign n5989 = ~n5980 & ~n5988;
  assign n5990 = ~n5979 & n5989;
  assign n5991 = n5931 & n5990;
  assign n5992 = ~n5931 & ~n5990;
  assign po0202 = n5991 | n5992;
  assign n5994 = ~pi1001 & ~n5980;
  assign n5995 = ~n5472 & ~n5980;
  assign n5996 = ~n5929 & n5930;
  assign n5997 = ~n5995 & ~n5996;
  assign n5998 = ~n5994 & n5997;
  assign n5999 = ~n5930 & ~n5932;
  assign n6000 = ~n5933 & n5981;
  assign n6001 = ~n5986 & ~n6000;
  assign n6002 = n5999 & ~n6001;
  assign n6003 = ~n5998 & ~n6002;
  assign n6004 = ~n5933 & ~n5974;
  assign n6005 = n5999 & n6004;
  assign n6006 = n5962 & ~n5975;
  assign n6007 = ~n5982 & ~n6006;
  assign n6008 = ~n5935 & n5966;
  assign n6009 = ~n5963 & ~n6008;
  assign n6010 = ~n5934 & ~n5975;
  assign n6011 = ~n6009 & n6010;
  assign n6012 = n6007 & ~n6011;
  assign n6013 = ~n5935 & ~n5936;
  assign n6014 = n6010 & n6013;
  assign n6015 = ~n5937 & ~n5942;
  assign n6016 = ~n5943 & n5951;
  assign n6017 = n6015 & ~n6016;
  assign n6018 = ~n5948 & ~n5956;
  assign n6019 = ~n5947 & ~n6018;
  assign n6020 = ~n5943 & ~n5946;
  assign n6021 = ~n6019 & n6020;
  assign n6022 = n6017 & ~n6021;
  assign n6023 = ~n5937 & n5941;
  assign n6024 = ~n5967 & ~n6023;
  assign n6025 = ~n6022 & n6024;
  assign n6026 = n6014 & ~n6025;
  assign n6027 = n6012 & ~n6026;
  assign n6028 = n6005 & ~n6027;
  assign n6029 = n6003 & ~n6028;
  assign n6030 = pi1002 & ~n6029;
  assign n6031 = ~pi1002 & n6029;
  assign po0203 = n6030 | n6031;
  assign n6033 = pi0092 & n5900;
  assign n6034 = n4138 & n5454;
  assign n6035 = pi0092 & n5236;
  assign n6036 = n5238 & ~n6035;
  assign n6037 = n4133 & ~n6036;
  assign n6038 = n6034 & n6037;
  assign n6039 = pi0092 & ~n4138;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = n5252 & ~n6040;
  assign n6042 = ~n6033 & ~n6041;
  assign po0204 = n5416 & ~n6042;
  assign n6044 = ~pi0138 & n4152;
  assign n6045 = n4157 & n6044;
  assign n6046 = n4138 & n5231;
  assign n6047 = ~n4139 & ~n6046;
  assign n6048 = n4148 & ~n6047;
  assign n6049 = ~n6045 & ~n6048;
  assign po0205 = n4162 | ~n6049;
  assign n6051 = ~pi0806 & ~pi0808;
  assign n6052 = ~pi0750 & ~pi0804;
  assign n6053 = n4699 & n4733;
  assign n6054 = n6052 & n6053;
  assign n6055 = n6051 & n6054;
  assign n6056 = ~pi0859 & n6055;
  assign n6057 = ~n5238 & n6056;
  assign n6058 = ~pi0809 & n6057;
  assign n6059 = ~pi0877 & n6058;
  assign n6060 = n4133 & ~n5231;
  assign n6061 = ~n4149 & n6060;
  assign n6062 = n4138 & n6061;
  assign n6063 = n4147 & n6062;
  assign po0206 = n6059 & n6063;
  assign n6065 = pi0111 & n5277;
  assign n6066 = ~pi0112 & n6065;
  assign n6067 = n4165 & n5273;
  assign n6068 = ~n6066 & ~n6067;
  assign n6069 = pi0095 & pi1251;
  assign n6070 = pi0799 & ~pi0800;
  assign n6071 = ~pi1251 & n6070;
  assign n6072 = ~n6069 & ~n6071;
  assign n6073 = n5899 & ~n6072;
  assign n6074 = n6068 & ~n6073;
  assign n6075 = ~pi0095 & ~n5260;
  assign n6076 = n5267 & ~n6075;
  assign n6077 = ~pi1417 & n6076;
  assign n6078 = pi0095 & n5252;
  assign n6079 = ~n4138 & n6078;
  assign n6080 = ~n6077 & ~n6079;
  assign n6081 = n6074 & n6080;
  assign po0207 = n5416 & ~n6081;
  assign n6083 = ~n5236 & n5238;
  assign po0208 = n6063 & n6083;
  assign n6085 = ~n4182 & ~n4183;
  assign n6086 = po0244 & n6085;
  assign n6087 = ~n4228 & ~n6086;
  assign po0209 = n4227 | ~n6087;
  assign n6089 = po0243 & n6085;
  assign n6090 = ~n4213 & ~n6089;
  assign po0210 = n4212 | ~n6090;
  assign n6092 = po0245 & n6085;
  assign n6093 = ~n4220 & ~n6092;
  assign po0211 = n4219 | ~n6093;
  assign n6095 = po0246 & n6085;
  assign n6096 = ~n4196 & ~n6095;
  assign po0212 = n4200 | ~n6096;
  assign n6098 = ~n5974 & ~n5981;
  assign n6099 = n6027 & n6098;
  assign n6100 = ~n6027 & ~n6098;
  assign po0213 = n6099 | n6100;
  assign n6102 = ~n4183 & po0298;
  assign n6103 = ~n4268 & ~n6102;
  assign n6104 = ~n4182 & ~n6103;
  assign po0214 = n4266 | n6104;
  assign n6106 = ~n4183 & po0259;
  assign n6107 = ~n4274 & ~n6106;
  assign n6108 = ~n4182 & ~n6107;
  assign po0215 = n4273 | n6108;
  assign n6110 = ~n4183 & po0261;
  assign n6111 = ~n4245 & ~n6110;
  assign n6112 = ~n4182 & ~n6111;
  assign po0216 = n4244 | n6112;
  assign n6114 = ~n4183 & po0260;
  assign n6115 = ~n4258 & ~n6114;
  assign n6116 = ~n4182 & ~n6115;
  assign po0217 = n4262 | n6116;
  assign n6118 = ~n4183 & po0262;
  assign n6119 = ~n4235 & ~n6118;
  assign n6120 = ~n4182 & ~n6119;
  assign po0218 = n4234 | n6120;
  assign n6122 = ~n4138 & n5252;
  assign n6123 = pi0108 & n6122;
  assign n6124 = ~n5260 & n5267;
  assign n6125 = pi0108 & ~pi1417;
  assign n6126 = n6124 & n6125;
  assign n6127 = ~pi1251 & ~n6070;
  assign n6128 = pi0108 & pi1251;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = n5899 & ~n6129;
  assign n6131 = ~n6126 & ~n6130;
  assign n6132 = ~n6123 & n6131;
  assign po0219 = n5416 & ~n6132;
  assign n6134 = pi0109 & n6122;
  assign n6135 = po1526 & ~n6070;
  assign n6136 = pi0109 & ~po1526;
  assign n6137 = ~n6135 & ~n6136;
  assign n6138 = n5913 & ~n6137;
  assign n6139 = pi0109 & pi1251;
  assign n6140 = n5899 & n6139;
  assign n6141 = ~n6138 & ~n6140;
  assign n6142 = ~n6134 & n6141;
  assign po0220 = n5416 & ~n6142;
  assign n6144 = ~pi0138 & n5282;
  assign n6145 = pi0110 & n6122;
  assign n6146 = ~n6144 & ~n6145;
  assign po0221 = n5416 & ~n6146;
  assign n6148 = pi0111 & n6122;
  assign n6149 = ~pi0111 & ~po1526;
  assign n6150 = ~n6135 & ~n6149;
  assign n6151 = n5913 & n6150;
  assign n6152 = pi0111 & pi1251;
  assign n6153 = n5899 & n6152;
  assign n6154 = ~n6151 & ~n6153;
  assign n6155 = ~n6148 & n6154;
  assign po0222 = n5416 & ~n6155;
  assign n6157 = pi0112 & n6122;
  assign n6158 = n5264 & n5271;
  assign n6159 = pi0095 & n6158;
  assign n6160 = ~pi0110 & n6159;
  assign n6161 = ~n6157 & ~n6160;
  assign po0223 = n5416 & ~n6161;
  assign n6163 = ~n5932 & ~n5980;
  assign n6164 = n6013 & n6015;
  assign n6165 = n5946 & ~n5951;
  assign n6166 = ~n5943 & ~n6165;
  assign n6167 = ~n5951 & ~n6018;
  assign n6168 = ~n5947 & n6167;
  assign n6169 = n6166 & ~n6168;
  assign n6170 = n6004 & ~n6169;
  assign n6171 = n6164 & n6170;
  assign n6172 = n6010 & n6171;
  assign n6173 = n6013 & ~n6024;
  assign n6174 = n6009 & ~n6173;
  assign n6175 = n6010 & ~n6174;
  assign n6176 = n6007 & ~n6175;
  assign n6177 = n6004 & ~n6176;
  assign n6178 = n6001 & ~n6177;
  assign n6179 = ~n6172 & n6178;
  assign n6180 = n6163 & n6179;
  assign n6181 = ~n6163 & ~n6179;
  assign po0224 = n6180 | n6181;
  assign n6183 = pi0198 & pi1459;
  assign n6184 = ~pi0114 & ~n6183;
  assign n6185 = pi1439 & pi1747;
  assign po0225 = ~n6184 & n6185;
  assign n6187 = pi0198 & pi1480;
  assign n6188 = ~pi0115 & ~n6187;
  assign n6189 = pi1473 & pi1747;
  assign po0226 = ~n6188 & n6189;
  assign n6191 = pi0198 & pi1430;
  assign n6192 = ~pi0116 & ~n6191;
  assign n6193 = pi1440 & pi1747;
  assign po0227 = ~n6192 & n6193;
  assign n6195 = ~n4183 & po0299;
  assign n6196 = ~n4251 & ~n6195;
  assign n6197 = ~n4182 & ~n6196;
  assign po0228 = n4255 | n6197;
  assign n6199 = pi0198 & pi1447;
  assign n6200 = ~pi0118 & ~n6199;
  assign n6201 = pi1437 & pi1747;
  assign po0229 = ~n6200 & n6201;
  assign n6203 = ~n4183 & po0300;
  assign n6204 = ~n4190 & ~n6203;
  assign n6205 = ~n4182 & ~n6204;
  assign po0230 = n4189 | n6205;
  assign n6207 = ~n5975 & ~n5982;
  assign n6208 = n5973 & n6207;
  assign n6209 = ~n5973 & ~n6207;
  assign po0231 = n6208 | n6209;
  assign n6211 = ~n5933 & ~n5986;
  assign n6212 = n5938 & n5970;
  assign n6213 = ~n5947 & n5956;
  assign n6214 = n5950 & ~n6213;
  assign n6215 = n5976 & ~n6214;
  assign n6216 = n5952 & n6215;
  assign n6217 = n6212 & n6216;
  assign n6218 = n5938 & ~n5945;
  assign n6219 = n5969 & ~n6218;
  assign n6220 = n5970 & ~n6219;
  assign n6221 = n5965 & ~n6220;
  assign n6222 = n5976 & ~n6221;
  assign n6223 = n5984 & ~n6222;
  assign n6224 = ~n6217 & n6223;
  assign n6225 = n6211 & n6224;
  assign n6226 = ~n6211 & ~n6224;
  assign po0233 = n6225 | n6226;
  assign n6228 = ~n4183 & po0303;
  assign po0234 = ~n4182 & n6228;
  assign n6230 = ~pi0218 & ~pi1099;
  assign n6231 = pi0236 & pi1099;
  assign po0235 = n6230 | n6231;
  assign n6233 = ~pi1148 & ~pi1317;
  assign n6234 = pi1148 & pi1317;
  assign n6235 = ~n6233 & ~n6234;
  assign n6236 = ~pi1253 & ~pi1313;
  assign n6237 = pi1253 & pi1313;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = ~pi1044 & ~pi1146;
  assign n6240 = pi1044 & pi1146;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = ~pi1147 & ~pi1318;
  assign n6243 = pi1147 & pi1318;
  assign n6244 = ~n6242 & ~n6243;
  assign n6245 = ~n6241 & ~n6244;
  assign n6246 = ~n6238 & n6245;
  assign po1567 = ~n6235 & n6246;
  assign n6248 = ~pi1116 & ~pi1313;
  assign n6249 = pi1116 & pi1313;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~pi1117 & ~pi1317;
  assign n6252 = pi1117 & pi1317;
  assign n6253 = ~n6251 & ~n6252;
  assign n6254 = ~pi1044 & ~pi1115;
  assign n6255 = pi1044 & pi1115;
  assign n6256 = ~n6254 & ~n6255;
  assign n6257 = ~pi1070 & ~pi1318;
  assign n6258 = pi1070 & pi1318;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = ~n6256 & ~n6259;
  assign n6261 = ~n6253 & n6260;
  assign po1588 = ~n6250 & n6261;
  assign n6263 = ~pi1262 & ~pi1318;
  assign n6264 = pi1262 & pi1318;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = ~pi1260 & ~pi1313;
  assign n6267 = pi1260 & pi1313;
  assign n6268 = ~n6266 & ~n6267;
  assign n6269 = ~pi1026 & ~pi1044;
  assign n6270 = pi1026 & pi1044;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = ~pi1123 & ~pi1317;
  assign n6273 = pi1123 & pi1317;
  assign n6274 = ~n6272 & ~n6273;
  assign n6275 = ~n6271 & ~n6274;
  assign n6276 = ~n6268 & n6275;
  assign po1538 = ~n6265 & n6276;
  assign n6278 = ~pi1135 & ~pi1317;
  assign n6279 = pi1135 & pi1317;
  assign n6280 = ~n6278 & ~n6279;
  assign n6281 = ~pi1134 & ~pi1313;
  assign n6282 = pi1134 & pi1313;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = ~pi1044 & ~pi1054;
  assign n6285 = pi1044 & pi1054;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~pi1136 & ~pi1318;
  assign n6288 = pi1136 & pi1318;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~n6286 & ~n6289;
  assign n6291 = ~n6283 & n6290;
  assign po1555 = ~n6280 & n6291;
  assign n6293 = ~po1538 & ~po1555;
  assign n6294 = ~po1588 & n6293;
  assign po1343 = po1567 | ~n6294;
  assign n6296 = pi0125 & ~po1343;
  assign n6297 = pi0264 & po1538;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = po1567 & n6293;
  assign n6300 = ~pi0265 & n6299;
  assign n6301 = po1588 & n6293;
  assign n6302 = ~po1567 & n6301;
  assign n6303 = pi0266 & n6302;
  assign n6304 = ~n6300 & ~n6303;
  assign n6305 = ~po1538 & po1555;
  assign n6306 = pi0249 & n6305;
  assign n6307 = n6304 & ~n6306;
  assign po0236 = ~n6298 | ~n6307;
  assign n6309 = ~n4183 & po0301;
  assign po0237 = ~n4182 & n6309;
  assign n6311 = ~n4183 & po0302;
  assign po0238 = ~n4182 & n6311;
  assign n6313 = pi0259 & pi1459;
  assign n6314 = ~pi0128 & ~n6313;
  assign po0239 = n6185 & ~n6314;
  assign n6316 = pi0259 & pi1480;
  assign n6317 = ~pi0129 & ~n6316;
  assign po0240 = n6189 & ~n6317;
  assign n6319 = pi0259 & pi1430;
  assign n6320 = ~pi0130 & ~n6319;
  assign po0241 = n6193 & ~n6320;
  assign n6322 = pi0259 & pi1447;
  assign n6323 = ~pi0131 & ~n6322;
  assign po0242 = n6201 & ~n6323;
  assign n6325 = pi1424 & pi1747;
  assign n6326 = ~pi0136 & pi0222;
  assign po0247 = n6325 & ~n6326;
  assign n6328 = pi0618 & pi1637;
  assign n6329 = ~pi0506 & ~pi1678;
  assign n6330 = ~pi0618 & ~pi1637;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = ~n6328 & ~n6331;
  assign n6333 = pi0587 & pi0622;
  assign n6334 = pi1482 & pi1489;
  assign n6335 = pi0622 & pi1489;
  assign n6336 = pi0587 & pi1482;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~n6334 & n6337;
  assign n6339 = ~n6333 & n6338;
  assign n6340 = ~n6332 & ~n6339;
  assign n6341 = pi1489 & n6333;
  assign n6342 = pi0587 & n6334;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = pi0622 & pi1482;
  assign n6345 = pi0483 & pi0485;
  assign n6346 = pi1454 & pi1490;
  assign n6347 = pi0485 & pi1454;
  assign n6348 = pi0483 & pi1490;
  assign n6349 = ~n6347 & ~n6348;
  assign n6350 = ~n6346 & n6349;
  assign n6351 = ~n6345 & n6350;
  assign n6352 = pi1513 & ~n6351;
  assign n6353 = pi0549 & n6352;
  assign n6354 = pi0549 & pi0567;
  assign n6355 = pi0567 & pi1513;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = pi1488 & ~n6356;
  assign n6358 = ~n6351 & n6357;
  assign n6359 = pi1490 & n6345;
  assign n6360 = pi0485 & n6346;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = pi0468 & pi0562;
  assign n6363 = pi0562 & pi1421;
  assign n6364 = pi0468 & pi1456;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = pi1421 & pi1456;
  assign n6367 = n6365 & ~n6366;
  assign n6368 = ~n6362 & n6367;
  assign n6369 = pi1468 & ~n6368;
  assign n6370 = pi0380 & n6369;
  assign n6371 = pi0380 & pi0533;
  assign n6372 = pi0533 & pi1468;
  assign n6373 = ~n6371 & ~n6372;
  assign n6374 = pi1455 & ~n6373;
  assign n6375 = ~n6368 & n6374;
  assign n6376 = pi1456 & n6362;
  assign n6377 = pi0562 & n6366;
  assign n6378 = ~n6376 & ~n6377;
  assign n6379 = pi0468 & pi1421;
  assign n6380 = n6378 & ~n6379;
  assign n6381 = ~n6375 & n6380;
  assign n6382 = ~n6370 & n6381;
  assign n6383 = pi0483 & pi1454;
  assign n6384 = n6382 & ~n6383;
  assign n6385 = n6361 & n6384;
  assign n6386 = ~n6358 & n6385;
  assign n6387 = ~n6353 & n6386;
  assign n6388 = ~pi0380 & ~pi1468;
  assign n6389 = pi1455 & ~n6388;
  assign n6390 = ~n6371 & ~n6389;
  assign n6391 = ~n6372 & n6390;
  assign n6392 = ~n6368 & ~n6391;
  assign n6393 = n6382 & ~n6392;
  assign n6394 = ~n6387 & ~n6393;
  assign n6395 = ~n6344 & ~n6394;
  assign n6396 = n6343 & n6395;
  assign n6397 = ~n6340 & n6396;
  assign n6398 = ~pi0549 & ~pi1513;
  assign n6399 = pi1488 & ~n6398;
  assign n6400 = n6356 & ~n6399;
  assign n6401 = ~n6351 & ~n6368;
  assign n6402 = ~n6391 & n6401;
  assign n6403 = ~n6400 & n6402;
  assign n6404 = ~n6394 & ~n6403;
  assign po0248 = n6397 | n6404;
  assign n6406 = ~pi0092 & n4143;
  assign n6407 = n4144 & n5251;
  assign n6408 = n6406 & n6407;
  assign n6409 = ~pi0109 & n6408;
  assign n6410 = po0462 & ~n6409;
  assign n6411 = pi0352 & pi0725;
  assign n6412 = ~n6410 & ~n6411;
  assign po0249 = ~pi0244 | ~n6412;
  assign n6414 = ~n5934 & ~n5962;
  assign n6415 = n6164 & ~n6169;
  assign n6416 = n6174 & ~n6415;
  assign n6417 = ~n6414 & ~n6416;
  assign n6418 = n6414 & n6416;
  assign po0250 = n6417 | n6418;
  assign n6420 = ~n5936 & ~n5966;
  assign n6421 = ~n6025 & ~n6420;
  assign n6422 = n6025 & n6420;
  assign po0251 = n6421 | n6422;
  assign n6424 = pi0213 & ~pi0261;
  assign n6425 = pi0141 & pi0261;
  assign po0252 = n6424 | n6425;
  assign n6427 = pi0662 & pi1567;
  assign n6428 = ~pi0586 & ~pi1703;
  assign n6429 = ~pi0662 & ~pi1567;
  assign n6430 = ~n6428 & ~n6429;
  assign n6431 = ~n6427 & ~n6430;
  assign n6432 = pi0653 & pi0654;
  assign n6433 = pi1525 & pi1536;
  assign n6434 = pi0654 & pi1536;
  assign n6435 = pi0653 & pi1525;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = ~n6433 & n6436;
  assign n6438 = ~n6432 & n6437;
  assign n6439 = ~n6431 & ~n6438;
  assign n6440 = pi1536 & n6432;
  assign n6441 = pi0653 & n6433;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = pi0654 & pi1525;
  assign n6444 = pi0566 & pi0569;
  assign n6445 = pi1475 & pi1484;
  assign n6446 = pi0569 & pi1484;
  assign n6447 = pi0566 & pi1475;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = ~n6445 & n6448;
  assign n6450 = ~n6444 & n6449;
  assign n6451 = pi1515 & ~n6450;
  assign n6452 = pi0648 & n6451;
  assign n6453 = pi0648 & pi0650;
  assign n6454 = pi0650 & pi1515;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = pi1535 & ~n6455;
  assign n6457 = ~n6450 & n6456;
  assign n6458 = pi1475 & n6444;
  assign n6459 = pi0569 & n6445;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = pi0621 & pi0645;
  assign n6462 = pi0645 & pi1449;
  assign n6463 = pi0621 & pi1441;
  assign n6464 = ~n6462 & ~n6463;
  assign n6465 = pi1441 & pi1449;
  assign n6466 = n6464 & ~n6465;
  assign n6467 = ~n6461 & n6466;
  assign n6468 = pi1436 & ~n6467;
  assign n6469 = pi0358 & n6468;
  assign n6470 = pi0358 & pi0623;
  assign n6471 = pi0623 & pi1436;
  assign n6472 = ~n6470 & ~n6471;
  assign n6473 = pi1486 & ~n6472;
  assign n6474 = ~n6467 & n6473;
  assign n6475 = pi1441 & n6461;
  assign n6476 = pi0645 & n6465;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = pi0621 & pi1449;
  assign n6479 = n6477 & ~n6478;
  assign n6480 = ~n6474 & n6479;
  assign n6481 = ~n6469 & n6480;
  assign n6482 = pi0566 & pi1484;
  assign n6483 = n6481 & ~n6482;
  assign n6484 = n6460 & n6483;
  assign n6485 = ~n6457 & n6484;
  assign n6486 = ~n6452 & n6485;
  assign n6487 = ~pi0358 & ~pi1436;
  assign n6488 = pi1486 & ~n6487;
  assign n6489 = ~n6470 & ~n6488;
  assign n6490 = ~n6471 & n6489;
  assign n6491 = ~n6467 & ~n6490;
  assign n6492 = n6481 & ~n6491;
  assign n6493 = ~n6486 & ~n6492;
  assign n6494 = ~n6443 & ~n6493;
  assign n6495 = n6442 & n6494;
  assign n6496 = ~n6439 & n6495;
  assign n6497 = ~pi0648 & ~pi1515;
  assign n6498 = pi1535 & ~n6497;
  assign n6499 = n6455 & ~n6498;
  assign n6500 = ~n6450 & ~n6467;
  assign n6501 = ~n6490 & n6500;
  assign n6502 = ~n6499 & n6501;
  assign n6503 = ~n6493 & ~n6502;
  assign po0253 = n6496 | n6503;
  assign n6505 = pi0507 & pi1565;
  assign n6506 = ~pi0408 & ~pi1702;
  assign n6507 = ~pi0507 & ~pi1565;
  assign n6508 = ~n6506 & ~n6507;
  assign n6509 = ~n6505 & ~n6508;
  assign n6510 = pi0508 & pi0509;
  assign n6511 = pi1497 & pi1509;
  assign n6512 = pi0509 & pi1509;
  assign n6513 = pi0508 & pi1497;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = ~n6511 & n6514;
  assign n6516 = ~n6510 & n6515;
  assign n6517 = ~n6509 & ~n6516;
  assign n6518 = pi1509 & n6510;
  assign n6519 = pi0508 & n6511;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = pi0509 & pi1497;
  assign n6522 = pi0386 & pi0387;
  assign n6523 = pi1461 & pi1474;
  assign n6524 = pi0387 & pi1461;
  assign n6525 = pi0386 & pi1474;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = ~n6523 & n6526;
  assign n6528 = ~n6522 & n6527;
  assign n6529 = pi1512 & ~n6528;
  assign n6530 = pi0480 & n6529;
  assign n6531 = pi0480 & pi0484;
  assign n6532 = pi0484 & pi1512;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = pi1507 & ~n6533;
  assign n6535 = ~n6528 & n6534;
  assign n6536 = pi1474 & n6522;
  assign n6537 = pi0387 & n6523;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = pi0381 & pi0470;
  assign n6540 = pi0470 & pi1434;
  assign n6541 = pi0381 & pi1438;
  assign n6542 = ~n6540 & ~n6541;
  assign n6543 = pi1434 & pi1438;
  assign n6544 = n6542 & ~n6543;
  assign n6545 = ~n6539 & n6544;
  assign n6546 = pi1435 & ~n6545;
  assign n6547 = pi0379 & n6546;
  assign n6548 = pi0379 & pi0466;
  assign n6549 = pi0466 & pi1435;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = pi1462 & ~n6550;
  assign n6552 = ~n6545 & n6551;
  assign n6553 = pi1438 & n6539;
  assign n6554 = pi0470 & n6543;
  assign n6555 = ~n6553 & ~n6554;
  assign n6556 = pi0381 & pi1434;
  assign n6557 = n6555 & ~n6556;
  assign n6558 = ~n6552 & n6557;
  assign n6559 = ~n6547 & n6558;
  assign n6560 = pi0386 & pi1461;
  assign n6561 = n6559 & ~n6560;
  assign n6562 = n6538 & n6561;
  assign n6563 = ~n6535 & n6562;
  assign n6564 = ~n6530 & n6563;
  assign n6565 = ~pi0379 & ~pi1435;
  assign n6566 = pi1462 & ~n6565;
  assign n6567 = ~n6548 & ~n6566;
  assign n6568 = ~n6549 & n6567;
  assign n6569 = ~n6545 & ~n6568;
  assign n6570 = n6559 & ~n6569;
  assign n6571 = ~n6564 & ~n6570;
  assign n6572 = ~n6521 & ~n6571;
  assign n6573 = n6520 & n6572;
  assign n6574 = ~n6517 & n6573;
  assign n6575 = ~pi0480 & ~pi1512;
  assign n6576 = pi1507 & ~n6575;
  assign n6577 = n6533 & ~n6576;
  assign n6578 = ~n6528 & ~n6545;
  assign n6579 = ~n6568 & n6578;
  assign n6580 = ~n6577 & n6579;
  assign n6581 = ~n6571 & ~n6580;
  assign po0254 = n6574 | n6581;
  assign n6583 = pi0232 & ~pi0261;
  assign n6584 = pi0144 & pi0261;
  assign po0255 = n6583 | n6584;
  assign n6586 = pi0211 & ~pi0261;
  assign n6587 = pi0145 & pi0261;
  assign po0256 = n6586 | n6587;
  assign n6589 = pi0230 & ~pi0261;
  assign n6590 = pi0146 & pi0261;
  assign po0257 = n6589 | n6590;
  assign n6592 = pi0220 & ~pi0261;
  assign n6593 = pi0147 & pi0261;
  assign po0258 = n6592 | n6593;
  assign n6595 = pi0997 & ~n4820;
  assign n6596 = n3953 & n4820;
  assign n6597 = ~n6595 & ~n6596;
  assign po0263 = pi1747 & ~n6597;
  assign n6599 = pi0429 & ~pi0706;
  assign n6600 = pi1747 & ~n6599;
  assign n6601 = pi0153 & pi0429;
  assign n6602 = ~pi0153 & pi0186;
  assign n6603 = pi0153 & ~pi0186;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = ~pi0429 & ~n6604;
  assign n6606 = ~n6601 & ~n6605;
  assign po0264 = n6600 & ~n6606;
  assign n6608 = ~pi0353 & ~pi1099;
  assign n6609 = pi0224 & pi1099;
  assign po0265 = n6608 | n6609;
  assign n6611 = pi0243 & pi1099;
  assign n6612 = ~pi0280 & ~pi1099;
  assign po0266 = n6611 | n6612;
  assign n6614 = pi0229 & ~pi0261;
  assign n6615 = pi0156 & pi0261;
  assign po0267 = n6614 | n6615;
  assign n6617 = pi0201 & ~pi0261;
  assign n6618 = pi0157 & pi0261;
  assign po0268 = n6617 | n6618;
  assign n6620 = pi0197 & ~pi0261;
  assign n6621 = pi0158 & pi0261;
  assign po0269 = n6620 | n6621;
  assign n6623 = pi0202 & ~pi0261;
  assign n6624 = pi0159 & pi0261;
  assign po0270 = n6623 | n6624;
  assign n6626 = pi0203 & ~pi0261;
  assign n6627 = pi0160 & pi0261;
  assign po0271 = n6626 | n6627;
  assign n6629 = pi0204 & ~pi0261;
  assign n6630 = pi0161 & pi0261;
  assign po0272 = n6629 | n6630;
  assign n6632 = pi0205 & ~pi0261;
  assign n6633 = pi0162 & pi0261;
  assign po0273 = n6632 | n6633;
  assign n6635 = pi0206 & ~pi0261;
  assign n6636 = pi0163 & pi0261;
  assign po0274 = n6635 | n6636;
  assign n6638 = pi0225 & ~pi0261;
  assign n6639 = pi0164 & pi0261;
  assign po0275 = n6638 | n6639;
  assign n6641 = pi0219 & ~pi0261;
  assign n6642 = pi0165 & pi0261;
  assign po0276 = n6641 | n6642;
  assign n6644 = pi0226 & ~pi0261;
  assign n6645 = pi0166 & pi0261;
  assign po0277 = n6644 | n6645;
  assign n6647 = pi0227 & ~pi0261;
  assign n6648 = pi0167 & pi0261;
  assign po0278 = n6647 | n6648;
  assign n6650 = pi0246 & ~pi0261;
  assign n6651 = pi0168 & pi0261;
  assign po0279 = n6650 | n6651;
  assign n6653 = pi0207 & ~pi0261;
  assign n6654 = pi0169 & pi0261;
  assign po0280 = n6653 | n6654;
  assign n6656 = pi0209 & ~pi0261;
  assign n6657 = pi0170 & pi0261;
  assign po0281 = n6656 | n6657;
  assign n6659 = pi0208 & ~pi0261;
  assign n6660 = pi0171 & pi0261;
  assign po0282 = n6659 | n6660;
  assign n6662 = pi0210 & ~pi0261;
  assign n6663 = pi0172 & pi0261;
  assign po0283 = n6662 | n6663;
  assign n6665 = pi0217 & ~pi0261;
  assign n6666 = pi0173 & pi0261;
  assign po0284 = n6665 | n6666;
  assign n6668 = pi0212 & ~pi0261;
  assign n6669 = pi0174 & pi0261;
  assign po0285 = n6668 | n6669;
  assign n6671 = pi0247 & ~pi0261;
  assign n6672 = pi0175 & pi0261;
  assign po0286 = n6671 | n6672;
  assign n6674 = pi0214 & ~pi0261;
  assign n6675 = pi0176 & pi0261;
  assign po0287 = n6674 | n6675;
  assign n6677 = pi0235 & ~pi0261;
  assign n6678 = pi0177 & pi0261;
  assign po0288 = n6677 | n6678;
  assign n6680 = pi0231 & ~pi0261;
  assign n6681 = pi0178 & pi0261;
  assign po0289 = n6680 | n6681;
  assign n6683 = pi0233 & ~pi0261;
  assign n6684 = pi0179 & pi0261;
  assign po0290 = n6683 | n6684;
  assign n6686 = pi0234 & ~pi0261;
  assign n6687 = pi0180 & pi0261;
  assign po0291 = n6686 | n6687;
  assign n6689 = pi0248 & ~pi0261;
  assign n6690 = pi0181 & pi0261;
  assign po0292 = n6689 | n6690;
  assign n6692 = pi0228 & ~pi0261;
  assign n6693 = pi0182 & pi0261;
  assign po0293 = n6692 | n6693;
  assign n6695 = pi0284 & pi0306;
  assign n6696 = ~pi0916 & pi1046;
  assign n6697 = ~pi1677 & n6696;
  assign po1775 = pi0984 | pi1045;
  assign n6699 = ~pi0954 & ~pi1050;
  assign n6700 = ~po1775 & n6699;
  assign n6701 = ~pi0760 & ~pi1021;
  assign n6702 = ~pi0773 & ~pi0937;
  assign n6703 = n6701 & n6702;
  assign n6704 = ~pi0971 & ~pi0995;
  assign n6705 = ~pi0966 & ~pi1019;
  assign n6706 = n6704 & n6705;
  assign n6707 = n6703 & n6706;
  assign n6708 = n6700 & n6707;
  assign n6709 = n6697 & n6708;
  assign n6710 = pi0954 & ~pi1050;
  assign n6711 = ~pi0916 & ~pi1046;
  assign n6712 = ~pi1677 & n6711;
  assign n6713 = n6703 & n6712;
  assign n6714 = ~po1775 & n6713;
  assign n6715 = n6706 & n6714;
  assign n6716 = n6710 & n6715;
  assign n6717 = n6700 & n6713;
  assign n6718 = pi0971 & ~pi0995;
  assign n6719 = n6717 & n6718;
  assign n6720 = n6705 & n6719;
  assign n6721 = ~n6716 & ~n6720;
  assign n6722 = ~n6709 & n6721;
  assign n6723 = ~pi0966 & pi1019;
  assign n6724 = n6700 & n6723;
  assign n6725 = n6713 & n6724;
  assign n6726 = n6704 & n6725;
  assign n6727 = pi0966 & ~pi1019;
  assign n6728 = n6704 & n6713;
  assign n6729 = n6700 & n6728;
  assign n6730 = n6727 & n6729;
  assign n6731 = ~n6716 & ~n6730;
  assign n6732 = ~n6726 & n6731;
  assign n6733 = pi0916 & ~pi1046;
  assign n6734 = n6708 & n6733;
  assign n6735 = ~pi1677 & n6734;
  assign n6736 = ~n6726 & ~n6735;
  assign n6737 = ~n6720 & n6736;
  assign n6738 = pi0785 & pi1479;
  assign n6739 = pi0785 & ~pi1479;
  assign n6740 = n6738 & ~n6739;
  assign n6741 = pi0960 & ~pi1345;
  assign n6742 = ~pi1479 & n6741;
  assign n6743 = pi0724 & n6742;
  assign n6744 = ~n6740 & ~n6743;
  assign n6745 = ~n6737 & ~n6744;
  assign n6746 = n6732 & n6745;
  assign n6747 = ~n6732 & ~n6737;
  assign n6748 = pi0262 & n6747;
  assign n6749 = ~n6746 & ~n6748;
  assign n6750 = n6722 & ~n6749;
  assign n6751 = ~n6722 & ~n6737;
  assign po1737 = pi1737 & ~pi1739;
  assign n6753 = pi1629 & po1737;
  assign n6754 = pi0724 & n6753;
  assign n6755 = n6751 & n6754;
  assign n6756 = n6732 & n6755;
  assign n6757 = ~n6750 & ~n6756;
  assign n6758 = ~n6722 & n6737;
  assign n6759 = pi0276 & n6753;
  assign n6760 = n6732 & n6759;
  assign n6761 = n6758 & n6760;
  assign n6762 = n6722 & n6737;
  assign n6763 = ~n6751 & ~n6762;
  assign n6764 = pi1677 & n6711;
  assign n6765 = n6708 & n6764;
  assign n6766 = ~n6730 & n6737;
  assign n6767 = ~n6716 & n6766;
  assign n6768 = ~n6765 & n6767;
  assign n6769 = ~n6709 & n6768;
  assign n6770 = ~n6732 & n6737;
  assign n6771 = n6732 & ~n6737;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~n6769 & n6772;
  assign n6774 = ~n6763 & n6773;
  assign n6775 = ~n6761 & ~n6774;
  assign n6776 = pi0277 & n6758;
  assign n6777 = po1737 & n6762;
  assign n6778 = ~n6776 & ~n6777;
  assign n6779 = ~n6732 & ~n6778;
  assign n6780 = n6775 & ~n6779;
  assign n6781 = n6757 & n6780;
  assign n6782 = ~pi0300 & ~pi0302;
  assign n6783 = n6781 & n6782;
  assign n6784 = pi0303 & n6783;
  assign n6785 = n6695 & n6784;
  assign n6786 = ~pi0301 & n6785;
  assign n6787 = ~pi0304 & n6786;
  assign po0294 = ~pi0305 & n6787;
  assign n6789 = pi0718 & pi1566;
  assign n6790 = ~pi0697 & ~pi1704;
  assign n6791 = ~pi0718 & ~pi1566;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = ~n6789 & ~n6792;
  assign n6794 = pi0708 & pi0719;
  assign n6795 = pi1524 & pi1545;
  assign n6796 = pi0708 & pi1545;
  assign n6797 = pi0719 & pi1524;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = ~n6795 & n6798;
  assign n6800 = ~n6794 & n6799;
  assign n6801 = ~n6793 & ~n6800;
  assign n6802 = pi1545 & n6794;
  assign n6803 = pi0719 & n6795;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = pi0708 & pi1524;
  assign n6806 = pi0675 & pi0678;
  assign n6807 = pi1483 & pi1514;
  assign n6808 = pi0678 & pi1483;
  assign n6809 = pi0675 & pi1514;
  assign n6810 = ~n6808 & ~n6809;
  assign n6811 = ~n6807 & n6810;
  assign n6812 = ~n6806 & n6811;
  assign n6813 = pi1537 & ~n6812;
  assign n6814 = pi0714 & n6813;
  assign n6815 = pi0714 & pi0717;
  assign n6816 = pi0717 & pi1537;
  assign n6817 = ~n6815 & ~n6816;
  assign n6818 = pi1533 & ~n6817;
  assign n6819 = ~n6812 & n6818;
  assign n6820 = pi1514 & n6806;
  assign n6821 = pi0678 & n6807;
  assign n6822 = ~n6820 & ~n6821;
  assign n6823 = pi0664 & pi0665;
  assign n6824 = pi0664 & pi1448;
  assign n6825 = pi0665 & pi1469;
  assign n6826 = ~n6824 & ~n6825;
  assign n6827 = pi1448 & pi1469;
  assign n6828 = n6826 & ~n6827;
  assign n6829 = ~n6823 & n6828;
  assign n6830 = pi1467 & ~n6829;
  assign n6831 = pi0359 & n6830;
  assign n6832 = pi0359 & pi0712;
  assign n6833 = pi0712 & pi1467;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = pi1485 & ~n6834;
  assign n6836 = ~n6829 & n6835;
  assign n6837 = pi1469 & n6823;
  assign n6838 = pi0664 & n6827;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = pi0665 & pi1448;
  assign n6841 = n6839 & ~n6840;
  assign n6842 = ~n6836 & n6841;
  assign n6843 = ~n6831 & n6842;
  assign n6844 = pi0675 & pi1483;
  assign n6845 = n6843 & ~n6844;
  assign n6846 = n6822 & n6845;
  assign n6847 = ~n6819 & n6846;
  assign n6848 = ~n6814 & n6847;
  assign n6849 = ~pi0359 & ~pi1467;
  assign n6850 = pi1485 & ~n6849;
  assign n6851 = ~n6832 & ~n6850;
  assign n6852 = ~n6833 & n6851;
  assign n6853 = ~n6829 & ~n6852;
  assign n6854 = n6843 & ~n6853;
  assign n6855 = ~n6848 & ~n6854;
  assign n6856 = ~n6805 & ~n6855;
  assign n6857 = n6804 & n6856;
  assign n6858 = ~n6801 & n6857;
  assign n6859 = ~pi0714 & ~pi1537;
  assign n6860 = pi1533 & ~n6859;
  assign n6861 = n6817 & ~n6860;
  assign n6862 = ~n6812 & ~n6829;
  assign n6863 = ~n6852 & n6862;
  assign n6864 = ~n6861 & n6863;
  assign n6865 = ~n6855 & ~n6864;
  assign po0295 = n6858 | n6865;
  assign n6867 = pi0153 & pi0186;
  assign n6868 = pi0195 & n6867;
  assign n6869 = pi0185 & ~n6868;
  assign n6870 = ~pi0185 & n6868;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = ~pi0429 & ~n6871;
  assign n6873 = pi0185 & pi0429;
  assign n6874 = ~n6872 & ~n6873;
  assign po0296 = n6600 & ~n6874;
  assign n6876 = pi0186 & ~pi0429;
  assign n6877 = ~pi0186 & pi0429;
  assign n6878 = ~n6876 & ~n6877;
  assign po0297 = n6600 & n6878;
  assign n6880 = n3974 & n4820;
  assign n6881 = ~n5032 & ~n6880;
  assign po0304 = pi1747 & ~n6881;
  assign po0305 = ~pi0281 & ~pi1099;
  assign n6884 = pi0195 & ~n6867;
  assign n6885 = ~pi0195 & n6867;
  assign n6886 = ~n6884 & ~n6885;
  assign n6887 = ~pi0429 & ~n6886;
  assign n6888 = pi0195 & pi0429;
  assign n6889 = ~n6887 & ~n6888;
  assign po0306 = n6600 & ~n6889;
  assign po0307 = ~pi0196 & ~pi0261;
  assign n6892 = ~pi1579 & pi1818;
  assign n6893 = ~pi1709 & n3967;
  assign n6894 = pi0197 & ~n3967;
  assign n6895 = ~n6893 & ~n6894;
  assign n6896 = pi0874 & ~n6895;
  assign n6897 = pi0197 & ~pi0874;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = pi1579 & ~n6898;
  assign po0308 = n6892 | n6899;
  assign n6901 = pi1582 & n4128;
  assign n6902 = pi1568 & n6901;
  assign n6903 = pi1570 & n4126;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = pi1570 & pi1580;
  assign n6906 = pi1568 & n6905;
  assign n6907 = n4122 & n6906;
  assign n6908 = pi1582 & n6907;
  assign n6909 = n6904 & ~n6908;
  assign po0309 = n4136 & ~n6909;
  assign n6911 = ~pi0998 & ~n4820;
  assign n6912 = ~n3977 & n4820;
  assign n6913 = ~n6911 & ~n6912;
  assign po0310 = pi1747 & n6913;
  assign n6915 = ~n5821 & ~n5830;
  assign n6916 = n5839 & ~n5867;
  assign n6917 = n5876 & n6916;
  assign n6918 = n5857 & n6917;
  assign n6919 = ~n5872 & n5875;
  assign n6920 = n5852 & ~n6919;
  assign n6921 = n5847 & ~n6920;
  assign n6922 = n5845 & ~n6921;
  assign n6923 = n5839 & ~n6922;
  assign n6924 = n5828 & ~n6923;
  assign n6925 = ~n6918 & n6924;
  assign n6926 = n6915 & n6925;
  assign n6927 = ~n6915 & ~n6925;
  assign po0311 = n6926 | n6927;
  assign n6929 = ~pi1579 & pi1816;
  assign n6930 = ~pi1713 & n3967;
  assign n6931 = pi0201 & ~n3967;
  assign n6932 = ~n6930 & ~n6931;
  assign n6933 = pi0874 & ~n6932;
  assign n6934 = pi0201 & ~pi0874;
  assign n6935 = ~n6933 & ~n6934;
  assign n6936 = pi1579 & ~n6935;
  assign po0312 = n6929 | n6936;
  assign n6938 = ~pi1579 & pi1817;
  assign n6939 = ~pi1714 & n3967;
  assign n6940 = pi0202 & ~n3967;
  assign n6941 = ~n6939 & ~n6940;
  assign n6942 = pi0874 & ~n6941;
  assign n6943 = pi0202 & ~pi0874;
  assign n6944 = ~n6942 & ~n6943;
  assign n6945 = pi1579 & ~n6944;
  assign po0313 = n6938 | n6945;
  assign n6947 = ~pi1579 & pi1819;
  assign n6948 = ~pi1717 & n3967;
  assign n6949 = pi0203 & ~n3967;
  assign n6950 = ~n6948 & ~n6949;
  assign n6951 = pi0874 & ~n6950;
  assign n6952 = pi0203 & ~pi0874;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = pi1579 & ~n6953;
  assign po0314 = n6947 | n6954;
  assign n6956 = ~pi1579 & pi1820;
  assign n6957 = ~pi1718 & n3967;
  assign n6958 = pi0204 & ~n3967;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = pi0874 & ~n6959;
  assign n6961 = pi0204 & ~pi0874;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = pi1579 & ~n6962;
  assign po0315 = n6956 | n6963;
  assign n6965 = ~pi1579 & pi1821;
  assign n6966 = ~pi1711 & n3967;
  assign n6967 = pi0205 & ~n3967;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = pi0874 & ~n6968;
  assign n6970 = pi0205 & ~pi0874;
  assign n6971 = ~n6969 & ~n6970;
  assign n6972 = pi1579 & ~n6971;
  assign po0316 = n6965 | n6972;
  assign n6974 = ~pi1579 & pi1823;
  assign n6975 = ~pi1716 & n3965;
  assign n6976 = pi0206 & ~n3965;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = pi0874 & ~n6977;
  assign n6979 = pi0206 & ~pi0874;
  assign n6980 = ~n6978 & ~n6979;
  assign n6981 = pi1579 & ~n6980;
  assign po0317 = n6974 | n6981;
  assign n6983 = ~pi1579 & pi1829;
  assign n6984 = pi0207 & ~n3965;
  assign n6985 = ~pi1711 & n3965;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 = pi0874 & ~n6986;
  assign n6988 = pi0207 & ~pi0874;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = pi1579 & ~n6989;
  assign po0318 = n6983 | n6990;
  assign n6992 = ~pi1579 & pi1831;
  assign n6993 = ~pi1716 & n3958;
  assign n6994 = pi0208 & ~n3958;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = pi0874 & ~n6995;
  assign n6997 = pi0208 & ~pi0874;
  assign n6998 = ~n6996 & ~n6997;
  assign n6999 = pi1579 & ~n6998;
  assign po0319 = n6992 | n6999;
  assign n7001 = ~pi1579 & pi1830;
  assign n7002 = ~pi1712 & n3958;
  assign n7003 = pi0209 & ~n3958;
  assign n7004 = ~n7002 & ~n7003;
  assign n7005 = pi0874 & ~n7004;
  assign n7006 = pi0209 & ~pi0874;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 = pi1579 & ~n7007;
  assign po0320 = n7001 | n7008;
  assign n7010 = ~pi1579 & pi1832;
  assign n7011 = ~pi1713 & n3958;
  assign n7012 = pi0210 & ~n3958;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = pi0874 & ~n7013;
  assign n7015 = pi0210 & ~pi0874;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = pi1579 & ~n7016;
  assign po0321 = n7010 | n7017;
  assign n7019 = ~pi1579 & pi1833;
  assign n7020 = ~pi1714 & n3958;
  assign n7021 = pi0211 & ~n3958;
  assign n7022 = ~n7020 & ~n7021;
  assign n7023 = pi0874 & ~n7022;
  assign n7024 = pi0211 & ~pi0874;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = pi1579 & ~n7025;
  assign po0322 = n7019 | n7026;
  assign n7028 = ~pi1579 & pi1835;
  assign n7029 = ~pi1717 & n3958;
  assign n7030 = pi0212 & ~n3958;
  assign n7031 = ~n7029 & ~n7030;
  assign n7032 = pi0874 & ~n7031;
  assign n7033 = pi0212 & ~pi0874;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = pi1579 & ~n7034;
  assign po0323 = n7028 | n7035;
  assign n7037 = ~pi1579 & pi1836;
  assign n7038 = ~pi1718 & n3958;
  assign n7039 = pi0213 & ~n3958;
  assign n7040 = ~n7038 & ~n7039;
  assign n7041 = pi0874 & ~n7040;
  assign n7042 = pi0213 & ~pi0874;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = pi1579 & ~n7043;
  assign po0324 = n7037 | n7044;
  assign n7046 = ~pi1579 & pi1837;
  assign n7047 = ~pi1711 & n3958;
  assign n7048 = pi0214 & ~n3958;
  assign n7049 = ~n7047 & ~n7048;
  assign n7050 = pi0874 & ~n7049;
  assign n7051 = pi0214 & ~pi0874;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = pi1579 & ~n7052;
  assign po0325 = n7046 | n7053;
  assign n7055 = ~n5941 & ~n5942;
  assign n7056 = n6169 & n7055;
  assign n7057 = ~n6169 & ~n7055;
  assign po0326 = n7056 | n7057;
  assign n7059 = ~n5937 & ~n5967;
  assign n7060 = n5960 & n7059;
  assign n7061 = ~n5960 & ~n7059;
  assign po0327 = n7060 | n7061;
  assign n7063 = ~pi1579 & pi1834;
  assign n7064 = ~pi1709 & n3958;
  assign n7065 = pi0217 & ~n3958;
  assign n7066 = ~n7064 & ~n7065;
  assign n7067 = pi0874 & ~n7066;
  assign n7068 = pi0217 & ~pi0874;
  assign n7069 = ~n7067 & ~n7068;
  assign n7070 = pi1579 & ~n7069;
  assign po0328 = n7063 | n7070;
  assign n7072 = ~n5855 & ~n5861;
  assign n7073 = ~n5856 & ~n5874;
  assign n7074 = n7072 & n7073;
  assign n7075 = ~n5846 & ~n5849;
  assign n7076 = ~n5860 & ~n5864;
  assign n7077 = ~n5838 & ~n5842;
  assign n7078 = ~n7076 & n7077;
  assign n7079 = n7075 & n7078;
  assign n7080 = n7074 & n7079;
  assign n7081 = ~n5824 & ~n5827;
  assign n7082 = n7080 & ~n7081;
  assign n7083 = ~n5838 & n5841;
  assign n7084 = ~n5825 & ~n7083;
  assign n7085 = ~n5846 & n5848;
  assign n7086 = ~n5843 & ~n7085;
  assign n7087 = n5869 & ~n5874;
  assign n7088 = ~n5850 & ~n7087;
  assign n7089 = ~n5855 & n5863;
  assign n7090 = ~n5870 & ~n7089;
  assign n7091 = n7073 & ~n7090;
  assign n7092 = n7088 & ~n7091;
  assign n7093 = n7075 & ~n7092;
  assign n7094 = n7086 & ~n7093;
  assign n7095 = n7077 & ~n7094;
  assign n7096 = n7084 & ~n7095;
  assign n7097 = ~n7081 & ~n7096;
  assign n7098 = ~n7082 & ~n7097;
  assign n7099 = ~n7080 & n7081;
  assign n7100 = n7096 & n7099;
  assign po0329 = ~n7098 | n7100;
  assign n7102 = ~pi1579 & pi1825;
  assign n7103 = ~pi1714 & n3965;
  assign n7104 = pi0219 & ~n3965;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = pi0874 & ~n7105;
  assign n7107 = pi0219 & ~pi0874;
  assign n7108 = ~n7106 & ~n7107;
  assign n7109 = pi1579 & ~n7108;
  assign po0330 = n7102 | n7109;
  assign n7111 = ~pi1579 & pi1822;
  assign n7112 = ~pi1712 & n3965;
  assign n7113 = pi0220 & ~n3965;
  assign n7114 = ~n7112 & ~n7113;
  assign n7115 = pi0874 & ~n7114;
  assign n7116 = pi0220 & ~pi0874;
  assign n7117 = ~n7115 & ~n7116;
  assign n7118 = pi1579 & ~n7117;
  assign po0331 = n7111 | n7118;
  assign n7120 = pi0239 & pi0240;
  assign n7121 = pi0237 & pi0238;
  assign n7122 = n7120 & n7121;
  assign n7123 = pi0257 & n7122;
  assign n7124 = pi0221 & n7123;
  assign n7125 = ~pi0221 & ~n7123;
  assign n7126 = ~n7124 & ~n7125;
  assign n7127 = pi0874 & n7126;
  assign n7128 = pi0221 & ~pi0874;
  assign n7129 = ~n7127 & ~n7128;
  assign n7130 = ~pi0097 & pi1747;
  assign po0332 = ~n7129 & n7130;
  assign n7132 = pi0242 & pi1099;
  assign n7133 = ~pi0355 & ~pi1099;
  assign po0334 = n7132 | n7133;
  assign n7135 = pi0221 & pi0241;
  assign n7136 = pi0237 & pi0257;
  assign n7137 = pi0238 & n7136;
  assign n7138 = pi0239 & n7137;
  assign n7139 = pi0240 & n7138;
  assign n7140 = pi0242 & n7139;
  assign n7141 = n7135 & n7140;
  assign n7142 = pi0224 & n7141;
  assign n7143 = ~pi0224 & ~n7141;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = pi0874 & n7144;
  assign n7146 = pi0224 & ~pi0874;
  assign n7147 = ~n7145 & ~n7146;
  assign po0335 = n7130 & ~n7147;
  assign n7149 = ~pi1579 & pi1824;
  assign n7150 = ~pi1713 & n3965;
  assign n7151 = pi0225 & ~n3965;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = pi0874 & ~n7152;
  assign n7154 = pi0225 & ~pi0874;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = pi1579 & ~n7155;
  assign po0336 = n7149 | n7156;
  assign n7158 = ~pi1579 & pi1826;
  assign n7159 = ~pi1709 & n3965;
  assign n7160 = pi0226 & ~n3965;
  assign n7161 = ~n7159 & ~n7160;
  assign n7162 = pi0874 & ~n7161;
  assign n7163 = pi0226 & ~pi0874;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = pi1579 & ~n7164;
  assign po0337 = n7158 | n7165;
  assign n7167 = ~pi1579 & pi1827;
  assign n7168 = ~pi1717 & n3965;
  assign n7169 = pi0227 & ~n3965;
  assign n7170 = ~n7168 & ~n7169;
  assign n7171 = pi0874 & ~n7170;
  assign n7172 = pi0227 & ~pi0874;
  assign n7173 = ~n7171 & ~n7172;
  assign n7174 = pi1579 & ~n7173;
  assign po0338 = n7167 | n7174;
  assign n7176 = ~pi1579 & pi1815;
  assign n7177 = pi0228 & ~n3967;
  assign n7178 = ~pi1716 & n3967;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = pi0874 & ~n7179;
  assign n7181 = pi0228 & ~pi0874;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = pi1579 & ~n7182;
  assign po0339 = n7176 | n7183;
  assign n7185 = ~pi0152 & ~pi0199;
  assign n7186 = pi0229 & ~n7185;
  assign n7187 = ~pi1712 & n7185;
  assign n7188 = ~n7186 & ~n7187;
  assign n7189 = pi0874 & ~n7188;
  assign n7190 = pi0229 & ~pi0874;
  assign n7191 = ~n7189 & ~n7190;
  assign n7192 = pi1579 & ~n7191;
  assign n7193 = ~pi1579 & pi1806;
  assign po0340 = n7192 | n7193;
  assign n7195 = pi0230 & ~n7185;
  assign n7196 = ~pi1716 & n7185;
  assign n7197 = ~n7195 & ~n7196;
  assign n7198 = pi0874 & ~n7197;
  assign n7199 = pi0230 & ~pi0874;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201 = pi1579 & ~n7200;
  assign n7202 = ~pi1579 & pi1807;
  assign po0341 = n7201 | n7202;
  assign n7204 = pi0231 & ~n7185;
  assign n7205 = ~pi1709 & n7185;
  assign n7206 = ~n7204 & ~n7205;
  assign n7207 = pi0874 & ~n7206;
  assign n7208 = pi0231 & ~pi0874;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = pi1579 & ~n7209;
  assign n7211 = ~pi1579 & pi1810;
  assign po0342 = n7210 | n7211;
  assign n7213 = pi0232 & ~n7185;
  assign n7214 = ~pi1717 & n7185;
  assign n7215 = ~n7213 & ~n7214;
  assign n7216 = pi0874 & ~n7215;
  assign n7217 = pi0232 & ~pi0874;
  assign n7218 = ~n7216 & ~n7217;
  assign n7219 = pi1579 & ~n7218;
  assign n7220 = ~pi1579 & pi1811;
  assign po0343 = n7219 | n7220;
  assign n7222 = pi0233 & ~n7185;
  assign n7223 = ~pi1718 & n7185;
  assign n7224 = ~n7222 & ~n7223;
  assign n7225 = pi0874 & ~n7224;
  assign n7226 = pi0233 & ~pi0874;
  assign n7227 = ~n7225 & ~n7226;
  assign n7228 = pi1579 & ~n7227;
  assign n7229 = ~pi1579 & pi1812;
  assign po0344 = n7228 | n7229;
  assign n7231 = pi0234 & ~n7185;
  assign n7232 = ~pi1711 & n7185;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = pi0874 & ~n7233;
  assign n7235 = pi0234 & ~pi0874;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = pi1579 & ~n7236;
  assign n7238 = ~pi1579 & pi1813;
  assign po0345 = n7237 | n7238;
  assign n7240 = pi0235 & ~n7185;
  assign n7241 = ~pi1714 & n7185;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = pi0874 & ~n7242;
  assign n7244 = pi0235 & ~pi0874;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = pi1579 & ~n7245;
  assign n7247 = ~pi1579 & pi1809;
  assign po0346 = n7246 | n7247;
  assign n7249 = pi0224 & pi0242;
  assign n7250 = n7120 & n7137;
  assign n7251 = pi0221 & n7250;
  assign n7252 = pi0241 & n7251;
  assign n7253 = n7249 & n7252;
  assign n7254 = pi0243 & n7253;
  assign n7255 = pi0236 & n7254;
  assign n7256 = ~pi0236 & ~n7254;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = pi0874 & n7257;
  assign n7259 = pi0236 & ~pi0874;
  assign n7260 = ~n7258 & ~n7259;
  assign po0347 = n7130 & ~n7260;
  assign n7262 = pi0237 & ~pi0874;
  assign n7263 = pi0237 & ~pi0257;
  assign n7264 = ~pi0237 & pi0257;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = pi0874 & ~n7265;
  assign n7267 = ~n7262 & ~n7266;
  assign po0348 = n7130 & ~n7267;
  assign n7269 = ~pi0238 & ~n7136;
  assign n7270 = ~n7137 & ~n7269;
  assign n7271 = pi0874 & n7270;
  assign n7272 = pi0238 & ~pi0874;
  assign n7273 = ~n7271 & ~n7272;
  assign po0349 = n7130 & ~n7273;
  assign n7275 = ~pi0239 & ~n7137;
  assign n7276 = ~n7138 & ~n7275;
  assign n7277 = pi0874 & n7276;
  assign n7278 = pi0239 & ~pi0874;
  assign n7279 = ~n7277 & ~n7278;
  assign po0350 = n7130 & ~n7279;
  assign n7281 = ~pi0240 & ~n7138;
  assign n7282 = ~n7139 & ~n7281;
  assign n7283 = pi0874 & n7282;
  assign n7284 = pi0240 & ~pi0874;
  assign n7285 = ~n7283 & ~n7284;
  assign po0351 = n7130 & ~n7285;
  assign n7287 = ~pi0241 & ~n7251;
  assign n7288 = ~n7252 & ~n7287;
  assign n7289 = pi0874 & n7288;
  assign n7290 = pi0241 & ~pi0874;
  assign n7291 = ~n7289 & ~n7290;
  assign po0352 = n7130 & ~n7291;
  assign n7293 = n7135 & n7250;
  assign n7294 = pi0242 & n7293;
  assign n7295 = ~pi0242 & ~n7293;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = pi0874 & n7296;
  assign n7298 = pi0242 & ~pi0874;
  assign n7299 = ~n7297 & ~n7298;
  assign po0353 = n7130 & ~n7299;
  assign n7301 = pi0241 & n7122;
  assign n7302 = pi0221 & n7301;
  assign n7303 = pi0257 & n7302;
  assign n7304 = n7249 & n7303;
  assign n7305 = pi0243 & n7304;
  assign n7306 = ~pi0243 & ~n7304;
  assign n7307 = ~n7305 & ~n7306;
  assign n7308 = pi0874 & n7307;
  assign n7309 = pi0243 & ~pi0874;
  assign n7310 = ~n7308 & ~n7309;
  assign po0354 = n7130 & ~n7310;
  assign n7312 = ~pi0221 & ~n5488;
  assign n7313 = ~pi0221 & ~n5491;
  assign n7314 = ~pi0240 & ~n5488;
  assign n7315 = ~pi0221 & ~pi0240;
  assign n7316 = ~n5492 & ~n7315;
  assign n7317 = ~n7314 & n7316;
  assign n7318 = ~n7313 & n7317;
  assign n7319 = pi0237 & n5528;
  assign n7320 = n5524 & ~n7319;
  assign n7321 = ~n5528 & ~n7136;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = ~pi0237 & ~pi0257;
  assign n7324 = n7322 & ~n7323;
  assign n7325 = ~pi0239 & ~n5512;
  assign n7326 = ~pi0238 & ~n5503;
  assign n7327 = ~pi0238 & ~pi0239;
  assign n7328 = ~n5518 & ~n7327;
  assign n7329 = ~n7326 & n7328;
  assign n7330 = ~n7325 & n7329;
  assign n7331 = ~n7324 & ~n7330;
  assign n7332 = ~n7318 & n7331;
  assign n7333 = pi0236 & n5463;
  assign n7334 = ~n5464 & ~n7333;
  assign n7335 = ~pi0224 & n5552;
  assign n7336 = ~pi0224 & ~pi0243;
  assign n7337 = ~n5551 & n7336;
  assign n7338 = ~n7335 & ~n7337;
  assign n7339 = ~pi0243 & ~n5482;
  assign n7340 = ~pi0241 & ~pi0242;
  assign n7341 = ~n5539 & n7340;
  assign n7342 = ~n5539 & ~n5545;
  assign n7343 = ~pi0241 & n7342;
  assign n7344 = ~n7341 & ~n7343;
  assign n7345 = ~pi0243 & ~n5551;
  assign n7346 = ~pi0224 & ~n5482;
  assign n7347 = ~n5552 & ~n7336;
  assign n7348 = ~n7346 & n7347;
  assign n7349 = ~n7345 & n7348;
  assign n7350 = ~n7344 & ~n7349;
  assign n7351 = ~pi0242 & ~n5545;
  assign n7352 = ~n7349 & n7351;
  assign n7353 = ~n7350 & ~n7352;
  assign n7354 = ~n7339 & n7353;
  assign n7355 = n7338 & n7354;
  assign n7356 = pi0236 & n5460;
  assign n7357 = ~n7355 & ~n7356;
  assign n7358 = ~n7334 & ~n7357;
  assign n7359 = pi0974 & n7358;
  assign n7360 = n5473 & n7359;
  assign n7361 = ~n5491 & n7315;
  assign n7362 = ~pi0240 & n5492;
  assign n7363 = ~n7361 & ~n7362;
  assign n7364 = ~pi0239 & ~n5503;
  assign n7365 = ~pi0238 & n5518;
  assign n7366 = ~n5512 & n7327;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = ~n7364 & n7367;
  assign n7369 = ~n7318 & ~n7368;
  assign n7370 = n7363 & ~n7369;
  assign n7371 = n7360 & n7370;
  assign n7372 = ~n7332 & n7371;
  assign n7373 = ~n7312 & n7372;
  assign n7374 = ~pi0242 & ~n5539;
  assign n7375 = ~pi0241 & ~n5545;
  assign n7376 = ~n7340 & ~n7342;
  assign n7377 = ~n7375 & n7376;
  assign n7378 = ~n7374 & n7377;
  assign n7379 = ~n7349 & ~n7378;
  assign n7380 = ~n7356 & n7379;
  assign n7381 = n7360 & ~n7380;
  assign po0355 = n7373 | n7381;
  assign n7383 = ~n5935 & ~n5963;
  assign n7384 = n5938 & n5952;
  assign n7385 = ~n6214 & n7384;
  assign n7386 = n6219 & ~n7385;
  assign n7387 = ~n7383 & ~n7386;
  assign n7388 = n7383 & n7386;
  assign po0356 = n7387 | n7388;
  assign n7390 = ~pi1579 & pi1828;
  assign n7391 = ~pi1718 & n3965;
  assign n7392 = pi0246 & ~n3965;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 = pi0874 & ~n7393;
  assign n7395 = pi0246 & ~pi0874;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = pi1579 & ~n7396;
  assign po0357 = n7390 | n7397;
  assign n7399 = pi0247 & ~n7185;
  assign n7400 = ~pi1713 & n7185;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = pi0874 & ~n7401;
  assign n7403 = pi0247 & ~pi0874;
  assign n7404 = ~n7402 & ~n7403;
  assign n7405 = pi1579 & ~n7404;
  assign n7406 = ~pi1579 & pi1808;
  assign po0358 = n7405 | n7406;
  assign n7408 = ~pi1579 & pi1814;
  assign n7409 = pi0248 & ~n3967;
  assign n7410 = ~pi1712 & n3967;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = pi0874 & ~n7411;
  assign n7413 = pi0248 & ~pi0874;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = pi1579 & ~n7414;
  assign po0359 = n7408 | n7415;
  assign n7417 = ~pi1127 & ~pi1308;
  assign n7418 = pi1127 & pi1308;
  assign n7419 = ~pi1076 & pi1420;
  assign n7420 = ~pi1029 & pi1444;
  assign n7421 = ~pi1029 & ~pi1076;
  assign n7422 = pi1420 & pi1444;
  assign n7423 = ~n7421 & ~n7422;
  assign n7424 = ~n7420 & n7423;
  assign n7425 = ~n7419 & n7424;
  assign n7426 = ~pi1130 & ~pi1452;
  assign n7427 = ~n7425 & n7426;
  assign n7428 = ~pi1083 & ~pi1130;
  assign n7429 = ~pi1500 & n7428;
  assign n7430 = ~pi1452 & ~pi1500;
  assign n7431 = ~pi1083 & n7430;
  assign n7432 = ~n7429 & ~n7431;
  assign n7433 = ~n7425 & ~n7432;
  assign n7434 = ~n7427 & ~n7433;
  assign n7435 = ~pi1076 & n7422;
  assign n7436 = pi1444 & n7421;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~pi1029 & pi1420;
  assign n7439 = n7437 & ~n7438;
  assign n7440 = n7434 & n7439;
  assign n7441 = ~n7418 & ~n7440;
  assign n7442 = ~n7417 & ~n7441;
  assign n7443 = ~pi1083 & ~pi1452;
  assign n7444 = ~pi1130 & ~pi1500;
  assign n7445 = ~n7428 & ~n7430;
  assign n7446 = ~n7444 & n7445;
  assign n7447 = ~n7443 & n7446;
  assign n7448 = ~pi1129 & ~pi1530;
  assign n7449 = ~pi1028 & pi1552;
  assign n7450 = ~pi1028 & ~pi1129;
  assign n7451 = ~pi1530 & pi1552;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = ~n7449 & n7452;
  assign n7454 = ~n7448 & n7453;
  assign n7455 = ~pi1310 & ~pi1558;
  assign n7456 = pi1027 & pi1630;
  assign n7457 = pi1310 & pi1558;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = ~n7455 & ~n7458;
  assign n7460 = ~n7454 & ~n7459;
  assign n7461 = ~pi1129 & n7451;
  assign n7462 = pi1552 & n7450;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = ~pi1028 & ~pi1530;
  assign n7465 = n7463 & ~n7464;
  assign n7466 = ~n7460 & n7465;
  assign n7467 = ~n7418 & ~n7425;
  assign n7468 = ~n7466 & n7467;
  assign n7469 = ~n7447 & n7468;
  assign n7470 = ~pi0949 & ~pi0980;
  assign n7471 = ~n7469 & n7470;
  assign n7472 = pi1341 & n7471;
  assign po0360 = ~n7442 | ~n7472;
  assign n7474 = ~pi0706 & pi1318;
  assign n7475 = pi0250 & pi0706;
  assign n7476 = ~n7474 & ~n7475;
  assign po0361 = pi1747 & ~n7476;
  assign n7478 = ~pi0706 & pi1042;
  assign n7479 = pi0251 & pi0706;
  assign n7480 = ~n7478 & ~n7479;
  assign po0362 = pi1747 & ~n7480;
  assign n7482 = ~pi0706 & pi1044;
  assign n7483 = pi0252 & pi0706;
  assign n7484 = ~n7482 & ~n7483;
  assign po0363 = pi1747 & ~n7484;
  assign n7486 = ~pi0706 & pi1313;
  assign n7487 = pi0253 & pi0706;
  assign n7488 = ~n7486 & ~n7487;
  assign po0364 = pi1747 & ~n7488;
  assign n7490 = pi0241 & pi1099;
  assign n7491 = ~pi0431 & ~pi1099;
  assign po0365 = n7490 | n7491;
  assign n7493 = ~pi0706 & pi1317;
  assign n7494 = pi0255 & pi0706;
  assign n7495 = ~n7493 & ~n7494;
  assign po0366 = pi1747 & ~n7495;
  assign n7497 = ~pi0256 & pi0630;
  assign po0367 = pi0354 & n7497;
  assign n7499 = ~pi0257 & ~pi0874;
  assign n7500 = pi0257 & pi0874;
  assign n7501 = ~n7499 & ~n7500;
  assign po0368 = n7130 & n7501;
  assign n7503 = ~pi0874 & ~n7185;
  assign n7504 = n3710 & n3715;
  assign n7505 = ~pi0336 & n7504;
  assign n7506 = pi0660 & n7505;
  assign n7507 = pi1409 & n7506;
  assign n7508 = ~pi0138 & n7507;
  assign n7509 = n3711 & n3715;
  assign n7510 = pi0336 & n7509;
  assign n7511 = ~n7506 & n7510;
  assign n7512 = ~n7508 & ~n7511;
  assign po0369 = n7503 & ~n7512;
  assign n7514 = n5442 & n6070;
  assign n7515 = pi0625 & n7514;
  assign n7516 = po1526 & n7515;
  assign po0370 = pi0089 & n7516;
  assign n7518 = ~n5946 & ~n5947;
  assign n7519 = ~n6018 & ~n7518;
  assign n7520 = n6018 & n7518;
  assign po0371 = n7519 | n7520;
  assign n7522 = pi0874 & n3958;
  assign po0372 = pi0258 | n7522;
  assign n7524 = pi0300 & pi0301;
  assign n7525 = ~pi0302 & ~n7524;
  assign n7526 = pi0303 & ~n7525;
  assign n7527 = n6781 & n7526;
  assign n7528 = pi0304 & pi0305;
  assign n7529 = n6695 & n7528;
  assign n7530 = n6781 & ~n7529;
  assign po0373 = n7527 | n7530;
  assign n7532 = ~pi0706 & pi1043;
  assign n7533 = pi0263 & pi0706;
  assign n7534 = ~n7532 & ~n7533;
  assign po0374 = pi1747 & ~n7534;
  assign n7536 = ~pi1119 & ~pi1307;
  assign n7537 = pi1119 & pi1307;
  assign n7538 = ~pi1270 & pi1432;
  assign n7539 = ~pi1267 & pi1443;
  assign n7540 = ~pi1267 & ~pi1270;
  assign n7541 = pi1432 & pi1443;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = ~n7539 & n7542;
  assign n7544 = ~n7538 & n7543;
  assign n7545 = ~pi1450 & ~pi1499;
  assign n7546 = ~pi1121 & n7545;
  assign n7547 = ~pi1121 & ~pi1274;
  assign n7548 = ~pi1499 & n7547;
  assign n7549 = ~n7546 & ~n7548;
  assign n7550 = ~n7544 & ~n7549;
  assign n7551 = ~pi1274 & ~pi1450;
  assign n7552 = ~n7544 & n7551;
  assign n7553 = ~n7550 & ~n7552;
  assign n7554 = ~pi1270 & n7541;
  assign n7555 = pi1443 & n7540;
  assign n7556 = ~n7554 & ~n7555;
  assign n7557 = ~pi1267 & pi1432;
  assign n7558 = n7556 & ~n7557;
  assign n7559 = n7553 & n7558;
  assign n7560 = ~n7537 & ~n7559;
  assign n7561 = ~n7536 & ~n7560;
  assign n7562 = ~pi1121 & ~pi1450;
  assign n7563 = ~pi1274 & ~pi1499;
  assign n7564 = ~n7545 & ~n7547;
  assign n7565 = ~n7563 & n7564;
  assign n7566 = ~n7562 & n7565;
  assign n7567 = ~pi1023 & ~pi1529;
  assign n7568 = ~pi1272 & pi1553;
  assign n7569 = ~pi1023 & ~pi1272;
  assign n7570 = ~pi1529 & pi1553;
  assign n7571 = ~n7569 & ~n7570;
  assign n7572 = ~n7568 & n7571;
  assign n7573 = ~n7567 & n7572;
  assign n7574 = ~pi1277 & ~pi1559;
  assign n7575 = pi1022 & pi1624;
  assign n7576 = pi1277 & pi1559;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = ~n7574 & ~n7577;
  assign n7579 = ~n7573 & ~n7578;
  assign n7580 = ~pi1023 & n7570;
  assign n7581 = pi1553 & n7569;
  assign n7582 = ~n7580 & ~n7581;
  assign n7583 = ~pi1272 & ~pi1529;
  assign n7584 = n7582 & ~n7583;
  assign n7585 = ~n7579 & n7584;
  assign n7586 = ~n7537 & ~n7544;
  assign n7587 = ~n7585 & n7586;
  assign n7588 = ~n7566 & n7587;
  assign n7589 = ~pi0948 & ~pi0979;
  assign n7590 = ~n7588 & n7589;
  assign n7591 = pi1340 & n7590;
  assign po0375 = ~n7561 | ~n7591;
  assign n7593 = ~pi1139 & ~pi1309;
  assign n7594 = pi1139 & pi1309;
  assign n7595 = ~pi1265 & pi1433;
  assign n7596 = ~pi1034 & pi1446;
  assign n7597 = ~pi1034 & ~pi1265;
  assign n7598 = pi1433 & pi1446;
  assign n7599 = ~n7597 & ~n7598;
  assign n7600 = ~n7596 & n7599;
  assign n7601 = ~n7595 & n7600;
  assign n7602 = ~pi1142 & ~pi1453;
  assign n7603 = ~n7601 & n7602;
  assign n7604 = ~pi1033 & ~pi1142;
  assign n7605 = ~pi1501 & n7604;
  assign n7606 = ~pi1453 & ~pi1501;
  assign n7607 = ~pi1033 & n7606;
  assign n7608 = ~n7605 & ~n7607;
  assign n7609 = ~n7601 & ~n7608;
  assign n7610 = ~n7603 & ~n7609;
  assign n7611 = ~pi1265 & n7598;
  assign n7612 = pi1446 & n7597;
  assign n7613 = ~n7611 & ~n7612;
  assign n7614 = ~pi1034 & pi1433;
  assign n7615 = n7613 & ~n7614;
  assign n7616 = n7610 & n7615;
  assign n7617 = ~n7594 & ~n7616;
  assign n7618 = ~n7593 & ~n7617;
  assign n7619 = ~pi1033 & ~pi1453;
  assign n7620 = ~pi1142 & ~pi1501;
  assign n7621 = ~n7604 & ~n7606;
  assign n7622 = ~n7620 & n7621;
  assign n7623 = ~n7619 & n7622;
  assign n7624 = ~pi1141 & ~pi1531;
  assign n7625 = ~pi1258 & pi1555;
  assign n7626 = ~pi1141 & ~pi1258;
  assign n7627 = ~pi1531 & pi1555;
  assign n7628 = ~n7626 & ~n7627;
  assign n7629 = ~n7625 & n7628;
  assign n7630 = ~n7624 & n7629;
  assign n7631 = ~pi1342 & ~pi1557;
  assign n7632 = pi1032 & pi1623;
  assign n7633 = pi1342 & pi1557;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = ~n7631 & ~n7634;
  assign n7636 = ~n7630 & ~n7635;
  assign n7637 = ~pi1141 & n7627;
  assign n7638 = pi1555 & n7626;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = ~pi1258 & ~pi1531;
  assign n7641 = n7639 & ~n7640;
  assign n7642 = ~n7636 & n7641;
  assign n7643 = ~n7594 & ~n7601;
  assign n7644 = ~n7642 & n7643;
  assign n7645 = ~n7623 & n7644;
  assign n7646 = ~pi0950 & ~pi0981;
  assign n7647 = ~n7645 & n7646;
  assign n7648 = pi1399 & n7647;
  assign po0376 = ~n7618 | ~n7648;
  assign n7650 = ~pi1102 & ~pi1306;
  assign n7651 = pi1102 & pi1306;
  assign n7652 = ~pi1109 & pi1431;
  assign n7653 = ~pi1110 & pi1442;
  assign n7654 = ~pi1109 & ~pi1110;
  assign n7655 = pi1431 & pi1442;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = ~n7653 & n7656;
  assign n7658 = ~n7652 & n7657;
  assign n7659 = ~pi1081 & ~pi1451;
  assign n7660 = ~n7658 & n7659;
  assign n7661 = ~pi1081 & ~pi1108;
  assign n7662 = ~pi1498 & n7661;
  assign n7663 = ~pi1451 & ~pi1498;
  assign n7664 = ~pi1108 & n7663;
  assign n7665 = ~n7662 & ~n7664;
  assign n7666 = ~n7658 & ~n7665;
  assign n7667 = ~n7660 & ~n7666;
  assign n7668 = ~pi1109 & n7655;
  assign n7669 = pi1442 & n7654;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~pi1110 & pi1431;
  assign n7672 = n7670 & ~n7671;
  assign n7673 = n7667 & n7672;
  assign n7674 = ~n7651 & ~n7673;
  assign n7675 = ~n7650 & ~n7674;
  assign n7676 = ~pi1108 & ~pi1451;
  assign n7677 = ~pi1081 & ~pi1498;
  assign n7678 = ~n7661 & ~n7663;
  assign n7679 = ~n7677 & n7678;
  assign n7680 = ~n7676 & n7679;
  assign n7681 = ~pi1106 & ~pi1528;
  assign n7682 = ~pi1107 & pi1554;
  assign n7683 = ~pi1106 & ~pi1107;
  assign n7684 = ~pi1528 & pi1554;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = ~n7682 & n7685;
  assign n7687 = ~n7681 & n7686;
  assign n7688 = ~pi1338 & ~pi1560;
  assign n7689 = pi1105 & pi1622;
  assign n7690 = pi1338 & pi1560;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~n7688 & ~n7691;
  assign n7693 = ~n7687 & ~n7692;
  assign n7694 = ~pi1106 & n7684;
  assign n7695 = pi1554 & n7683;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = ~pi1107 & ~pi1528;
  assign n7698 = n7696 & ~n7697;
  assign n7699 = ~n7693 & n7698;
  assign n7700 = ~n7651 & ~n7658;
  assign n7701 = ~n7699 & n7700;
  assign n7702 = ~n7680 & n7701;
  assign n7703 = ~pi0947 & ~pi0978;
  assign n7704 = ~n7702 & n7703;
  assign n7705 = pi1398 & n7704;
  assign po0377 = ~n7675 | ~n7705;
  assign n7707 = pi1233 & ~po0462;
  assign n7708 = ~po1678 & n5234;
  assign po0378 = n7707 & ~n7708;
  assign n7710 = ~pi0268 & pi0331;
  assign n7711 = pi0268 & ~pi0331;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = pi0706 & ~pi1671;
  assign n7714 = pi1747 & n7713;
  assign po0379 = ~n7712 & n7714;
  assign n7716 = ~pi0706 & pi1039;
  assign n7717 = pi0269 & pi0706;
  assign n7718 = ~n7716 & ~n7717;
  assign po0380 = pi1747 & ~n7718;
  assign n7720 = ~pi0706 & pi1041;
  assign n7721 = pi0270 & pi0706;
  assign n7722 = ~n7720 & ~n7721;
  assign po0381 = pi1747 & ~n7722;
  assign n7724 = ~pi0706 & pi1040;
  assign n7725 = pi0271 & pi0706;
  assign n7726 = ~n7724 & ~n7725;
  assign po0382 = pi1747 & ~n7726;
  assign n7728 = ~pi0706 & pi1049;
  assign n7729 = pi0272 & pi0706;
  assign n7730 = ~n7728 & ~n7729;
  assign po0383 = pi1747 & ~n7730;
  assign n7732 = ~pi0706 & pi1017;
  assign n7733 = pi0273 & pi0706;
  assign n7734 = ~n7732 & ~n7733;
  assign po0384 = pi1747 & ~n7734;
  assign n7736 = pi0268 & pi0331;
  assign n7737 = pi0274 & ~n7736;
  assign n7738 = ~pi0274 & n7736;
  assign n7739 = ~n7737 & ~n7738;
  assign po0385 = n7714 & ~n7739;
  assign n7741 = pi0274 & n7736;
  assign n7742 = pi0275 & ~n7741;
  assign n7743 = ~pi0275 & n7741;
  assign n7744 = ~n7742 & ~n7743;
  assign po0386 = n7714 & ~n7744;
  assign n7746 = pi0292 & pi0293;
  assign n7747 = pi0283 & n7746;
  assign n7748 = pi0291 & n7746;
  assign n7749 = pi0287 & pi0288;
  assign n7750 = pi0289 & n7749;
  assign n7751 = pi0290 & ~n7750;
  assign n7752 = n7748 & ~n7751;
  assign n7753 = n6781 & ~n7752;
  assign po0387 = ~n7747 & n7753;
  assign n7755 = ~pi0303 & n7525;
  assign n7756 = n6781 & ~n7755;
  assign po0388 = n7530 | n7756;
  assign n7758 = ~pi0279 & pi0294;
  assign n7759 = pi0279 & ~pi0294;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~pi1621 & n6781;
  assign po0389 = ~n7760 & n7761;
  assign n7763 = ~n5825 & ~n5838;
  assign n7764 = ~n5878 & ~n7763;
  assign n7765 = n5878 & n7763;
  assign po0390 = n7764 | n7765;
  assign n7767 = ~n5822 & ~n5833;
  assign n7768 = n7073 & n7075;
  assign n7769 = n7072 & ~n7076;
  assign n7770 = n7090 & ~n7769;
  assign n7771 = ~n5821 & ~n5824;
  assign n7772 = n7077 & n7771;
  assign n7773 = ~n7770 & n7772;
  assign n7774 = n7768 & n7773;
  assign n7775 = ~n5824 & ~n7084;
  assign n7776 = ~n5827 & ~n7775;
  assign n7777 = ~n5821 & ~n7776;
  assign n7778 = n7075 & ~n7088;
  assign n7779 = n7086 & ~n7778;
  assign n7780 = n7772 & ~n7779;
  assign n7781 = ~n7777 & ~n7780;
  assign n7782 = ~n7774 & n7781;
  assign n7783 = ~n5830 & n7782;
  assign n7784 = n7767 & n7783;
  assign n7785 = ~n7767 & ~n7783;
  assign po0391 = n7784 | n7785;
  assign n7787 = ~n5943 & ~n5951;
  assign n7788 = n6214 & n7787;
  assign n7789 = ~n6214 & ~n7787;
  assign po0392 = n7788 | n7789;
  assign n7791 = ~pi0283 & ~pi1621;
  assign n7792 = pi0290 & ~pi0291;
  assign n7793 = ~pi0289 & n7792;
  assign n7794 = ~pi0287 & ~pi0288;
  assign n7795 = n7793 & n7794;
  assign n7796 = ~pi0283 & ~n7795;
  assign n7797 = pi0283 & n7795;
  assign n7798 = ~n7796 & ~n7797;
  assign n7799 = pi1621 & ~n7798;
  assign n7800 = ~n7791 & ~n7799;
  assign n7801 = ~pi1534 & n6781;
  assign po0393 = ~n7800 & n7801;
  assign n7803 = pi0183 & pi1534;
  assign n7804 = pi0302 & n7524;
  assign n7805 = pi0303 & n7804;
  assign n7806 = ~pi0284 & n7805;
  assign n7807 = pi0284 & ~n7805;
  assign n7808 = ~n7806 & ~n7807;
  assign n7809 = n7803 & n7808;
  assign n7810 = ~pi0284 & ~n7803;
  assign n7811 = ~n7809 & ~n7810;
  assign po0394 = n6781 & ~n7811;
  assign n7813 = pi0275 & n7741;
  assign n7814 = pi0285 & n7813;
  assign n7815 = ~pi0285 & ~n7813;
  assign n7816 = ~n7814 & ~n7815;
  assign po0395 = n7714 & n7816;
  assign n7818 = pi0620 & ~pi1099;
  assign n7819 = pi0240 & pi1099;
  assign po0396 = n7818 | n7819;
  assign n7821 = ~pi0287 & ~pi1621;
  assign n7822 = pi0287 & pi1621;
  assign n7823 = ~n7821 & ~n7822;
  assign po0397 = n7801 & ~n7823;
  assign n7825 = ~pi0288 & ~pi1621;
  assign n7826 = ~pi0287 & pi0288;
  assign n7827 = pi0287 & ~pi0288;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = pi1621 & ~n7828;
  assign n7830 = ~n7825 & ~n7829;
  assign po0398 = n7801 & ~n7830;
  assign n7832 = ~pi0289 & ~pi1621;
  assign n7833 = ~pi0289 & ~n7794;
  assign n7834 = pi0289 & n7794;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = pi1621 & ~n7835;
  assign n7837 = ~n7832 & ~n7836;
  assign po0399 = n7801 & ~n7837;
  assign n7839 = pi0290 & ~pi1621;
  assign n7840 = ~pi0289 & n7794;
  assign n7841 = pi0290 & ~n7840;
  assign n7842 = ~pi0290 & n7840;
  assign n7843 = ~n7841 & ~n7842;
  assign n7844 = pi1621 & ~n7843;
  assign n7845 = ~n7839 & ~n7844;
  assign po0400 = n7801 & ~n7845;
  assign n7847 = ~pi0291 & ~pi1621;
  assign n7848 = pi0290 & n7840;
  assign n7849 = ~pi0291 & ~n7848;
  assign n7850 = pi0291 & n7848;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = pi1621 & ~n7851;
  assign n7853 = ~n7847 & ~n7852;
  assign po0401 = n7801 & ~n7853;
  assign n7855 = ~pi0292 & ~pi1621;
  assign n7856 = ~pi0283 & n7848;
  assign n7857 = ~pi0291 & n7856;
  assign n7858 = ~pi0292 & ~n7857;
  assign n7859 = pi0292 & n7857;
  assign n7860 = ~n7858 & ~n7859;
  assign n7861 = pi1621 & ~n7860;
  assign n7862 = ~n7855 & ~n7861;
  assign po0402 = n7801 & ~n7862;
  assign n7864 = ~pi0293 & ~pi1621;
  assign n7865 = n7792 & n7840;
  assign n7866 = ~pi0292 & n7865;
  assign n7867 = ~pi0283 & n7866;
  assign n7868 = ~pi0293 & ~n7867;
  assign n7869 = pi0293 & n7867;
  assign n7870 = ~n7868 & ~n7869;
  assign n7871 = pi1621 & ~n7870;
  assign n7872 = ~n7864 & ~n7871;
  assign po0403 = n7801 & ~n7872;
  assign po0404 = pi0294 & n7761;
  assign n7875 = ~pi0279 & ~pi0294;
  assign n7876 = ~pi0295 & n7875;
  assign n7877 = pi0295 & ~n7875;
  assign n7878 = ~n7876 & ~n7877;
  assign po0405 = n7761 & n7878;
  assign n7880 = ~pi0307 & n7876;
  assign n7881 = ~pi0296 & n7880;
  assign n7882 = pi0296 & ~n7880;
  assign n7883 = ~n7881 & ~n7882;
  assign po0406 = n7761 & n7883;
  assign n7885 = ~pi0296 & ~pi0307;
  assign n7886 = n7876 & n7885;
  assign n7887 = ~pi0297 & n7886;
  assign n7888 = pi0297 & ~n7886;
  assign n7889 = ~n7887 & ~n7888;
  assign po0407 = n7761 & n7889;
  assign n7891 = ~pi0297 & n7880;
  assign n7892 = ~pi0296 & n7891;
  assign n7893 = ~pi0298 & n7892;
  assign n7894 = pi0298 & ~n7892;
  assign n7895 = ~n7893 & ~n7894;
  assign po0408 = n7761 & n7895;
  assign n7897 = pi0239 & pi1099;
  assign n7898 = ~pi0545 & ~pi1099;
  assign po0409 = n7897 | n7898;
  assign n7900 = pi0300 & n7803;
  assign n7901 = ~pi0300 & ~n7803;
  assign n7902 = ~n7900 & ~n7901;
  assign po0410 = n6781 & n7902;
  assign n7904 = pi0301 & ~n7803;
  assign n7905 = pi0300 & ~pi0301;
  assign n7906 = ~pi0300 & pi0301;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = n7803 & ~n7907;
  assign n7909 = ~n7904 & ~n7908;
  assign po0411 = n6781 & ~n7909;
  assign n7911 = ~n7525 & ~n7804;
  assign n7912 = n7803 & n7911;
  assign n7913 = pi0302 & ~n7803;
  assign n7914 = ~n7912 & ~n7913;
  assign po0412 = n6781 & ~n7914;
  assign n7916 = ~pi0303 & ~n7804;
  assign n7917 = ~n7805 & ~n7916;
  assign n7918 = n7803 & n7917;
  assign n7919 = pi0303 & ~n7803;
  assign n7920 = ~n7918 & ~n7919;
  assign po0413 = n6781 & ~n7920;
  assign n7922 = ~pi0306 & n7805;
  assign n7923 = ~pi0284 & n7922;
  assign n7924 = ~pi0304 & n7923;
  assign n7925 = pi0304 & ~n7923;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = n7803 & n7926;
  assign n7928 = ~pi0304 & ~n7803;
  assign n7929 = ~n7927 & ~n7928;
  assign po0414 = n6781 & ~n7929;
  assign n7931 = ~pi0284 & pi0303;
  assign n7932 = n7804 & n7931;
  assign n7933 = ~pi0304 & n7932;
  assign n7934 = ~pi0306 & n7933;
  assign n7935 = ~pi0305 & n7934;
  assign n7936 = pi0305 & ~n7934;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = n7803 & n7937;
  assign n7939 = ~pi0305 & ~n7803;
  assign n7940 = ~n7938 & ~n7939;
  assign po0415 = n6781 & ~n7940;
  assign n7942 = ~pi0306 & n7932;
  assign n7943 = pi0306 & ~n7932;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n7803 & n7944;
  assign n7946 = ~pi0306 & ~n7803;
  assign n7947 = ~n7945 & ~n7946;
  assign po0416 = n6781 & ~n7947;
  assign n7949 = pi0307 & ~n7876;
  assign n7950 = ~n7880 & ~n7949;
  assign po0417 = n7761 & n7950;
  assign n7952 = ~pi0298 & n7886;
  assign n7953 = ~pi0297 & n7952;
  assign n7954 = ~pi0308 & n7953;
  assign n7955 = pi0308 & ~n7953;
  assign n7956 = ~n7954 & ~n7955;
  assign po0418 = n7761 & n7956;
  assign n7958 = ~pi1088 & ~pi1370;
  assign n7959 = n3721 & n7958;
  assign n7960 = pi0409 & n7959;
  assign n7961 = ~pi0309 & ~pi1101;
  assign n7962 = n7960 & ~n7961;
  assign n7963 = pi0309 & ~pi1409;
  assign n7964 = ~pi0138 & ~n7963;
  assign n7965 = n7506 & ~n7964;
  assign n7966 = ~n7962 & ~n7965;
  assign n7967 = pi0309 & n3712;
  assign n7968 = ~pi1090 & n7967;
  assign n7969 = pi0121 & ~pi0138;
  assign n7970 = ~pi0096 & n7969;
  assign n7971 = n7968 & ~n7970;
  assign n7972 = pi0097 & ~pi0138;
  assign n7973 = n7971 & ~n7972;
  assign n7974 = pi0309 & n7973;
  assign n7975 = pi0309 & ~pi1101;
  assign n7976 = ~pi0138 & ~n7975;
  assign n7977 = n3714 & ~n7976;
  assign n7978 = ~n7974 & ~n7977;
  assign n7979 = ~pi0309 & pi1250;
  assign n7980 = ~pi0258 & ~n7979;
  assign n7981 = ~pi0138 & ~n7980;
  assign n7982 = n7510 & ~n7981;
  assign n7983 = ~n3725 & ~n7976;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = n7978 & n7984;
  assign n7986 = ~pi0138 & ~pi1547;
  assign n7987 = n3955 & n3958;
  assign n7988 = pi0309 & ~n7987;
  assign n7989 = n7986 & ~n7988;
  assign n7990 = n3709 & n3721;
  assign n7991 = pi1370 & n7990;
  assign n7992 = ~n7989 & n7991;
  assign n7993 = n7985 & ~n7992;
  assign n7994 = pi1747 & n7993;
  assign po0419 = ~n7966 | ~n7994;
  assign n7996 = ~pi0726 & ~pi1099;
  assign n7997 = pi0237 & pi1099;
  assign po0420 = n7996 | n7997;
  assign n7999 = ~pi1758 & pi1759;
  assign n8000 = ~pi1761 & pi1762;
  assign n8001 = ~pi1763 & ~pi1764;
  assign n8002 = ~pi1760 & n8001;
  assign n8003 = n8000 & n8002;
  assign n8004 = ~pi1773 & n3738;
  assign n8005 = n3855 & n8004;
  assign n8006 = n8003 & n8005;
  assign n8007 = n7999 & n8006;
  assign n8008 = pi1802 & n8007;
  assign n8009 = pi1430 & pi1526;
  assign n8010 = pi1082 & n8009;
  assign n8011 = pi1047 & pi1430;
  assign n8012 = ~pi0311 & ~n8011;
  assign n8013 = ~pi1672 & n8011;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~n8009 & ~n8014;
  assign n8016 = ~n8010 & ~n8015;
  assign n8017 = ~n8007 & ~n8016;
  assign n8018 = pi1747 & ~n8017;
  assign po0421 = n8008 | ~n8018;
  assign n8020 = pi1805 & n8007;
  assign n8021 = ~pi1075 & n8009;
  assign n8022 = ~pi0312 & ~n8011;
  assign n8023 = ~pi1666 & n8011;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = ~n8009 & ~n8024;
  assign n8026 = ~n8021 & ~n8025;
  assign n8027 = ~n8007 & ~n8026;
  assign n8028 = pi1747 & ~n8027;
  assign po0422 = n8020 | ~n8028;
  assign n8030 = pi1783 & n8007;
  assign n8031 = ~pi1182 & n8009;
  assign n8032 = pi0022 & n8011;
  assign n8033 = ~pi0313 & ~n8011;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 = ~n8009 & ~n8034;
  assign n8036 = ~n8031 & ~n8035;
  assign n8037 = ~n8007 & ~n8036;
  assign n8038 = pi1747 & ~n8037;
  assign po0423 = n8030 | ~n8038;
  assign n8040 = pi1801 & n8007;
  assign n8041 = pi1176 & n8009;
  assign n8042 = pi0124 & n8011;
  assign n8043 = ~pi0314 & ~n8011;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = ~n8009 & ~n8044;
  assign n8046 = ~n8041 & ~n8045;
  assign n8047 = ~n8007 & ~n8046;
  assign n8048 = pi1747 & ~n8047;
  assign po0424 = n8040 | ~n8048;
  assign n8050 = pi1788 & n8007;
  assign n8051 = ~pi1169 & n8009;
  assign n8052 = pi0011 & n8011;
  assign n8053 = ~pi0315 & ~n8011;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = ~n8009 & ~n8054;
  assign n8056 = ~n8051 & ~n8055;
  assign n8057 = ~n8007 & ~n8056;
  assign n8058 = pi1747 & ~n8057;
  assign po0425 = n8050 | ~n8058;
  assign n8060 = pi1784 & n8007;
  assign n8061 = ~pi1166 & n8009;
  assign n8062 = pi0016 & n8011;
  assign n8063 = ~pi0316 & ~n8011;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = ~n8009 & ~n8064;
  assign n8066 = ~n8061 & ~n8065;
  assign n8067 = ~n8007 & ~n8066;
  assign n8068 = pi1747 & ~n8067;
  assign po0426 = n8060 | ~n8068;
  assign n8070 = pi1787 & n8007;
  assign n8071 = ~pi1239 & n8009;
  assign n8072 = pi0007 & n8011;
  assign n8073 = ~pi0317 & ~n8011;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = ~n8009 & ~n8074;
  assign n8076 = ~n8071 & ~n8075;
  assign n8077 = ~n8007 & ~n8076;
  assign n8078 = pi1747 & ~n8077;
  assign po0427 = n8070 | ~n8078;
  assign n8080 = pi1758 & pi1759;
  assign n8081 = n8006 & n8080;
  assign n8082 = pi1430 & pi1729;
  assign n8083 = pi0996 & pi1430;
  assign n8084 = ~n8082 & ~n8083;
  assign n8085 = pi0011 & ~n8084;
  assign n8086 = ~pi0318 & n8084;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = ~n8081 & ~n8087;
  assign n8089 = pi1788 & n8081;
  assign n8090 = ~n8088 & ~n8089;
  assign po0428 = ~pi1747 | ~n8090;
  assign n8092 = pi1785 & n8007;
  assign n8093 = ~pi1167 & n8009;
  assign n8094 = pi0019 & n8011;
  assign n8095 = ~pi0319 & ~n8011;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = ~n8009 & ~n8096;
  assign n8098 = ~n8093 & ~n8097;
  assign n8099 = ~n8007 & ~n8098;
  assign n8100 = pi1747 & ~n8099;
  assign po0429 = n8092 | ~n8100;
  assign n8102 = pi1789 & n8007;
  assign n8103 = ~pi1246 & n8009;
  assign n8104 = pi0018 & n8011;
  assign n8105 = ~pi0320 & ~n8011;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = ~n8009 & ~n8106;
  assign n8108 = ~n8103 & ~n8107;
  assign n8109 = ~n8007 & ~n8108;
  assign n8110 = pi1747 & ~n8109;
  assign po0430 = n8102 | ~n8110;
  assign n8112 = pi1780 & n8007;
  assign n8113 = ~pi1073 & n8009;
  assign n8114 = pi0023 & n8011;
  assign n8115 = ~pi0321 & ~n8011;
  assign n8116 = ~n8114 & ~n8115;
  assign n8117 = ~n8009 & ~n8116;
  assign n8118 = ~n8113 & ~n8117;
  assign n8119 = ~n8007 & ~n8118;
  assign n8120 = pi1747 & ~n8119;
  assign po0431 = n8112 | ~n8120;
  assign n8122 = pi0016 & ~n8084;
  assign n8123 = ~pi0322 & n8084;
  assign n8124 = ~n8122 & ~n8123;
  assign n8125 = ~n8081 & ~n8124;
  assign n8126 = pi1784 & n8081;
  assign n8127 = ~n8125 & ~n8126;
  assign po0432 = ~pi1747 | ~n8127;
  assign n8129 = pi0007 & ~n8084;
  assign n8130 = ~pi0323 & n8084;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = ~n8081 & ~n8131;
  assign n8133 = pi1787 & n8081;
  assign n8134 = ~n8132 & ~n8133;
  assign po0433 = ~pi1747 | ~n8134;
  assign n8136 = pi1781 & n8007;
  assign n8137 = ~pi1053 & n8009;
  assign n8138 = pi0030 & n8011;
  assign n8139 = ~pi0324 & ~n8011;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n8009 & ~n8140;
  assign n8142 = ~n8137 & ~n8141;
  assign n8143 = ~n8007 & ~n8142;
  assign n8144 = ~n8136 & ~n8143;
  assign po0434 = ~pi1747 | ~n8144;
  assign n8146 = pi0019 & ~n8084;
  assign n8147 = ~pi0325 & n8084;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = ~n8081 & ~n8148;
  assign n8150 = pi1785 & n8081;
  assign n8151 = ~n8149 & ~n8150;
  assign po0435 = ~pi1747 | ~n8151;
  assign n8153 = pi0018 & ~n8084;
  assign n8154 = ~pi0326 & n8084;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = ~n8081 & ~n8155;
  assign n8157 = pi1789 & n8081;
  assign n8158 = ~n8156 & ~n8157;
  assign po0436 = ~pi1747 | ~n8158;
  assign n8160 = pi0023 & ~n8084;
  assign n8161 = ~pi0327 & n8084;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~n8081 & ~n8162;
  assign n8164 = pi1780 & n8081;
  assign n8165 = ~n8163 & ~n8164;
  assign po0437 = ~pi1747 | ~n8165;
  assign n8167 = pi0046 & ~n8084;
  assign n8168 = ~pi0328 & n8084;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = ~n8081 & ~n8169;
  assign n8171 = pi1778 & n8081;
  assign n8172 = ~n8170 & ~n8171;
  assign po0438 = ~pi1747 | ~n8172;
  assign n8174 = pi0028 & ~n8084;
  assign n8175 = ~pi0329 & n8084;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8081 & ~n8176;
  assign n8178 = pi1779 & n8081;
  assign n8179 = ~n8177 & ~n8178;
  assign po0439 = ~pi1747 | ~n8179;
  assign n8181 = pi0030 & ~n8084;
  assign n8182 = ~pi0330 & n8084;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = ~n8081 & ~n8183;
  assign n8185 = pi1781 & n8081;
  assign n8186 = ~n8184 & ~n8185;
  assign po0440 = ~pi1747 | ~n8186;
  assign n8188 = ~pi0331 & n7713;
  assign po0441 = pi1747 & n8188;
  assign n8190 = pi0238 & pi1099;
  assign n8191 = ~pi0673 & ~pi1099;
  assign po0442 = n8190 | n8191;
  assign n8193 = ~n5850 & ~n5874;
  assign n8194 = n5873 & n8193;
  assign n8195 = ~n5873 & ~n8193;
  assign po0443 = n8194 | n8195;
  assign n8197 = ~pi1672 & ~n8084;
  assign n8198 = ~pi0334 & n8084;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = ~n8081 & ~n8199;
  assign n8201 = pi1802 & n8081;
  assign n8202 = ~n8200 & ~n8201;
  assign po0444 = ~pi1747 | ~n8202;
  assign n8204 = ~pi1666 & ~n8084;
  assign n8205 = ~pi0335 & n8084;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = ~n8081 & ~n8206;
  assign n8208 = pi1805 & n8081;
  assign n8209 = ~n8207 & ~n8208;
  assign po0445 = ~pi1747 | ~n8209;
  assign n8211 = ~pi0138 & ~pi1101;
  assign n8212 = ~n3725 & n8211;
  assign n8213 = pi0336 & n8212;
  assign n8214 = ~pi0138 & pi0336;
  assign n8215 = n7510 & n8214;
  assign n8216 = ~pi0258 & pi1250;
  assign n8217 = n8215 & n8216;
  assign n8218 = n7506 & n8214;
  assign n8219 = ~n7508 & ~n8218;
  assign n8220 = ~n8217 & n8219;
  assign n8221 = ~n8213 & n8220;
  assign po0446 = pi1747 & ~n8221;
  assign n8223 = pi1774 & n8007;
  assign n8224 = ~pi1254 & n8009;
  assign n8225 = pi0064 & n8011;
  assign n8226 = ~pi0337 & ~n8011;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~n8009 & ~n8227;
  assign n8229 = ~n8224 & ~n8228;
  assign n8230 = ~n8007 & ~n8229;
  assign n8231 = pi1747 & ~n8230;
  assign po0447 = n8223 | ~n8231;
  assign n8233 = pi1792 & n8007;
  assign n8234 = ~pi1171 & n8009;
  assign n8235 = pi0310 & n8011;
  assign n8236 = ~pi0338 & ~n8011;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = ~n8009 & ~n8237;
  assign n8239 = ~n8234 & ~n8238;
  assign n8240 = ~n8007 & ~n8239;
  assign n8241 = pi1747 & ~n8240;
  assign po0448 = n8233 | ~n8241;
  assign n8243 = pi1793 & n8007;
  assign n8244 = pi1241 & n8009;
  assign n8245 = pi0332 & n8011;
  assign n8246 = ~pi0339 & ~n8011;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = ~n8009 & ~n8247;
  assign n8249 = ~n8244 & ~n8248;
  assign n8250 = ~n8007 & ~n8249;
  assign n8251 = pi1747 & ~n8250;
  assign po0449 = n8243 | ~n8251;
  assign n8253 = pi1775 & n8007;
  assign n8254 = ~pi1172 & n8009;
  assign n8255 = pi0057 & n8011;
  assign n8256 = ~pi0340 & ~n8011;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = ~n8009 & ~n8257;
  assign n8259 = ~n8254 & ~n8258;
  assign n8260 = ~n8007 & ~n8259;
  assign n8261 = pi1747 & ~n8260;
  assign po0450 = n8253 | ~n8261;
  assign n8263 = pi1794 & n8007;
  assign n8264 = pi1077 & n8009;
  assign n8265 = pi0299 & n8011;
  assign n8266 = ~pi0341 & ~n8011;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~n8009 & ~n8267;
  assign n8269 = ~n8264 & ~n8268;
  assign n8270 = ~n8007 & ~n8269;
  assign n8271 = pi1747 & ~n8270;
  assign po0451 = n8263 | ~n8271;
  assign n8273 = pi1795 & n8007;
  assign n8274 = pi1173 & n8009;
  assign n8275 = pi0286 & n8011;
  assign n8276 = ~pi0342 & ~n8011;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = ~n8009 & ~n8277;
  assign n8279 = ~n8274 & ~n8278;
  assign n8280 = ~n8007 & ~n8279;
  assign n8281 = pi1747 & ~n8280;
  assign po0452 = n8273 | ~n8281;
  assign n8283 = pi1797 & n8007;
  assign n8284 = pi1174 & n8009;
  assign n8285 = pi0254 & n8011;
  assign n8286 = ~pi0343 & ~n8011;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~n8009 & ~n8287;
  assign n8289 = ~n8284 & ~n8288;
  assign n8290 = ~n8007 & ~n8289;
  assign n8291 = pi1747 & ~n8290;
  assign po0453 = n8283 | ~n8291;
  assign n8293 = pi1798 & n8007;
  assign n8294 = pi1093 & n8009;
  assign n8295 = pi0223 & n8011;
  assign n8296 = ~pi0344 & ~n8011;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = ~n8009 & ~n8297;
  assign n8299 = ~n8294 & ~n8298;
  assign n8300 = ~n8007 & ~n8299;
  assign n8301 = pi1747 & ~n8300;
  assign po0454 = n8293 | ~n8301;
  assign n8303 = pi1799 & n8007;
  assign n8304 = pi1175 & n8009;
  assign n8305 = pi0154 & n8011;
  assign n8306 = ~pi0345 & ~n8011;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = ~n8009 & ~n8307;
  assign n8309 = ~n8304 & ~n8308;
  assign n8310 = ~n8007 & ~n8309;
  assign n8311 = pi1747 & ~n8310;
  assign po0455 = n8303 | ~n8311;
  assign n8313 = pi1800 & n8007;
  assign n8314 = pi1089 & n8009;
  assign n8315 = pi0155 & n8011;
  assign n8316 = ~pi0346 & ~n8011;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = ~n8009 & ~n8317;
  assign n8319 = ~n8314 & ~n8318;
  assign n8320 = ~n8007 & ~n8319;
  assign n8321 = pi1747 & ~n8320;
  assign po0456 = n8313 | ~n8321;
  assign n8323 = pi1804 & n8007;
  assign n8324 = pi1179 & n8009;
  assign n8325 = pi0063 & n8011;
  assign n8326 = ~pi0347 & ~n8011;
  assign n8327 = ~n8325 & ~n8326;
  assign n8328 = ~n8009 & ~n8327;
  assign n8329 = ~n8324 & ~n8328;
  assign n8330 = ~n8007 & ~n8329;
  assign n8331 = pi1747 & ~n8330;
  assign po0457 = n8323 | ~n8331;
  assign n8333 = pi1777 & n8007;
  assign n8334 = ~pi1180 & n8009;
  assign n8335 = pi0049 & n8011;
  assign n8336 = ~pi0348 & ~n8011;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~n8009 & ~n8337;
  assign n8339 = ~n8334 & ~n8338;
  assign n8340 = ~n8007 & ~n8339;
  assign n8341 = pi1747 & ~n8340;
  assign po0458 = n8333 | ~n8341;
  assign n8343 = pi1782 & n8007;
  assign n8344 = ~pi1055 & n8009;
  assign n8345 = pi0027 & n8011;
  assign n8346 = ~pi0349 & ~n8011;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = ~n8009 & ~n8347;
  assign n8349 = ~n8344 & ~n8348;
  assign n8350 = ~n8007 & ~n8349;
  assign n8351 = pi1747 & ~n8350;
  assign po0459 = n8343 | ~n8351;
  assign n8353 = pi1760 & n8001;
  assign n8354 = n8000 & n8353;
  assign n8355 = n8005 & n8354;
  assign n8356 = n7999 & n8355;
  assign n8357 = pi1802 & n8356;
  assign n8358 = pi1447 & pi1526;
  assign n8359 = pi1249 & n8358;
  assign n8360 = pi1047 & pi1447;
  assign n8361 = ~pi0350 & ~n8360;
  assign n8362 = ~pi1672 & n8360;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n8358 & ~n8363;
  assign n8365 = ~n8359 & ~n8364;
  assign n8366 = ~n8356 & ~n8365;
  assign n8367 = pi1747 & ~n8366;
  assign po0460 = n8357 | ~n8367;
  assign n8369 = pi1805 & n8356;
  assign n8370 = ~pi1238 & n8358;
  assign n8371 = ~pi0351 & ~n8360;
  assign n8372 = ~pi1666 & n8360;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n8358 & ~n8373;
  assign n8375 = ~n8370 & ~n8374;
  assign n8376 = ~n8356 & ~n8375;
  assign n8377 = pi1747 & ~n8376;
  assign po0461 = n8369 | ~n8377;
  assign n8379 = ~n5841 & ~n5842;
  assign n8380 = n7768 & ~n7770;
  assign n8381 = n7779 & ~n8380;
  assign n8382 = ~n8379 & ~n8381;
  assign n8383 = n8379 & n8381;
  assign po0463 = n8382 | n8383;
  assign n8385 = ~n5843 & ~n5846;
  assign n8386 = n5857 & n5875;
  assign n8387 = ~n5867 & n8386;
  assign n8388 = n6920 & ~n8387;
  assign n8389 = ~n8385 & ~n8388;
  assign n8390 = n8385 & n8388;
  assign po0465 = n8389 | n8390;
  assign n8392 = pi1782 & n8356;
  assign n8393 = ~pi1245 & n8358;
  assign n8394 = pi0027 & n8360;
  assign n8395 = ~pi0356 & ~n8360;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~n8358 & ~n8396;
  assign n8398 = ~n8393 & ~n8397;
  assign n8399 = ~n8356 & ~n8398;
  assign n8400 = pi1747 & ~n8399;
  assign po0466 = n8392 | ~n8400;
  assign n8402 = n8080 & n8355;
  assign n8403 = pi1447 & pi1729;
  assign n8404 = pi0996 & pi1447;
  assign n8405 = ~n8403 & ~n8404;
  assign n8406 = pi0023 & ~n8405;
  assign n8407 = ~pi0357 & n8405;
  assign n8408 = ~n8406 & ~n8407;
  assign n8409 = ~n8402 & ~n8408;
  assign n8410 = pi1780 & n8402;
  assign n8411 = ~n8409 & ~n8410;
  assign po0467 = ~pi1747 | ~n8411;
  assign n8413 = pi1047 & pi1459;
  assign n8414 = pi1459 & pi1526;
  assign n8415 = pi1459 & pi1569;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~n8413 & n8416;
  assign n8418 = pi0358 & n8417;
  assign n8419 = pi0623 & ~pi1139;
  assign n8420 = ~pi0623 & pi1139;
  assign n8421 = pi0566 & ~pi1034;
  assign n8422 = ~n8420 & n8421;
  assign n8423 = ~n8419 & ~n8422;
  assign n8424 = ~pi0566 & pi1034;
  assign n8425 = ~n8420 & ~n8424;
  assign n8426 = pi0569 & ~pi1265;
  assign n8427 = ~pi0569 & pi1265;
  assign n8428 = pi0648 & ~pi1142;
  assign n8429 = ~n8427 & n8428;
  assign n8430 = ~n8426 & ~n8429;
  assign n8431 = ~pi0648 & pi1142;
  assign n8432 = ~n8427 & ~n8431;
  assign n8433 = ~pi0650 & pi1033;
  assign n8434 = ~pi0654 & pi1258;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = pi0650 & ~pi1033;
  assign n8437 = n8433 & ~n8436;
  assign n8438 = ~n8435 & n8437;
  assign n8439 = pi0654 & ~pi1258;
  assign n8440 = ~n8436 & ~n8439;
  assign n8441 = pi0653 & ~pi1141;
  assign n8442 = ~pi0653 & pi1141;
  assign n8443 = pi0662 & ~pi1342;
  assign n8444 = ~n8442 & n8443;
  assign n8445 = ~n8441 & ~n8444;
  assign n8446 = n8435 & ~n8445;
  assign n8447 = n8440 & ~n8446;
  assign n8448 = ~n8438 & ~n8447;
  assign n8449 = n8437 & n8445;
  assign n8450 = n8448 & ~n8449;
  assign n8451 = n8432 & n8450;
  assign n8452 = n8430 & ~n8451;
  assign n8453 = n8425 & ~n8452;
  assign n8454 = n8423 & ~n8453;
  assign n8455 = n8425 & n8432;
  assign n8456 = ~pi0662 & pi1342;
  assign n8457 = ~n8442 & ~n8456;
  assign n8458 = n8435 & n8457;
  assign n8459 = ~pi0586 & pi1032;
  assign n8460 = n8458 & ~n8459;
  assign n8461 = n8455 & n8460;
  assign n8462 = n8454 & ~n8461;
  assign n8463 = pi0358 & ~n8462;
  assign n8464 = ~pi0358 & n8462;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = ~n8417 & ~n8465;
  assign n8467 = ~n8418 & ~n8466;
  assign n8468 = pi1697 & ~n8467;
  assign n8469 = pi0648 & n6444;
  assign n8470 = pi0653 & pi0662;
  assign n8471 = pi0650 & pi0654;
  assign n8472 = n8470 & n8471;
  assign n8473 = n8469 & n8472;
  assign n8474 = pi0586 & n8473;
  assign n8475 = pi0623 & n8474;
  assign n8476 = pi0358 & n8475;
  assign n8477 = ~pi0358 & ~n8475;
  assign n8478 = ~n8476 & ~n8477;
  assign n8479 = ~pi1697 & n8478;
  assign n8480 = ~n8468 & ~n8479;
  assign po0468 = pi1143 & ~n8480;
  assign n8482 = pi1047 & pi1480;
  assign n8483 = pi1480 & pi1526;
  assign n8484 = pi1480 & pi1594;
  assign n8485 = ~n8483 & ~n8484;
  assign n8486 = ~n8482 & n8485;
  assign n8487 = pi0359 & n8486;
  assign n8488 = pi0712 & ~pi1102;
  assign n8489 = ~pi0712 & pi1102;
  assign n8490 = pi0675 & ~pi1110;
  assign n8491 = ~n8489 & n8490;
  assign n8492 = ~n8488 & ~n8491;
  assign n8493 = ~pi0675 & pi1110;
  assign n8494 = ~n8489 & ~n8493;
  assign n8495 = pi0678 & ~pi1109;
  assign n8496 = ~pi0678 & pi1109;
  assign n8497 = pi0714 & ~pi1081;
  assign n8498 = ~n8496 & n8497;
  assign n8499 = ~n8495 & ~n8498;
  assign n8500 = ~pi0714 & pi1081;
  assign n8501 = ~n8496 & ~n8500;
  assign n8502 = ~pi0717 & pi1108;
  assign n8503 = ~pi0708 & pi1107;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = pi0717 & ~pi1108;
  assign n8506 = n8502 & ~n8505;
  assign n8507 = ~n8504 & n8506;
  assign n8508 = pi0708 & ~pi1107;
  assign n8509 = ~n8505 & ~n8508;
  assign n8510 = pi0719 & ~pi1106;
  assign n8511 = ~pi0719 & pi1106;
  assign n8512 = pi0718 & ~pi1338;
  assign n8513 = ~n8511 & n8512;
  assign n8514 = ~n8510 & ~n8513;
  assign n8515 = n8504 & ~n8514;
  assign n8516 = n8509 & ~n8515;
  assign n8517 = ~n8507 & ~n8516;
  assign n8518 = n8506 & n8514;
  assign n8519 = n8517 & ~n8518;
  assign n8520 = n8501 & n8519;
  assign n8521 = n8499 & ~n8520;
  assign n8522 = n8494 & ~n8521;
  assign n8523 = n8492 & ~n8522;
  assign n8524 = n8494 & n8501;
  assign n8525 = ~pi0718 & pi1338;
  assign n8526 = ~n8511 & ~n8525;
  assign n8527 = n8504 & n8526;
  assign n8528 = ~pi0697 & pi1105;
  assign n8529 = n8527 & ~n8528;
  assign n8530 = n8524 & n8529;
  assign n8531 = n8523 & ~n8530;
  assign n8532 = pi0359 & ~n8531;
  assign n8533 = ~pi0359 & n8531;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = ~n8486 & ~n8534;
  assign n8536 = ~n8487 & ~n8535;
  assign n8537 = pi1699 & ~n8536;
  assign n8538 = pi0714 & n6806;
  assign n8539 = pi0718 & pi0719;
  assign n8540 = pi0708 & pi0717;
  assign n8541 = n8539 & n8540;
  assign n8542 = n8538 & n8541;
  assign n8543 = pi0697 & n8542;
  assign n8544 = pi0712 & n8543;
  assign n8545 = pi0359 & n8544;
  assign n8546 = ~pi0359 & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = ~pi1699 & n8547;
  assign n8549 = ~n8537 & ~n8548;
  assign po0469 = pi1111 & ~n8549;
  assign n8551 = ~pi0360 & n8084;
  assign n8552 = pi0049 & ~n8084;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 = ~n8081 & ~n8553;
  assign n8555 = pi1777 & n8081;
  assign n8556 = ~n8554 & ~n8555;
  assign po0470 = ~pi1747 | ~n8556;
  assign n8558 = ~n5948 & ~n5955;
  assign n8559 = ~n5954 & n8558;
  assign n8560 = n5954 & ~n8558;
  assign po0471 = n8559 | n8560;
  assign n8562 = pi1780 & n8356;
  assign n8563 = ~pi1244 & n8358;
  assign n8564 = pi0023 & n8360;
  assign n8565 = ~pi0362 & ~n8360;
  assign n8566 = ~n8564 & ~n8565;
  assign n8567 = ~n8358 & ~n8566;
  assign n8568 = ~n8563 & ~n8567;
  assign n8569 = ~n8356 & ~n8568;
  assign n8570 = pi1747 & ~n8569;
  assign po0472 = n8562 | ~n8570;
  assign n8572 = pi1788 & n8356;
  assign n8573 = ~pi1188 & n8358;
  assign n8574 = pi0011 & n8360;
  assign n8575 = ~pi0363 & ~n8360;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~n8358 & ~n8576;
  assign n8578 = ~n8573 & ~n8577;
  assign n8579 = ~n8356 & ~n8578;
  assign n8580 = pi1747 & ~n8579;
  assign po0473 = n8572 | ~n8580;
  assign n8582 = pi1784 & n8356;
  assign n8583 = ~pi1185 & n8358;
  assign n8584 = pi0016 & n8360;
  assign n8585 = ~pi0364 & ~n8360;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = ~n8358 & ~n8586;
  assign n8588 = ~n8583 & ~n8587;
  assign n8589 = ~n8356 & ~n8588;
  assign n8590 = pi1747 & ~n8589;
  assign po0474 = n8582 | ~n8590;
  assign n8592 = pi1787 & n8356;
  assign n8593 = ~pi1063 & n8358;
  assign n8594 = pi0007 & n8360;
  assign n8595 = ~pi0365 & ~n8360;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~n8358 & ~n8596;
  assign n8598 = ~n8593 & ~n8597;
  assign n8599 = ~n8356 & ~n8598;
  assign n8600 = pi1747 & ~n8599;
  assign po0475 = n8592 | ~n8600;
  assign n8602 = pi0011 & ~n8405;
  assign n8603 = ~pi0366 & n8405;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8402 & ~n8604;
  assign n8606 = pi1788 & n8402;
  assign n8607 = ~n8605 & ~n8606;
  assign po0476 = ~pi1747 | ~n8607;
  assign n8609 = pi1785 & n8356;
  assign n8610 = ~pi1186 & n8358;
  assign n8611 = pi0019 & n8360;
  assign n8612 = ~pi0367 & ~n8360;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = ~n8358 & ~n8613;
  assign n8615 = ~n8610 & ~n8614;
  assign n8616 = ~n8356 & ~n8615;
  assign n8617 = pi1747 & ~n8616;
  assign po0477 = n8609 | ~n8617;
  assign n8619 = pi1789 & n8356;
  assign n8620 = ~pi1189 & n8358;
  assign n8621 = pi0018 & n8360;
  assign n8622 = ~pi0368 & ~n8360;
  assign n8623 = ~n8621 & ~n8622;
  assign n8624 = ~n8358 & ~n8623;
  assign n8625 = ~n8620 & ~n8624;
  assign n8626 = ~n8356 & ~n8625;
  assign n8627 = pi1747 & ~n8626;
  assign po0478 = n8619 | ~n8627;
  assign n8629 = pi0016 & ~n8405;
  assign n8630 = ~pi0369 & n8405;
  assign n8631 = ~n8629 & ~n8630;
  assign n8632 = ~n8402 & ~n8631;
  assign n8633 = pi1784 & n8402;
  assign n8634 = ~n8632 & ~n8633;
  assign po0479 = ~pi1747 | ~n8634;
  assign n8636 = pi0007 & ~n8405;
  assign n8637 = ~pi0370 & n8405;
  assign n8638 = ~n8636 & ~n8637;
  assign n8639 = ~n8402 & ~n8638;
  assign n8640 = pi1787 & n8402;
  assign n8641 = ~n8639 & ~n8640;
  assign po0480 = ~pi1747 | ~n8641;
  assign n8643 = pi1781 & n8356;
  assign n8644 = ~pi1205 & n8358;
  assign n8645 = pi0030 & n8360;
  assign n8646 = ~pi0371 & ~n8360;
  assign n8647 = ~n8645 & ~n8646;
  assign n8648 = ~n8358 & ~n8647;
  assign n8649 = ~n8644 & ~n8648;
  assign n8650 = ~n8356 & ~n8649;
  assign n8651 = pi1747 & ~n8650;
  assign po0481 = n8643 | ~n8651;
  assign n8653 = pi0019 & ~n8405;
  assign n8654 = ~pi0372 & n8405;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = ~n8402 & ~n8655;
  assign n8657 = pi1785 & n8402;
  assign n8658 = ~n8656 & ~n8657;
  assign po0482 = ~pi1747 | ~n8658;
  assign n8660 = pi0018 & ~n8405;
  assign n8661 = ~pi0373 & n8405;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = ~n8402 & ~n8662;
  assign n8664 = pi1789 & n8402;
  assign n8665 = ~n8663 & ~n8664;
  assign po0483 = ~pi1747 | ~n8665;
  assign n8667 = pi0046 & ~n8405;
  assign n8668 = ~pi0374 & n8405;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = ~n8402 & ~n8669;
  assign n8671 = pi1778 & n8402;
  assign n8672 = ~n8670 & ~n8671;
  assign po0484 = ~pi1747 | ~n8672;
  assign n8674 = pi0030 & ~n8405;
  assign n8675 = ~pi0375 & n8405;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = ~n8402 & ~n8676;
  assign n8678 = pi1781 & n8402;
  assign n8679 = ~n8677 & ~n8678;
  assign po0485 = ~pi1747 | ~n8679;
  assign n8681 = pi0028 & ~n8405;
  assign n8682 = ~pi0376 & n8405;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = ~n8402 & ~n8683;
  assign n8685 = pi1779 & n8402;
  assign n8686 = ~n8684 & ~n8685;
  assign po0486 = ~pi1747 | ~n8686;
  assign n8688 = ~pi0377 & n8084;
  assign n8689 = pi0194 & ~n8084;
  assign n8690 = ~n8688 & ~n8689;
  assign n8691 = ~n8081 & ~n8690;
  assign n8692 = pi1803 & n8081;
  assign n8693 = ~n8691 & ~n8692;
  assign po0487 = ~pi1747 | ~n8693;
  assign n8695 = ~pi0378 & n8084;
  assign n8696 = pi0286 & ~n8084;
  assign n8697 = ~n8695 & ~n8696;
  assign n8698 = ~n8081 & ~n8697;
  assign n8699 = pi1795 & n8081;
  assign n8700 = ~n8698 & ~n8699;
  assign po0488 = ~pi1747 | ~n8700;
  assign n8702 = pi1430 & pi1571;
  assign n8703 = ~n8009 & ~n8702;
  assign n8704 = ~n8011 & n8703;
  assign n8705 = pi0379 & n8704;
  assign n8706 = pi0466 & ~pi1119;
  assign n8707 = ~pi0466 & pi1119;
  assign n8708 = pi0386 & ~pi1267;
  assign n8709 = ~n8707 & n8708;
  assign n8710 = ~n8706 & ~n8709;
  assign n8711 = ~pi0386 & pi1267;
  assign n8712 = ~n8707 & ~n8711;
  assign n8713 = pi0387 & ~pi1270;
  assign n8714 = ~pi0387 & pi1270;
  assign n8715 = pi0480 & ~pi1274;
  assign n8716 = ~n8714 & n8715;
  assign n8717 = ~n8713 & ~n8716;
  assign n8718 = ~pi0480 & pi1274;
  assign n8719 = ~n8714 & ~n8718;
  assign n8720 = ~pi0484 & pi1121;
  assign n8721 = ~pi0509 & pi1272;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = pi0484 & ~pi1121;
  assign n8724 = n8720 & ~n8723;
  assign n8725 = ~n8722 & n8724;
  assign n8726 = pi0509 & ~pi1272;
  assign n8727 = ~n8723 & ~n8726;
  assign n8728 = pi0508 & ~pi1023;
  assign n8729 = ~pi0508 & pi1023;
  assign n8730 = pi0507 & ~pi1277;
  assign n8731 = ~n8729 & n8730;
  assign n8732 = ~n8728 & ~n8731;
  assign n8733 = n8722 & ~n8732;
  assign n8734 = n8727 & ~n8733;
  assign n8735 = ~n8725 & ~n8734;
  assign n8736 = n8724 & n8732;
  assign n8737 = n8735 & ~n8736;
  assign n8738 = n8719 & n8737;
  assign n8739 = n8717 & ~n8738;
  assign n8740 = n8712 & ~n8739;
  assign n8741 = n8710 & ~n8740;
  assign n8742 = n8712 & n8719;
  assign n8743 = ~pi0507 & pi1277;
  assign n8744 = ~n8729 & ~n8743;
  assign n8745 = n8722 & n8744;
  assign n8746 = ~pi0408 & pi1022;
  assign n8747 = n8745 & ~n8746;
  assign n8748 = n8742 & n8747;
  assign n8749 = n8741 & ~n8748;
  assign n8750 = pi0379 & ~n8749;
  assign n8751 = ~pi0379 & n8749;
  assign n8752 = ~n8750 & ~n8751;
  assign n8753 = ~n8704 & ~n8752;
  assign n8754 = ~n8705 & ~n8753;
  assign n8755 = pi1690 & ~n8754;
  assign n8756 = pi0480 & n6522;
  assign n8757 = pi0507 & pi0508;
  assign n8758 = pi0484 & pi0509;
  assign n8759 = n8757 & n8758;
  assign n8760 = n8756 & n8759;
  assign n8761 = pi0408 & n8760;
  assign n8762 = pi0466 & n8761;
  assign n8763 = pi0379 & n8762;
  assign n8764 = ~pi0379 & ~n8762;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = ~pi1690 & n8765;
  assign n8767 = ~n8755 & ~n8766;
  assign po0489 = pi1122 & ~n8767;
  assign n8769 = pi1447 & pi1572;
  assign n8770 = ~n8358 & ~n8769;
  assign n8771 = ~n8360 & n8770;
  assign n8772 = pi0380 & n8771;
  assign n8773 = pi0533 & ~pi1127;
  assign n8774 = ~pi0533 & pi1127;
  assign n8775 = pi0483 & ~pi1029;
  assign n8776 = ~n8774 & n8775;
  assign n8777 = ~n8773 & ~n8776;
  assign n8778 = ~pi0483 & pi1029;
  assign n8779 = ~n8774 & ~n8778;
  assign n8780 = pi0485 & ~pi1076;
  assign n8781 = ~pi0485 & pi1076;
  assign n8782 = pi0549 & ~pi1130;
  assign n8783 = ~n8781 & n8782;
  assign n8784 = ~n8780 & ~n8783;
  assign n8785 = ~pi0549 & pi1130;
  assign n8786 = ~n8781 & ~n8785;
  assign n8787 = ~pi0567 & pi1083;
  assign n8788 = ~pi0622 & pi1028;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = pi0622 & ~pi1028;
  assign n8791 = pi0567 & ~pi1083;
  assign n8792 = ~n8790 & ~n8791;
  assign n8793 = ~n8789 & n8792;
  assign n8794 = n8787 & ~n8791;
  assign n8795 = pi0587 & ~pi1129;
  assign n8796 = ~pi0587 & pi1129;
  assign n8797 = pi0618 & ~pi1310;
  assign n8798 = ~n8796 & n8797;
  assign n8799 = ~n8795 & ~n8798;
  assign n8800 = n8789 & ~n8799;
  assign n8801 = n8794 & ~n8800;
  assign n8802 = ~n8793 & ~n8801;
  assign n8803 = n8792 & n8799;
  assign n8804 = n8802 & ~n8803;
  assign n8805 = n8786 & n8804;
  assign n8806 = n8784 & ~n8805;
  assign n8807 = n8779 & ~n8806;
  assign n8808 = n8777 & ~n8807;
  assign n8809 = n8779 & n8786;
  assign n8810 = ~pi0618 & pi1310;
  assign n8811 = ~n8796 & ~n8810;
  assign n8812 = n8789 & n8811;
  assign n8813 = ~pi0506 & pi1027;
  assign n8814 = n8812 & ~n8813;
  assign n8815 = n8809 & n8814;
  assign n8816 = n8808 & ~n8815;
  assign n8817 = pi0380 & ~n8816;
  assign n8818 = ~pi0380 & n8816;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~n8771 & ~n8819;
  assign n8821 = ~n8772 & ~n8820;
  assign n8822 = pi1679 & ~n8821;
  assign n8823 = pi0549 & n6345;
  assign n8824 = pi0587 & pi0618;
  assign n8825 = pi0567 & pi0622;
  assign n8826 = n8824 & n8825;
  assign n8827 = n8823 & n8826;
  assign n8828 = pi0506 & n8827;
  assign n8829 = pi0533 & n8828;
  assign n8830 = pi0380 & n8829;
  assign n8831 = ~pi0380 & ~n8829;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = ~pi1679 & n8832;
  assign n8834 = ~n8822 & ~n8833;
  assign po0490 = pi1131 & ~n8834;
  assign n8836 = pi0381 & n8704;
  assign n8837 = n8719 & ~n8724;
  assign n8838 = ~n8727 & n8837;
  assign n8839 = n8717 & ~n8838;
  assign n8840 = n8712 & ~n8839;
  assign n8841 = n8744 & ~n8746;
  assign n8842 = n8732 & ~n8841;
  assign n8843 = n8719 & n8722;
  assign n8844 = ~n8842 & n8843;
  assign n8845 = n8712 & n8844;
  assign n8846 = ~pi0379 & ~pi0470;
  assign n8847 = ~n8845 & n8846;
  assign n8848 = n8710 & n8847;
  assign n8849 = ~n8840 & n8848;
  assign n8850 = pi0381 & ~n8849;
  assign n8851 = ~pi0381 & n8849;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = ~n8704 & ~n8852;
  assign n8854 = ~n8836 & ~n8853;
  assign n8855 = pi1690 & ~n8854;
  assign n8856 = pi0408 & pi0507;
  assign n8857 = pi0508 & n8856;
  assign n8858 = pi0509 & n8857;
  assign n8859 = n6531 & n8858;
  assign n8860 = pi0387 & n8859;
  assign n8861 = n6548 & n8860;
  assign n8862 = pi0470 & n8861;
  assign n8863 = pi0386 & n8862;
  assign n8864 = pi0381 & n8863;
  assign n8865 = ~pi0381 & ~n8863;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = ~pi1690 & n8866;
  assign n8868 = ~n8855 & ~n8867;
  assign po0491 = pi1122 & ~n8868;
  assign n8870 = pi0696 & n5420;
  assign n8871 = ~pi0647 & n8870;
  assign n8872 = ~pi1627 & n5259;
  assign n8873 = ~pi1626 & pi1628;
  assign n8874 = ~pi1627 & n8873;
  assign n8875 = ~po1678 & ~n4135;
  assign n8876 = ~po1690 & ~po1688;
  assign n8877 = ~po1676 & n8876;
  assign n8878 = n8875 & n8877;
  assign n8879 = n8874 & ~n8878;
  assign n8880 = ~n8872 & n8879;
  assign n8881 = pi1227 & pi1228;
  assign n8882 = n4134 & n8881;
  assign n8883 = n4114 & n8881;
  assign n8884 = n4118 & n8881;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = ~n8882 & n8885;
  assign n8887 = n5232 & n8881;
  assign n8888 = n8886 & ~n8887;
  assign n8889 = pi1628 & n8888;
  assign n8890 = n8878 & n8889;
  assign n8891 = n5423 & ~n8890;
  assign n8892 = pi0382 & n8891;
  assign n8893 = pi0382 & ~pi1626;
  assign n8894 = ~n8891 & n8893;
  assign n8895 = ~n8892 & ~n8894;
  assign n8896 = n8874 & ~n8888;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = ~n8872 & n8897;
  assign n8899 = ~n8880 & ~n8898;
  assign n8900 = n8871 & ~n8899;
  assign n8901 = n8871 & n8872;
  assign n8902 = n8893 & n8901;
  assign n8903 = ~n8900 & ~n8902;
  assign n8904 = pi0382 & ~n8873;
  assign n8905 = ~pi0647 & ~pi0696;
  assign n8906 = ~pi0382 & n8905;
  assign n8907 = pi0695 & n8906;
  assign n8908 = n8904 & n8907;
  assign n8909 = n8903 & ~n8908;
  assign n8910 = pi0382 & n8905;
  assign n8911 = ~pi0695 & n8910;
  assign n8912 = ~n8874 & n8911;
  assign n8913 = ~n5422 & ~n8912;
  assign n8914 = ~n5423 & n8893;
  assign n8915 = pi0382 & n5423;
  assign n8916 = ~n8914 & ~n8915;
  assign n8917 = ~n8913 & ~n8916;
  assign n8918 = n8909 & ~n8917;
  assign po0492 = pi1747 & ~n8918;
  assign n8920 = pi0383 & n8704;
  assign n8921 = pi0384 & pi0481;
  assign n8922 = ~pi0482 & ~pi1267;
  assign n8923 = ~pi0441 & ~pi1119;
  assign n8924 = ~n8922 & ~n8923;
  assign n8925 = n8921 & n8924;
  assign n8926 = ~pi0510 & ~pi1274;
  assign n8927 = ~pi0388 & ~pi1270;
  assign n8928 = ~n8926 & ~n8927;
  assign n8929 = pi0442 & pi1121;
  assign n8930 = ~pi0442 & ~pi1121;
  assign n8931 = pi0413 & pi1272;
  assign n8932 = ~n8930 & n8931;
  assign n8933 = ~n8929 & ~n8932;
  assign n8934 = n8928 & ~n8933;
  assign n8935 = pi0388 & pi1270;
  assign n8936 = pi0510 & pi1274;
  assign n8937 = ~n8927 & n8936;
  assign n8938 = ~n8935 & ~n8937;
  assign n8939 = ~n8934 & n8938;
  assign n8940 = n8925 & ~n8939;
  assign n8941 = pi0441 & pi1119;
  assign n8942 = pi0482 & pi1267;
  assign n8943 = ~n8923 & n8942;
  assign n8944 = ~n8941 & ~n8943;
  assign n8945 = n8921 & ~n8944;
  assign n8946 = ~n8940 & ~n8945;
  assign n8947 = ~pi0413 & ~pi1272;
  assign n8948 = ~n8930 & ~n8947;
  assign n8949 = n8928 & n8948;
  assign n8950 = n8925 & n8949;
  assign n8951 = pi0412 & pi1023;
  assign n8952 = ~pi0412 & ~pi1023;
  assign n8953 = pi0411 & pi1277;
  assign n8954 = ~n8952 & n8953;
  assign n8955 = ~n8951 & ~n8954;
  assign n8956 = ~pi0411 & ~pi1277;
  assign n8957 = ~n8952 & ~n8956;
  assign n8958 = pi0410 & pi1022;
  assign n8959 = n8957 & n8958;
  assign n8960 = n8955 & ~n8959;
  assign n8961 = n8950 & ~n8960;
  assign n8962 = n8946 & ~n8961;
  assign n8963 = pi0383 & n8962;
  assign n8964 = ~pi0383 & ~n8962;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = ~n8704 & ~n8965;
  assign n8967 = ~n8920 & ~n8966;
  assign n8968 = pi1690 & ~n8967;
  assign n8969 = ~pi0384 & ~pi0441;
  assign n8970 = ~pi0481 & ~pi0482;
  assign n8971 = ~pi0410 & ~pi0411;
  assign n8972 = ~pi0412 & n8971;
  assign n8973 = ~pi0413 & n8972;
  assign n8974 = ~pi0442 & ~pi0510;
  assign n8975 = ~pi0388 & n8974;
  assign n8976 = n8973 & n8975;
  assign n8977 = n8970 & n8976;
  assign n8978 = n8969 & n8977;
  assign n8979 = pi0383 & n8978;
  assign n8980 = ~pi0383 & ~n8978;
  assign n8981 = ~n8979 & ~n8980;
  assign n8982 = ~pi1690 & n8981;
  assign n8983 = ~n8968 & ~n8982;
  assign po0493 = pi1122 & ~n8983;
  assign n8985 = pi0384 & n8704;
  assign n8986 = n8948 & ~n8955;
  assign n8987 = n8933 & ~n8986;
  assign n8988 = n8928 & ~n8987;
  assign n8989 = n8938 & ~n8988;
  assign n8990 = n8924 & ~n8989;
  assign n8991 = n8944 & ~n8990;
  assign n8992 = n8924 & n8928;
  assign n8993 = ~n8952 & n8958;
  assign n8994 = n8948 & n8993;
  assign n8995 = ~n8956 & n8994;
  assign n8996 = n8992 & n8995;
  assign n8997 = n8991 & ~n8996;
  assign n8998 = pi0384 & n8997;
  assign n8999 = ~pi0384 & ~n8997;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = ~n8704 & ~n9000;
  assign n9002 = ~n8985 & ~n9001;
  assign n9003 = pi1690 & ~n9002;
  assign n9004 = ~pi0482 & ~pi0510;
  assign n9005 = ~pi0410 & ~pi0442;
  assign n9006 = ~pi0412 & ~pi0413;
  assign n9007 = ~pi0411 & n9006;
  assign n9008 = n9005 & n9007;
  assign n9009 = ~pi0441 & n9008;
  assign n9010 = ~pi0388 & n9009;
  assign n9011 = n9004 & n9010;
  assign n9012 = pi0384 & n9011;
  assign n9013 = ~pi0384 & ~n9011;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~pi1690 & n9014;
  assign n9016 = ~n9003 & ~n9015;
  assign po0494 = pi1122 & ~n9016;
  assign n9018 = pi0385 & ~po1343;
  assign n9019 = pi0897 & po1538;
  assign n9020 = ~n9018 & ~n9019;
  assign n9021 = ~pi0899 & n6299;
  assign n9022 = pi0898 & n6302;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = pi0896 & n6305;
  assign n9025 = n9023 & ~n9024;
  assign po0495 = ~n9020 | ~n9025;
  assign n9027 = pi0386 & n8704;
  assign n9028 = ~n8708 & ~n8711;
  assign n9029 = n8839 & ~n8844;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = n9028 & n9029;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = ~n8704 & ~n9032;
  assign n9034 = ~n9027 & ~n9033;
  assign n9035 = pi1690 & ~n9034;
  assign n9036 = pi0386 & n8860;
  assign n9037 = ~pi0386 & ~n8860;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~pi1690 & n9038;
  assign n9040 = ~n9035 & ~n9039;
  assign po0496 = pi1122 & ~n9040;
  assign n9042 = pi0387 & n8704;
  assign n9043 = ~n8713 & ~n8714;
  assign n9044 = ~n8721 & n8728;
  assign n9045 = ~n8726 & ~n9044;
  assign n9046 = ~n8718 & ~n8720;
  assign n9047 = ~n9045 & n9046;
  assign n9048 = ~n8718 & n8723;
  assign n9049 = ~n8715 & ~n9048;
  assign n9050 = ~n9047 & n9049;
  assign n9051 = ~n8721 & ~n8729;
  assign n9052 = n9046 & n9051;
  assign n9053 = ~n8743 & ~n8746;
  assign n9054 = ~n8730 & ~n9053;
  assign n9055 = n9052 & ~n9054;
  assign n9056 = n9050 & ~n9055;
  assign n9057 = ~n9043 & ~n9056;
  assign n9058 = n9043 & n9056;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = ~n8704 & ~n9059;
  assign n9061 = ~n9042 & ~n9060;
  assign n9062 = pi1690 & ~n9061;
  assign n9063 = ~pi0387 & ~n8859;
  assign n9064 = ~n8860 & ~n9063;
  assign n9065 = ~pi1690 & n9064;
  assign n9066 = ~n9062 & ~n9065;
  assign po0497 = pi1122 & ~n9066;
  assign n9068 = pi0388 & n8704;
  assign n9069 = ~n8927 & ~n8935;
  assign n9070 = ~n8926 & ~n8930;
  assign n9071 = ~n8947 & n8951;
  assign n9072 = ~n8931 & ~n9071;
  assign n9073 = n9070 & ~n9072;
  assign n9074 = ~n8926 & n8929;
  assign n9075 = ~n8936 & ~n9074;
  assign n9076 = ~n9073 & n9075;
  assign n9077 = ~n8956 & n8958;
  assign n9078 = ~n8953 & ~n9077;
  assign n9079 = ~n8947 & ~n8952;
  assign n9080 = n9070 & n9079;
  assign n9081 = ~n9078 & n9080;
  assign n9082 = n9076 & ~n9081;
  assign n9083 = n9069 & n9082;
  assign n9084 = ~n9069 & ~n9082;
  assign n9085 = ~n9083 & ~n9084;
  assign n9086 = ~n8704 & ~n9085;
  assign n9087 = ~n9068 & ~n9086;
  assign n9088 = pi1690 & ~n9087;
  assign n9089 = n8971 & n8974;
  assign n9090 = n9006 & n9089;
  assign n9091 = pi0388 & n9090;
  assign n9092 = ~pi0388 & ~n9090;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = ~pi1690 & n9093;
  assign n9095 = ~n9088 & ~n9094;
  assign po0498 = pi1122 & ~n9095;
  assign n9097 = ~pi0389 & n8084;
  assign n9098 = pi0064 & ~n8084;
  assign n9099 = ~n9097 & ~n9098;
  assign n9100 = ~n8081 & ~n9099;
  assign n9101 = pi1774 & n8081;
  assign n9102 = ~n9100 & ~n9101;
  assign po0499 = ~pi1747 | ~n9102;
  assign n9104 = ~pi0390 & n8084;
  assign n9105 = pi0014 & ~n8084;
  assign n9106 = ~n9104 & ~n9105;
  assign n9107 = ~n8081 & ~n9106;
  assign n9108 = pi1786 & n8081;
  assign n9109 = ~n9107 & ~n9108;
  assign po0500 = ~pi1747 | ~n9109;
  assign n9111 = ~pi0391 & n8084;
  assign n9112 = pi0015 & ~n8084;
  assign n9113 = ~n9111 & ~n9112;
  assign n9114 = ~n8081 & ~n9113;
  assign n9115 = pi1790 & n8081;
  assign n9116 = ~n9114 & ~n9115;
  assign po0501 = ~pi1747 | ~n9116;
  assign n9118 = ~pi0392 & n8084;
  assign n9119 = pi0953 & ~n8084;
  assign n9120 = ~n9118 & ~n9119;
  assign n9121 = ~n8081 & ~n9120;
  assign n9122 = pi1791 & n8081;
  assign n9123 = ~n9121 & ~n9122;
  assign po0502 = ~pi1747 | ~n9123;
  assign n9125 = ~pi0393 & n8084;
  assign n9126 = pi0332 & ~n8084;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = ~n8081 & ~n9127;
  assign n9129 = pi1793 & n8081;
  assign n9130 = ~n9128 & ~n9129;
  assign po0503 = ~pi1747 | ~n9130;
  assign n9132 = ~pi0394 & n8084;
  assign n9133 = pi0057 & ~n8084;
  assign n9134 = ~n9132 & ~n9133;
  assign n9135 = ~n8081 & ~n9134;
  assign n9136 = pi1775 & n8081;
  assign n9137 = ~n9135 & ~n9136;
  assign po0504 = ~pi1747 | ~n9137;
  assign n9139 = ~pi0395 & n8084;
  assign n9140 = pi0299 & ~n8084;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = ~n8081 & ~n9141;
  assign n9143 = pi1794 & n8081;
  assign n9144 = ~n9142 & ~n9143;
  assign po0505 = ~pi1747 | ~n9144;
  assign n9146 = ~pi0396 & n8084;
  assign n9147 = pi1481 & ~n8084;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n8081 & ~n9148;
  assign n9150 = pi1796 & n8081;
  assign n9151 = ~n9149 & ~n9150;
  assign po0506 = ~pi1747 | ~n9151;
  assign n9153 = ~pi0397 & n8084;
  assign n9154 = pi0223 & ~n8084;
  assign n9155 = ~n9153 & ~n9154;
  assign n9156 = ~n8081 & ~n9155;
  assign n9157 = pi1798 & n8081;
  assign n9158 = ~n9156 & ~n9157;
  assign po0507 = ~pi1747 | ~n9158;
  assign n9160 = ~pi0398 & n8084;
  assign n9161 = pi0154 & ~n8084;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = ~n8081 & ~n9162;
  assign n9164 = pi1799 & n8081;
  assign n9165 = ~n9163 & ~n9164;
  assign po0508 = ~pi1747 | ~n9165;
  assign n9167 = ~pi0399 & n8084;
  assign n9168 = pi0254 & ~n8084;
  assign n9169 = ~n9167 & ~n9168;
  assign n9170 = ~n8081 & ~n9169;
  assign n9171 = pi1797 & n8081;
  assign n9172 = ~n9170 & ~n9171;
  assign po0509 = ~pi1747 | ~n9172;
  assign n9174 = ~pi0400 & n8084;
  assign n9175 = pi0124 & ~n8084;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = ~n8081 & ~n9176;
  assign n9178 = pi1801 & n8081;
  assign n9179 = ~n9177 & ~n9178;
  assign po0510 = ~pi1747 | ~n9179;
  assign n9181 = ~pi0401 & n8084;
  assign n9182 = pi0155 & ~n8084;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = ~n8081 & ~n9183;
  assign n9185 = pi1800 & n8081;
  assign n9186 = ~n9184 & ~n9185;
  assign po0511 = ~pi1747 | ~n9186;
  assign n9188 = ~pi0402 & n8084;
  assign n9189 = pi0056 & ~n8084;
  assign n9190 = ~n9188 & ~n9189;
  assign n9191 = ~n8081 & ~n9190;
  assign n9192 = pi1776 & n8081;
  assign n9193 = ~n9191 & ~n9192;
  assign po0512 = ~pi1747 | ~n9193;
  assign n9195 = ~pi0403 & n8084;
  assign n9196 = pi0063 & ~n8084;
  assign n9197 = ~n9195 & ~n9196;
  assign n9198 = ~n8081 & ~n9197;
  assign n9199 = pi1804 & n8081;
  assign n9200 = ~n9198 & ~n9199;
  assign po0513 = ~pi1747 | ~n9200;
  assign n9202 = ~pi0404 & n8084;
  assign n9203 = pi0027 & ~n8084;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = ~n8081 & ~n9204;
  assign n9206 = pi1782 & n8081;
  assign n9207 = ~n9205 & ~n9206;
  assign po0514 = ~pi1747 | ~n9207;
  assign n9209 = ~pi0405 & n8084;
  assign n9210 = pi0022 & ~n8084;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = ~n8081 & ~n9211;
  assign n9213 = pi1783 & n8081;
  assign n9214 = ~n9212 & ~n9213;
  assign po0515 = ~pi1747 | ~n9214;
  assign n9216 = ~pi1672 & ~n8405;
  assign n9217 = ~pi0406 & n8405;
  assign n9218 = ~n9216 & ~n9217;
  assign n9219 = ~n8402 & ~n9218;
  assign n9220 = pi1802 & n8402;
  assign n9221 = ~n9219 & ~n9220;
  assign po0516 = ~pi1747 | ~n9221;
  assign n9223 = ~pi1666 & ~n8405;
  assign n9224 = ~pi0407 & n8405;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n8402 & ~n9225;
  assign n9227 = pi1805 & n8402;
  assign n9228 = ~n9226 & ~n9227;
  assign po0517 = ~pi1747 | ~n9228;
  assign n9230 = pi0408 & n8704;
  assign n9231 = pi0408 & ~pi1022;
  assign n9232 = ~n8746 & ~n9231;
  assign n9233 = ~n8704 & ~n9232;
  assign n9234 = ~n9230 & ~n9233;
  assign n9235 = pi1690 & ~n9234;
  assign n9236 = ~pi0408 & ~pi1690;
  assign n9237 = ~n9235 & ~n9236;
  assign po0518 = pi1122 & ~n9237;
  assign n9239 = pi0409 & pi1250;
  assign n9240 = ~pi0258 & ~n9239;
  assign n9241 = n7510 & ~n9240;
  assign n9242 = ~pi0138 & n9241;
  assign n9243 = ~pi1101 & n7960;
  assign n9244 = ~n8212 & ~n9243;
  assign n9245 = pi0409 & ~n9244;
  assign n9246 = ~n9242 & ~n9245;
  assign po0519 = pi1747 & ~n9246;
  assign n9248 = pi0410 & n8704;
  assign n9249 = ~pi0410 & pi1022;
  assign n9250 = pi0410 & ~pi1022;
  assign n9251 = ~n9249 & ~n9250;
  assign n9252 = ~n8704 & ~n9251;
  assign n9253 = ~n9248 & ~n9252;
  assign n9254 = pi1690 & ~n9253;
  assign n9255 = ~pi0410 & ~pi1690;
  assign n9256 = ~n9254 & ~n9255;
  assign po0520 = pi1122 & ~n9256;
  assign n9258 = pi0411 & n8704;
  assign n9259 = ~n8953 & ~n8956;
  assign n9260 = n8958 & ~n9259;
  assign n9261 = ~n8958 & n9259;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~n8704 & ~n9262;
  assign n9264 = ~n9258 & ~n9263;
  assign n9265 = pi1690 & ~n9264;
  assign n9266 = pi0410 & pi0411;
  assign n9267 = ~n8971 & ~n9266;
  assign n9268 = ~pi1690 & ~n9267;
  assign n9269 = ~n9265 & ~n9268;
  assign po0521 = pi1122 & ~n9269;
  assign n9271 = pi0412 & n8704;
  assign n9272 = ~n8951 & ~n8952;
  assign n9273 = ~n9078 & ~n9272;
  assign n9274 = n9078 & n9272;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = ~n8704 & ~n9275;
  assign n9277 = ~n9271 & ~n9276;
  assign n9278 = pi1690 & ~n9277;
  assign n9279 = pi0412 & ~n8971;
  assign n9280 = ~n8972 & ~n9279;
  assign n9281 = ~pi1690 & ~n9280;
  assign n9282 = ~n9278 & ~n9281;
  assign po0522 = pi1122 & ~n9282;
  assign n9284 = pi0413 & n8704;
  assign n9285 = ~n8931 & ~n8947;
  assign n9286 = ~n8960 & ~n9285;
  assign n9287 = n8960 & n9285;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = ~n8704 & ~n9288;
  assign n9290 = ~n9284 & ~n9289;
  assign n9291 = pi1690 & ~n9290;
  assign n9292 = pi0413 & ~n8972;
  assign n9293 = ~n8973 & ~n9292;
  assign n9294 = ~pi1690 & ~n9293;
  assign n9295 = ~n9291 & ~n9294;
  assign po0523 = pi1122 & ~n9295;
  assign n9297 = pi1790 & n8356;
  assign n9298 = ~pi1190 & n8358;
  assign n9299 = pi0015 & n8360;
  assign n9300 = ~pi0414 & ~n8360;
  assign n9301 = ~n9299 & ~n9300;
  assign n9302 = ~n8358 & ~n9301;
  assign n9303 = ~n9298 & ~n9302;
  assign n9304 = ~n8356 & ~n9303;
  assign n9305 = pi1747 & ~n9304;
  assign po0524 = n9297 | ~n9305;
  assign n9307 = pi1792 & n8356;
  assign n9308 = ~pi1191 & n8358;
  assign n9309 = pi0310 & n8360;
  assign n9310 = ~pi0415 & ~n8360;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = ~n8358 & ~n9311;
  assign n9313 = ~n9308 & ~n9312;
  assign n9314 = ~n8356 & ~n9313;
  assign n9315 = pi1747 & ~n9314;
  assign po0525 = n9307 | ~n9315;
  assign n9317 = pi1793 & n8356;
  assign n9318 = pi1192 & n8358;
  assign n9319 = pi0332 & n8360;
  assign n9320 = ~pi0416 & ~n8360;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = ~n8358 & ~n9321;
  assign n9323 = ~n9318 & ~n9322;
  assign n9324 = ~n8356 & ~n9323;
  assign n9325 = pi1747 & ~n9324;
  assign po0526 = n9317 | ~n9325;
  assign n9327 = pi1775 & n8356;
  assign n9328 = ~pi1193 & n8358;
  assign n9329 = pi0057 & n8360;
  assign n9330 = ~pi0417 & ~n8360;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~n8358 & ~n9331;
  assign n9333 = ~n9328 & ~n9332;
  assign n9334 = ~n8356 & ~n9333;
  assign n9335 = pi1747 & ~n9334;
  assign po0527 = n9327 | ~n9335;
  assign n9337 = pi1794 & n8356;
  assign n9338 = pi1276 & n8358;
  assign n9339 = pi0299 & n8360;
  assign n9340 = ~pi0418 & ~n8360;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n8358 & ~n9341;
  assign n9343 = ~n9338 & ~n9342;
  assign n9344 = ~n8356 & ~n9343;
  assign n9345 = pi1747 & ~n9344;
  assign po0528 = n9337 | ~n9345;
  assign n9347 = pi1795 & n8356;
  assign n9348 = pi1194 & n8358;
  assign n9349 = pi0286 & n8360;
  assign n9350 = ~pi0419 & ~n8360;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n8358 & ~n9351;
  assign n9353 = ~n9348 & ~n9352;
  assign n9354 = ~n8356 & ~n9353;
  assign n9355 = pi1747 & ~n9354;
  assign po0529 = n9347 | ~n9355;
  assign n9357 = pi1797 & n8356;
  assign n9358 = pi1196 & n8358;
  assign n9359 = pi0254 & n8360;
  assign n9360 = ~pi0420 & ~n8360;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n8358 & ~n9361;
  assign n9363 = ~n9358 & ~n9362;
  assign n9364 = ~n8356 & ~n9363;
  assign n9365 = pi1747 & ~n9364;
  assign po0530 = n9357 | ~n9365;
  assign n9367 = pi1798 & n8356;
  assign n9368 = pi1264 & n8358;
  assign n9369 = pi0223 & n8360;
  assign n9370 = ~pi0421 & ~n8360;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n8358 & ~n9371;
  assign n9373 = ~n9368 & ~n9372;
  assign n9374 = ~n8356 & ~n9373;
  assign n9375 = pi1747 & ~n9374;
  assign po0531 = n9367 | ~n9375;
  assign n9377 = pi1799 & n8356;
  assign n9378 = pi1197 & n8358;
  assign n9379 = pi0154 & n8360;
  assign n9380 = ~pi0422 & ~n8360;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = ~n8358 & ~n9381;
  assign n9383 = ~n9378 & ~n9382;
  assign n9384 = ~n8356 & ~n9383;
  assign n9385 = pi1747 & ~n9384;
  assign po0532 = n9377 | ~n9385;
  assign n9387 = pi1801 & n8356;
  assign n9388 = pi1199 & n8358;
  assign n9389 = pi0124 & n8360;
  assign n9390 = ~pi0423 & ~n8360;
  assign n9391 = ~n9389 & ~n9390;
  assign n9392 = ~n8358 & ~n9391;
  assign n9393 = ~n9388 & ~n9392;
  assign n9394 = ~n8356 & ~n9393;
  assign n9395 = pi1747 & ~n9394;
  assign po0533 = n9387 | ~n9395;
  assign n9397 = pi1804 & n8356;
  assign n9398 = pi1036 & n8358;
  assign n9399 = pi0063 & n8360;
  assign n9400 = ~pi0424 & ~n8360;
  assign n9401 = ~n9399 & ~n9400;
  assign n9402 = ~n8358 & ~n9401;
  assign n9403 = ~n9398 & ~n9402;
  assign n9404 = ~n8356 & ~n9403;
  assign n9405 = pi1747 & ~n9404;
  assign po0534 = n9397 | ~n9405;
  assign n9407 = pi1777 & n8356;
  assign n9408 = ~pi1202 & n8358;
  assign n9409 = pi0049 & n8360;
  assign n9410 = ~pi0425 & ~n8360;
  assign n9411 = ~n9409 & ~n9410;
  assign n9412 = ~n8358 & ~n9411;
  assign n9413 = ~n9408 & ~n9412;
  assign n9414 = ~n8356 & ~n9413;
  assign n9415 = pi1747 & ~n9414;
  assign po0535 = n9407 | ~n9415;
  assign n9417 = pi1783 & n8356;
  assign n9418 = ~pi1240 & n8358;
  assign n9419 = pi0022 & n8360;
  assign n9420 = ~pi0426 & ~n8360;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n8358 & ~n9421;
  assign n9423 = ~n9418 & ~n9422;
  assign n9424 = ~n8356 & ~n9423;
  assign n9425 = pi1747 & ~n9424;
  assign po0536 = n9417 | ~n9425;
  assign n9427 = pi1761 & pi1762;
  assign n9428 = n8002 & n9427;
  assign n9429 = n8005 & n9428;
  assign n9430 = n7999 & n9429;
  assign n9431 = pi1802 & n9430;
  assign n9432 = pi1057 & n8414;
  assign n9433 = ~pi0427 & ~n8413;
  assign n9434 = ~pi1672 & n8413;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = ~n8414 & ~n9435;
  assign n9437 = ~n9432 & ~n9436;
  assign n9438 = ~n9430 & ~n9437;
  assign n9439 = pi1747 & ~n9438;
  assign po0537 = n9431 | ~n9439;
  assign n9441 = pi1805 & n9430;
  assign n9442 = ~pi1221 & n8414;
  assign n9443 = ~pi0428 & ~n8413;
  assign n9444 = ~pi1666 & n8413;
  assign n9445 = ~n9443 & ~n9444;
  assign n9446 = ~n8414 & ~n9445;
  assign n9447 = ~n9442 & ~n9446;
  assign n9448 = ~n9430 & ~n9447;
  assign n9449 = pi1747 & ~n9448;
  assign po0538 = n9441 | ~n9449;
  assign n9451 = pi0269 & ~pi1039;
  assign n9452 = ~pi0269 & pi1039;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = pi0271 & ~pi1040;
  assign n9455 = ~pi0271 & pi1040;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = pi0270 & ~pi1041;
  assign n9458 = ~pi0270 & pi1041;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = pi0272 & ~pi1049;
  assign n9461 = ~pi0272 & pi1049;
  assign n9462 = ~n9460 & ~n9461;
  assign n9463 = n9459 & n9462;
  assign n9464 = n9456 & n9463;
  assign n9465 = n9453 & n9464;
  assign n9466 = pi0250 & ~pi1318;
  assign n9467 = ~pi0250 & pi1318;
  assign n9468 = ~n9466 & ~n9467;
  assign n9469 = n9465 & n9468;
  assign n9470 = pi0255 & ~pi1317;
  assign n9471 = ~pi0255 & pi1317;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = pi0253 & ~pi1313;
  assign n9474 = ~pi0253 & pi1313;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = n9472 & n9475;
  assign n9477 = pi0251 & ~pi1042;
  assign n9478 = ~pi0251 & pi1042;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = pi0263 & ~pi1043;
  assign n9481 = ~pi0263 & pi1043;
  assign n9482 = ~n9480 & ~n9481;
  assign n9483 = n9479 & n9482;
  assign n9484 = pi0273 & ~pi1017;
  assign n9485 = ~pi0273 & pi1017;
  assign n9486 = ~n9484 & ~n9485;
  assign n9487 = n9483 & n9486;
  assign n9488 = pi1233 & n4135;
  assign po0815 = ~po1002 & n9488;
  assign n9490 = pi0252 & ~pi1044;
  assign n9491 = ~pi0252 & pi1044;
  assign n9492 = ~n9490 & ~n9491;
  assign n9493 = po0815 & n9492;
  assign n9494 = n9487 & n9493;
  assign n9495 = n9476 & n9494;
  assign po0539 = n9469 & n9495;
  assign n9497 = ~pi0430 & n8084;
  assign n9498 = pi0310 & ~n8084;
  assign n9499 = ~n9497 & ~n9498;
  assign n9500 = ~n8081 & ~n9499;
  assign n9501 = pi1792 & n8081;
  assign n9502 = ~n9500 & ~n9501;
  assign po0540 = ~pi1747 | ~n9502;
  assign n9504 = ~n5848 & ~n5849;
  assign n9505 = n7074 & ~n7076;
  assign n9506 = n7092 & ~n9505;
  assign n9507 = ~n9504 & ~n9506;
  assign n9508 = n9504 & n9506;
  assign po0541 = n9507 | n9508;
  assign n9510 = pi1800 & n8356;
  assign n9511 = pi1198 & n8358;
  assign n9512 = pi0155 & n8360;
  assign n9513 = ~pi0432 & ~n8360;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = ~n8358 & ~n9514;
  assign n9516 = ~n9511 & ~n9515;
  assign n9517 = ~n8356 & ~n9516;
  assign n9518 = pi1747 & ~n9517;
  assign po0542 = n9510 | ~n9518;
  assign n9520 = pi0469 & pi0474;
  assign n9521 = pi0433 & ~n9520;
  assign n9522 = ~pi0433 & n9520;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = pi1671 & ~n9523;
  assign n9525 = pi0433 & ~pi1671;
  assign n9526 = ~n9524 & ~n9525;
  assign po0543 = ~pi0705 & ~n9526;
  assign n9528 = pi1776 & n8007;
  assign n9529 = ~pi1178 & n8009;
  assign n9530 = pi0056 & n8011;
  assign n9531 = ~pi0435 & ~n8011;
  assign n9532 = ~n9530 & ~n9531;
  assign n9533 = ~n8009 & ~n9532;
  assign n9534 = ~n9529 & ~n9533;
  assign n9535 = ~n8007 & ~n9534;
  assign n9536 = pi1747 & ~n9535;
  assign po0545 = n9528 | ~n9536;
  assign n9538 = pi1782 & n9430;
  assign n9539 = ~pi1279 & n8414;
  assign n9540 = pi0027 & n8413;
  assign n9541 = ~pi0436 & ~n8413;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = ~n8414 & ~n9542;
  assign n9544 = ~n9539 & ~n9543;
  assign n9545 = ~n9430 & ~n9544;
  assign n9546 = pi1747 & ~n9545;
  assign po0546 = n9538 | ~n9546;
  assign n9548 = n8353 & n9427;
  assign n9549 = n8005 & n9548;
  assign n9550 = n7999 & n9549;
  assign n9551 = pi1805 & n9550;
  assign n9552 = ~pi1161 & n8483;
  assign n9553 = ~pi0437 & ~n8482;
  assign n9554 = ~pi1666 & n8482;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = ~n8483 & ~n9555;
  assign n9557 = ~n9552 & ~n9556;
  assign n9558 = ~n9550 & ~n9557;
  assign n9559 = pi1747 & ~n9558;
  assign po0547 = n9551 | ~n9559;
  assign n9561 = pi1796 & n8007;
  assign n9562 = pi1087 & n8009;
  assign n9563 = pi1481 & n8011;
  assign n9564 = ~pi0438 & ~n8011;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = ~n8009 & ~n9565;
  assign n9567 = ~n9562 & ~n9566;
  assign n9568 = ~n8007 & ~n9567;
  assign n9569 = pi1747 & ~n9568;
  assign po0548 = n9561 | ~n9569;
  assign n9571 = pi1786 & n9430;
  assign n9572 = ~pi1086 & n8414;
  assign n9573 = pi0014 & n8413;
  assign n9574 = ~pi0439 & ~n8413;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = ~n8414 & ~n9575;
  assign n9577 = ~n9572 & ~n9576;
  assign n9578 = ~n9430 & ~n9577;
  assign n9579 = pi1747 & ~n9578;
  assign po0549 = n9571 | ~n9579;
  assign n9581 = ~pi0440 & n8405;
  assign n9582 = pi0057 & ~n8405;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = ~n8402 & ~n9583;
  assign n9585 = pi1775 & n8402;
  assign n9586 = ~n9584 & ~n9585;
  assign po0550 = ~pi1747 | ~n9586;
  assign n9588 = ~pi0388 & ~pi0482;
  assign n9589 = n8974 & n9588;
  assign n9590 = n8973 & n9589;
  assign n9591 = pi0441 & ~n9590;
  assign n9592 = ~pi0441 & n9590;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = ~pi1690 & ~n9593;
  assign n9595 = pi0441 & n8704;
  assign n9596 = ~n8923 & ~n8941;
  assign n9597 = ~n8922 & n8935;
  assign n9598 = ~n8942 & ~n9597;
  assign n9599 = ~n9078 & n9079;
  assign n9600 = n9072 & ~n9599;
  assign n9601 = n9070 & ~n9600;
  assign n9602 = n9075 & ~n9601;
  assign n9603 = ~n8922 & ~n8927;
  assign n9604 = ~n9602 & n9603;
  assign n9605 = n9598 & ~n9604;
  assign n9606 = ~n9596 & ~n9605;
  assign n9607 = n9596 & n9605;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~n8704 & ~n9608;
  assign n9610 = ~n9595 & ~n9609;
  assign n9611 = pi1690 & ~n9610;
  assign n9612 = ~n9594 & ~n9611;
  assign po0551 = pi1122 & ~n9612;
  assign n9614 = pi0442 & ~n8973;
  assign n9615 = ~pi0442 & n8973;
  assign n9616 = ~n9614 & ~n9615;
  assign n9617 = ~pi1690 & ~n9616;
  assign n9618 = pi0442 & n8704;
  assign n9619 = ~n8929 & ~n8930;
  assign n9620 = ~n9600 & ~n9619;
  assign n9621 = n9600 & n9619;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = ~n8704 & ~n9622;
  assign n9624 = ~n9618 & ~n9623;
  assign n9625 = pi1690 & ~n9624;
  assign n9626 = ~n9617 & ~n9625;
  assign po0552 = pi1122 & ~n9626;
  assign n9628 = ~pi0443 & n8405;
  assign n9629 = pi0022 & ~n8405;
  assign n9630 = ~n9628 & ~n9629;
  assign n9631 = ~n8402 & ~n9630;
  assign n9632 = pi1783 & n8402;
  assign n9633 = ~n9631 & ~n9632;
  assign po0553 = ~pi1747 | ~n9633;
  assign n9635 = pi1793 & n9430;
  assign n9636 = pi1213 & n8414;
  assign n9637 = pi0332 & n8413;
  assign n9638 = ~pi0444 & ~n8413;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = ~n8414 & ~n9639;
  assign n9641 = ~n9636 & ~n9640;
  assign n9642 = ~n9430 & ~n9641;
  assign n9643 = pi1747 & ~n9642;
  assign po0554 = n9635 | ~n9643;
  assign n9645 = ~pi0445 & n8405;
  assign n9646 = pi0124 & ~n8405;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = ~n8402 & ~n9647;
  assign n9649 = pi1801 & n8402;
  assign n9650 = ~n9648 & ~n9649;
  assign po0555 = ~pi1747 | ~n9650;
  assign n9652 = ~pi0446 & n8405;
  assign n9653 = pi0254 & ~n8405;
  assign n9654 = ~n9652 & ~n9653;
  assign n9655 = ~n8402 & ~n9654;
  assign n9656 = pi1797 & n8402;
  assign n9657 = ~n9655 & ~n9656;
  assign po0556 = ~pi1747 | ~n9657;
  assign n9659 = pi1779 & n8007;
  assign n9660 = ~pi1181 & n8009;
  assign n9661 = pi0028 & n8011;
  assign n9662 = ~pi0447 & ~n8011;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = ~n8009 & ~n9663;
  assign n9665 = ~n9660 & ~n9664;
  assign n9666 = ~n8007 & ~n9665;
  assign n9667 = pi1747 & ~n9666;
  assign po0557 = n9659 | ~n9667;
  assign n9669 = pi0476 & pi0477;
  assign n9670 = pi0475 & n9669;
  assign n9671 = pi0433 & n9520;
  assign n9672 = n9670 & n9671;
  assign n9673 = pi0448 & ~n9672;
  assign n9674 = ~pi0448 & n9672;
  assign n9675 = ~n9673 & ~n9674;
  assign n9676 = pi1671 & ~n9675;
  assign n9677 = pi0448 & ~pi1671;
  assign n9678 = ~n9676 & ~n9677;
  assign po0558 = ~pi0705 & ~n9678;
  assign n9680 = pi1780 & n9430;
  assign n9681 = ~pi1278 & n8414;
  assign n9682 = pi0023 & n8413;
  assign n9683 = ~pi0449 & ~n8413;
  assign n9684 = ~n9682 & ~n9683;
  assign n9685 = ~n8414 & ~n9684;
  assign n9686 = ~n9681 & ~n9685;
  assign n9687 = ~n9430 & ~n9686;
  assign n9688 = pi1747 & ~n9687;
  assign po0559 = n9680 | ~n9688;
  assign n9690 = pi1785 & n9430;
  assign n9691 = ~pi1208 & n8414;
  assign n9692 = pi0019 & n8413;
  assign n9693 = ~pi0450 & ~n8413;
  assign n9694 = ~n9692 & ~n9693;
  assign n9695 = ~n8414 & ~n9694;
  assign n9696 = ~n9691 & ~n9695;
  assign n9697 = ~n9430 & ~n9696;
  assign n9698 = pi1747 & ~n9697;
  assign po0560 = n9690 | ~n9698;
  assign n9700 = pi1784 & n9430;
  assign n9701 = ~pi1085 & n8414;
  assign n9702 = pi0016 & n8413;
  assign n9703 = ~pi0451 & ~n8413;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = ~n8414 & ~n9704;
  assign n9706 = ~n9701 & ~n9705;
  assign n9707 = ~n9430 & ~n9706;
  assign n9708 = pi1747 & ~n9707;
  assign po0561 = n9700 | ~n9708;
  assign n9710 = pi1788 & n9430;
  assign n9711 = ~pi1062 & n8414;
  assign n9712 = pi0011 & n8413;
  assign n9713 = ~pi0452 & ~n8413;
  assign n9714 = ~n9712 & ~n9713;
  assign n9715 = ~n8414 & ~n9714;
  assign n9716 = ~n9711 & ~n9715;
  assign n9717 = ~n9430 & ~n9716;
  assign n9718 = pi1747 & ~n9717;
  assign po0562 = n9710 | ~n9718;
  assign n9720 = pi1787 & n9430;
  assign n9721 = ~pi1209 & n8414;
  assign n9722 = pi0007 & n8413;
  assign n9723 = ~pi0453 & ~n8413;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = ~n8414 & ~n9724;
  assign n9726 = ~n9721 & ~n9725;
  assign n9727 = ~n9430 & ~n9726;
  assign n9728 = pi1747 & ~n9727;
  assign po0563 = n9720 | ~n9728;
  assign n9730 = n8080 & n9429;
  assign n9731 = pi1459 & pi1729;
  assign n9732 = pi0996 & pi1459;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = pi0011 & ~n9733;
  assign n9735 = ~pi0454 & n9733;
  assign n9736 = ~n9734 & ~n9735;
  assign n9737 = ~n9730 & ~n9736;
  assign n9738 = pi1788 & n9730;
  assign n9739 = ~n9737 & ~n9738;
  assign po0564 = ~pi1747 | ~n9739;
  assign n9741 = pi1789 & n9430;
  assign n9742 = ~pi1210 & n8414;
  assign n9743 = pi0018 & n8413;
  assign n9744 = ~pi0455 & ~n8413;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = ~n8414 & ~n9745;
  assign n9747 = ~n9742 & ~n9746;
  assign n9748 = ~n9430 & ~n9747;
  assign n9749 = pi1747 & ~n9748;
  assign po0565 = n9741 | ~n9749;
  assign n9751 = pi0016 & ~n9733;
  assign n9752 = ~pi0456 & n9733;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~n9730 & ~n9753;
  assign n9755 = pi1784 & n9730;
  assign n9756 = ~n9754 & ~n9755;
  assign po0566 = ~pi1747 | ~n9756;
  assign n9758 = pi0007 & ~n9733;
  assign n9759 = ~pi0457 & n9733;
  assign n9760 = ~n9758 & ~n9759;
  assign n9761 = ~n9730 & ~n9760;
  assign n9762 = pi1787 & n9730;
  assign n9763 = ~n9761 & ~n9762;
  assign po0567 = ~pi1747 | ~n9763;
  assign n9765 = pi1778 & n8007;
  assign n9766 = ~pi1067 & n8009;
  assign n9767 = pi0046 & n8011;
  assign n9768 = ~pi0458 & ~n8011;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = ~n8009 & ~n9769;
  assign n9771 = ~n9766 & ~n9770;
  assign n9772 = ~n8007 & ~n9771;
  assign n9773 = pi1747 & ~n9772;
  assign po0568 = n9765 | ~n9773;
  assign n9775 = pi1781 & n9430;
  assign n9776 = ~pi1223 & n8414;
  assign n9777 = pi0030 & n8413;
  assign n9778 = ~pi0459 & ~n8413;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = ~n8414 & ~n9779;
  assign n9781 = ~n9776 & ~n9780;
  assign n9782 = ~n9430 & ~n9781;
  assign n9783 = pi1747 & ~n9782;
  assign po0569 = n9775 | ~n9783;
  assign n9785 = pi0019 & ~n9733;
  assign n9786 = ~pi0460 & n9733;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = ~n9730 & ~n9787;
  assign n9789 = pi1785 & n9730;
  assign n9790 = ~n9788 & ~n9789;
  assign po0570 = ~pi1747 | ~n9790;
  assign n9792 = pi0023 & ~n9733;
  assign n9793 = ~pi0461 & n9733;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = ~n9730 & ~n9794;
  assign n9796 = pi1780 & n9730;
  assign n9797 = ~n9795 & ~n9796;
  assign po0571 = ~pi1747 | ~n9797;
  assign n9799 = pi0046 & ~n9733;
  assign n9800 = ~pi0462 & n9733;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = ~n9730 & ~n9801;
  assign n9803 = pi1778 & n9730;
  assign n9804 = ~n9802 & ~n9803;
  assign po0572 = ~pi1747 | ~n9804;
  assign n9806 = pi0028 & ~n9733;
  assign n9807 = ~pi0463 & n9733;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = ~n9730 & ~n9808;
  assign n9810 = pi1779 & n9730;
  assign n9811 = ~n9809 & ~n9810;
  assign po0573 = ~pi1747 | ~n9811;
  assign n9813 = pi0030 & ~n9733;
  assign n9814 = ~pi0464 & n9733;
  assign n9815 = ~n9813 & ~n9814;
  assign n9816 = ~n9730 & ~n9815;
  assign n9817 = pi1781 & n9730;
  assign n9818 = ~n9816 & ~n9817;
  assign po0574 = ~pi1747 | ~n9818;
  assign n9820 = pi0465 & ~pi1671;
  assign n9821 = pi0475 & n9671;
  assign n9822 = pi0476 & n9821;
  assign n9823 = pi0448 & n9822;
  assign n9824 = pi0477 & n9823;
  assign n9825 = pi0478 & pi0479;
  assign n9826 = n9824 & n9825;
  assign n9827 = pi0473 & n9826;
  assign n9828 = pi0467 & n9827;
  assign n9829 = ~pi0465 & n9828;
  assign n9830 = pi0465 & ~n9828;
  assign n9831 = ~n9829 & ~n9830;
  assign n9832 = pi1671 & ~n9831;
  assign n9833 = ~n9820 & ~n9832;
  assign po0575 = ~pi0705 & n9833;
  assign n9835 = n6522 & n6531;
  assign n9836 = n8858 & n9835;
  assign n9837 = pi0466 & ~n9836;
  assign n9838 = ~pi0466 & n9836;
  assign n9839 = ~n9837 & ~n9838;
  assign n9840 = ~pi1690 & ~n9839;
  assign n9841 = pi0466 & n8704;
  assign n9842 = ~n8706 & ~n8707;
  assign n9843 = ~n8711 & n8713;
  assign n9844 = ~n8708 & ~n9843;
  assign n9845 = n9051 & ~n9054;
  assign n9846 = n9045 & ~n9845;
  assign n9847 = n9046 & ~n9846;
  assign n9848 = n9049 & ~n9847;
  assign n9849 = ~n8711 & ~n8714;
  assign n9850 = ~n9848 & n9849;
  assign n9851 = n9844 & ~n9850;
  assign n9852 = n9842 & n9851;
  assign n9853 = ~n9842 & ~n9851;
  assign n9854 = ~n9852 & ~n9853;
  assign n9855 = ~n8704 & ~n9854;
  assign n9856 = ~n9841 & ~n9855;
  assign n9857 = pi1690 & ~n9856;
  assign n9858 = ~n9840 & ~n9857;
  assign po0576 = pi1122 & ~n9858;
  assign n9860 = pi0467 & ~n9824;
  assign n9861 = ~pi0467 & n9824;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = pi1671 & ~n9862;
  assign n9864 = pi0467 & ~pi1671;
  assign n9865 = ~n9863 & ~n9864;
  assign po0577 = ~pi0705 & ~n9865;
  assign n9867 = pi0468 & n8771;
  assign n9868 = n8786 & ~n8792;
  assign n9869 = ~n8794 & n9868;
  assign n9870 = n8784 & ~n9869;
  assign n9871 = n8779 & ~n9870;
  assign n9872 = n8811 & ~n8813;
  assign n9873 = n8799 & ~n9872;
  assign n9874 = n8786 & n8789;
  assign n9875 = ~n9873 & n9874;
  assign n9876 = n8779 & n9875;
  assign n9877 = ~pi0380 & ~pi0562;
  assign n9878 = ~n9876 & n9877;
  assign n9879 = n8777 & n9878;
  assign n9880 = ~n9871 & n9879;
  assign n9881 = pi0468 & ~n9880;
  assign n9882 = ~pi0468 & n9880;
  assign n9883 = ~n9881 & ~n9882;
  assign n9884 = ~n8771 & ~n9883;
  assign n9885 = ~n9867 & ~n9884;
  assign n9886 = pi1679 & ~n9885;
  assign n9887 = pi0506 & pi0618;
  assign n9888 = pi0587 & n9887;
  assign n9889 = pi0622 & n9888;
  assign n9890 = n6354 & n9889;
  assign n9891 = pi0485 & n9890;
  assign n9892 = n6371 & n9891;
  assign n9893 = pi0562 & n9892;
  assign n9894 = pi0483 & n9893;
  assign n9895 = pi0468 & n9894;
  assign n9896 = ~pi0468 & ~n9894;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~pi1679 & n9897;
  assign n9899 = ~n9886 & ~n9898;
  assign po0578 = pi1131 & ~n9899;
  assign n9901 = pi0469 & ~pi1671;
  assign n9902 = ~pi0469 & pi1671;
  assign n9903 = ~n9901 & ~n9902;
  assign po0579 = ~pi0705 & ~n9903;
  assign n9905 = n6522 & n6548;
  assign n9906 = n8859 & n9905;
  assign n9907 = pi0470 & ~n9906;
  assign n9908 = ~pi0470 & n9906;
  assign n9909 = ~n9907 & ~n9908;
  assign n9910 = ~pi1690 & ~n9909;
  assign n9911 = pi0470 & n8704;
  assign n9912 = ~n9050 & n9849;
  assign n9913 = n9844 & ~n9912;
  assign n9914 = ~n8707 & ~n9913;
  assign n9915 = ~pi0379 & ~n8706;
  assign n9916 = ~n9914 & n9915;
  assign n9917 = ~n8707 & n9849;
  assign n9918 = n9055 & n9917;
  assign n9919 = n9916 & ~n9918;
  assign n9920 = pi0470 & ~n9919;
  assign n9921 = ~pi0470 & n9919;
  assign n9922 = ~n9920 & ~n9921;
  assign n9923 = ~n8704 & ~n9922;
  assign n9924 = ~n9911 & ~n9923;
  assign n9925 = pi1690 & ~n9924;
  assign n9926 = ~n9910 & ~n9925;
  assign po0580 = pi1122 & ~n9926;
  assign n9928 = pi0471 & n8771;
  assign n9929 = pi0472 & pi0564;
  assign n9930 = ~pi0565 & ~pi1029;
  assign n9931 = ~pi0560 & ~pi1127;
  assign n9932 = ~n9930 & ~n9931;
  assign n9933 = n9929 & n9932;
  assign n9934 = ~pi0588 & ~pi1130;
  assign n9935 = ~pi0486 & ~pi1076;
  assign n9936 = ~n9934 & ~n9935;
  assign n9937 = pi0541 & pi1083;
  assign n9938 = ~pi0541 & ~pi1083;
  assign n9939 = pi0514 & pi1028;
  assign n9940 = ~n9938 & n9939;
  assign n9941 = ~n9937 & ~n9940;
  assign n9942 = n9936 & ~n9941;
  assign n9943 = pi0486 & pi1076;
  assign n9944 = pi0588 & pi1130;
  assign n9945 = ~n9935 & n9944;
  assign n9946 = ~n9943 & ~n9945;
  assign n9947 = ~n9942 & n9946;
  assign n9948 = n9933 & ~n9947;
  assign n9949 = pi0560 & pi1127;
  assign n9950 = pi0565 & pi1029;
  assign n9951 = ~n9931 & n9950;
  assign n9952 = ~n9949 & ~n9951;
  assign n9953 = n9929 & ~n9952;
  assign n9954 = ~n9948 & ~n9953;
  assign n9955 = ~pi0514 & ~pi1028;
  assign n9956 = ~n9938 & ~n9955;
  assign n9957 = n9936 & n9956;
  assign n9958 = n9933 & n9957;
  assign n9959 = pi0513 & pi1129;
  assign n9960 = ~pi0513 & ~pi1129;
  assign n9961 = pi0512 & pi1310;
  assign n9962 = ~n9960 & n9961;
  assign n9963 = ~n9959 & ~n9962;
  assign n9964 = ~pi0512 & ~pi1310;
  assign n9965 = ~n9960 & ~n9964;
  assign n9966 = pi0511 & pi1027;
  assign n9967 = n9965 & n9966;
  assign n9968 = n9963 & ~n9967;
  assign n9969 = n9958 & ~n9968;
  assign n9970 = n9954 & ~n9969;
  assign n9971 = pi0471 & n9970;
  assign n9972 = ~pi0471 & ~n9970;
  assign n9973 = ~n9971 & ~n9972;
  assign n9974 = ~n8771 & ~n9973;
  assign n9975 = ~n9928 & ~n9974;
  assign n9976 = pi1679 & ~n9975;
  assign n9977 = ~pi0472 & ~pi0560;
  assign n9978 = ~pi0564 & ~pi0565;
  assign n9979 = ~pi0511 & ~pi0512;
  assign n9980 = ~pi0513 & n9979;
  assign n9981 = ~pi0514 & n9980;
  assign n9982 = ~pi0541 & ~pi0588;
  assign n9983 = ~pi0486 & n9982;
  assign n9984 = n9981 & n9983;
  assign n9985 = n9978 & n9984;
  assign n9986 = n9977 & n9985;
  assign n9987 = pi0471 & n9986;
  assign n9988 = ~pi0471 & ~n9986;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = ~pi1679 & n9989;
  assign n9991 = ~n9976 & ~n9990;
  assign po0581 = pi1131 & ~n9991;
  assign n9993 = pi0472 & n8771;
  assign n9994 = n9956 & ~n9963;
  assign n9995 = n9941 & ~n9994;
  assign n9996 = n9936 & ~n9995;
  assign n9997 = n9946 & ~n9996;
  assign n9998 = n9932 & ~n9997;
  assign n9999 = n9952 & ~n9998;
  assign n10000 = n9932 & n9936;
  assign n10001 = ~n9960 & n9966;
  assign n10002 = n9956 & n10001;
  assign n10003 = ~n9964 & n10002;
  assign n10004 = n10000 & n10003;
  assign n10005 = n9999 & ~n10004;
  assign n10006 = pi0472 & n10005;
  assign n10007 = ~pi0472 & ~n10005;
  assign n10008 = ~n10006 & ~n10007;
  assign n10009 = ~n8771 & ~n10008;
  assign n10010 = ~n9993 & ~n10009;
  assign n10011 = pi1679 & ~n10010;
  assign n10012 = ~pi0565 & ~pi0588;
  assign n10013 = ~pi0511 & ~pi0541;
  assign n10014 = ~pi0513 & ~pi0514;
  assign n10015 = ~pi0512 & n10014;
  assign n10016 = n10013 & n10015;
  assign n10017 = ~pi0560 & n10016;
  assign n10018 = ~pi0486 & n10017;
  assign n10019 = n10012 & n10018;
  assign n10020 = pi0472 & n10019;
  assign n10021 = ~pi0472 & ~n10019;
  assign n10022 = ~n10020 & ~n10021;
  assign n10023 = ~pi1679 & n10022;
  assign n10024 = ~n10011 & ~n10023;
  assign po0582 = pi1131 & ~n10024;
  assign n10026 = pi0448 & pi0467;
  assign n10027 = n9825 & n10026;
  assign n10028 = n9672 & n10027;
  assign n10029 = pi0473 & ~n10028;
  assign n10030 = ~pi0473 & n10028;
  assign n10031 = ~n10029 & ~n10030;
  assign n10032 = pi1671 & ~n10031;
  assign n10033 = pi0473 & ~pi1671;
  assign n10034 = ~n10032 & ~n10033;
  assign po0583 = ~pi0705 & ~n10034;
  assign n10036 = pi0469 & ~pi0474;
  assign n10037 = ~pi0469 & pi0474;
  assign n10038 = ~n10036 & ~n10037;
  assign n10039 = pi1671 & ~n10038;
  assign n10040 = pi0474 & ~pi1671;
  assign n10041 = ~n10039 & ~n10040;
  assign po0584 = ~pi0705 & ~n10041;
  assign n10043 = pi0475 & ~n9671;
  assign n10044 = ~pi0475 & n9671;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = pi1671 & ~n10045;
  assign n10047 = pi0475 & ~pi1671;
  assign n10048 = ~n10046 & ~n10047;
  assign po0585 = ~pi0705 & ~n10048;
  assign n10050 = pi0476 & ~n9821;
  assign n10051 = ~pi0476 & n9821;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = pi1671 & ~n10052;
  assign n10054 = pi0476 & ~pi1671;
  assign n10055 = ~n10053 & ~n10054;
  assign po0586 = ~pi0705 & ~n10055;
  assign n10057 = pi0433 & pi0474;
  assign n10058 = pi0476 & n10057;
  assign n10059 = pi0475 & n10058;
  assign n10060 = pi0469 & n10059;
  assign n10061 = pi0477 & ~n10060;
  assign n10062 = ~pi0477 & n10060;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = pi1671 & ~n10063;
  assign n10065 = pi0477 & ~pi1671;
  assign n10066 = ~n10064 & ~n10065;
  assign po0587 = ~pi0705 & ~n10066;
  assign n10068 = pi0469 & pi0477;
  assign n10069 = n10059 & n10068;
  assign n10070 = pi0448 & n10069;
  assign n10071 = pi0479 & n10070;
  assign n10072 = pi0467 & n10071;
  assign n10073 = pi0478 & ~n10072;
  assign n10074 = ~pi0478 & n10072;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076 = pi1671 & ~n10075;
  assign n10077 = pi0478 & ~pi1671;
  assign n10078 = ~n10076 & ~n10077;
  assign po0588 = ~pi0705 & ~n10078;
  assign n10080 = n9669 & n10026;
  assign n10081 = n9821 & n10080;
  assign n10082 = pi0479 & ~n10081;
  assign n10083 = ~pi0479 & n10081;
  assign n10084 = ~n10082 & ~n10083;
  assign n10085 = pi1671 & ~n10084;
  assign n10086 = pi0479 & ~pi1671;
  assign n10087 = ~n10085 & ~n10086;
  assign po0589 = ~pi0705 & ~n10087;
  assign n10089 = pi0408 & n8759;
  assign n10090 = pi0480 & ~n10089;
  assign n10091 = ~pi0480 & n10089;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = ~pi1690 & ~n10092;
  assign n10094 = pi0480 & n8704;
  assign n10095 = ~n8715 & ~n8718;
  assign n10096 = ~n8737 & ~n8747;
  assign n10097 = n10095 & n10096;
  assign n10098 = ~n10095 & ~n10096;
  assign n10099 = ~n10097 & ~n10098;
  assign n10100 = ~n8704 & ~n10099;
  assign n10101 = ~n10094 & ~n10100;
  assign n10102 = pi1690 & ~n10101;
  assign n10103 = ~n10093 & ~n10102;
  assign po0590 = pi1122 & ~n10103;
  assign n10105 = n8969 & n9588;
  assign n10106 = n9090 & n10105;
  assign n10107 = pi0481 & ~n10106;
  assign n10108 = ~pi0481 & n10106;
  assign n10109 = ~n10107 & ~n10108;
  assign n10110 = ~pi1690 & ~n10109;
  assign n10111 = pi0481 & n8704;
  assign n10112 = pi0384 & ~n8923;
  assign n10113 = n9603 & n10112;
  assign n10114 = ~n9076 & n10113;
  assign n10115 = n9080 & n10113;
  assign n10116 = ~n9078 & n10115;
  assign n10117 = pi0384 & n8941;
  assign n10118 = ~n9598 & n10112;
  assign n10119 = ~n10117 & ~n10118;
  assign n10120 = ~n10116 & n10119;
  assign n10121 = ~n10114 & n10120;
  assign n10122 = pi0481 & n10121;
  assign n10123 = ~pi0481 & ~n10121;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = ~n8704 & ~n10124;
  assign n10126 = ~n10111 & ~n10125;
  assign n10127 = pi1690 & ~n10126;
  assign n10128 = ~n10110 & ~n10127;
  assign po0591 = pi1122 & ~n10128;
  assign n10130 = pi0482 & ~n8976;
  assign n10131 = ~pi0482 & n8976;
  assign n10132 = ~n10130 & ~n10131;
  assign n10133 = ~pi1690 & ~n10132;
  assign n10134 = pi0482 & n8704;
  assign n10135 = ~n8922 & ~n8942;
  assign n10136 = n8949 & ~n8960;
  assign n10137 = n8939 & ~n10136;
  assign n10138 = n10135 & n10137;
  assign n10139 = ~n10135 & ~n10137;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = ~n8704 & ~n10140;
  assign n10142 = ~n10134 & ~n10141;
  assign n10143 = pi1690 & ~n10142;
  assign n10144 = ~n10133 & ~n10143;
  assign po0592 = pi1122 & ~n10144;
  assign n10146 = pi0483 & n8771;
  assign n10147 = ~n8775 & ~n8778;
  assign n10148 = n9870 & ~n9875;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = n10147 & n10148;
  assign n10151 = ~n10149 & ~n10150;
  assign n10152 = ~n8771 & ~n10151;
  assign n10153 = ~n10146 & ~n10152;
  assign n10154 = pi1679 & ~n10153;
  assign n10155 = pi0483 & n9891;
  assign n10156 = ~pi0483 & ~n9891;
  assign n10157 = ~n10155 & ~n10156;
  assign n10158 = ~pi1679 & n10157;
  assign n10159 = ~n10154 & ~n10158;
  assign po0593 = pi1131 & ~n10159;
  assign n10161 = pi0484 & ~n8858;
  assign n10162 = ~pi0484 & n8858;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = ~pi1690 & ~n10163;
  assign n10165 = pi0484 & n8704;
  assign n10166 = ~n8720 & ~n8723;
  assign n10167 = n9846 & n10166;
  assign n10168 = ~n9846 & ~n10166;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = ~n8704 & ~n10169;
  assign n10171 = ~n10165 & ~n10170;
  assign n10172 = pi1690 & ~n10171;
  assign n10173 = ~n10164 & ~n10172;
  assign po0594 = pi1122 & ~n10173;
  assign n10175 = pi0485 & n8771;
  assign n10176 = ~n8780 & ~n8781;
  assign n10177 = ~n8788 & n8795;
  assign n10178 = ~n8790 & ~n10177;
  assign n10179 = ~n8785 & ~n8787;
  assign n10180 = ~n10178 & n10179;
  assign n10181 = ~n8785 & n8791;
  assign n10182 = ~n8782 & ~n10181;
  assign n10183 = ~n10180 & n10182;
  assign n10184 = ~n8788 & ~n8796;
  assign n10185 = n10179 & n10184;
  assign n10186 = ~n8810 & ~n8813;
  assign n10187 = ~n8797 & ~n10186;
  assign n10188 = n10185 & ~n10187;
  assign n10189 = n10183 & ~n10188;
  assign n10190 = ~n10176 & ~n10189;
  assign n10191 = n10176 & n10189;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = ~n8771 & ~n10192;
  assign n10194 = ~n10175 & ~n10193;
  assign n10195 = pi1679 & ~n10194;
  assign n10196 = ~pi0485 & ~n9890;
  assign n10197 = ~n9891 & ~n10196;
  assign n10198 = ~pi1679 & n10197;
  assign n10199 = ~n10195 & ~n10198;
  assign po0595 = pi1131 & ~n10199;
  assign n10201 = pi0486 & n8771;
  assign n10202 = ~n9935 & ~n9943;
  assign n10203 = ~n9934 & ~n9938;
  assign n10204 = ~n9955 & n9959;
  assign n10205 = ~n9939 & ~n10204;
  assign n10206 = n10203 & ~n10205;
  assign n10207 = ~n9934 & n9937;
  assign n10208 = ~n9944 & ~n10207;
  assign n10209 = ~n10206 & n10208;
  assign n10210 = ~n9964 & n9966;
  assign n10211 = ~n9961 & ~n10210;
  assign n10212 = ~n9955 & ~n9960;
  assign n10213 = n10203 & n10212;
  assign n10214 = ~n10211 & n10213;
  assign n10215 = n10209 & ~n10214;
  assign n10216 = n10202 & n10215;
  assign n10217 = ~n10202 & ~n10215;
  assign n10218 = ~n10216 & ~n10217;
  assign n10219 = ~n8771 & ~n10218;
  assign n10220 = ~n10201 & ~n10219;
  assign n10221 = pi1679 & ~n10220;
  assign n10222 = n9979 & n9982;
  assign n10223 = n10014 & n10222;
  assign n10224 = pi0486 & n10223;
  assign n10225 = ~pi0486 & ~n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = ~pi1679 & n10226;
  assign n10228 = ~n10221 & ~n10227;
  assign po0596 = pi1131 & ~n10228;
  assign n10230 = ~pi0487 & n8405;
  assign n10231 = pi0064 & ~n8405;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = ~n8402 & ~n10232;
  assign n10234 = pi1774 & n8402;
  assign n10235 = ~n10233 & ~n10234;
  assign po0597 = ~pi1747 | ~n10235;
  assign n10237 = ~pi0488 & n8405;
  assign n10238 = pi0014 & ~n8405;
  assign n10239 = ~n10237 & ~n10238;
  assign n10240 = ~n8402 & ~n10239;
  assign n10241 = pi1786 & n8402;
  assign n10242 = ~n10240 & ~n10241;
  assign po0598 = ~pi1747 | ~n10242;
  assign n10244 = ~pi0489 & n8405;
  assign n10245 = pi0015 & ~n8405;
  assign n10246 = ~n10244 & ~n10245;
  assign n10247 = ~n8402 & ~n10246;
  assign n10248 = pi1790 & n8402;
  assign n10249 = ~n10247 & ~n10248;
  assign po0599 = ~pi1747 | ~n10249;
  assign n10251 = ~pi0490 & n8405;
  assign n10252 = pi0953 & ~n8405;
  assign n10253 = ~n10251 & ~n10252;
  assign n10254 = ~n8402 & ~n10253;
  assign n10255 = pi1791 & n8402;
  assign n10256 = ~n10254 & ~n10255;
  assign po0600 = ~pi1747 | ~n10256;
  assign n10258 = ~pi0491 & n8405;
  assign n10259 = pi0310 & ~n8405;
  assign n10260 = ~n10258 & ~n10259;
  assign n10261 = ~n8402 & ~n10260;
  assign n10262 = pi1792 & n8402;
  assign n10263 = ~n10261 & ~n10262;
  assign po0601 = ~pi1747 | ~n10263;
  assign n10265 = ~pi0492 & n8405;
  assign n10266 = pi0332 & ~n8405;
  assign n10267 = ~n10265 & ~n10266;
  assign n10268 = ~n8402 & ~n10267;
  assign n10269 = pi1793 & n8402;
  assign n10270 = ~n10268 & ~n10269;
  assign po0602 = ~pi1747 | ~n10270;
  assign n10272 = ~pi0493 & n8405;
  assign n10273 = pi0299 & ~n8405;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = ~n8402 & ~n10274;
  assign n10276 = pi1794 & n8402;
  assign n10277 = ~n10275 & ~n10276;
  assign po0603 = ~pi1747 | ~n10277;
  assign n10279 = ~pi0494 & n8405;
  assign n10280 = pi0286 & ~n8405;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = ~n8402 & ~n10281;
  assign n10283 = pi1795 & n8402;
  assign n10284 = ~n10282 & ~n10283;
  assign po0604 = ~pi1747 | ~n10284;
  assign n10286 = ~pi0495 & n8405;
  assign n10287 = pi1481 & ~n8405;
  assign n10288 = ~n10286 & ~n10287;
  assign n10289 = ~n8402 & ~n10288;
  assign n10290 = pi1796 & n8402;
  assign n10291 = ~n10289 & ~n10290;
  assign po0605 = ~pi1747 | ~n10291;
  assign n10293 = ~pi0496 & n8405;
  assign n10294 = pi0223 & ~n8405;
  assign n10295 = ~n10293 & ~n10294;
  assign n10296 = ~n8402 & ~n10295;
  assign n10297 = pi1798 & n8402;
  assign n10298 = ~n10296 & ~n10297;
  assign po0606 = ~pi1747 | ~n10298;
  assign n10300 = ~pi0497 & n8405;
  assign n10301 = pi0154 & ~n8405;
  assign n10302 = ~n10300 & ~n10301;
  assign n10303 = ~n8402 & ~n10302;
  assign n10304 = pi1799 & n8402;
  assign n10305 = ~n10303 & ~n10304;
  assign po0607 = ~pi1747 | ~n10305;
  assign n10307 = ~pi0498 & n8405;
  assign n10308 = pi0155 & ~n8405;
  assign n10309 = ~n10307 & ~n10308;
  assign n10310 = ~n8402 & ~n10309;
  assign n10311 = pi1800 & n8402;
  assign n10312 = ~n10310 & ~n10311;
  assign po0608 = ~pi1747 | ~n10312;
  assign n10314 = ~pi0499 & n8405;
  assign n10315 = pi0056 & ~n8405;
  assign n10316 = ~n10314 & ~n10315;
  assign n10317 = ~n8402 & ~n10316;
  assign n10318 = pi1776 & n8402;
  assign n10319 = ~n10317 & ~n10318;
  assign po0609 = ~pi1747 | ~n10319;
  assign n10321 = ~pi0500 & n8405;
  assign n10322 = pi0063 & ~n8405;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n8402 & ~n10323;
  assign n10325 = pi1804 & n8402;
  assign n10326 = ~n10324 & ~n10325;
  assign po0610 = ~pi1747 | ~n10326;
  assign n10328 = ~pi0501 & n8405;
  assign n10329 = pi0194 & ~n8405;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = ~n8402 & ~n10330;
  assign n10332 = pi1803 & n8402;
  assign n10333 = ~n10331 & ~n10332;
  assign po0611 = ~pi1747 | ~n10333;
  assign n10335 = ~pi0502 & n8405;
  assign n10336 = pi0049 & ~n8405;
  assign n10337 = ~n10335 & ~n10336;
  assign n10338 = ~n8402 & ~n10337;
  assign n10339 = pi1777 & n8402;
  assign n10340 = ~n10338 & ~n10339;
  assign po0612 = ~pi1747 | ~n10340;
  assign n10342 = ~pi0503 & n8405;
  assign n10343 = pi0027 & ~n8405;
  assign n10344 = ~n10342 & ~n10343;
  assign n10345 = ~n8402 & ~n10344;
  assign n10346 = pi1782 & n8402;
  assign n10347 = ~n10345 & ~n10346;
  assign po0613 = ~pi1747 | ~n10347;
  assign n10349 = ~pi1672 & ~n9733;
  assign n10350 = ~pi0504 & n9733;
  assign n10351 = ~n10349 & ~n10350;
  assign n10352 = ~n9730 & ~n10351;
  assign n10353 = pi1802 & n9730;
  assign n10354 = ~n10352 & ~n10353;
  assign po0614 = ~pi1747 | ~n10354;
  assign n10356 = ~pi1666 & ~n9733;
  assign n10357 = ~pi0505 & n9733;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n9730 & ~n10358;
  assign n10360 = pi1805 & n9730;
  assign n10361 = ~n10359 & ~n10360;
  assign po0615 = ~pi1747 | ~n10361;
  assign n10363 = pi0506 & n8771;
  assign n10364 = pi0506 & ~pi1027;
  assign n10365 = ~n8813 & ~n10364;
  assign n10366 = ~n8771 & ~n10365;
  assign n10367 = ~n10363 & ~n10366;
  assign n10368 = pi1679 & ~n10367;
  assign n10369 = ~pi0506 & ~pi1679;
  assign n10370 = ~n10368 & ~n10369;
  assign po0616 = pi1131 & ~n10370;
  assign n10372 = pi0408 & ~pi0507;
  assign n10373 = ~pi0408 & pi0507;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = ~pi1690 & ~n10374;
  assign n10376 = pi0507 & n8704;
  assign n10377 = ~n8730 & ~n8743;
  assign n10378 = ~n8746 & ~n10377;
  assign n10379 = n8746 & n10377;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = ~n8704 & ~n10380;
  assign n10382 = ~n10376 & ~n10381;
  assign n10383 = pi1690 & ~n10382;
  assign n10384 = ~n10375 & ~n10383;
  assign po0617 = pi1122 & ~n10384;
  assign n10386 = ~pi0508 & n8856;
  assign n10387 = pi0508 & ~n8856;
  assign n10388 = ~n10386 & ~n10387;
  assign n10389 = ~pi1690 & ~n10388;
  assign n10390 = pi0508 & n8704;
  assign n10391 = ~n8728 & ~n8729;
  assign n10392 = ~n9054 & ~n10391;
  assign n10393 = n9054 & n10391;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = ~n8704 & ~n10394;
  assign n10396 = ~n10390 & ~n10395;
  assign n10397 = pi1690 & ~n10396;
  assign n10398 = ~n10389 & ~n10397;
  assign po0618 = pi1122 & ~n10398;
  assign n10400 = pi0509 & ~n8857;
  assign n10401 = ~pi0509 & n8857;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = ~pi1690 & ~n10402;
  assign n10404 = pi0509 & n8704;
  assign n10405 = ~n8721 & ~n8726;
  assign n10406 = n8842 & n10405;
  assign n10407 = ~n8842 & ~n10405;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = ~n8704 & ~n10408;
  assign n10410 = ~n10404 & ~n10409;
  assign n10411 = pi1690 & ~n10410;
  assign n10412 = ~n10403 & ~n10411;
  assign po0619 = pi1122 & ~n10412;
  assign n10414 = pi0510 & ~n9008;
  assign n10415 = ~pi0510 & n9008;
  assign n10416 = ~n10414 & ~n10415;
  assign n10417 = ~pi1690 & ~n10416;
  assign n10418 = pi0510 & n8704;
  assign n10419 = ~n8926 & ~n8936;
  assign n10420 = n8987 & ~n8995;
  assign n10421 = n10419 & n10420;
  assign n10422 = ~n10419 & ~n10420;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = ~n8704 & ~n10423;
  assign n10425 = ~n10418 & ~n10424;
  assign n10426 = pi1690 & ~n10425;
  assign n10427 = ~n10417 & ~n10426;
  assign po0620 = pi1122 & ~n10427;
  assign n10429 = pi0511 & n8771;
  assign n10430 = ~pi0511 & pi1027;
  assign n10431 = pi0511 & ~pi1027;
  assign n10432 = ~n10430 & ~n10431;
  assign n10433 = ~n8771 & ~n10432;
  assign n10434 = ~n10429 & ~n10433;
  assign n10435 = pi1679 & ~n10434;
  assign n10436 = ~pi0511 & ~pi1679;
  assign n10437 = ~n10435 & ~n10436;
  assign po0621 = pi1131 & ~n10437;
  assign n10439 = pi0512 & n8771;
  assign n10440 = ~n9961 & ~n9964;
  assign n10441 = n9966 & ~n10440;
  assign n10442 = ~n9966 & n10440;
  assign n10443 = ~n10441 & ~n10442;
  assign n10444 = ~n8771 & ~n10443;
  assign n10445 = ~n10439 & ~n10444;
  assign n10446 = pi1679 & ~n10445;
  assign n10447 = pi0511 & pi0512;
  assign n10448 = ~n9979 & ~n10447;
  assign n10449 = ~pi1679 & ~n10448;
  assign n10450 = ~n10446 & ~n10449;
  assign po0622 = pi1131 & ~n10450;
  assign n10452 = pi0513 & n8771;
  assign n10453 = ~n9959 & ~n9960;
  assign n10454 = ~n10211 & ~n10453;
  assign n10455 = n10211 & n10453;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = ~n8771 & ~n10456;
  assign n10458 = ~n10452 & ~n10457;
  assign n10459 = pi1679 & ~n10458;
  assign n10460 = pi0513 & ~n9979;
  assign n10461 = ~n9980 & ~n10460;
  assign n10462 = ~pi1679 & ~n10461;
  assign n10463 = ~n10459 & ~n10462;
  assign po0623 = pi1131 & ~n10463;
  assign n10465 = pi0514 & n8771;
  assign n10466 = ~n9939 & ~n9955;
  assign n10467 = ~n9968 & ~n10466;
  assign n10468 = n9968 & n10466;
  assign n10469 = ~n10467 & ~n10468;
  assign n10470 = ~n8771 & ~n10469;
  assign n10471 = ~n10465 & ~n10470;
  assign n10472 = pi1679 & ~n10471;
  assign n10473 = pi0514 & ~n9980;
  assign n10474 = ~n9981 & ~n10473;
  assign n10475 = ~pi1679 & ~n10474;
  assign n10476 = ~n10472 & ~n10475;
  assign po0624 = pi1131 & ~n10476;
  assign n10478 = pi1802 & n9550;
  assign n10479 = pi1159 & n8483;
  assign n10480 = ~pi0515 & ~n8482;
  assign n10481 = ~pi1672 & n8482;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = ~n8483 & ~n10482;
  assign n10484 = ~n10479 & ~n10483;
  assign n10485 = ~n9550 & ~n10484;
  assign n10486 = pi1747 & ~n10485;
  assign po0625 = n10478 | ~n10486;
  assign n10488 = pi1786 & n8007;
  assign n10489 = ~pi1168 & n8009;
  assign n10490 = pi0014 & n8011;
  assign n10491 = ~pi0516 & ~n8011;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = ~n8009 & ~n10492;
  assign n10494 = ~n10489 & ~n10493;
  assign n10495 = ~n8007 & ~n10494;
  assign n10496 = pi1747 & ~n10495;
  assign po0626 = n10488 | ~n10496;
  assign n10498 = pi1790 & n8007;
  assign n10499 = ~pi1170 & n8009;
  assign n10500 = pi0015 & n8011;
  assign n10501 = ~pi0517 & ~n8011;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = ~n8009 & ~n10502;
  assign n10504 = ~n10499 & ~n10503;
  assign n10505 = ~n8007 & ~n10504;
  assign n10506 = pi1747 & ~n10505;
  assign po0627 = n10498 | ~n10506;
  assign n10508 = pi1791 & n8007;
  assign n10509 = ~pi1247 & n8009;
  assign n10510 = pi0953 & n8011;
  assign n10511 = ~pi0518 & ~n8011;
  assign n10512 = ~n10510 & ~n10511;
  assign n10513 = ~n8009 & ~n10512;
  assign n10514 = ~n10509 & ~n10513;
  assign n10515 = ~n8007 & ~n10514;
  assign n10516 = pi1747 & ~n10515;
  assign po0628 = n10508 | ~n10516;
  assign n10518 = pi1803 & n8007;
  assign n10519 = pi1177 & n8009;
  assign n10520 = pi0194 & n8011;
  assign n10521 = ~pi0519 & ~n8011;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = ~n8009 & ~n10522;
  assign n10524 = ~n10519 & ~n10523;
  assign n10525 = ~n8007 & ~n10524;
  assign n10526 = pi1747 & ~n10525;
  assign po0629 = n10518 | ~n10526;
  assign n10528 = pi1774 & n9430;
  assign n10529 = ~pi1207 & n8414;
  assign n10530 = pi0064 & n8413;
  assign n10531 = ~pi0520 & ~n8413;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = ~n8414 & ~n10532;
  assign n10534 = ~n10529 & ~n10533;
  assign n10535 = ~n9430 & ~n10534;
  assign n10536 = pi1747 & ~n10535;
  assign po0630 = n10528 | ~n10536;
  assign n10538 = pi1790 & n9430;
  assign n10539 = ~pi1071 & n8414;
  assign n10540 = pi0015 & n8413;
  assign n10541 = ~pi0521 & ~n8413;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = ~n8414 & ~n10542;
  assign n10544 = ~n10539 & ~n10543;
  assign n10545 = ~n9430 & ~n10544;
  assign n10546 = pi1747 & ~n10545;
  assign po0631 = n10538 | ~n10546;
  assign n10548 = pi1791 & n9430;
  assign n10549 = ~pi1211 & n8414;
  assign n10550 = pi0953 & n8413;
  assign n10551 = ~pi0522 & ~n8413;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = ~n8414 & ~n10552;
  assign n10554 = ~n10549 & ~n10553;
  assign n10555 = ~n9430 & ~n10554;
  assign n10556 = pi1747 & ~n10555;
  assign po0632 = n10548 | ~n10556;
  assign n10558 = pi1792 & n9430;
  assign n10559 = ~pi1212 & n8414;
  assign n10560 = pi0310 & n8413;
  assign n10561 = ~pi0523 & ~n8413;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = ~n8414 & ~n10562;
  assign n10564 = ~n10559 & ~n10563;
  assign n10565 = ~n9430 & ~n10564;
  assign n10566 = pi1747 & ~n10565;
  assign po0633 = n10558 | ~n10566;
  assign n10568 = pi1794 & n9430;
  assign n10569 = pi1214 & n8414;
  assign n10570 = pi0299 & n8413;
  assign n10571 = ~pi0524 & ~n8413;
  assign n10572 = ~n10570 & ~n10571;
  assign n10573 = ~n8414 & ~n10572;
  assign n10574 = ~n10569 & ~n10573;
  assign n10575 = ~n9430 & ~n10574;
  assign n10576 = pi1747 & ~n10575;
  assign po0634 = n10568 | ~n10576;
  assign n10578 = pi1796 & n9430;
  assign n10579 = pi1216 & n8414;
  assign n10580 = pi1481 & n8413;
  assign n10581 = ~pi0525 & ~n8413;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = ~n8414 & ~n10582;
  assign n10584 = ~n10579 & ~n10583;
  assign n10585 = ~n9430 & ~n10584;
  assign n10586 = pi1747 & ~n10585;
  assign po0635 = n10578 | ~n10586;
  assign n10588 = pi1798 & n9430;
  assign n10589 = pi1217 & n8414;
  assign n10590 = pi0223 & n8413;
  assign n10591 = ~pi0526 & ~n8413;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = ~n8414 & ~n10592;
  assign n10594 = ~n10589 & ~n10593;
  assign n10595 = ~n9430 & ~n10594;
  assign n10596 = pi1747 & ~n10595;
  assign po0636 = n10588 | ~n10596;
  assign n10598 = pi1799 & n9430;
  assign n10599 = pi1218 & n8414;
  assign n10600 = pi0154 & n8413;
  assign n10601 = ~pi0527 & ~n8413;
  assign n10602 = ~n10600 & ~n10601;
  assign n10603 = ~n8414 & ~n10602;
  assign n10604 = ~n10599 & ~n10603;
  assign n10605 = ~n9430 & ~n10604;
  assign n10606 = pi1747 & ~n10605;
  assign po0637 = n10598 | ~n10606;
  assign n10608 = pi1803 & n9430;
  assign n10609 = pi1232 & n8414;
  assign n10610 = pi0194 & n8413;
  assign n10611 = ~pi0528 & ~n8413;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = ~n8414 & ~n10612;
  assign n10614 = ~n10609 & ~n10613;
  assign n10615 = ~n9430 & ~n10614;
  assign n10616 = pi1747 & ~n10615;
  assign po0638 = n10608 | ~n10616;
  assign n10618 = pi1775 & n9430;
  assign n10619 = ~pi1064 & n8414;
  assign n10620 = pi0057 & n8413;
  assign n10621 = ~pi0529 & ~n8413;
  assign n10622 = ~n10620 & ~n10621;
  assign n10623 = ~n8414 & ~n10622;
  assign n10624 = ~n10619 & ~n10623;
  assign n10625 = ~n9430 & ~n10624;
  assign n10626 = pi1747 & ~n10625;
  assign po0639 = n10618 | ~n10626;
  assign n10628 = pi1804 & n9430;
  assign n10629 = pi1266 & n8414;
  assign n10630 = pi0063 & n8413;
  assign n10631 = ~pi0530 & ~n8413;
  assign n10632 = ~n10630 & ~n10631;
  assign n10633 = ~n8414 & ~n10632;
  assign n10634 = ~n10629 & ~n10633;
  assign n10635 = ~n9430 & ~n10634;
  assign n10636 = pi1747 & ~n10635;
  assign po0640 = n10628 | ~n10636;
  assign n10638 = pi1777 & n9430;
  assign n10639 = ~pi1282 & n8414;
  assign n10640 = pi0049 & n8413;
  assign n10641 = ~pi0531 & ~n8413;
  assign n10642 = ~n10640 & ~n10641;
  assign n10643 = ~n8414 & ~n10642;
  assign n10644 = ~n10639 & ~n10643;
  assign n10645 = ~n9430 & ~n10644;
  assign n10646 = pi1747 & ~n10645;
  assign po0641 = n10638 | ~n10646;
  assign n10648 = pi0018 & ~n9733;
  assign n10649 = ~pi0532 & n9733;
  assign n10650 = ~n10648 & ~n10649;
  assign n10651 = ~n9730 & ~n10650;
  assign n10652 = pi1789 & n9730;
  assign n10653 = ~n10651 & ~n10652;
  assign po0642 = ~pi1747 | ~n10653;
  assign n10655 = n6345 & n6354;
  assign n10656 = n9889 & n10655;
  assign n10657 = pi0533 & ~n10656;
  assign n10658 = ~pi0533 & n10656;
  assign n10659 = ~n10657 & ~n10658;
  assign n10660 = ~pi1679 & ~n10659;
  assign n10661 = pi0533 & n8771;
  assign n10662 = ~n8773 & ~n8774;
  assign n10663 = ~n8778 & n8780;
  assign n10664 = ~n8775 & ~n10663;
  assign n10665 = n10184 & ~n10187;
  assign n10666 = n10178 & ~n10665;
  assign n10667 = n10179 & ~n10666;
  assign n10668 = n10182 & ~n10667;
  assign n10669 = ~n8778 & ~n8781;
  assign n10670 = ~n10668 & n10669;
  assign n10671 = n10664 & ~n10670;
  assign n10672 = n10662 & n10671;
  assign n10673 = ~n10662 & ~n10671;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = ~n8771 & ~n10674;
  assign n10676 = ~n10661 & ~n10675;
  assign n10677 = pi1679 & ~n10676;
  assign n10678 = ~n10660 & ~n10677;
  assign po0643 = pi1131 & ~n10678;
  assign n10680 = pi1776 & n8356;
  assign n10681 = ~pi1200 & n8358;
  assign n10682 = pi0056 & n8360;
  assign n10683 = ~pi0534 & ~n8360;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = ~n8358 & ~n10684;
  assign n10686 = ~n10681 & ~n10685;
  assign n10687 = ~n8356 & ~n10686;
  assign n10688 = pi1747 & ~n10687;
  assign po0644 = n10680 | ~n10688;
  assign n10690 = ~pi0089 & n5266;
  assign n10691 = pi1417 & n10690;
  assign n10692 = n6406 & n10691;
  assign n10693 = ~pi1416 & n5445;
  assign n10694 = n6406 & n10693;
  assign n10695 = pi0089 & n10694;
  assign n10696 = ~n10692 & ~n10695;
  assign n10697 = pi1480 & ~n10696;
  assign n10698 = ~pi0535 & ~n10697;
  assign po0645 = n6189 & ~n10698;
  assign n10700 = pi1796 & n8356;
  assign n10701 = pi1195 & n8358;
  assign n10702 = pi1481 & n8360;
  assign n10703 = ~pi0536 & ~n8360;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n8358 & ~n10704;
  assign n10706 = ~n10701 & ~n10705;
  assign n10707 = ~n8356 & ~n10706;
  assign n10708 = pi1747 & ~n10707;
  assign po0646 = n10700 | ~n10708;
  assign n10710 = ~pi0537 & n9733;
  assign n10711 = pi0049 & ~n9733;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~n9730 & ~n10712;
  assign n10714 = pi1777 & n9730;
  assign n10715 = ~n10713 & ~n10714;
  assign po0647 = ~pi1747 | ~n10715;
  assign n10717 = ~pi0538 & n9733;
  assign n10718 = pi0299 & ~n9733;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 = ~n9730 & ~n10719;
  assign n10721 = pi1794 & n9730;
  assign n10722 = ~n10720 & ~n10721;
  assign po0648 = ~pi1747 | ~n10722;
  assign n10724 = ~pi0539 & n9733;
  assign n10725 = pi0124 & ~n9733;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = ~n9730 & ~n10726;
  assign n10728 = pi1801 & n9730;
  assign n10729 = ~n10727 & ~n10728;
  assign po0649 = ~pi1747 | ~n10729;
  assign n10731 = ~pi0540 & n9733;
  assign n10732 = pi0223 & ~n9733;
  assign n10733 = ~n10731 & ~n10732;
  assign n10734 = ~n9730 & ~n10733;
  assign n10735 = pi1798 & n9730;
  assign n10736 = ~n10734 & ~n10735;
  assign po0650 = ~pi1747 | ~n10736;
  assign n10738 = pi0541 & ~n9981;
  assign n10739 = ~pi0541 & n9981;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~pi1679 & ~n10740;
  assign n10742 = pi0541 & n8771;
  assign n10743 = ~n9937 & ~n9938;
  assign n10744 = ~n10211 & n10212;
  assign n10745 = n10205 & ~n10744;
  assign n10746 = ~n10743 & ~n10745;
  assign n10747 = n10743 & n10745;
  assign n10748 = ~n10746 & ~n10747;
  assign n10749 = ~n8771 & ~n10748;
  assign n10750 = ~n10742 & ~n10749;
  assign n10751 = pi1679 & ~n10750;
  assign n10752 = ~n10741 & ~n10751;
  assign po0651 = pi1131 & ~n10752;
  assign n10754 = pi1803 & n9550;
  assign n10755 = pi1269 & n8483;
  assign n10756 = pi0194 & n8482;
  assign n10757 = ~pi0542 & ~n8482;
  assign n10758 = ~n10756 & ~n10757;
  assign n10759 = ~n8483 & ~n10758;
  assign n10760 = ~n10755 & ~n10759;
  assign n10761 = ~n9550 & ~n10760;
  assign n10762 = pi1747 & ~n10761;
  assign po0652 = n10754 | ~n10762;
  assign n10764 = ~pi0543 & n9733;
  assign n10765 = pi0953 & ~n9733;
  assign n10766 = ~n10764 & ~n10765;
  assign n10767 = ~n9730 & ~n10766;
  assign n10768 = pi1791 & n9730;
  assign n10769 = ~n10767 & ~n10768;
  assign po0653 = ~pi1747 | ~n10769;
  assign n10771 = pi1799 & n9550;
  assign n10772 = pi1275 & n8483;
  assign n10773 = pi0154 & n8482;
  assign n10774 = ~pi0544 & ~n8482;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~n8483 & ~n10775;
  assign n10777 = ~n10772 & ~n10776;
  assign n10778 = ~n9550 & ~n10777;
  assign n10779 = pi1747 & ~n10778;
  assign po0654 = n10771 | ~n10779;
  assign n10781 = ~n5855 & ~n5870;
  assign n10782 = n5867 & n10781;
  assign n10783 = ~n5867 & ~n10781;
  assign po0655 = n10782 | n10783;
  assign n10785 = pi1795 & n9550;
  assign n10786 = pi1154 & n8483;
  assign n10787 = pi0286 & n8482;
  assign n10788 = ~pi0546 & ~n8482;
  assign n10789 = ~n10787 & ~n10788;
  assign n10790 = ~n8483 & ~n10789;
  assign n10791 = ~n10786 & ~n10790;
  assign n10792 = ~n9550 & ~n10791;
  assign n10793 = pi1747 & ~n10792;
  assign po0656 = n10785 | ~n10793;
  assign n10795 = pi1779 & n9550;
  assign n10796 = ~pi1162 & n8483;
  assign n10797 = pi0028 & n8482;
  assign n10798 = ~pi0547 & ~n8482;
  assign n10799 = ~n10797 & ~n10798;
  assign n10800 = ~n8483 & ~n10799;
  assign n10801 = ~n10796 & ~n10800;
  assign n10802 = ~n9550 & ~n10801;
  assign n10803 = pi1747 & ~n10802;
  assign po0657 = n10795 | ~n10803;
  assign n10805 = pi1779 & n8356;
  assign n10806 = ~pi1204 & n8358;
  assign n10807 = pi0028 & n8360;
  assign n10808 = ~pi0548 & ~n8360;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = ~n8358 & ~n10809;
  assign n10811 = ~n10806 & ~n10810;
  assign n10812 = ~n8356 & ~n10811;
  assign n10813 = pi1747 & ~n10812;
  assign po0658 = n10805 | ~n10813;
  assign n10815 = pi0506 & n8826;
  assign n10816 = pi0549 & ~n10815;
  assign n10817 = ~pi0549 & n10815;
  assign n10818 = ~n10816 & ~n10817;
  assign n10819 = ~pi1679 & ~n10818;
  assign n10820 = pi0549 & n8771;
  assign n10821 = ~n8782 & ~n8785;
  assign n10822 = ~n8804 & ~n8814;
  assign n10823 = n10821 & n10822;
  assign n10824 = ~n10821 & ~n10822;
  assign n10825 = ~n10823 & ~n10824;
  assign n10826 = ~n8771 & ~n10825;
  assign n10827 = ~n10820 & ~n10826;
  assign n10828 = pi1679 & ~n10827;
  assign n10829 = ~n10819 & ~n10828;
  assign po0659 = pi1131 & ~n10829;
  assign n10831 = pi1780 & n9550;
  assign n10832 = ~pi1343 & n8483;
  assign n10833 = pi0023 & n8482;
  assign n10834 = ~pi0550 & ~n8482;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = ~n8483 & ~n10835;
  assign n10837 = ~n10832 & ~n10836;
  assign n10838 = ~n9550 & ~n10837;
  assign n10839 = pi1747 & ~n10838;
  assign po0660 = n10831 | ~n10839;
  assign n10841 = pi1784 & n9550;
  assign n10842 = ~pi1316 & n8483;
  assign n10843 = pi0016 & n8482;
  assign n10844 = ~pi0551 & ~n8482;
  assign n10845 = ~n10843 & ~n10844;
  assign n10846 = ~n8483 & ~n10845;
  assign n10847 = ~n10842 & ~n10846;
  assign n10848 = ~n9550 & ~n10847;
  assign n10849 = pi1747 & ~n10848;
  assign po0661 = n10841 | ~n10849;
  assign n10851 = pi0552 & n8417;
  assign n10852 = pi0642 & pi1139;
  assign n10853 = ~pi0642 & ~pi1139;
  assign n10854 = pi0631 & pi1034;
  assign n10855 = ~n10853 & n10854;
  assign n10856 = ~n10852 & ~n10855;
  assign n10857 = ~pi0631 & ~pi1034;
  assign n10858 = ~n10853 & ~n10857;
  assign n10859 = pi0568 & pi1265;
  assign n10860 = ~pi0568 & ~pi1265;
  assign n10861 = pi0655 & pi1142;
  assign n10862 = ~n10860 & n10861;
  assign n10863 = ~n10859 & ~n10862;
  assign n10864 = ~pi0655 & ~pi1142;
  assign n10865 = ~n10860 & ~n10864;
  assign n10866 = pi0627 & pi1033;
  assign n10867 = ~pi0627 & ~pi1033;
  assign n10868 = pi0591 & pi1258;
  assign n10869 = ~n10867 & n10868;
  assign n10870 = ~n10866 & ~n10869;
  assign n10871 = ~pi0591 & ~pi1258;
  assign n10872 = ~n10867 & ~n10871;
  assign n10873 = pi0590 & pi1141;
  assign n10874 = ~pi0590 & ~pi1141;
  assign n10875 = pi0589 & pi1342;
  assign n10876 = ~n10874 & n10875;
  assign n10877 = ~n10873 & ~n10876;
  assign n10878 = n10872 & ~n10877;
  assign n10879 = n10870 & ~n10878;
  assign n10880 = n10865 & ~n10879;
  assign n10881 = n10863 & ~n10880;
  assign n10882 = n10858 & ~n10881;
  assign n10883 = n10856 & ~n10882;
  assign n10884 = n10858 & n10865;
  assign n10885 = ~pi0589 & ~pi1342;
  assign n10886 = pi0594 & pi1032;
  assign n10887 = ~n10874 & n10886;
  assign n10888 = n10872 & n10887;
  assign n10889 = ~n10885 & n10888;
  assign n10890 = n10884 & n10889;
  assign n10891 = n10883 & ~n10890;
  assign n10892 = pi0552 & n10891;
  assign n10893 = ~pi0552 & ~n10891;
  assign n10894 = ~n10892 & ~n10893;
  assign n10895 = ~n8417 & ~n10894;
  assign n10896 = ~n10851 & ~n10895;
  assign n10897 = pi1697 & ~n10896;
  assign n10898 = ~pi0631 & ~pi0655;
  assign n10899 = ~pi0594 & ~pi0627;
  assign n10900 = ~pi0590 & ~pi0591;
  assign n10901 = ~pi0589 & n10900;
  assign n10902 = n10899 & n10901;
  assign n10903 = ~pi0642 & n10902;
  assign n10904 = ~pi0568 & n10903;
  assign n10905 = n10898 & n10904;
  assign n10906 = pi0552 & n10905;
  assign n10907 = ~pi0552 & ~n10905;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = ~pi1697 & n10908;
  assign n10910 = ~n10897 & ~n10909;
  assign po0662 = pi1143 & ~n10910;
  assign n10912 = pi1788 & n9550;
  assign n10913 = ~pi1151 & n8483;
  assign n10914 = pi0011 & n8482;
  assign n10915 = ~pi0553 & ~n8482;
  assign n10916 = ~n10914 & ~n10915;
  assign n10917 = ~n8483 & ~n10916;
  assign n10918 = ~n10913 & ~n10917;
  assign n10919 = ~n9550 & ~n10918;
  assign n10920 = pi1747 & ~n10919;
  assign po0663 = n10912 | ~n10920;
  assign n10922 = pi1787 & n9550;
  assign n10923 = ~pi1312 & n8483;
  assign n10924 = pi0007 & n8482;
  assign n10925 = ~pi0554 & ~n8482;
  assign n10926 = ~n10924 & ~n10925;
  assign n10927 = ~n8483 & ~n10926;
  assign n10928 = ~n10923 & ~n10927;
  assign n10929 = ~n9550 & ~n10928;
  assign n10930 = pi1747 & ~n10929;
  assign po0664 = n10922 | ~n10930;
  assign n10932 = pi1785 & n9550;
  assign n10933 = ~pi1311 & n8483;
  assign n10934 = pi0019 & n8482;
  assign n10935 = ~pi0555 & ~n8482;
  assign n10936 = ~n10934 & ~n10935;
  assign n10937 = ~n8483 & ~n10936;
  assign n10938 = ~n10933 & ~n10937;
  assign n10939 = ~n9550 & ~n10938;
  assign n10940 = pi1747 & ~n10939;
  assign po0665 = n10932 | ~n10940;
  assign n10942 = pi1789 & n9550;
  assign n10943 = ~pi1152 & n8483;
  assign n10944 = pi0018 & n8482;
  assign n10945 = ~pi0556 & ~n8482;
  assign n10946 = ~n10944 & ~n10945;
  assign n10947 = ~n8483 & ~n10946;
  assign n10948 = ~n10943 & ~n10947;
  assign n10949 = ~n9550 & ~n10948;
  assign n10950 = pi1747 & ~n10949;
  assign po0666 = n10942 | ~n10950;
  assign n10952 = pi1778 & n9550;
  assign n10953 = ~pi1332 & n8483;
  assign n10954 = pi0046 & n8482;
  assign n10955 = ~pi0557 & ~n8482;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = ~n8483 & ~n10956;
  assign n10958 = ~n10953 & ~n10957;
  assign n10959 = ~n9550 & ~n10958;
  assign n10960 = pi1747 & ~n10959;
  assign po0667 = n10952 | ~n10960;
  assign n10962 = pi1781 & n9550;
  assign n10963 = ~pi1333 & n8483;
  assign n10964 = pi0030 & n8482;
  assign n10965 = ~pi0558 & ~n8482;
  assign n10966 = ~n10964 & ~n10965;
  assign n10967 = ~n8483 & ~n10966;
  assign n10968 = ~n10963 & ~n10967;
  assign n10969 = ~n9550 & ~n10968;
  assign n10970 = pi1747 & ~n10969;
  assign po0668 = n10962 | ~n10970;
  assign n10972 = pi1778 & n8356;
  assign n10973 = ~pi1203 & n8358;
  assign n10974 = pi0046 & n8360;
  assign n10975 = ~pi0559 & ~n8360;
  assign n10976 = ~n10974 & ~n10975;
  assign n10977 = ~n8358 & ~n10976;
  assign n10978 = ~n10973 & ~n10977;
  assign n10979 = ~n8356 & ~n10978;
  assign n10980 = pi1747 & ~n10979;
  assign po0669 = n10972 | ~n10980;
  assign n10982 = ~pi0486 & ~pi0565;
  assign n10983 = n9982 & n10982;
  assign n10984 = n9981 & n10983;
  assign n10985 = pi0560 & ~n10984;
  assign n10986 = ~pi0560 & n10984;
  assign n10987 = ~n10985 & ~n10986;
  assign n10988 = ~pi1679 & ~n10987;
  assign n10989 = pi0560 & n8771;
  assign n10990 = ~n9931 & ~n9949;
  assign n10991 = ~n9930 & n9943;
  assign n10992 = ~n9950 & ~n10991;
  assign n10993 = n10203 & ~n10745;
  assign n10994 = n10208 & ~n10993;
  assign n10995 = ~n9930 & ~n9935;
  assign n10996 = ~n10994 & n10995;
  assign n10997 = n10992 & ~n10996;
  assign n10998 = ~n10990 & ~n10997;
  assign n10999 = n10990 & n10997;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n8771 & ~n11000;
  assign n11002 = ~n10989 & ~n11001;
  assign n11003 = pi1679 & ~n11002;
  assign n11004 = ~n10988 & ~n11003;
  assign po0670 = pi1131 & ~n11004;
  assign n11006 = pi0753 & ~pi1773;
  assign n11007 = pi1773 & pi1807;
  assign po0671 = n11006 | n11007;
  assign n11009 = n6345 & n6371;
  assign n11010 = n9890 & n11009;
  assign n11011 = pi0562 & ~n11010;
  assign n11012 = ~pi0562 & n11010;
  assign n11013 = ~n11011 & ~n11012;
  assign n11014 = ~pi1679 & ~n11013;
  assign n11015 = pi0562 & n8771;
  assign n11016 = ~n10183 & n10669;
  assign n11017 = n10664 & ~n11016;
  assign n11018 = ~n8774 & ~n11017;
  assign n11019 = ~pi0380 & ~n8773;
  assign n11020 = ~n11018 & n11019;
  assign n11021 = ~n8774 & n10669;
  assign n11022 = n10188 & n11021;
  assign n11023 = n11020 & ~n11022;
  assign n11024 = pi0562 & ~n11023;
  assign n11025 = ~pi0562 & n11023;
  assign n11026 = ~n11024 & ~n11025;
  assign n11027 = ~n8771 & ~n11026;
  assign n11028 = ~n11015 & ~n11027;
  assign n11029 = pi1679 & ~n11028;
  assign n11030 = ~n11014 & ~n11029;
  assign po0672 = pi1131 & ~n11030;
  assign n11032 = pi0563 & n8417;
  assign n11033 = pi0552 & pi0649;
  assign n11034 = n10858 & n11033;
  assign n11035 = n10865 & ~n10870;
  assign n11036 = n10863 & ~n11035;
  assign n11037 = n11034 & ~n11036;
  assign n11038 = ~n10856 & n11033;
  assign n11039 = ~n11037 & ~n11038;
  assign n11040 = n10865 & n10872;
  assign n11041 = n11034 & n11040;
  assign n11042 = ~n10874 & ~n10885;
  assign n11043 = n10886 & n11042;
  assign n11044 = n10877 & ~n11043;
  assign n11045 = n11041 & ~n11044;
  assign n11046 = n11039 & ~n11045;
  assign n11047 = pi0563 & n11046;
  assign n11048 = ~pi0563 & ~n11046;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = ~n8417 & ~n11049;
  assign n11051 = ~n11032 & ~n11050;
  assign n11052 = pi1697 & ~n11051;
  assign n11053 = ~pi0552 & ~pi0642;
  assign n11054 = ~pi0631 & ~pi0649;
  assign n11055 = ~pi0589 & ~pi0594;
  assign n11056 = ~pi0590 & n11055;
  assign n11057 = ~pi0591 & n11056;
  assign n11058 = ~pi0627 & ~pi0655;
  assign n11059 = ~pi0568 & n11058;
  assign n11060 = n11057 & n11059;
  assign n11061 = n11054 & n11060;
  assign n11062 = n11053 & n11061;
  assign n11063 = pi0563 & n11062;
  assign n11064 = ~pi0563 & ~n11062;
  assign n11065 = ~n11063 & ~n11064;
  assign n11066 = ~pi1697 & n11065;
  assign n11067 = ~n11052 & ~n11066;
  assign po0673 = pi1143 & ~n11067;
  assign n11069 = n9977 & n10982;
  assign n11070 = n10223 & n11069;
  assign n11071 = pi0564 & ~n11070;
  assign n11072 = ~pi0564 & n11070;
  assign n11073 = ~n11071 & ~n11072;
  assign n11074 = ~pi1679 & ~n11073;
  assign n11075 = pi0564 & n8771;
  assign n11076 = pi0472 & ~n9931;
  assign n11077 = n10995 & n11076;
  assign n11078 = ~n10209 & n11077;
  assign n11079 = n10213 & n11077;
  assign n11080 = ~n10211 & n11079;
  assign n11081 = pi0472 & n9949;
  assign n11082 = ~n10992 & n11076;
  assign n11083 = ~n11081 & ~n11082;
  assign n11084 = ~n11080 & n11083;
  assign n11085 = ~n11078 & n11084;
  assign n11086 = pi0564 & n11085;
  assign n11087 = ~pi0564 & ~n11085;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = ~n8771 & ~n11088;
  assign n11090 = ~n11075 & ~n11089;
  assign n11091 = pi1679 & ~n11090;
  assign n11092 = ~n11074 & ~n11091;
  assign po0674 = pi1131 & ~n11092;
  assign n11094 = pi0565 & ~n9984;
  assign n11095 = ~pi0565 & n9984;
  assign n11096 = ~n11094 & ~n11095;
  assign n11097 = ~pi1679 & ~n11096;
  assign n11098 = pi0565 & n8771;
  assign n11099 = ~n9930 & ~n9950;
  assign n11100 = n9957 & ~n9968;
  assign n11101 = n9947 & ~n11100;
  assign n11102 = n11099 & n11101;
  assign n11103 = ~n11099 & ~n11101;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = ~n8771 & ~n11104;
  assign n11106 = ~n11098 & ~n11105;
  assign n11107 = pi1679 & ~n11106;
  assign n11108 = ~n11097 & ~n11107;
  assign po0675 = pi1131 & ~n11108;
  assign n11110 = pi0566 & n8417;
  assign n11111 = ~n8421 & ~n8424;
  assign n11112 = n8432 & ~n8437;
  assign n11113 = ~n8440 & n11112;
  assign n11114 = n8430 & ~n11113;
  assign n11115 = n8457 & ~n8459;
  assign n11116 = n8445 & ~n11115;
  assign n11117 = n8432 & n8435;
  assign n11118 = ~n11116 & n11117;
  assign n11119 = n11114 & ~n11118;
  assign n11120 = ~n11111 & ~n11119;
  assign n11121 = n11111 & n11119;
  assign n11122 = ~n11120 & ~n11121;
  assign n11123 = ~n8417 & ~n11122;
  assign n11124 = ~n11110 & ~n11123;
  assign n11125 = pi1697 & ~n11124;
  assign n11126 = pi0586 & pi0662;
  assign n11127 = pi0653 & n11126;
  assign n11128 = pi0654 & n11127;
  assign n11129 = n6453 & n11128;
  assign n11130 = pi0569 & n11129;
  assign n11131 = pi0566 & n11130;
  assign n11132 = ~pi0566 & ~n11130;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~pi1697 & n11133;
  assign n11135 = ~n11125 & ~n11134;
  assign po0676 = pi1143 & ~n11135;
  assign n11137 = pi0567 & ~n9889;
  assign n11138 = ~pi0567 & n9889;
  assign n11139 = ~n11137 & ~n11138;
  assign n11140 = ~pi1679 & ~n11139;
  assign n11141 = pi0567 & n8771;
  assign n11142 = ~n8787 & ~n8791;
  assign n11143 = n10666 & n11142;
  assign n11144 = ~n10666 & ~n11142;
  assign n11145 = ~n11143 & ~n11144;
  assign n11146 = ~n8771 & ~n11145;
  assign n11147 = ~n11141 & ~n11146;
  assign n11148 = pi1679 & ~n11147;
  assign n11149 = ~n11140 & ~n11148;
  assign po0677 = pi1131 & ~n11149;
  assign n11151 = pi0568 & n8417;
  assign n11152 = ~n10859 & ~n10860;
  assign n11153 = ~n10864 & ~n10867;
  assign n11154 = ~n10871 & n10873;
  assign n11155 = ~n10868 & ~n11154;
  assign n11156 = n11153 & ~n11155;
  assign n11157 = ~n10864 & n10866;
  assign n11158 = ~n10861 & ~n11157;
  assign n11159 = ~n11156 & n11158;
  assign n11160 = ~n10885 & n10886;
  assign n11161 = ~n10875 & ~n11160;
  assign n11162 = ~n10871 & ~n10874;
  assign n11163 = n11153 & n11162;
  assign n11164 = ~n11161 & n11163;
  assign n11165 = n11159 & ~n11164;
  assign n11166 = n11152 & n11165;
  assign n11167 = ~n11152 & ~n11165;
  assign n11168 = ~n11166 & ~n11167;
  assign n11169 = ~n8417 & ~n11168;
  assign n11170 = ~n11151 & ~n11169;
  assign n11171 = pi1697 & ~n11170;
  assign n11172 = n11055 & n11058;
  assign n11173 = n10900 & n11172;
  assign n11174 = pi0568 & n11173;
  assign n11175 = ~pi0568 & ~n11173;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = ~pi1697 & n11176;
  assign n11178 = ~n11171 & ~n11177;
  assign po0678 = pi1143 & ~n11178;
  assign n11180 = pi0569 & n8417;
  assign n11181 = ~n8426 & ~n8427;
  assign n11182 = ~n8434 & n8441;
  assign n11183 = ~n8439 & ~n11182;
  assign n11184 = ~n8431 & ~n8433;
  assign n11185 = ~n11183 & n11184;
  assign n11186 = ~n8431 & n8436;
  assign n11187 = ~n8428 & ~n11186;
  assign n11188 = ~n11185 & n11187;
  assign n11189 = ~n8434 & ~n8442;
  assign n11190 = n11184 & n11189;
  assign n11191 = ~n8456 & ~n8459;
  assign n11192 = ~n8443 & ~n11191;
  assign n11193 = n11190 & ~n11192;
  assign n11194 = n11188 & ~n11193;
  assign n11195 = ~n11181 & ~n11194;
  assign n11196 = n11181 & n11194;
  assign n11197 = ~n11195 & ~n11196;
  assign n11198 = ~n8417 & ~n11197;
  assign n11199 = ~n11180 & ~n11198;
  assign n11200 = pi1697 & ~n11199;
  assign n11201 = ~pi0569 & ~n11129;
  assign n11202 = ~n11130 & ~n11201;
  assign n11203 = ~pi1697 & n11202;
  assign n11204 = ~n11200 & ~n11203;
  assign po0679 = pi1143 & ~n11204;
  assign n11206 = ~pi0570 & n9733;
  assign n11207 = pi0064 & ~n9733;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = ~n9730 & ~n11208;
  assign n11210 = pi1774 & n9730;
  assign n11211 = ~n11209 & ~n11210;
  assign po0680 = ~pi1747 | ~n11211;
  assign n11213 = ~pi0571 & n9733;
  assign n11214 = pi0014 & ~n9733;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = ~n9730 & ~n11215;
  assign n11217 = pi1786 & n9730;
  assign n11218 = ~n11216 & ~n11217;
  assign po0681 = ~pi1747 | ~n11218;
  assign n11220 = ~pi0572 & n9733;
  assign n11221 = pi0015 & ~n9733;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = ~n9730 & ~n11222;
  assign n11224 = pi1790 & n9730;
  assign n11225 = ~n11223 & ~n11224;
  assign po0682 = ~pi1747 | ~n11225;
  assign n11227 = ~pi0573 & n9733;
  assign n11228 = pi0310 & ~n9733;
  assign n11229 = ~n11227 & ~n11228;
  assign n11230 = ~n9730 & ~n11229;
  assign n11231 = pi1792 & n9730;
  assign n11232 = ~n11230 & ~n11231;
  assign po0683 = ~pi1747 | ~n11232;
  assign n11234 = ~pi0574 & n9733;
  assign n11235 = pi0332 & ~n9733;
  assign n11236 = ~n11234 & ~n11235;
  assign n11237 = ~n9730 & ~n11236;
  assign n11238 = pi1793 & n9730;
  assign n11239 = ~n11237 & ~n11238;
  assign po0684 = ~pi1747 | ~n11239;
  assign n11241 = ~pi0575 & n9733;
  assign n11242 = pi0057 & ~n9733;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = ~n9730 & ~n11243;
  assign n11245 = pi1775 & n9730;
  assign n11246 = ~n11244 & ~n11245;
  assign po0685 = ~pi1747 | ~n11246;
  assign n11248 = ~pi0576 & n9733;
  assign n11249 = pi1481 & ~n9733;
  assign n11250 = ~n11248 & ~n11249;
  assign n11251 = ~n9730 & ~n11250;
  assign n11252 = pi1796 & n9730;
  assign n11253 = ~n11251 & ~n11252;
  assign po0686 = ~pi1747 | ~n11253;
  assign n11255 = ~pi0577 & n9733;
  assign n11256 = pi0254 & ~n9733;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~n9730 & ~n11257;
  assign n11259 = pi1797 & n9730;
  assign n11260 = ~n11258 & ~n11259;
  assign po0687 = ~pi1747 | ~n11260;
  assign n11262 = ~pi0578 & n9733;
  assign n11263 = pi0286 & ~n9733;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = ~n9730 & ~n11264;
  assign n11266 = pi1795 & n9730;
  assign n11267 = ~n11265 & ~n11266;
  assign po0688 = ~pi1747 | ~n11267;
  assign n11269 = ~pi0579 & n9733;
  assign n11270 = pi0155 & ~n9733;
  assign n11271 = ~n11269 & ~n11270;
  assign n11272 = ~n9730 & ~n11271;
  assign n11273 = pi1800 & n9730;
  assign n11274 = ~n11272 & ~n11273;
  assign po0689 = ~pi1747 | ~n11274;
  assign n11276 = ~pi0580 & n9733;
  assign n11277 = pi0154 & ~n9733;
  assign n11278 = ~n11276 & ~n11277;
  assign n11279 = ~n9730 & ~n11278;
  assign n11280 = pi1799 & n9730;
  assign n11281 = ~n11279 & ~n11280;
  assign po0690 = ~pi1747 | ~n11281;
  assign n11283 = ~pi0581 & n9733;
  assign n11284 = pi0194 & ~n9733;
  assign n11285 = ~n11283 & ~n11284;
  assign n11286 = ~n9730 & ~n11285;
  assign n11287 = pi1803 & n9730;
  assign n11288 = ~n11286 & ~n11287;
  assign po0691 = ~pi1747 | ~n11288;
  assign n11290 = ~pi0582 & n9733;
  assign n11291 = pi0056 & ~n9733;
  assign n11292 = ~n11290 & ~n11291;
  assign n11293 = ~n9730 & ~n11292;
  assign n11294 = pi1776 & n9730;
  assign n11295 = ~n11293 & ~n11294;
  assign po0692 = ~pi1747 | ~n11295;
  assign n11297 = ~pi0583 & n9733;
  assign n11298 = pi0063 & ~n9733;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n9730 & ~n11299;
  assign n11301 = pi1804 & n9730;
  assign n11302 = ~n11300 & ~n11301;
  assign po0693 = ~pi1747 | ~n11302;
  assign n11304 = ~pi0584 & n9733;
  assign n11305 = pi0027 & ~n9733;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = ~n9730 & ~n11306;
  assign n11308 = pi1782 & n9730;
  assign n11309 = ~n11307 & ~n11308;
  assign po0694 = ~pi1747 | ~n11309;
  assign n11311 = ~pi0585 & n9733;
  assign n11312 = pi0022 & ~n9733;
  assign n11313 = ~n11311 & ~n11312;
  assign n11314 = ~n9730 & ~n11313;
  assign n11315 = pi1783 & n9730;
  assign n11316 = ~n11314 & ~n11315;
  assign po0695 = ~pi1747 | ~n11316;
  assign n11318 = pi0586 & n8417;
  assign n11319 = pi0586 & ~pi1032;
  assign n11320 = ~n8459 & ~n11319;
  assign n11321 = ~n8417 & ~n11320;
  assign n11322 = ~n11318 & ~n11321;
  assign n11323 = pi1697 & ~n11322;
  assign n11324 = ~pi0586 & ~pi1697;
  assign n11325 = ~n11323 & ~n11324;
  assign po0696 = pi1143 & ~n11325;
  assign n11327 = ~pi0587 & n9887;
  assign n11328 = pi0587 & ~n9887;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~pi1679 & ~n11329;
  assign n11331 = pi0587 & n8771;
  assign n11332 = ~n8795 & ~n8796;
  assign n11333 = ~n10187 & ~n11332;
  assign n11334 = n10187 & n11332;
  assign n11335 = ~n11333 & ~n11334;
  assign n11336 = ~n8771 & ~n11335;
  assign n11337 = ~n11331 & ~n11336;
  assign n11338 = pi1679 & ~n11337;
  assign n11339 = ~n11330 & ~n11338;
  assign po0697 = pi1131 & ~n11339;
  assign n11341 = pi0588 & ~n10016;
  assign n11342 = ~pi0588 & n10016;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = ~pi1679 & ~n11343;
  assign n11345 = pi0588 & n8771;
  assign n11346 = ~n9934 & ~n9944;
  assign n11347 = n9995 & ~n10003;
  assign n11348 = n11346 & n11347;
  assign n11349 = ~n11346 & ~n11347;
  assign n11350 = ~n11348 & ~n11349;
  assign n11351 = ~n8771 & ~n11350;
  assign n11352 = ~n11345 & ~n11351;
  assign n11353 = pi1679 & ~n11352;
  assign n11354 = ~n11344 & ~n11353;
  assign po0698 = pi1131 & ~n11354;
  assign n11356 = pi0589 & n8417;
  assign n11357 = ~n10875 & ~n10885;
  assign n11358 = n10886 & ~n11357;
  assign n11359 = ~n10886 & n11357;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = ~n8417 & ~n11360;
  assign n11362 = ~n11356 & ~n11361;
  assign n11363 = pi1697 & ~n11362;
  assign n11364 = pi0589 & pi0594;
  assign n11365 = ~n11055 & ~n11364;
  assign n11366 = ~pi1697 & ~n11365;
  assign n11367 = ~n11363 & ~n11366;
  assign po0699 = pi1143 & ~n11367;
  assign n11369 = pi0590 & n8417;
  assign n11370 = ~n10873 & ~n10874;
  assign n11371 = ~n11161 & ~n11370;
  assign n11372 = n11161 & n11370;
  assign n11373 = ~n11371 & ~n11372;
  assign n11374 = ~n8417 & ~n11373;
  assign n11375 = ~n11369 & ~n11374;
  assign n11376 = pi1697 & ~n11375;
  assign n11377 = pi0590 & ~n11055;
  assign n11378 = ~n11056 & ~n11377;
  assign n11379 = ~pi1697 & ~n11378;
  assign n11380 = ~n11376 & ~n11379;
  assign po0700 = pi1143 & ~n11380;
  assign n11382 = pi0591 & n8417;
  assign n11383 = ~n10868 & ~n10871;
  assign n11384 = ~n11044 & ~n11383;
  assign n11385 = n11044 & n11383;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = ~n8417 & ~n11386;
  assign n11388 = ~n11382 & ~n11387;
  assign n11389 = pi1697 & ~n11388;
  assign n11390 = pi0591 & ~n11056;
  assign n11391 = ~n11057 & ~n11390;
  assign n11392 = ~pi1697 & ~n11391;
  assign n11393 = ~n11389 & ~n11392;
  assign po0701 = pi1143 & ~n11393;
  assign n11395 = pi1459 & ~n10696;
  assign n11396 = ~pi0592 & ~n11395;
  assign po0702 = n6185 & ~n11396;
  assign n11398 = pi1774 & n9550;
  assign n11399 = ~pi1149 & n8483;
  assign n11400 = pi0064 & n8482;
  assign n11401 = ~pi0593 & ~n8482;
  assign n11402 = ~n11400 & ~n11401;
  assign n11403 = ~n8483 & ~n11402;
  assign n11404 = ~n11399 & ~n11403;
  assign n11405 = ~n9550 & ~n11404;
  assign n11406 = pi1747 & ~n11405;
  assign po0703 = n11398 | ~n11406;
  assign n11408 = pi0594 & n8417;
  assign n11409 = ~pi0594 & pi1032;
  assign n11410 = pi0594 & ~pi1032;
  assign n11411 = ~n11409 & ~n11410;
  assign n11412 = ~n8417 & ~n11411;
  assign n11413 = ~n11408 & ~n11412;
  assign n11414 = pi1697 & ~n11413;
  assign n11415 = ~pi0594 & ~pi1697;
  assign n11416 = ~n11414 & ~n11415;
  assign po0704 = pi1143 & ~n11416;
  assign n11418 = pi1790 & n9550;
  assign n11419 = ~pi1153 & n8483;
  assign n11420 = pi0015 & n8482;
  assign n11421 = ~pi0595 & ~n8482;
  assign n11422 = ~n11420 & ~n11421;
  assign n11423 = ~n8483 & ~n11422;
  assign n11424 = ~n11419 & ~n11423;
  assign n11425 = ~n9550 & ~n11424;
  assign n11426 = pi1747 & ~n11425;
  assign po0705 = n11418 | ~n11426;
  assign n11428 = pi1791 & n9550;
  assign n11429 = ~pi1305 & n8483;
  assign n11430 = pi0953 & n8482;
  assign n11431 = ~pi0596 & ~n8482;
  assign n11432 = ~n11430 & ~n11431;
  assign n11433 = ~n8483 & ~n11432;
  assign n11434 = ~n11429 & ~n11433;
  assign n11435 = ~n9550 & ~n11434;
  assign n11436 = pi1747 & ~n11435;
  assign po0706 = n11428 | ~n11436;
  assign n11438 = pi1792 & n9550;
  assign n11439 = ~pi1284 & n8483;
  assign n11440 = pi0310 & n8482;
  assign n11441 = ~pi0597 & ~n8482;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = ~n8483 & ~n11442;
  assign n11444 = ~n11439 & ~n11443;
  assign n11445 = ~n9550 & ~n11444;
  assign n11446 = pi1747 & ~n11445;
  assign po0707 = n11438 | ~n11446;
  assign n11448 = pi1793 & n9550;
  assign n11449 = pi1331 & n8483;
  assign n11450 = pi0332 & n8482;
  assign n11451 = ~pi0598 & ~n8482;
  assign n11452 = ~n11450 & ~n11451;
  assign n11453 = ~n8483 & ~n11452;
  assign n11454 = ~n11449 & ~n11453;
  assign n11455 = ~n9550 & ~n11454;
  assign n11456 = pi1747 & ~n11455;
  assign po0708 = n11448 | ~n11456;
  assign n11458 = pi1775 & n9550;
  assign n11459 = ~pi1292 & n8483;
  assign n11460 = pi0057 & n8482;
  assign n11461 = ~pi0599 & ~n8482;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = ~n8483 & ~n11462;
  assign n11464 = ~n11459 & ~n11463;
  assign n11465 = ~n9550 & ~n11464;
  assign n11466 = pi1747 & ~n11465;
  assign po0709 = n11458 | ~n11466;
  assign n11468 = pi1794 & n9550;
  assign n11469 = pi1283 & n8483;
  assign n11470 = pi0299 & n8482;
  assign n11471 = ~pi0600 & ~n8482;
  assign n11472 = ~n11470 & ~n11471;
  assign n11473 = ~n8483 & ~n11472;
  assign n11474 = ~n11469 & ~n11473;
  assign n11475 = ~n9550 & ~n11474;
  assign n11476 = pi1747 & ~n11475;
  assign po0710 = n11468 | ~n11476;
  assign n11478 = pi1786 & n9550;
  assign n11479 = ~pi1150 & n8483;
  assign n11480 = pi0014 & n8482;
  assign n11481 = ~pi0601 & ~n8482;
  assign n11482 = ~n11480 & ~n11481;
  assign n11483 = ~n8483 & ~n11482;
  assign n11484 = ~n11479 & ~n11483;
  assign n11485 = ~n9550 & ~n11484;
  assign n11486 = pi1747 & ~n11485;
  assign po0711 = n11478 | ~n11486;
  assign n11488 = pi1797 & n9550;
  assign n11489 = pi1156 & n8483;
  assign n11490 = pi0254 & n8482;
  assign n11491 = ~pi0602 & ~n8482;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = ~n8483 & ~n11492;
  assign n11494 = ~n11489 & ~n11493;
  assign n11495 = ~n9550 & ~n11494;
  assign n11496 = pi1747 & ~n11495;
  assign po0712 = n11488 | ~n11496;
  assign n11498 = pi1798 & n9550;
  assign n11499 = pi1157 & n8483;
  assign n11500 = pi0223 & n8482;
  assign n11501 = ~pi0603 & ~n8482;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = ~n8483 & ~n11502;
  assign n11504 = ~n11499 & ~n11503;
  assign n11505 = ~n9550 & ~n11504;
  assign n11506 = pi1747 & ~n11505;
  assign po0713 = n11498 | ~n11506;
  assign n11508 = pi1796 & n9550;
  assign n11509 = pi1155 & n8483;
  assign n11510 = pi1481 & n8482;
  assign n11511 = ~pi0604 & ~n8482;
  assign n11512 = ~n11510 & ~n11511;
  assign n11513 = ~n8483 & ~n11512;
  assign n11514 = ~n11509 & ~n11513;
  assign n11515 = ~n9550 & ~n11514;
  assign n11516 = pi1747 & ~n11515;
  assign po0714 = n11508 | ~n11516;
  assign n11518 = pi1801 & n9550;
  assign n11519 = pi1346 & n8483;
  assign n11520 = pi0124 & n8482;
  assign n11521 = ~pi0605 & ~n8482;
  assign n11522 = ~n11520 & ~n11521;
  assign n11523 = ~n8483 & ~n11522;
  assign n11524 = ~n11519 & ~n11523;
  assign n11525 = ~n9550 & ~n11524;
  assign n11526 = pi1747 & ~n11525;
  assign po0715 = n11518 | ~n11526;
  assign n11528 = pi1800 & n9550;
  assign n11529 = pi1158 & n8483;
  assign n11530 = pi0155 & n8482;
  assign n11531 = ~pi0606 & ~n8482;
  assign n11532 = ~n11530 & ~n11531;
  assign n11533 = ~n8483 & ~n11532;
  assign n11534 = ~n11529 & ~n11533;
  assign n11535 = ~n9550 & ~n11534;
  assign n11536 = pi1747 & ~n11535;
  assign po0716 = n11528 | ~n11536;
  assign n11538 = pi1776 & n9550;
  assign n11539 = ~pi1344 & n8483;
  assign n11540 = pi0056 & n8482;
  assign n11541 = ~pi0607 & ~n8482;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = ~n8483 & ~n11542;
  assign n11544 = ~n11539 & ~n11543;
  assign n11545 = ~n9550 & ~n11544;
  assign n11546 = pi1747 & ~n11545;
  assign po0717 = n11538 | ~n11546;
  assign n11548 = pi1804 & n9550;
  assign n11549 = pi1160 & n8483;
  assign n11550 = pi0063 & n8482;
  assign n11551 = ~pi0608 & ~n8482;
  assign n11552 = ~n11550 & ~n11551;
  assign n11553 = ~n8483 & ~n11552;
  assign n11554 = ~n11549 & ~n11553;
  assign n11555 = ~n9550 & ~n11554;
  assign n11556 = pi1747 & ~n11555;
  assign po0718 = n11548 | ~n11556;
  assign n11558 = pi1777 & n9550;
  assign n11559 = ~pi1263 & n8483;
  assign n11560 = pi0049 & n8482;
  assign n11561 = ~pi0609 & ~n8482;
  assign n11562 = ~n11560 & ~n11561;
  assign n11563 = ~n8483 & ~n11562;
  assign n11564 = ~n11559 & ~n11563;
  assign n11565 = ~n9550 & ~n11564;
  assign n11566 = pi1747 & ~n11565;
  assign po0719 = n11558 | ~n11566;
  assign n11568 = pi1782 & n9550;
  assign n11569 = ~pi1163 & n8483;
  assign n11570 = pi0027 & n8482;
  assign n11571 = ~pi0610 & ~n8482;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = ~n8483 & ~n11572;
  assign n11574 = ~n11569 & ~n11573;
  assign n11575 = ~n9550 & ~n11574;
  assign n11576 = pi1747 & ~n11575;
  assign po0720 = n11568 | ~n11576;
  assign n11578 = pi1783 & n9550;
  assign n11579 = ~pi1183 & n8483;
  assign n11580 = pi0022 & n8482;
  assign n11581 = ~pi0611 & ~n8482;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = ~n8483 & ~n11582;
  assign n11584 = ~n11579 & ~n11583;
  assign n11585 = ~n9550 & ~n11584;
  assign n11586 = pi1747 & ~n11585;
  assign po0721 = n11578 | ~n11586;
  assign n11588 = pi1774 & n8356;
  assign n11589 = ~pi1065 & n8358;
  assign n11590 = pi0064 & n8360;
  assign n11591 = ~pi0612 & ~n8360;
  assign n11592 = ~n11590 & ~n11591;
  assign n11593 = ~n8358 & ~n11592;
  assign n11594 = ~n11589 & ~n11593;
  assign n11595 = ~n8356 & ~n11594;
  assign n11596 = pi1747 & ~n11595;
  assign po0722 = n11588 | ~n11596;
  assign n11598 = pi1786 & n8356;
  assign n11599 = ~pi1187 & n8358;
  assign n11600 = pi0014 & n8360;
  assign n11601 = ~pi0613 & ~n8360;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = ~n8358 & ~n11602;
  assign n11604 = ~n11599 & ~n11603;
  assign n11605 = ~n8356 & ~n11604;
  assign n11606 = pi1747 & ~n11605;
  assign po0723 = n11598 | ~n11606;
  assign n11608 = pi1791 & n8356;
  assign n11609 = ~pi1248 & n8358;
  assign n11610 = pi0953 & n8360;
  assign n11611 = ~pi0614 & ~n8360;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = ~n8358 & ~n11612;
  assign n11614 = ~n11609 & ~n11613;
  assign n11615 = ~n8356 & ~n11614;
  assign n11616 = pi1747 & ~n11615;
  assign po0724 = n11608 | ~n11616;
  assign n11618 = pi1430 & ~n10696;
  assign n11619 = ~pi0615 & ~n11618;
  assign po0725 = n6193 & ~n11619;
  assign n11621 = pi1803 & n8356;
  assign n11622 = pi1201 & n8358;
  assign n11623 = pi0194 & n8360;
  assign n11624 = ~pi0616 & ~n8360;
  assign n11625 = ~n11623 & ~n11624;
  assign n11626 = ~n8358 & ~n11625;
  assign n11627 = ~n11622 & ~n11626;
  assign n11628 = ~n8356 & ~n11627;
  assign n11629 = pi1747 & ~n11628;
  assign po0726 = n11621 | ~n11629;
  assign n11631 = pi1447 & ~n10696;
  assign n11632 = ~pi0617 & ~n11631;
  assign po0727 = n6201 & ~n11632;
  assign n11634 = pi0506 & ~pi0618;
  assign n11635 = ~pi0506 & pi0618;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = ~pi1679 & ~n11636;
  assign n11638 = pi0618 & n8771;
  assign n11639 = ~n8797 & ~n8810;
  assign n11640 = ~n8813 & ~n11639;
  assign n11641 = n8813 & n11639;
  assign n11642 = ~n11640 & ~n11641;
  assign n11643 = ~n8771 & ~n11642;
  assign n11644 = ~n11638 & ~n11643;
  assign n11645 = pi1679 & ~n11644;
  assign n11646 = ~n11637 & ~n11645;
  assign po0728 = pi1131 & ~n11646;
  assign n11648 = pi0619 & n3751;
  assign n11649 = ~pi1773 & n3740;
  assign n11650 = pi0619 & n3742;
  assign n11651 = n3746 & n11650;
  assign n11652 = ~n11649 & n11651;
  assign n11653 = ~n8004 & n11652;
  assign n11654 = ~pi0716 & n3734;
  assign n11655 = ~pi0677 & n11654;
  assign n11656 = ~pi1401 & n11655;
  assign n11657 = pi0634 & n11656;
  assign n11658 = pi1747 & ~n11657;
  assign n11659 = ~n11653 & n11658;
  assign po0729 = n11648 | ~n11659;
  assign n11661 = ~n5856 & ~n5869;
  assign n11662 = n7770 & n11661;
  assign n11663 = ~n7770 & ~n11661;
  assign po0730 = n11662 | n11663;
  assign n11665 = pi0621 & n8417;
  assign n11666 = n8425 & ~n11114;
  assign n11667 = n8425 & n11118;
  assign n11668 = ~pi0358 & ~pi0645;
  assign n11669 = ~n11667 & n11668;
  assign n11670 = n8423 & n11669;
  assign n11671 = ~n11666 & n11670;
  assign n11672 = pi0621 & ~n11671;
  assign n11673 = ~pi0621 & n11671;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n8417 & ~n11674;
  assign n11676 = ~n11665 & ~n11675;
  assign n11677 = pi1697 & ~n11676;
  assign n11678 = n6470 & n11130;
  assign n11679 = pi0645 & n11678;
  assign n11680 = pi0566 & n11679;
  assign n11681 = pi0621 & n11680;
  assign n11682 = ~pi0621 & ~n11680;
  assign n11683 = ~n11681 & ~n11682;
  assign n11684 = ~pi1697 & n11683;
  assign n11685 = ~n11677 & ~n11684;
  assign po0731 = pi1143 & ~n11685;
  assign n11687 = pi0622 & ~n9888;
  assign n11688 = ~pi0622 & n9888;
  assign n11689 = ~n11687 & ~n11688;
  assign n11690 = ~pi1679 & ~n11689;
  assign n11691 = pi0622 & n8771;
  assign n11692 = ~n8788 & ~n8790;
  assign n11693 = n9873 & n11692;
  assign n11694 = ~n9873 & ~n11692;
  assign n11695 = ~n11693 & ~n11694;
  assign n11696 = ~n8771 & ~n11695;
  assign n11697 = ~n11691 & ~n11696;
  assign n11698 = pi1679 & ~n11697;
  assign n11699 = ~n11690 & ~n11698;
  assign po0732 = pi1131 & ~n11699;
  assign n11701 = n6444 & n6453;
  assign n11702 = n11128 & n11701;
  assign n11703 = pi0623 & ~n11702;
  assign n11704 = ~pi0623 & n11702;
  assign n11705 = ~n11703 & ~n11704;
  assign n11706 = ~pi1697 & ~n11705;
  assign n11707 = pi0623 & n8417;
  assign n11708 = ~n8419 & ~n8420;
  assign n11709 = ~n8424 & n8426;
  assign n11710 = ~n8421 & ~n11709;
  assign n11711 = n11189 & ~n11192;
  assign n11712 = n11183 & ~n11711;
  assign n11713 = n11184 & ~n11712;
  assign n11714 = n11187 & ~n11713;
  assign n11715 = ~n8424 & ~n8427;
  assign n11716 = ~n11714 & n11715;
  assign n11717 = n11710 & ~n11716;
  assign n11718 = n11708 & n11717;
  assign n11719 = ~n11708 & ~n11717;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 = ~n8417 & ~n11720;
  assign n11722 = ~n11707 & ~n11721;
  assign n11723 = pi1697 & ~n11722;
  assign n11724 = ~n11706 & ~n11723;
  assign po0733 = pi1143 & ~n11724;
  assign n11726 = n8080 & n9549;
  assign n11727 = pi0996 & pi1480;
  assign n11728 = pi1480 & pi1729;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = pi0030 & ~n11729;
  assign n11731 = ~pi0624 & n11729;
  assign n11732 = ~n11730 & ~n11731;
  assign n11733 = ~n11726 & ~n11732;
  assign n11734 = pi1781 & n11726;
  assign n11735 = ~n11733 & ~n11734;
  assign po0734 = ~pi1747 | ~n11735;
  assign n11737 = ~pi1016 & n8884;
  assign n11738 = pi1016 & n8887;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = pi0982 & ~n11739;
  assign n11741 = ~pi1016 & n8883;
  assign n11742 = pi1016 & n8882;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = ~pi0982 & ~n11743;
  assign po0735 = ~n11740 & ~n11744;
  assign n11746 = pi1776 & n9430;
  assign n11747 = ~pi1220 & n8414;
  assign n11748 = pi0056 & n8413;
  assign n11749 = ~pi0626 & ~n8413;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = ~n8414 & ~n11750;
  assign n11752 = ~n11747 & ~n11751;
  assign n11753 = ~n9430 & ~n11752;
  assign n11754 = pi1747 & ~n11753;
  assign po0736 = n11746 | ~n11754;
  assign n11756 = pi0627 & ~n11057;
  assign n11757 = ~pi0627 & n11057;
  assign n11758 = ~n11756 & ~n11757;
  assign n11759 = ~pi1697 & ~n11758;
  assign n11760 = pi0627 & n8417;
  assign n11761 = ~n10866 & ~n10867;
  assign n11762 = ~n11161 & n11162;
  assign n11763 = n11155 & ~n11762;
  assign n11764 = ~n11761 & ~n11763;
  assign n11765 = n11761 & n11763;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = ~n8417 & ~n11766;
  assign n11768 = ~n11760 & ~n11767;
  assign n11769 = pi1697 & ~n11768;
  assign n11770 = ~n11759 & ~n11769;
  assign po0737 = pi1143 & ~n11770;
  assign n11772 = pi0028 & ~n11729;
  assign n11773 = ~pi0628 & n11729;
  assign n11774 = ~n11772 & ~n11773;
  assign n11775 = ~n11726 & ~n11774;
  assign n11776 = pi1779 & n11726;
  assign n11777 = ~n11775 & ~n11776;
  assign po0738 = ~pi1747 | ~n11777;
  assign n11779 = pi1800 & n9430;
  assign n11780 = pi1219 & n8414;
  assign n11781 = pi0155 & n8413;
  assign n11782 = ~pi0629 & ~n8413;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = ~n8414 & ~n11783;
  assign n11785 = ~n11780 & ~n11784;
  assign n11786 = ~n9430 & ~n11785;
  assign n11787 = pi1747 & ~n11786;
  assign po0739 = n11779 | ~n11787;
  assign n11789 = pi0702 & pi0716;
  assign n11790 = ~n3854 & ~n11789;
  assign n11791 = n3732 & n3854;
  assign n11792 = ~n11790 & n11791;
  assign n11793 = ~pi0619 & n11792;
  assign n11794 = pi1401 & n11793;
  assign n11795 = ~pi0702 & n3731;
  assign n11796 = pi0716 & n11795;
  assign n11797 = pi0702 & n3731;
  assign n11798 = ~pi0716 & n11797;
  assign n11799 = ~n11796 & ~n11798;
  assign po0740 = n11794 | ~n11799;
  assign n11801 = pi0631 & ~n11060;
  assign n11802 = ~pi0631 & n11060;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = ~pi1697 & ~n11803;
  assign n11805 = pi0631 & n8417;
  assign n11806 = ~n10854 & ~n10857;
  assign n11807 = n11040 & ~n11044;
  assign n11808 = n11036 & ~n11807;
  assign n11809 = n11806 & n11808;
  assign n11810 = ~n11806 & ~n11808;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = ~n8417 & ~n11811;
  assign n11813 = ~n11805 & ~n11812;
  assign n11814 = pi1697 & ~n11813;
  assign n11815 = ~n11804 & ~n11814;
  assign po0741 = pi1143 & ~n11815;
  assign n11817 = pi1778 & n9430;
  assign n11818 = ~pi1222 & n8414;
  assign n11819 = pi0046 & n8413;
  assign n11820 = ~pi0632 & ~n8413;
  assign n11821 = ~n11819 & ~n11820;
  assign n11822 = ~n8414 & ~n11821;
  assign n11823 = ~n11818 & ~n11822;
  assign n11824 = ~n9430 & ~n11823;
  assign n11825 = pi1747 & ~n11824;
  assign po0742 = n11817 | ~n11825;
  assign n11827 = pi0023 & ~n11729;
  assign n11828 = ~pi0633 & n11729;
  assign n11829 = ~n11827 & ~n11828;
  assign n11830 = ~n11726 & ~n11829;
  assign n11831 = pi1780 & n11726;
  assign n11832 = ~n11830 & ~n11831;
  assign po0743 = ~pi1747 | ~n11832;
  assign n11834 = pi0634 & n3751;
  assign n11835 = ~pi0634 & ~pi1401;
  assign n11836 = n11654 & n11835;
  assign n11837 = pi0677 & n11836;
  assign n11838 = ~n11834 & ~n11837;
  assign po0744 = pi1747 & ~n11838;
  assign n11840 = pi0011 & ~n11729;
  assign n11841 = ~pi0635 & n11729;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11726 & ~n11842;
  assign n11844 = pi1788 & n11726;
  assign n11845 = ~n11843 & ~n11844;
  assign po0745 = ~pi1747 | ~n11845;
  assign n11847 = pi0016 & ~n11729;
  assign n11848 = ~pi0636 & n11729;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = ~n11726 & ~n11849;
  assign n11851 = pi1784 & n11726;
  assign n11852 = ~n11850 & ~n11851;
  assign po0746 = ~pi1747 | ~n11852;
  assign n11854 = pi0007 & ~n11729;
  assign n11855 = ~pi0637 & n11729;
  assign n11856 = ~n11854 & ~n11855;
  assign n11857 = ~n11726 & ~n11856;
  assign n11858 = pi1787 & n11726;
  assign n11859 = ~n11857 & ~n11858;
  assign po0747 = ~pi1747 | ~n11859;
  assign n11861 = pi0019 & ~n11729;
  assign n11862 = ~pi0638 & n11729;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = ~n11726 & ~n11863;
  assign n11865 = pi1785 & n11726;
  assign n11866 = ~n11864 & ~n11865;
  assign po0748 = ~pi1747 | ~n11866;
  assign n11868 = pi0018 & ~n11729;
  assign n11869 = ~pi0639 & n11729;
  assign n11870 = ~n11868 & ~n11869;
  assign n11871 = ~n11726 & ~n11870;
  assign n11872 = pi1789 & n11726;
  assign n11873 = ~n11871 & ~n11872;
  assign po0749 = ~pi1747 | ~n11873;
  assign n11875 = pi1779 & n9430;
  assign n11876 = ~pi1281 & n8414;
  assign n11877 = pi0028 & n8413;
  assign n11878 = ~pi0640 & ~n8413;
  assign n11879 = ~n11877 & ~n11878;
  assign n11880 = ~n8414 & ~n11879;
  assign n11881 = ~n11876 & ~n11880;
  assign n11882 = ~n9430 & ~n11881;
  assign n11883 = pi1747 & ~n11882;
  assign po0750 = n11875 | ~n11883;
  assign n11885 = pi0046 & ~n11729;
  assign n11886 = ~pi0641 & n11729;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11726 & ~n11887;
  assign n11889 = pi1778 & n11726;
  assign n11890 = ~n11888 & ~n11889;
  assign po0751 = ~pi1747 | ~n11890;
  assign n11892 = ~pi0568 & ~pi0631;
  assign n11893 = n11058 & n11892;
  assign n11894 = n11057 & n11893;
  assign n11895 = pi0642 & ~n11894;
  assign n11896 = ~pi0642 & n11894;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = ~pi1697 & ~n11897;
  assign n11899 = pi0642 & n8417;
  assign n11900 = ~n10852 & ~n10853;
  assign n11901 = ~n10857 & n10859;
  assign n11902 = ~n10854 & ~n11901;
  assign n11903 = n11153 & ~n11763;
  assign n11904 = n11158 & ~n11903;
  assign n11905 = ~n10857 & ~n10860;
  assign n11906 = ~n11904 & n11905;
  assign n11907 = n11902 & ~n11906;
  assign n11908 = ~n11900 & ~n11907;
  assign n11909 = n11900 & n11907;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = ~n8417 & ~n11910;
  assign n11912 = ~n11899 & ~n11911;
  assign n11913 = pi1697 & ~n11912;
  assign n11914 = ~n11898 & ~n11913;
  assign po0752 = pi1143 & ~n11914;
  assign n11916 = pi0886 & ~pi1773;
  assign n11917 = pi1773 & pi1809;
  assign po0753 = n11916 | n11917;
  assign n11919 = ~pi0644 & pi0893;
  assign po0754 = n6325 & ~n11919;
  assign n11921 = n6444 & n6470;
  assign n11922 = n11129 & n11921;
  assign n11923 = pi0645 & ~n11922;
  assign n11924 = ~pi0645 & n11922;
  assign n11925 = ~n11923 & ~n11924;
  assign n11926 = ~pi1697 & ~n11925;
  assign n11927 = pi0645 & n8417;
  assign n11928 = ~n11188 & n11715;
  assign n11929 = n11710 & ~n11928;
  assign n11930 = ~n8420 & ~n11929;
  assign n11931 = ~pi0358 & ~n8419;
  assign n11932 = ~n11930 & n11931;
  assign n11933 = ~n8420 & n11715;
  assign n11934 = n11193 & n11933;
  assign n11935 = n11932 & ~n11934;
  assign n11936 = pi0645 & ~n11935;
  assign n11937 = ~pi0645 & n11935;
  assign n11938 = ~n11936 & ~n11937;
  assign n11939 = ~n8417 & ~n11938;
  assign n11940 = ~n11927 & ~n11939;
  assign n11941 = pi1697 & ~n11940;
  assign n11942 = ~n11926 & ~n11941;
  assign po0755 = pi1143 & ~n11942;
  assign n11944 = ~po1210 & ~n3752;
  assign n11945 = pi1747 & n11944;
  assign po0756 = ~n3731 & n11945;
  assign n11947 = pi0647 & ~pi1626;
  assign n11948 = ~n5423 & n11947;
  assign n11949 = pi0647 & n5423;
  assign n11950 = ~n11948 & ~n11949;
  assign n11951 = ~n8913 & ~n11950;
  assign n11952 = n8901 & n11947;
  assign n11953 = pi0647 & ~n8873;
  assign n11954 = n8907 & n11953;
  assign n11955 = ~n11952 & ~n11954;
  assign n11956 = ~n8872 & ~n8879;
  assign n11957 = pi0647 & n8891;
  assign n11958 = ~n8891 & n11947;
  assign n11959 = ~n11957 & ~n11958;
  assign n11960 = ~n8896 & n11959;
  assign n11961 = n8871 & ~n11960;
  assign n11962 = n11956 & n11961;
  assign n11963 = n11955 & ~n11962;
  assign n11964 = ~n11951 & n11963;
  assign po0757 = pi1747 & ~n11964;
  assign n11966 = pi0586 & n8472;
  assign n11967 = pi0648 & ~n11966;
  assign n11968 = ~pi0648 & n11966;
  assign n11969 = ~n11967 & ~n11968;
  assign n11970 = ~pi1697 & ~n11969;
  assign n11971 = pi0648 & n8417;
  assign n11972 = ~n8428 & ~n8431;
  assign n11973 = ~n8450 & ~n8460;
  assign n11974 = n11972 & n11973;
  assign n11975 = ~n11972 & ~n11973;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = ~n8417 & ~n11976;
  assign n11978 = ~n11971 & ~n11977;
  assign n11979 = pi1697 & ~n11978;
  assign n11980 = ~n11970 & ~n11979;
  assign po0758 = pi1143 & ~n11980;
  assign n11982 = n11053 & n11892;
  assign n11983 = n11173 & n11982;
  assign n11984 = pi0649 & ~n11983;
  assign n11985 = ~pi0649 & n11983;
  assign n11986 = ~n11984 & ~n11985;
  assign n11987 = ~pi1697 & ~n11986;
  assign n11988 = pi0649 & n8417;
  assign n11989 = pi0552 & ~n10853;
  assign n11990 = n11905 & n11989;
  assign n11991 = ~n11159 & n11990;
  assign n11992 = n11163 & n11990;
  assign n11993 = ~n11161 & n11992;
  assign n11994 = pi0552 & n10852;
  assign n11995 = ~n11902 & n11989;
  assign n11996 = ~n11994 & ~n11995;
  assign n11997 = ~n11993 & n11996;
  assign n11998 = ~n11991 & n11997;
  assign n11999 = pi0649 & n11998;
  assign n12000 = ~pi0649 & ~n11998;
  assign n12001 = ~n11999 & ~n12000;
  assign n12002 = ~n8417 & ~n12001;
  assign n12003 = ~n11988 & ~n12002;
  assign n12004 = pi1697 & ~n12003;
  assign n12005 = ~n11987 & ~n12004;
  assign po0759 = pi1143 & ~n12005;
  assign n12007 = pi0650 & ~n11128;
  assign n12008 = ~pi0650 & n11128;
  assign n12009 = ~n12007 & ~n12008;
  assign n12010 = ~pi1697 & ~n12009;
  assign n12011 = pi0650 & n8417;
  assign n12012 = ~n8433 & ~n8436;
  assign n12013 = n11712 & n12012;
  assign n12014 = ~n11712 & ~n12012;
  assign n12015 = ~n12013 & ~n12014;
  assign n12016 = ~n8417 & ~n12015;
  assign n12017 = ~n12011 & ~n12016;
  assign n12018 = pi1697 & ~n12017;
  assign n12019 = ~n12010 & ~n12018;
  assign po0760 = pi1143 & ~n12019;
  assign n12021 = ~pi1672 & ~n11729;
  assign n12022 = ~pi0651 & n11729;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = ~n11726 & ~n12023;
  assign n12025 = pi1802 & n11726;
  assign n12026 = ~n12024 & ~n12025;
  assign po0761 = ~pi1747 | ~n12026;
  assign n12028 = ~pi1666 & ~n11729;
  assign n12029 = ~pi0652 & n11729;
  assign n12030 = ~n12028 & ~n12029;
  assign n12031 = ~n11726 & ~n12030;
  assign n12032 = pi1805 & n11726;
  assign n12033 = ~n12031 & ~n12032;
  assign po0762 = ~pi1747 | ~n12033;
  assign n12035 = ~pi0653 & n11126;
  assign n12036 = pi0653 & ~n11126;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = ~pi1697 & ~n12037;
  assign n12039 = pi0653 & n8417;
  assign n12040 = ~n8441 & ~n8442;
  assign n12041 = ~n11192 & ~n12040;
  assign n12042 = n11192 & n12040;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = ~n8417 & ~n12043;
  assign n12045 = ~n12039 & ~n12044;
  assign n12046 = pi1697 & ~n12045;
  assign n12047 = ~n12038 & ~n12046;
  assign po0763 = pi1143 & ~n12047;
  assign n12049 = ~pi0654 & n11127;
  assign n12050 = pi0654 & ~n11127;
  assign n12051 = ~n12049 & ~n12050;
  assign n12052 = ~pi1697 & ~n12051;
  assign n12053 = pi0654 & n8417;
  assign n12054 = ~n8434 & ~n8439;
  assign n12055 = n11116 & n12054;
  assign n12056 = ~n11116 & ~n12054;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = ~n8417 & ~n12057;
  assign n12059 = ~n12053 & ~n12058;
  assign n12060 = pi1697 & ~n12059;
  assign n12061 = ~n12052 & ~n12060;
  assign po0764 = pi1143 & ~n12061;
  assign n12063 = pi0655 & ~n10902;
  assign n12064 = ~pi0655 & n10902;
  assign n12065 = ~n12063 & ~n12064;
  assign n12066 = ~pi1697 & ~n12065;
  assign n12067 = pi0655 & n8417;
  assign n12068 = ~n10861 & ~n10864;
  assign n12069 = n10879 & ~n10889;
  assign n12070 = n12068 & n12069;
  assign n12071 = ~n12068 & ~n12069;
  assign n12072 = ~n12070 & ~n12071;
  assign n12073 = ~n8417 & ~n12072;
  assign n12074 = ~n12067 & ~n12073;
  assign n12075 = pi1697 & ~n12074;
  assign n12076 = ~n12066 & ~n12075;
  assign po0765 = pi1143 & ~n12076;
  assign n12078 = pi1795 & n9430;
  assign n12079 = pi1215 & n8414;
  assign n12080 = pi0286 & n8413;
  assign n12081 = ~pi0656 & ~n8413;
  assign n12082 = ~n12080 & ~n12081;
  assign n12083 = ~n8414 & ~n12082;
  assign n12084 = ~n12079 & ~n12083;
  assign n12085 = ~n9430 & ~n12084;
  assign n12086 = pi1747 & ~n12085;
  assign po0766 = n12078 | ~n12086;
  assign n12088 = pi1797 & n9430;
  assign n12089 = pi1066 & n8414;
  assign n12090 = pi0254 & n8413;
  assign n12091 = ~pi0657 & ~n8413;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = ~n8414 & ~n12092;
  assign n12094 = ~n12089 & ~n12093;
  assign n12095 = ~n9430 & ~n12094;
  assign n12096 = pi1747 & ~n12095;
  assign po0767 = n12088 | ~n12096;
  assign n12098 = pi1801 & n9430;
  assign n12099 = pi1056 & n8414;
  assign n12100 = pi0124 & n8413;
  assign n12101 = ~pi0658 & ~n8413;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = ~n8414 & ~n12102;
  assign n12104 = ~n12099 & ~n12103;
  assign n12105 = ~n9430 & ~n12104;
  assign n12106 = pi1747 & ~n12105;
  assign po0768 = n12098 | ~n12106;
  assign n12108 = pi1783 & n9430;
  assign n12109 = ~pi1224 & n8414;
  assign n12110 = pi0022 & n8413;
  assign n12111 = ~pi0659 & ~n8413;
  assign n12112 = ~n12110 & ~n12111;
  assign n12113 = ~n8414 & ~n12112;
  assign n12114 = ~n12109 & ~n12113;
  assign n12115 = ~n9430 & ~n12114;
  assign n12116 = pi1747 & ~n12115;
  assign po0769 = n12108 | ~n12116;
  assign n12118 = ~pi0138 & pi0660;
  assign n12119 = ~pi0138 & pi1101;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = n3714 & ~n12120;
  assign n12122 = pi0660 & n8212;
  assign n12123 = ~pi1409 & n12118;
  assign n12124 = n7506 & n12123;
  assign n12125 = ~n12122 & ~n12124;
  assign n12126 = ~n12121 & n12125;
  assign po0770 = pi1747 & ~n12126;
  assign n12128 = pi0883 & ~pi1773;
  assign n12129 = pi1773 & pi1806;
  assign po0771 = n12128 | n12129;
  assign n12131 = pi0586 & ~pi0662;
  assign n12132 = ~pi0586 & pi0662;
  assign n12133 = ~n12131 & ~n12132;
  assign n12134 = ~pi1697 & ~n12133;
  assign n12135 = pi0662 & n8417;
  assign n12136 = ~n8443 & ~n8456;
  assign n12137 = ~n8459 & ~n12136;
  assign n12138 = n8459 & n12136;
  assign n12139 = ~n12137 & ~n12138;
  assign n12140 = ~n8417 & ~n12139;
  assign n12141 = ~n12135 & ~n12140;
  assign n12142 = pi1697 & ~n12141;
  assign n12143 = ~n12134 & ~n12142;
  assign po0772 = pi1143 & ~n12143;
  assign n12145 = pi0663 & n8486;
  assign n12146 = pi0709 & pi1102;
  assign n12147 = ~pi0709 & ~pi1102;
  assign n12148 = pi0720 & pi1110;
  assign n12149 = ~n12147 & n12148;
  assign n12150 = ~n12146 & ~n12149;
  assign n12151 = ~pi0720 & ~pi1110;
  assign n12152 = ~n12147 & ~n12151;
  assign n12153 = pi0679 & pi1109;
  assign n12154 = ~pi0679 & ~pi1109;
  assign n12155 = pi0707 & pi1081;
  assign n12156 = ~n12154 & n12155;
  assign n12157 = ~n12153 & ~n12156;
  assign n12158 = ~pi0707 & ~pi1081;
  assign n12159 = ~n12154 & ~n12158;
  assign n12160 = pi0710 & pi1108;
  assign n12161 = ~pi0710 & ~pi1108;
  assign n12162 = pi0669 & pi1107;
  assign n12163 = ~n12161 & n12162;
  assign n12164 = ~n12160 & ~n12163;
  assign n12165 = ~pi0669 & ~pi1107;
  assign n12166 = ~n12161 & ~n12165;
  assign n12167 = pi0699 & pi1106;
  assign n12168 = ~pi0699 & ~pi1106;
  assign n12169 = pi0698 & pi1338;
  assign n12170 = ~n12168 & n12169;
  assign n12171 = ~n12167 & ~n12170;
  assign n12172 = n12166 & ~n12171;
  assign n12173 = n12164 & ~n12172;
  assign n12174 = n12159 & ~n12173;
  assign n12175 = n12157 & ~n12174;
  assign n12176 = n12152 & ~n12175;
  assign n12177 = n12150 & ~n12176;
  assign n12178 = n12152 & n12159;
  assign n12179 = ~pi0698 & ~pi1338;
  assign n12180 = pi0700 & pi1105;
  assign n12181 = ~n12168 & n12180;
  assign n12182 = n12166 & n12181;
  assign n12183 = ~n12179 & n12182;
  assign n12184 = n12178 & n12183;
  assign n12185 = n12177 & ~n12184;
  assign n12186 = pi0663 & n12185;
  assign n12187 = ~pi0663 & ~n12185;
  assign n12188 = ~n12186 & ~n12187;
  assign n12189 = ~n8486 & ~n12188;
  assign n12190 = ~n12145 & ~n12189;
  assign n12191 = pi1699 & ~n12190;
  assign n12192 = ~pi0707 & ~pi0720;
  assign n12193 = ~pi0700 & ~pi0710;
  assign n12194 = ~pi0669 & ~pi0699;
  assign n12195 = ~pi0698 & n12194;
  assign n12196 = n12193 & n12195;
  assign n12197 = ~pi0709 & n12196;
  assign n12198 = ~pi0679 & n12197;
  assign n12199 = n12192 & n12198;
  assign n12200 = pi0663 & n12199;
  assign n12201 = ~pi0663 & ~n12199;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = ~pi1699 & n12202;
  assign n12204 = ~n12191 & ~n12203;
  assign po0773 = pi1111 & ~n12204;
  assign n12206 = n6806 & n6832;
  assign n12207 = pi0697 & pi0718;
  assign n12208 = pi0719 & n12207;
  assign n12209 = pi0708 & n12208;
  assign n12210 = n6815 & n12209;
  assign n12211 = n12206 & n12210;
  assign n12212 = pi0664 & ~n12211;
  assign n12213 = ~pi0664 & n12211;
  assign n12214 = ~n12212 & ~n12213;
  assign n12215 = ~pi1699 & ~n12214;
  assign n12216 = pi0664 & n8486;
  assign n12217 = ~n8493 & ~n8496;
  assign n12218 = ~n8500 & ~n8502;
  assign n12219 = ~n8503 & n8510;
  assign n12220 = ~n8508 & ~n12219;
  assign n12221 = n12218 & ~n12220;
  assign n12222 = ~n8500 & n8505;
  assign n12223 = ~n8497 & ~n12222;
  assign n12224 = ~n12221 & n12223;
  assign n12225 = n12217 & ~n12224;
  assign n12226 = ~n8493 & n8495;
  assign n12227 = ~n8490 & ~n12226;
  assign n12228 = ~n12225 & n12227;
  assign n12229 = ~n8489 & ~n12228;
  assign n12230 = ~pi0359 & ~n8488;
  assign n12231 = ~n12229 & n12230;
  assign n12232 = ~n8489 & n12217;
  assign n12233 = ~n8503 & ~n8511;
  assign n12234 = n12218 & n12233;
  assign n12235 = ~n8525 & ~n8528;
  assign n12236 = ~n8512 & ~n12235;
  assign n12237 = n12234 & ~n12236;
  assign n12238 = n12232 & n12237;
  assign n12239 = n12231 & ~n12238;
  assign n12240 = pi0664 & ~n12239;
  assign n12241 = ~pi0664 & n12239;
  assign n12242 = ~n12240 & ~n12241;
  assign n12243 = ~n8486 & ~n12242;
  assign n12244 = ~n12216 & ~n12243;
  assign n12245 = pi1699 & ~n12244;
  assign n12246 = ~n12215 & ~n12245;
  assign po0774 = pi1111 & ~n12246;
  assign n12248 = pi0665 & n8486;
  assign n12249 = n8501 & ~n8506;
  assign n12250 = ~n8509 & n12249;
  assign n12251 = n8499 & ~n12250;
  assign n12252 = n8494 & ~n12251;
  assign n12253 = n8526 & ~n8528;
  assign n12254 = n8514 & ~n12253;
  assign n12255 = n8501 & n8504;
  assign n12256 = ~n12254 & n12255;
  assign n12257 = n8494 & n12256;
  assign n12258 = ~pi0359 & ~pi0664;
  assign n12259 = ~n12257 & n12258;
  assign n12260 = n8492 & n12259;
  assign n12261 = ~n12252 & n12260;
  assign n12262 = pi0665 & ~n12261;
  assign n12263 = ~pi0665 & n12261;
  assign n12264 = ~n12262 & ~n12263;
  assign n12265 = ~n8486 & ~n12264;
  assign n12266 = ~n12248 & ~n12265;
  assign n12267 = pi1699 & ~n12266;
  assign n12268 = pi0678 & n12210;
  assign n12269 = n6832 & n12268;
  assign n12270 = pi0664 & n12269;
  assign n12271 = pi0675 & n12270;
  assign n12272 = pi0665 & n12271;
  assign n12273 = ~pi0665 & ~n12271;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = ~pi1699 & n12274;
  assign n12276 = ~n12267 & ~n12275;
  assign po0775 = pi1111 & ~n12276;
  assign n12278 = pi0885 & ~pi1773;
  assign n12279 = pi1773 & pi1808;
  assign po0776 = n12278 | n12279;
  assign n12281 = ~pi0667 & n11729;
  assign n12282 = pi0154 & ~n11729;
  assign n12283 = ~n12281 & ~n12282;
  assign n12284 = ~n11726 & ~n12283;
  assign n12285 = pi1799 & n11726;
  assign n12286 = ~n12284 & ~n12285;
  assign po0777 = ~pi1747 | ~n12286;
  assign n12288 = ~pi0668 & n11729;
  assign n12289 = pi0286 & ~n11729;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n11726 & ~n12290;
  assign n12292 = pi1795 & n11726;
  assign n12293 = ~n12291 & ~n12292;
  assign po0778 = ~pi1747 | ~n12293;
  assign n12295 = pi0669 & n8486;
  assign n12296 = ~n12162 & ~n12165;
  assign n12297 = ~n12168 & ~n12179;
  assign n12298 = n12180 & n12297;
  assign n12299 = n12171 & ~n12298;
  assign n12300 = ~n12296 & ~n12299;
  assign n12301 = n12296 & n12299;
  assign n12302 = ~n12300 & ~n12301;
  assign n12303 = ~n8486 & ~n12302;
  assign n12304 = ~n12295 & ~n12303;
  assign n12305 = pi1699 & ~n12304;
  assign n12306 = ~pi0698 & ~pi0700;
  assign n12307 = ~pi0699 & n12306;
  assign n12308 = ~pi0669 & n12307;
  assign n12309 = pi0669 & ~n12307;
  assign n12310 = ~n12308 & ~n12309;
  assign n12311 = ~pi1699 & ~n12310;
  assign n12312 = ~n12305 & ~n12311;
  assign po0779 = pi1111 & ~n12312;
  assign n12314 = ~pi0670 & n11729;
  assign n12315 = pi0064 & ~n11729;
  assign n12316 = ~n12314 & ~n12315;
  assign n12317 = ~n11726 & ~n12316;
  assign n12318 = pi1774 & n11726;
  assign n12319 = ~n12317 & ~n12318;
  assign po0780 = ~pi1747 | ~n12319;
  assign n12321 = ~pi0671 & n11729;
  assign n12322 = pi0310 & ~n11729;
  assign n12323 = ~n12321 & ~n12322;
  assign n12324 = ~n11726 & ~n12323;
  assign n12325 = pi1792 & n11726;
  assign n12326 = ~n12324 & ~n12325;
  assign po0781 = ~pi1747 | ~n12326;
  assign n12328 = ~pi0749 & ~pi0852;
  assign n12329 = ~pi0849 & pi0877;
  assign n12330 = pi0748 & pi0848;
  assign n12331 = ~n4699 & ~n12330;
  assign n12332 = pi0748 & ~pi0759;
  assign n12333 = ~pi0810 & pi0848;
  assign n12334 = ~n12332 & ~n12333;
  assign n12335 = n12331 & n12334;
  assign n12336 = ~pi0809 & pi0847;
  assign n12337 = pi0846 & pi0847;
  assign n12338 = ~pi0808 & n12337;
  assign n12339 = pi0846 & n4707;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = ~n12336 & n12340;
  assign n12342 = ~n12335 & ~n12341;
  assign n12343 = ~pi0759 & pi0848;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = ~pi0810 & n12330;
  assign n12346 = pi0748 & n4699;
  assign n12347 = ~n12345 & ~n12346;
  assign n12348 = n12344 & n12347;
  assign n12349 = ~n12329 & ~n12348;
  assign n12350 = pi0849 & ~pi0877;
  assign n12351 = ~n12349 & ~n12350;
  assign n12352 = n12328 & n12351;
  assign n12353 = ~pi0850 & n12352;
  assign n12354 = ~n4707 & ~n12337;
  assign n12355 = ~pi0809 & pi0846;
  assign n12356 = ~pi0808 & pi0847;
  assign n12357 = ~n12355 & ~n12356;
  assign n12358 = n12354 & n12357;
  assign n12359 = ~n12335 & ~n12358;
  assign n12360 = ~n12329 & n12359;
  assign n12361 = n12353 & ~n12360;
  assign n12362 = pi0751 & ~pi0755;
  assign n12363 = ~pi0807 & pi0845;
  assign n12364 = ~n12362 & ~n12363;
  assign n12365 = pi0751 & pi0845;
  assign n12366 = n12364 & ~n12365;
  assign n12367 = ~n4733 & n12366;
  assign n12368 = ~pi0806 & pi0842;
  assign n12369 = ~pi0804 & pi0844;
  assign n12370 = ~n12368 & ~n12369;
  assign n12371 = pi0842 & pi0844;
  assign n12372 = n12370 & ~n12371;
  assign n12373 = ~n4737 & n12372;
  assign n12374 = pi0750 & ~pi0754;
  assign n12375 = pi0841 & ~n12374;
  assign n12376 = pi0754 & ~n4754;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = ~n4757 & n12377;
  assign n12379 = ~n12373 & ~n12378;
  assign n12380 = ~n12367 & n12379;
  assign n12381 = pi0751 & n4733;
  assign n12382 = ~pi0807 & n12365;
  assign n12383 = ~n12381 & ~n12382;
  assign n12384 = ~pi0804 & n12371;
  assign n12385 = pi0842 & n4737;
  assign n12386 = ~n12384 & ~n12385;
  assign n12387 = ~pi0806 & pi0844;
  assign n12388 = n12386 & ~n12387;
  assign n12389 = ~n12367 & ~n12388;
  assign n12390 = n12383 & ~n12389;
  assign n12391 = ~pi0755 & pi0845;
  assign n12392 = n12390 & ~n12391;
  assign n12393 = n12353 & n12392;
  assign n12394 = ~n12380 & n12393;
  assign po0782 = n12361 | n12394;
  assign n12396 = ~n5861 & ~n5863;
  assign n12397 = n7076 & n12396;
  assign n12398 = ~n7076 & ~n12396;
  assign po0783 = n12397 | n12398;
  assign n12400 = pi0674 & n8486;
  assign n12401 = pi0663 & pi0715;
  assign n12402 = n12152 & n12401;
  assign n12403 = n12159 & ~n12164;
  assign n12404 = n12157 & ~n12403;
  assign n12405 = n12402 & ~n12404;
  assign n12406 = ~n12150 & n12401;
  assign n12407 = ~n12405 & ~n12406;
  assign n12408 = n12159 & n12166;
  assign n12409 = n12402 & n12408;
  assign n12410 = ~n12299 & n12409;
  assign n12411 = n12407 & ~n12410;
  assign n12412 = pi0674 & n12411;
  assign n12413 = ~pi0674 & ~n12411;
  assign n12414 = ~n12412 & ~n12413;
  assign n12415 = ~n8486 & ~n12414;
  assign n12416 = ~n12400 & ~n12415;
  assign n12417 = pi1699 & ~n12416;
  assign n12418 = ~pi0663 & ~pi0709;
  assign n12419 = ~pi0715 & ~pi0720;
  assign n12420 = ~pi0707 & ~pi0710;
  assign n12421 = ~pi0679 & n12420;
  assign n12422 = n12308 & n12421;
  assign n12423 = n12419 & n12422;
  assign n12424 = n12418 & n12423;
  assign n12425 = pi0674 & n12424;
  assign n12426 = ~pi0674 & ~n12424;
  assign n12427 = ~n12425 & ~n12426;
  assign n12428 = ~pi1699 & n12427;
  assign n12429 = ~n12417 & ~n12428;
  assign po0784 = pi1111 & ~n12429;
  assign n12431 = pi0675 & n8486;
  assign n12432 = ~n8490 & ~n8493;
  assign n12433 = n12251 & ~n12256;
  assign n12434 = ~n12432 & ~n12433;
  assign n12435 = n12432 & n12433;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = ~n8486 & ~n12436;
  assign n12438 = ~n12431 & ~n12437;
  assign n12439 = pi1699 & ~n12438;
  assign n12440 = pi0675 & n12268;
  assign n12441 = ~pi0675 & ~n12268;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~pi1699 & n12442;
  assign n12444 = ~n12439 & ~n12443;
  assign po0785 = pi1111 & ~n12444;
  assign n12446 = ~pi0383 & ~pi0481;
  assign n12447 = n8969 & n12446;
  assign n12448 = n9589 & n12447;
  assign n12449 = n9007 & n12448;
  assign n12450 = ~pi0410 & n12449;
  assign n12451 = n5806 & ~n12450;
  assign n12452 = pi1122 & n12451;
  assign n12453 = ~pi1173 & n6510;
  assign n12454 = ~pi1087 & ~pi1173;
  assign n12455 = pi0508 & n12454;
  assign n12456 = ~n12453 & ~n12455;
  assign n12457 = ~pi0408 & pi1241;
  assign n12458 = ~pi0507 & pi1077;
  assign n12459 = ~n12457 & ~n12458;
  assign n12460 = pi0507 & ~pi1077;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~n6510 & ~n12454;
  assign n12463 = pi0508 & ~pi1087;
  assign n12464 = pi0509 & ~pi1173;
  assign n12465 = ~n12463 & ~n12464;
  assign n12466 = n12462 & n12465;
  assign n12467 = ~n12461 & ~n12466;
  assign n12468 = n12456 & ~n12467;
  assign n12469 = pi0509 & ~pi1087;
  assign n12470 = n12468 & ~n12469;
  assign n12471 = ~pi1093 & ~pi1174;
  assign n12472 = ~n6531 & ~n12471;
  assign n12473 = pi0480 & ~pi1174;
  assign n12474 = pi0484 & ~pi1093;
  assign n12475 = ~n12473 & ~n12474;
  assign n12476 = n12472 & n12475;
  assign n12477 = ~n12470 & ~n12476;
  assign n12478 = ~pi1082 & ~pi1176;
  assign n12479 = pi0466 & ~pi1082;
  assign n12480 = pi0379 & ~pi1176;
  assign n12481 = ~n12479 & ~n12480;
  assign n12482 = ~n6548 & n12481;
  assign n12483 = ~n12478 & n12482;
  assign n12484 = ~pi1177 & ~pi1179;
  assign n12485 = pi0470 & ~pi1179;
  assign n12486 = pi0381 & ~pi1177;
  assign n12487 = ~n12485 & ~n12486;
  assign n12488 = ~n6539 & n12487;
  assign n12489 = ~n12484 & n12488;
  assign n12490 = pi0387 & ~pi1089;
  assign n12491 = ~pi0386 & pi1089;
  assign n12492 = ~pi1175 & ~n12491;
  assign n12493 = ~n12490 & ~n12492;
  assign n12494 = ~n6522 & n12493;
  assign n12495 = ~n12489 & ~n12494;
  assign n12496 = ~n12483 & n12495;
  assign n12497 = n12477 & n12496;
  assign n12498 = pi0480 & ~n12494;
  assign n12499 = ~pi1093 & n12498;
  assign n12500 = ~n12471 & ~n12473;
  assign n12501 = ~n12494 & ~n12500;
  assign n12502 = pi0484 & n12501;
  assign n12503 = ~pi1176 & n6548;
  assign n12504 = pi0466 & n12478;
  assign n12505 = ~n12503 & ~n12504;
  assign n12506 = pi0379 & ~pi1082;
  assign n12507 = n12505 & ~n12506;
  assign n12508 = ~n12489 & ~n12507;
  assign n12509 = pi0381 & ~pi1179;
  assign n12510 = ~n12508 & ~n12509;
  assign n12511 = ~pi1177 & n6539;
  assign n12512 = pi0470 & n12484;
  assign n12513 = ~n12511 & ~n12512;
  assign n12514 = n12510 & n12513;
  assign n12515 = pi0386 & ~pi1089;
  assign n12516 = n12514 & ~n12515;
  assign n12517 = ~n6522 & ~n12490;
  assign n12518 = ~pi1175 & ~n12517;
  assign n12519 = n12516 & ~n12518;
  assign n12520 = ~n12502 & n12519;
  assign n12521 = ~n12499 & n12520;
  assign n12522 = ~n12483 & ~n12489;
  assign n12523 = n12514 & ~n12522;
  assign n12524 = ~n12521 & ~n12523;
  assign n12525 = pi1256 & ~pi1257;
  assign n12526 = pi1122 & n12525;
  assign n12527 = ~n12524 & n12526;
  assign n12528 = ~n12497 & n12527;
  assign n12529 = ~n12452 & ~n12528;
  assign n12530 = ~pi1607 & ~n12529;
  assign n12531 = pi1690 & ~pi1734;
  assign po0786 = n12530 & n12531;
  assign n12533 = n3732 & n11654;
  assign n12534 = pi1401 & n12533;
  assign n12535 = ~n3736 & ~n3750;
  assign n12536 = ~pi0677 & ~n3731;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~n12534 & ~n12537;
  assign po0787 = pi1747 & ~n12538;
  assign n12540 = pi0678 & n8486;
  assign n12541 = ~n8495 & ~n8496;
  assign n12542 = n12224 & ~n12237;
  assign n12543 = ~n12541 & ~n12542;
  assign n12544 = n12541 & n12542;
  assign n12545 = ~n12543 & ~n12544;
  assign n12546 = ~n8486 & ~n12545;
  assign n12547 = ~n12540 & ~n12546;
  assign n12548 = pi1699 & ~n12547;
  assign n12549 = ~pi0678 & ~n12210;
  assign n12550 = ~n12268 & ~n12549;
  assign n12551 = ~pi1699 & n12550;
  assign n12552 = ~n12548 & ~n12551;
  assign po0788 = pi1111 & ~n12552;
  assign n12554 = pi0679 & n8486;
  assign n12555 = ~n12153 & ~n12154;
  assign n12556 = ~n12158 & ~n12161;
  assign n12557 = ~n12165 & n12167;
  assign n12558 = ~n12162 & ~n12557;
  assign n12559 = n12556 & ~n12558;
  assign n12560 = ~n12158 & n12160;
  assign n12561 = ~n12155 & ~n12560;
  assign n12562 = ~n12559 & n12561;
  assign n12563 = ~n12179 & n12180;
  assign n12564 = ~n12169 & ~n12563;
  assign n12565 = ~n12165 & ~n12168;
  assign n12566 = n12556 & n12565;
  assign n12567 = ~n12564 & n12566;
  assign n12568 = n12562 & ~n12567;
  assign n12569 = n12555 & n12568;
  assign n12570 = ~n12555 & ~n12568;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = ~n8486 & ~n12571;
  assign n12573 = ~n12554 & ~n12572;
  assign n12574 = pi1699 & ~n12573;
  assign n12575 = n12306 & n12420;
  assign n12576 = n12194 & n12575;
  assign n12577 = pi0679 & n12576;
  assign n12578 = ~pi0679 & ~n12576;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = ~pi1699 & n12579;
  assign n12581 = ~n12574 & ~n12580;
  assign po0789 = pi1111 & ~n12581;
  assign n12583 = ~pi0680 & n11729;
  assign n12584 = pi0014 & ~n11729;
  assign n12585 = ~n12583 & ~n12584;
  assign n12586 = ~n11726 & ~n12585;
  assign n12587 = pi1786 & n11726;
  assign n12588 = ~n12586 & ~n12587;
  assign po0790 = ~pi1747 | ~n12588;
  assign n12590 = ~pi0681 & n11729;
  assign n12591 = pi0015 & ~n11729;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n11726 & ~n12592;
  assign n12594 = pi1790 & n11726;
  assign n12595 = ~n12593 & ~n12594;
  assign po0791 = ~pi1747 | ~n12595;
  assign n12597 = ~pi0682 & n11729;
  assign n12598 = pi0953 & ~n11729;
  assign n12599 = ~n12597 & ~n12598;
  assign n12600 = ~n11726 & ~n12599;
  assign n12601 = pi1791 & n11726;
  assign n12602 = ~n12600 & ~n12601;
  assign po0792 = ~pi1747 | ~n12602;
  assign n12604 = ~pi0683 & n11729;
  assign n12605 = pi0332 & ~n11729;
  assign n12606 = ~n12604 & ~n12605;
  assign n12607 = ~n11726 & ~n12606;
  assign n12608 = pi1793 & n11726;
  assign n12609 = ~n12607 & ~n12608;
  assign po0793 = ~pi1747 | ~n12609;
  assign n12611 = ~pi0684 & n11729;
  assign n12612 = pi0057 & ~n11729;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = ~n11726 & ~n12613;
  assign n12615 = pi1775 & n11726;
  assign n12616 = ~n12614 & ~n12615;
  assign po0794 = ~pi1747 | ~n12616;
  assign n12618 = ~pi0685 & n11729;
  assign n12619 = pi0299 & ~n11729;
  assign n12620 = ~n12618 & ~n12619;
  assign n12621 = ~n11726 & ~n12620;
  assign n12622 = pi1794 & n11726;
  assign n12623 = ~n12621 & ~n12622;
  assign po0795 = ~pi1747 | ~n12623;
  assign n12625 = ~pi0686 & n11729;
  assign n12626 = pi1481 & ~n11729;
  assign n12627 = ~n12625 & ~n12626;
  assign n12628 = ~n11726 & ~n12627;
  assign n12629 = pi1796 & n11726;
  assign n12630 = ~n12628 & ~n12629;
  assign po0796 = ~pi1747 | ~n12630;
  assign n12632 = ~pi0687 & n11729;
  assign n12633 = pi0254 & ~n11729;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = ~n11726 & ~n12634;
  assign n12636 = pi1797 & n11726;
  assign n12637 = ~n12635 & ~n12636;
  assign po0797 = ~pi1747 | ~n12637;
  assign n12639 = ~pi0688 & n11729;
  assign n12640 = pi0223 & ~n11729;
  assign n12641 = ~n12639 & ~n12640;
  assign n12642 = ~n11726 & ~n12641;
  assign n12643 = pi1798 & n11726;
  assign n12644 = ~n12642 & ~n12643;
  assign po0798 = ~pi1747 | ~n12644;
  assign n12646 = ~pi0689 & n11729;
  assign n12647 = pi0124 & ~n11729;
  assign n12648 = ~n12646 & ~n12647;
  assign n12649 = ~n11726 & ~n12648;
  assign n12650 = pi1801 & n11726;
  assign n12651 = ~n12649 & ~n12650;
  assign po0799 = ~pi1747 | ~n12651;
  assign n12653 = ~pi0690 & n11729;
  assign n12654 = pi0155 & ~n11729;
  assign n12655 = ~n12653 & ~n12654;
  assign n12656 = ~n11726 & ~n12655;
  assign n12657 = pi1800 & n11726;
  assign n12658 = ~n12656 & ~n12657;
  assign po0800 = ~pi1747 | ~n12658;
  assign n12660 = ~pi0691 & n11729;
  assign n12661 = pi0063 & ~n11729;
  assign n12662 = ~n12660 & ~n12661;
  assign n12663 = ~n11726 & ~n12662;
  assign n12664 = pi1804 & n11726;
  assign n12665 = ~n12663 & ~n12664;
  assign po0801 = ~pi1747 | ~n12665;
  assign n12667 = ~pi0692 & n11729;
  assign n12668 = pi0056 & ~n11729;
  assign n12669 = ~n12667 & ~n12668;
  assign n12670 = ~n11726 & ~n12669;
  assign n12671 = pi1776 & n11726;
  assign n12672 = ~n12670 & ~n12671;
  assign po0802 = ~pi1747 | ~n12672;
  assign n12674 = ~pi0693 & n11729;
  assign n12675 = pi0022 & ~n11729;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = ~n11726 & ~n12676;
  assign n12678 = pi1783 & n11726;
  assign n12679 = ~n12677 & ~n12678;
  assign po0803 = ~pi1747 | ~n12679;
  assign n12681 = ~pi0694 & n11729;
  assign n12682 = pi0027 & ~n11729;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~n11726 & ~n12683;
  assign n12685 = pi1782 & n11726;
  assign n12686 = ~n12684 & ~n12685;
  assign po0804 = ~pi1747 | ~n12686;
  assign n12688 = n8871 & ~n8872;
  assign n12689 = ~n8879 & n12688;
  assign n12690 = ~n8896 & n12689;
  assign n12691 = ~pi0695 & n8891;
  assign n12692 = ~pi0695 & ~pi1626;
  assign n12693 = ~n8891 & n12692;
  assign n12694 = ~n12691 & ~n12693;
  assign n12695 = n12690 & n12694;
  assign n12696 = pi0695 & ~n8873;
  assign n12697 = n8907 & n12696;
  assign n12698 = ~n5423 & ~n12692;
  assign n12699 = pi0695 & n5423;
  assign n12700 = ~n12698 & ~n12699;
  assign n12701 = n8911 & ~n12700;
  assign n12702 = ~n12697 & ~n12701;
  assign po1535 = n8874 & n8911;
  assign n12704 = n12702 & ~po1535;
  assign n12705 = n5422 & ~n12700;
  assign n12706 = n8901 & ~n12692;
  assign n12707 = ~n12705 & ~n12706;
  assign n12708 = pi1747 & n12707;
  assign n12709 = n12704 & n12708;
  assign po0805 = n12695 | ~n12709;
  assign n12711 = pi0696 & ~pi1626;
  assign n12712 = ~n5423 & n12711;
  assign n12713 = pi0696 & n5423;
  assign n12714 = ~n12712 & ~n12713;
  assign n12715 = ~n8913 & ~n12714;
  assign n12716 = n8901 & n12711;
  assign n12717 = ~pi0696 & ~n8873;
  assign n12718 = n8907 & ~n12717;
  assign n12719 = ~n12716 & ~n12718;
  assign n12720 = ~pi0696 & n8891;
  assign n12721 = ~n8891 & ~n12711;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = n12690 & n12722;
  assign n12724 = n12719 & ~n12723;
  assign n12725 = ~n12715 & n12724;
  assign po0806 = pi1747 & ~n12725;
  assign n12727 = pi0697 & n8486;
  assign n12728 = pi0697 & ~pi1105;
  assign n12729 = ~n8528 & ~n12728;
  assign n12730 = ~n8486 & ~n12729;
  assign n12731 = ~n12727 & ~n12730;
  assign n12732 = pi1699 & ~n12731;
  assign n12733 = ~pi0697 & ~pi1699;
  assign n12734 = ~n12732 & ~n12733;
  assign po0807 = pi1111 & ~n12734;
  assign n12736 = pi0698 & n8486;
  assign n12737 = ~n12169 & ~n12179;
  assign n12738 = n12180 & ~n12737;
  assign n12739 = ~n12180 & n12737;
  assign n12740 = ~n12738 & ~n12739;
  assign n12741 = ~n8486 & ~n12740;
  assign n12742 = ~n12736 & ~n12741;
  assign n12743 = pi1699 & ~n12742;
  assign n12744 = pi0698 & pi0700;
  assign n12745 = ~n12306 & ~n12744;
  assign n12746 = ~pi1699 & ~n12745;
  assign n12747 = ~n12743 & ~n12746;
  assign po0808 = pi1111 & ~n12747;
  assign n12749 = pi0699 & n8486;
  assign n12750 = ~n12167 & ~n12168;
  assign n12751 = ~n12564 & ~n12750;
  assign n12752 = n12564 & n12750;
  assign n12753 = ~n12751 & ~n12752;
  assign n12754 = ~n8486 & ~n12753;
  assign n12755 = ~n12749 & ~n12754;
  assign n12756 = pi1699 & ~n12755;
  assign n12757 = pi0699 & ~n12306;
  assign n12758 = ~n12307 & ~n12757;
  assign n12759 = ~pi1699 & ~n12758;
  assign n12760 = ~n12756 & ~n12759;
  assign po0809 = pi1111 & ~n12760;
  assign n12762 = pi0700 & n8486;
  assign n12763 = ~pi0700 & pi1105;
  assign n12764 = pi0700 & ~pi1105;
  assign n12765 = ~n12763 & ~n12764;
  assign n12766 = ~n8486 & ~n12765;
  assign n12767 = ~n12762 & ~n12766;
  assign n12768 = pi1699 & ~n12767;
  assign n12769 = ~pi0700 & ~pi1699;
  assign n12770 = ~n12768 & ~n12769;
  assign po0810 = pi1111 & ~n12770;
  assign n12772 = ~pi0997 & n5524;
  assign n12773 = pi0997 & ~n5524;
  assign po0811 = n12772 | n12773;
  assign n12775 = pi0702 & n3751;
  assign n12776 = pi1747 & n12775;
  assign n12777 = ~pi0702 & ~n3739;
  assign n12778 = n3746 & ~n12777;
  assign n12779 = ~n3741 & ~n11649;
  assign n12780 = ~n8004 & n12779;
  assign n12781 = n12778 & n12780;
  assign n12782 = pi1747 & n12781;
  assign po0812 = n12776 | n12782;
  assign n12784 = ~pi0703 & n11729;
  assign n12785 = pi0049 & ~n11729;
  assign n12786 = ~n12784 & ~n12785;
  assign n12787 = ~n11726 & ~n12786;
  assign n12788 = pi1777 & n11726;
  assign n12789 = ~n12787 & ~n12788;
  assign po0813 = ~pi1747 | ~n12789;
  assign n12791 = ~pi0704 & n11729;
  assign n12792 = pi0194 & ~n11729;
  assign n12793 = ~n12791 & ~n12792;
  assign n12794 = ~n11726 & ~n12793;
  assign n12795 = pi1803 & n11726;
  assign n12796 = ~n12794 & ~n12795;
  assign po0814 = ~pi1747 | ~n12796;
  assign n12798 = pi0707 & ~n12196;
  assign n12799 = ~pi0707 & n12196;
  assign n12800 = ~n12798 & ~n12799;
  assign n12801 = ~pi1699 & ~n12800;
  assign n12802 = pi0707 & n8486;
  assign n12803 = ~n12155 & ~n12158;
  assign n12804 = n12173 & ~n12183;
  assign n12805 = n12803 & n12804;
  assign n12806 = ~n12803 & ~n12804;
  assign n12807 = ~n12805 & ~n12806;
  assign n12808 = ~n8486 & ~n12807;
  assign n12809 = ~n12802 & ~n12808;
  assign n12810 = pi1699 & ~n12809;
  assign n12811 = ~n12801 & ~n12810;
  assign po0816 = pi1111 & ~n12811;
  assign n12813 = ~pi0708 & n12208;
  assign n12814 = pi0708 & ~n12208;
  assign n12815 = ~n12813 & ~n12814;
  assign n12816 = ~pi1699 & ~n12815;
  assign n12817 = pi0708 & n8486;
  assign n12818 = ~n8503 & ~n8508;
  assign n12819 = n12254 & n12818;
  assign n12820 = ~n12254 & ~n12818;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n8486 & ~n12821;
  assign n12823 = ~n12817 & ~n12822;
  assign n12824 = pi1699 & ~n12823;
  assign n12825 = ~n12816 & ~n12824;
  assign po0817 = pi1111 & ~n12825;
  assign n12827 = ~pi0679 & ~pi0720;
  assign n12828 = n12420 & n12827;
  assign n12829 = n12308 & n12828;
  assign n12830 = pi0709 & ~n12829;
  assign n12831 = ~pi0709 & n12829;
  assign n12832 = ~n12830 & ~n12831;
  assign n12833 = ~pi1699 & ~n12832;
  assign n12834 = pi0709 & n8486;
  assign n12835 = ~n12146 & ~n12147;
  assign n12836 = ~n12151 & n12153;
  assign n12837 = ~n12148 & ~n12836;
  assign n12838 = ~n12564 & n12565;
  assign n12839 = n12558 & ~n12838;
  assign n12840 = n12556 & ~n12839;
  assign n12841 = n12561 & ~n12840;
  assign n12842 = ~n12151 & ~n12154;
  assign n12843 = ~n12841 & n12842;
  assign n12844 = n12837 & ~n12843;
  assign n12845 = ~n12835 & ~n12844;
  assign n12846 = n12835 & n12844;
  assign n12847 = ~n12845 & ~n12846;
  assign n12848 = ~n8486 & ~n12847;
  assign n12849 = ~n12834 & ~n12848;
  assign n12850 = pi1699 & ~n12849;
  assign n12851 = ~n12833 & ~n12850;
  assign po0818 = pi1111 & ~n12851;
  assign n12853 = pi0710 & ~n12308;
  assign n12854 = ~pi0710 & n12308;
  assign n12855 = ~n12853 & ~n12854;
  assign n12856 = ~pi1699 & ~n12855;
  assign n12857 = pi0710 & n8486;
  assign n12858 = ~n12160 & ~n12161;
  assign n12859 = ~n12839 & ~n12858;
  assign n12860 = n12839 & n12858;
  assign n12861 = ~n12859 & ~n12860;
  assign n12862 = ~n8486 & ~n12861;
  assign n12863 = ~n12857 & ~n12862;
  assign n12864 = pi1699 & ~n12863;
  assign n12865 = ~n12856 & ~n12864;
  assign po0819 = pi1111 & ~n12865;
  assign n12867 = ~pi0471 & ~pi0564;
  assign n12868 = n9977 & n12867;
  assign n12869 = n10983 & n12868;
  assign n12870 = n10015 & n12869;
  assign n12871 = ~pi0511 & n12870;
  assign n12872 = n5631 & ~n12871;
  assign n12873 = pi1131 & n12872;
  assign n12874 = ~pi1194 & n6333;
  assign n12875 = ~pi1194 & ~pi1195;
  assign n12876 = pi0587 & n12875;
  assign n12877 = ~n12874 & ~n12876;
  assign n12878 = ~pi0506 & pi1192;
  assign n12879 = ~pi0618 & pi1276;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = pi0618 & ~pi1276;
  assign n12882 = ~n12880 & ~n12881;
  assign n12883 = ~n6333 & ~n12875;
  assign n12884 = pi0587 & ~pi1195;
  assign n12885 = pi0622 & ~pi1194;
  assign n12886 = ~n12884 & ~n12885;
  assign n12887 = n12883 & n12886;
  assign n12888 = ~n12882 & ~n12887;
  assign n12889 = n12877 & ~n12888;
  assign n12890 = pi0622 & ~pi1195;
  assign n12891 = n12889 & ~n12890;
  assign n12892 = ~pi1196 & ~pi1264;
  assign n12893 = ~n6354 & ~n12892;
  assign n12894 = pi0549 & ~pi1196;
  assign n12895 = pi0567 & ~pi1264;
  assign n12896 = ~n12894 & ~n12895;
  assign n12897 = n12893 & n12896;
  assign n12898 = ~n12891 & ~n12897;
  assign n12899 = ~pi1199 & ~pi1249;
  assign n12900 = pi0533 & ~pi1249;
  assign n12901 = pi0380 & ~pi1199;
  assign n12902 = ~n12900 & ~n12901;
  assign n12903 = ~n6371 & n12902;
  assign n12904 = ~n12899 & n12903;
  assign n12905 = ~pi1036 & ~pi1201;
  assign n12906 = pi0562 & ~pi1036;
  assign n12907 = pi0468 & ~pi1201;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = ~n6362 & n12908;
  assign n12910 = ~n12905 & n12909;
  assign n12911 = pi0485 & ~pi1198;
  assign n12912 = ~pi0483 & pi1198;
  assign n12913 = ~pi1197 & ~n12912;
  assign n12914 = ~n12911 & ~n12913;
  assign n12915 = ~n6345 & n12914;
  assign n12916 = ~n12910 & ~n12915;
  assign n12917 = ~n12904 & n12916;
  assign n12918 = n12898 & n12917;
  assign n12919 = pi0549 & ~n12915;
  assign n12920 = ~pi1264 & n12919;
  assign n12921 = ~n12892 & ~n12894;
  assign n12922 = ~n12915 & ~n12921;
  assign n12923 = pi0567 & n12922;
  assign n12924 = ~pi1199 & n6371;
  assign n12925 = pi0533 & n12899;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = pi0380 & ~pi1249;
  assign n12928 = n12926 & ~n12927;
  assign n12929 = ~n12910 & ~n12928;
  assign n12930 = pi0468 & ~pi1036;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = ~pi1201 & n6362;
  assign n12933 = pi0562 & n12905;
  assign n12934 = ~n12932 & ~n12933;
  assign n12935 = n12931 & n12934;
  assign n12936 = pi0483 & ~pi1198;
  assign n12937 = n12935 & ~n12936;
  assign n12938 = ~n6345 & ~n12911;
  assign n12939 = ~pi1197 & ~n12938;
  assign n12940 = n12937 & ~n12939;
  assign n12941 = ~n12923 & n12940;
  assign n12942 = ~n12920 & n12941;
  assign n12943 = ~n12904 & ~n12910;
  assign n12944 = n12935 & ~n12943;
  assign n12945 = ~n12942 & ~n12944;
  assign n12946 = pi1080 & ~pi1132;
  assign n12947 = pi1131 & n12946;
  assign n12948 = ~n12945 & n12947;
  assign n12949 = ~n12918 & n12948;
  assign n12950 = ~n12873 & ~n12949;
  assign n12951 = ~pi1608 & ~n12950;
  assign n12952 = pi1679 & ~pi1730;
  assign po0820 = n12951 & n12952;
  assign n12954 = n6806 & n6815;
  assign n12955 = n12209 & n12954;
  assign n12956 = pi0712 & ~n12955;
  assign n12957 = ~pi0712 & n12955;
  assign n12958 = ~n12956 & ~n12957;
  assign n12959 = ~pi1699 & ~n12958;
  assign n12960 = pi0712 & n8486;
  assign n12961 = ~n8488 & ~n8489;
  assign n12962 = n12233 & ~n12236;
  assign n12963 = n12220 & ~n12962;
  assign n12964 = n12218 & ~n12963;
  assign n12965 = n12223 & ~n12964;
  assign n12966 = n12217 & ~n12965;
  assign n12967 = n12227 & ~n12966;
  assign n12968 = n12961 & n12967;
  assign n12969 = ~n12961 & ~n12967;
  assign n12970 = ~n12968 & ~n12969;
  assign n12971 = ~n8486 & ~n12970;
  assign n12972 = ~n12960 & ~n12971;
  assign n12973 = pi1699 & ~n12972;
  assign n12974 = ~n12959 & ~n12973;
  assign po0821 = pi1111 & ~n12974;
  assign n12976 = ~pi0563 & ~pi0649;
  assign n12977 = n11053 & n12976;
  assign n12978 = n11893 & n12977;
  assign n12979 = n10901 & n12978;
  assign n12980 = ~pi0594 & n12979;
  assign n12981 = n5792 & ~n12980;
  assign n12982 = pi1143 & n12981;
  assign n12983 = ~pi0586 & pi1213;
  assign n12984 = ~pi0662 & pi1214;
  assign n12985 = ~n12983 & ~n12984;
  assign n12986 = pi0662 & ~pi1214;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~pi1215 & ~pi1216;
  assign n12989 = ~n6432 & ~n12988;
  assign n12990 = pi0653 & ~pi1216;
  assign n12991 = pi0654 & ~pi1215;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = n12989 & n12992;
  assign n12994 = ~n12987 & ~n12993;
  assign n12995 = pi0653 & n12988;
  assign n12996 = ~pi1215 & n6432;
  assign n12997 = ~n12995 & ~n12996;
  assign n12998 = ~n12994 & n12997;
  assign n12999 = pi0654 & ~pi1216;
  assign n13000 = n12998 & ~n12999;
  assign n13001 = ~pi1056 & ~pi1057;
  assign n13002 = pi0358 & ~pi1056;
  assign n13003 = pi0623 & ~pi1057;
  assign n13004 = ~n13002 & ~n13003;
  assign n13005 = ~n6470 & n13004;
  assign n13006 = ~n13001 & n13005;
  assign n13007 = ~pi1232 & ~pi1266;
  assign n13008 = pi0645 & ~pi1266;
  assign n13009 = pi0621 & ~pi1232;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~n6461 & n13010;
  assign n13012 = ~n13007 & n13011;
  assign n13013 = pi0569 & ~pi1219;
  assign n13014 = ~pi0566 & pi1219;
  assign n13015 = ~pi1218 & ~n13014;
  assign n13016 = ~n13013 & ~n13015;
  assign n13017 = ~n6444 & n13016;
  assign n13018 = ~n13012 & ~n13017;
  assign n13019 = ~pi1066 & ~pi1217;
  assign n13020 = pi0648 & ~pi1066;
  assign n13021 = pi0650 & ~pi1217;
  assign n13022 = ~n13020 & ~n13021;
  assign n13023 = ~n6453 & n13022;
  assign n13024 = ~n13019 & n13023;
  assign n13025 = n13018 & ~n13024;
  assign n13026 = ~n13006 & n13025;
  assign n13027 = ~n13000 & n13026;
  assign n13028 = pi0648 & ~n13017;
  assign n13029 = ~pi1217 & n13028;
  assign n13030 = ~n13019 & ~n13020;
  assign n13031 = ~n13017 & ~n13030;
  assign n13032 = pi0650 & n13031;
  assign n13033 = pi0358 & ~n13012;
  assign n13034 = ~pi1057 & n13033;
  assign n13035 = ~n13001 & ~n13002;
  assign n13036 = ~n13012 & ~n13035;
  assign n13037 = pi0623 & n13036;
  assign n13038 = ~pi1232 & n6461;
  assign n13039 = pi0645 & n13007;
  assign n13040 = ~n13038 & ~n13039;
  assign n13041 = pi0621 & ~pi1266;
  assign n13042 = n13040 & ~n13041;
  assign n13043 = ~n13037 & n13042;
  assign n13044 = ~n13034 & n13043;
  assign n13045 = pi0566 & ~pi1219;
  assign n13046 = n13044 & ~n13045;
  assign n13047 = ~n6444 & ~n13013;
  assign n13048 = ~pi1218 & ~n13047;
  assign n13049 = n13046 & ~n13048;
  assign n13050 = ~n13032 & n13049;
  assign n13051 = ~n13029 & n13050;
  assign n13052 = ~n13006 & ~n13012;
  assign n13053 = n13044 & ~n13052;
  assign n13054 = ~n13051 & ~n13053;
  assign n13055 = pi1144 & ~pi1259;
  assign n13056 = pi1143 & n13055;
  assign n13057 = ~n13054 & n13056;
  assign n13058 = ~n13027 & n13057;
  assign n13059 = ~n12982 & ~n13058;
  assign n13060 = ~pi1583 & ~n13059;
  assign n13061 = pi1697 & ~pi1743;
  assign po0822 = n13060 & n13061;
  assign n13063 = pi0697 & n8541;
  assign n13064 = pi0714 & ~n13063;
  assign n13065 = ~pi0714 & n13063;
  assign n13066 = ~n13064 & ~n13065;
  assign n13067 = ~pi1699 & ~n13066;
  assign n13068 = pi0714 & n8486;
  assign n13069 = ~n8497 & ~n8500;
  assign n13070 = ~n8519 & ~n8529;
  assign n13071 = n13069 & n13070;
  assign n13072 = ~n13069 & ~n13070;
  assign n13073 = ~n13071 & ~n13072;
  assign n13074 = ~n8486 & ~n13073;
  assign n13075 = ~n13068 & ~n13074;
  assign n13076 = pi1699 & ~n13075;
  assign n13077 = ~n13067 & ~n13076;
  assign po0823 = pi1111 & ~n13077;
  assign n13079 = n12418 & n12827;
  assign n13080 = n12576 & n13079;
  assign n13081 = pi0715 & ~n13080;
  assign n13082 = ~pi0715 & n13080;
  assign n13083 = ~n13081 & ~n13082;
  assign n13084 = ~pi1699 & ~n13083;
  assign n13085 = pi0715 & n8486;
  assign n13086 = pi0663 & ~n12147;
  assign n13087 = n12842 & n13086;
  assign n13088 = ~n12562 & n13087;
  assign n13089 = n12566 & n13087;
  assign n13090 = ~n12564 & n13089;
  assign n13091 = pi0663 & n12146;
  assign n13092 = ~n12837 & n13086;
  assign n13093 = ~n13091 & ~n13092;
  assign n13094 = ~n13090 & n13093;
  assign n13095 = ~n13088 & n13094;
  assign n13096 = pi0715 & n13095;
  assign n13097 = ~pi0715 & ~n13095;
  assign n13098 = ~n13096 & ~n13097;
  assign n13099 = ~n8486 & ~n13098;
  assign n13100 = ~n13085 & ~n13099;
  assign n13101 = pi1699 & ~n13100;
  assign n13102 = ~n13084 & ~n13101;
  assign po0824 = pi1111 & ~n13102;
  assign n13104 = n3746 & ~n8004;
  assign n13105 = pi0716 & ~n3739;
  assign n13106 = ~n3741 & ~n13105;
  assign n13107 = ~n11649 & ~n13106;
  assign n13108 = n13104 & n13107;
  assign n13109 = pi0716 & n3737;
  assign n13110 = ~n13108 & ~n13109;
  assign po0825 = pi1747 & ~n13110;
  assign n13112 = pi0717 & ~n12209;
  assign n13113 = ~pi0717 & n12209;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = ~pi1699 & ~n13114;
  assign n13116 = pi0717 & n8486;
  assign n13117 = ~n8502 & ~n8505;
  assign n13118 = n12963 & n13117;
  assign n13119 = ~n12963 & ~n13117;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = ~n8486 & ~n13120;
  assign n13122 = ~n13116 & ~n13121;
  assign n13123 = pi1699 & ~n13122;
  assign n13124 = ~n13115 & ~n13123;
  assign po0826 = pi1111 & ~n13124;
  assign n13126 = pi0697 & ~pi0718;
  assign n13127 = ~pi0697 & pi0718;
  assign n13128 = ~n13126 & ~n13127;
  assign n13129 = ~pi1699 & ~n13128;
  assign n13130 = pi0718 & n8486;
  assign n13131 = ~n8512 & ~n8525;
  assign n13132 = ~n8528 & ~n13131;
  assign n13133 = n8528 & n13131;
  assign n13134 = ~n13132 & ~n13133;
  assign n13135 = ~n8486 & ~n13134;
  assign n13136 = ~n13130 & ~n13135;
  assign n13137 = pi1699 & ~n13136;
  assign n13138 = ~n13129 & ~n13137;
  assign po0827 = pi1111 & ~n13138;
  assign n13140 = ~pi0719 & n12207;
  assign n13141 = pi0719 & ~n12207;
  assign n13142 = ~n13140 & ~n13141;
  assign n13143 = ~pi1699 & ~n13142;
  assign n13144 = pi0719 & n8486;
  assign n13145 = ~n8510 & ~n8511;
  assign n13146 = ~n12236 & ~n13145;
  assign n13147 = n12236 & n13145;
  assign n13148 = ~n13146 & ~n13147;
  assign n13149 = ~n8486 & ~n13148;
  assign n13150 = ~n13144 & ~n13149;
  assign n13151 = pi1699 & ~n13150;
  assign n13152 = ~n13143 & ~n13151;
  assign po0828 = pi1111 & ~n13152;
  assign n13154 = pi0720 & ~n12422;
  assign n13155 = ~pi0720 & n12422;
  assign n13156 = ~n13154 & ~n13155;
  assign n13157 = ~pi1699 & ~n13156;
  assign n13158 = pi0720 & n8486;
  assign n13159 = ~n12148 & ~n12151;
  assign n13160 = ~n12299 & n12408;
  assign n13161 = n12404 & ~n13160;
  assign n13162 = n13159 & n13161;
  assign n13163 = ~n13159 & ~n13161;
  assign n13164 = ~n13162 & ~n13163;
  assign n13165 = ~n8486 & ~n13164;
  assign n13166 = ~n13158 & ~n13165;
  assign n13167 = pi1699 & ~n13166;
  assign n13168 = ~n13157 & ~n13167;
  assign po0829 = pi1111 & ~n13168;
  assign n13170 = ~pi0674 & ~pi0715;
  assign n13171 = n12418 & n13170;
  assign n13172 = n12828 & n13171;
  assign n13173 = n12195 & n13172;
  assign n13174 = ~pi0700 & n13173;
  assign n13175 = n5886 & ~n13174;
  assign n13176 = pi1111 & n13175;
  assign n13177 = ~pi0697 & pi1331;
  assign n13178 = ~pi0718 & pi1283;
  assign n13179 = ~n13177 & ~n13178;
  assign n13180 = pi0718 & ~pi1283;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = ~pi1154 & ~pi1155;
  assign n13183 = ~n6794 & ~n13182;
  assign n13184 = pi0719 & ~pi1155;
  assign n13185 = pi0708 & ~pi1154;
  assign n13186 = ~n13184 & ~n13185;
  assign n13187 = n13183 & n13186;
  assign n13188 = ~n13181 & ~n13187;
  assign n13189 = pi0719 & n13182;
  assign n13190 = ~pi1154 & n6794;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n13188 & n13191;
  assign n13193 = pi0708 & ~pi1155;
  assign n13194 = n13192 & ~n13193;
  assign n13195 = ~pi1159 & ~pi1346;
  assign n13196 = pi0359 & ~pi1346;
  assign n13197 = pi0712 & ~pi1159;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = ~n6832 & n13198;
  assign n13200 = ~n13195 & n13199;
  assign n13201 = ~pi1160 & ~pi1269;
  assign n13202 = pi0664 & ~pi1160;
  assign n13203 = pi0665 & ~pi1269;
  assign n13204 = ~n13202 & ~n13203;
  assign n13205 = ~n6823 & n13204;
  assign n13206 = ~n13201 & n13205;
  assign n13207 = pi0678 & ~pi1158;
  assign n13208 = ~pi0675 & pi1158;
  assign n13209 = ~pi1275 & ~n13208;
  assign n13210 = ~n13207 & ~n13209;
  assign n13211 = ~n6806 & n13210;
  assign n13212 = ~n13206 & ~n13211;
  assign n13213 = ~pi1156 & ~pi1157;
  assign n13214 = pi0714 & ~pi1156;
  assign n13215 = pi0717 & ~pi1157;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = ~n6815 & n13216;
  assign n13218 = ~n13213 & n13217;
  assign n13219 = n13212 & ~n13218;
  assign n13220 = ~n13200 & n13219;
  assign n13221 = ~n13194 & n13220;
  assign n13222 = pi0714 & ~n13211;
  assign n13223 = ~pi1157 & n13222;
  assign n13224 = ~n13213 & ~n13214;
  assign n13225 = ~n13211 & ~n13224;
  assign n13226 = pi0717 & n13225;
  assign n13227 = pi0359 & ~n13206;
  assign n13228 = ~pi1159 & n13227;
  assign n13229 = ~n13195 & ~n13196;
  assign n13230 = ~n13206 & ~n13229;
  assign n13231 = pi0712 & n13230;
  assign n13232 = ~pi1269 & n6823;
  assign n13233 = pi0664 & n13201;
  assign n13234 = ~n13232 & ~n13233;
  assign n13235 = pi0665 & ~pi1160;
  assign n13236 = n13234 & ~n13235;
  assign n13237 = ~n13231 & n13236;
  assign n13238 = ~n13228 & n13237;
  assign n13239 = pi0675 & ~pi1158;
  assign n13240 = n13238 & ~n13239;
  assign n13241 = ~n6806 & ~n13207;
  assign n13242 = ~pi1275 & ~n13241;
  assign n13243 = n13240 & ~n13242;
  assign n13244 = ~n13226 & n13243;
  assign n13245 = ~n13223 & n13244;
  assign n13246 = ~n13200 & ~n13206;
  assign n13247 = n13238 & ~n13246;
  assign n13248 = ~n13245 & ~n13247;
  assign n13249 = pi1112 & ~pi1113;
  assign n13250 = pi1111 & n13249;
  assign n13251 = ~n13248 & n13250;
  assign n13252 = ~n13221 & n13251;
  assign n13253 = ~n13176 & ~n13252;
  assign n13254 = ~pi1604 & ~n13253;
  assign n13255 = pi1699 & ~pi1728;
  assign po0830 = n13254 & n13255;
  assign n13257 = n8896 & n12689;
  assign n13258 = n5422 & n8874;
  assign n13259 = ~n13257 & ~n13258;
  assign n13260 = pi0722 & n13259;
  assign n13261 = pi0723 & ~pi0730;
  assign n13262 = ~pi0723 & pi0730;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = pi0738 & n13263;
  assign n13265 = ~pi0738 & ~n13263;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = ~pi1735 & pi1740;
  assign n13268 = pi1735 & ~pi1740;
  assign n13269 = ~n13267 & ~n13268;
  assign n13270 = ~pi1738 & n13269;
  assign n13271 = pi1738 & ~n13269;
  assign n13272 = ~n13270 & ~n13271;
  assign n13273 = ~n13266 & n13272;
  assign n13274 = n13266 & ~n13272;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276 = ~pi0731 & pi0744;
  assign n13277 = pi0731 & ~pi0744;
  assign n13278 = ~n13276 & ~n13277;
  assign n13279 = pi0727 & ~pi0732;
  assign n13280 = ~pi0727 & pi0732;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = pi1733 & ~pi1741;
  assign n13283 = ~pi1733 & pi1741;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = pi1722 & ~pi1727;
  assign n13286 = ~pi1722 & pi1727;
  assign n13287 = ~n13285 & ~n13286;
  assign n13288 = ~n13284 & n13287;
  assign n13289 = n13284 & ~n13287;
  assign n13290 = ~n13288 & ~n13289;
  assign n13291 = ~n13281 & n13290;
  assign n13292 = n13281 & ~n13290;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = ~n13278 & n13293;
  assign n13295 = n13278 & ~n13293;
  assign n13296 = ~n13294 & ~n13295;
  assign n13297 = ~n13275 & n13296;
  assign n13298 = n13275 & ~n13296;
  assign n13299 = ~n13297 & ~n13298;
  assign n13300 = ~n13259 & ~n13299;
  assign n13301 = ~n13260 & ~n13300;
  assign n13302 = pi1496 & ~pi1626;
  assign po0831 = ~n13301 | n13302;
  assign n13304 = pi0723 & n13259;
  assign n13305 = pi0733 & ~n13259;
  assign n13306 = ~n13304 & ~n13305;
  assign po0832 = n13302 | ~n13306;
  assign n13308 = pi0764 & pi0790;
  assign n13309 = ~pi0765 & pi0766;
  assign n13310 = n13308 & n13309;
  assign n13311 = ~n6709 & n6735;
  assign n13312 = n6739 & ~n6743;
  assign n13313 = n13311 & n13312;
  assign n13314 = n6709 & ~n6735;
  assign n13315 = ~n13311 & ~n13314;
  assign n13316 = ~pi0954 & n6715;
  assign n13317 = pi1050 & n13316;
  assign n13318 = n13315 & n13317;
  assign n13319 = ~n13313 & ~n13318;
  assign po1776 = pi1737 & pi1739;
  assign n13321 = ~pi1668 & po1776;
  assign n13322 = pi0276 & n13321;
  assign n13323 = ~n6759 & n13322;
  assign n13324 = n6709 & n13323;
  assign n13325 = ~n6735 & n13324;
  assign n13326 = n13319 & ~n13325;
  assign n13327 = ~n13310 & n13326;
  assign n13328 = pi0761 & pi0787;
  assign n13329 = ~pi0788 & ~n13328;
  assign n13330 = pi0783 & ~n13329;
  assign n13331 = n13326 & n13330;
  assign po0833 = n13327 | n13331;
  assign n13333 = pi0238 & ~pi0804;
  assign n13334 = ~pi0237 & ~n13333;
  assign n13335 = pi0750 & n13334;
  assign n13336 = ~pi0238 & pi0804;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = pi0257 & ~pi0859;
  assign n13339 = pi0750 & ~n13333;
  assign n13340 = ~n13334 & ~n13339;
  assign n13341 = ~n13338 & ~n13340;
  assign n13342 = n13337 & ~n13341;
  assign n13343 = ~pi0236 & pi0877;
  assign n13344 = ~pi0236 & ~pi0243;
  assign n13345 = ~pi0243 & pi0877;
  assign n13346 = ~n13344 & ~n13345;
  assign n13347 = pi0759 & ~n13346;
  assign n13348 = pi0236 & ~pi0877;
  assign n13349 = pi0759 & ~n13348;
  assign n13350 = ~n13344 & ~n13349;
  assign n13351 = ~n13345 & n13350;
  assign n13352 = ~pi0224 & ~pi0242;
  assign n13353 = ~pi0242 & pi0810;
  assign n13354 = ~n13352 & ~n13353;
  assign n13355 = ~n13351 & ~n13354;
  assign n13356 = pi0809 & n13355;
  assign n13357 = ~pi0224 & pi0810;
  assign n13358 = ~n13351 & n13357;
  assign n13359 = ~n13356 & ~n13358;
  assign n13360 = ~n13347 & n13359;
  assign n13361 = ~n13343 & n13360;
  assign n13362 = pi0224 & ~pi0810;
  assign n13363 = pi0809 & ~n13362;
  assign n13364 = ~n13352 & ~n13363;
  assign n13365 = ~n13353 & n13364;
  assign n13366 = ~n13351 & ~n13365;
  assign n13367 = n13361 & ~n13366;
  assign n13368 = ~pi0241 & pi0808;
  assign n13369 = n13361 & ~n13368;
  assign n13370 = ~pi0221 & ~pi0241;
  assign n13371 = pi0241 & ~pi0808;
  assign n13372 = pi0755 & ~n13371;
  assign n13373 = ~n13370 & ~n13372;
  assign n13374 = ~pi0221 & pi0808;
  assign n13375 = n13373 & ~n13374;
  assign n13376 = ~pi0239 & ~pi0240;
  assign n13377 = ~pi0239 & pi0807;
  assign n13378 = ~n13376 & ~n13377;
  assign n13379 = pi0806 & ~n13378;
  assign n13380 = ~pi0240 & pi0807;
  assign n13381 = ~n13379 & ~n13380;
  assign n13382 = ~n13375 & ~n13381;
  assign n13383 = ~n13370 & ~n13374;
  assign n13384 = pi0755 & ~n13383;
  assign n13385 = ~n13382 & ~n13384;
  assign n13386 = n13369 & n13385;
  assign n13387 = ~n13367 & ~n13386;
  assign n13388 = pi0797 & ~n13387;
  assign n13389 = n13342 & n13388;
  assign n13390 = pi0240 & ~pi0807;
  assign n13391 = pi0806 & ~n13390;
  assign n13392 = ~n13376 & ~n13391;
  assign n13393 = ~n13377 & n13392;
  assign n13394 = ~n13351 & ~n13375;
  assign n13395 = ~n13393 & n13394;
  assign n13396 = ~n13365 & n13395;
  assign n13397 = ~n13387 & ~n13396;
  assign n13398 = pi0797 & n13397;
  assign po0834 = n13389 | n13398;
  assign n13400 = ~n5859 & ~n5864;
  assign n13401 = ~n5858 & ~n13400;
  assign n13402 = n5858 & n13400;
  assign po0835 = n13401 | n13402;
  assign n13404 = pi0727 & n13259;
  assign n13405 = n13269 & ~n13287;
  assign n13406 = ~n13269 & n13287;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = pi0736 & ~pi0737;
  assign n13409 = ~pi0736 & pi0737;
  assign n13410 = ~n13408 & ~n13409;
  assign n13411 = ~pi1725 & pi1738;
  assign n13412 = pi1725 & ~pi1738;
  assign n13413 = ~n13411 & ~n13412;
  assign n13414 = ~n13410 & n13413;
  assign n13415 = n13410 & ~n13413;
  assign n13416 = ~n13414 & ~n13415;
  assign n13417 = ~n13407 & n13416;
  assign n13418 = n13407 & ~n13416;
  assign n13419 = ~n13417 & ~n13418;
  assign n13420 = pi0723 & ~pi0731;
  assign n13421 = ~pi0723 & pi0731;
  assign n13422 = ~n13420 & ~n13421;
  assign n13423 = pi0730 & ~pi0738;
  assign n13424 = ~pi0730 & pi0738;
  assign n13425 = ~n13423 & ~n13424;
  assign n13426 = ~n13422 & n13425;
  assign n13427 = n13422 & ~n13425;
  assign n13428 = ~n13426 & ~n13427;
  assign n13429 = ~pi0732 & pi0744;
  assign n13430 = pi0732 & ~pi0744;
  assign n13431 = ~n13429 & ~n13430;
  assign n13432 = pi0727 & n13284;
  assign n13433 = ~pi0727 & ~n13284;
  assign n13434 = ~n13432 & ~n13433;
  assign n13435 = ~n13431 & n13434;
  assign n13436 = n13431 & ~n13434;
  assign n13437 = ~n13435 & ~n13436;
  assign n13438 = ~n13428 & n13437;
  assign n13439 = n13428 & ~n13437;
  assign n13440 = ~n13438 & ~n13439;
  assign n13441 = ~n13419 & n13440;
  assign n13442 = n13419 & ~n13440;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~n13259 & ~n13443;
  assign n13445 = ~n13404 & ~n13444;
  assign po0836 = n13302 | ~n13445;
  assign n13447 = pi0728 & pi1424;
  assign n13448 = pi1747 & n13447;
  assign n13449 = pi1676 & n6325;
  assign n13450 = pi1726 & n13449;
  assign po0837 = n13448 | n13450;
  assign n13452 = pi0729 & n13259;
  assign n13453 = pi0737 & ~pi0738;
  assign n13454 = ~pi0737 & pi0738;
  assign n13455 = ~n13453 & ~n13454;
  assign n13456 = n13263 & ~n13455;
  assign n13457 = ~n13263 & n13455;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = n13278 & ~n13281;
  assign n13460 = ~n13278 & n13281;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = ~n13458 & n13461;
  assign n13463 = n13458 & ~n13461;
  assign n13464 = ~n13462 & ~n13463;
  assign n13465 = n13269 & ~n13413;
  assign n13466 = ~n13269 & n13413;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = ~n13290 & n13467;
  assign n13469 = n13290 & ~n13467;
  assign n13470 = ~n13468 & ~n13469;
  assign n13471 = ~n13464 & n13470;
  assign n13472 = n13464 & ~n13470;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = ~n13259 & ~n13473;
  assign n13475 = ~n13452 & ~n13474;
  assign po0838 = n13302 | ~n13475;
  assign n13477 = pi0730 & n13259;
  assign n13478 = pi0746 & ~n13259;
  assign n13479 = ~n13477 & ~n13478;
  assign po0839 = n13302 | ~n13479;
  assign n13481 = pi0731 & n13259;
  assign n13482 = pi0734 & ~n13259;
  assign n13483 = ~n13481 & ~n13482;
  assign po0840 = n13302 | ~n13483;
  assign n13485 = pi0732 & n13259;
  assign n13486 = pi0745 & ~n13259;
  assign n13487 = ~n13485 & ~n13486;
  assign po0841 = n13302 | ~n13487;
  assign n13489 = pi0733 & n13259;
  assign n13490 = pi1735 & ~pi1738;
  assign n13491 = ~pi1735 & pi1738;
  assign n13492 = ~n13490 & ~n13491;
  assign n13493 = ~n13425 & n13492;
  assign n13494 = n13425 & ~n13492;
  assign n13495 = ~n13493 & ~n13494;
  assign n13496 = ~n13259 & ~n13495;
  assign n13497 = ~n13489 & ~n13496;
  assign po0842 = n13302 | ~n13497;
  assign n13499 = pi0734 & n13259;
  assign n13500 = ~n13263 & n13269;
  assign n13501 = n13263 & ~n13269;
  assign n13502 = ~n13500 & ~n13501;
  assign n13503 = ~n13259 & ~n13502;
  assign n13504 = ~n13499 & ~n13503;
  assign po0843 = n13302 | ~n13504;
  assign n13506 = pi0735 & n13259;
  assign n13507 = pi1727 & ~pi1740;
  assign n13508 = ~pi1727 & pi1740;
  assign n13509 = ~n13507 & ~n13508;
  assign n13510 = ~n13422 & n13509;
  assign n13511 = n13422 & ~n13509;
  assign n13512 = ~n13510 & ~n13511;
  assign n13513 = ~n13259 & ~n13512;
  assign n13514 = ~n13506 & ~n13513;
  assign po0844 = n13302 | ~n13514;
  assign n13516 = pi0736 & n13259;
  assign n13517 = ~pi1722 & pi1741;
  assign n13518 = pi1722 & ~pi1741;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = ~n13431 & n13519;
  assign n13521 = n13431 & ~n13519;
  assign n13522 = ~n13520 & ~n13521;
  assign n13523 = ~n13259 & ~n13522;
  assign n13524 = ~n13516 & ~n13523;
  assign po0845 = n13302 | ~n13524;
  assign n13526 = pi0737 & n13259;
  assign n13527 = pi0729 & ~pi0732;
  assign n13528 = ~pi0729 & pi0732;
  assign n13529 = ~n13527 & ~n13528;
  assign n13530 = n13434 & ~n13529;
  assign n13531 = ~n13434 & n13529;
  assign n13532 = ~n13530 & ~n13531;
  assign n13533 = ~n13259 & ~n13532;
  assign n13534 = ~n13526 & ~n13533;
  assign po0846 = n13302 | ~n13534;
  assign n13536 = pi0738 & n13259;
  assign n13537 = pi0722 & pi1733;
  assign n13538 = ~pi0722 & ~pi1733;
  assign n13539 = ~n13537 & ~n13538;
  assign n13540 = pi0727 & n13539;
  assign n13541 = ~pi0727 & ~n13539;
  assign n13542 = ~n13540 & ~n13541;
  assign n13543 = ~n13259 & ~n13542;
  assign n13544 = ~n13536 & ~n13543;
  assign po0847 = n13302 | ~n13544;
  assign n13546 = pi0236 & pi0243;
  assign n13547 = pi0243 & ~pi0877;
  assign n13548 = ~n13546 & ~n13547;
  assign n13549 = ~pi0759 & ~n13548;
  assign n13550 = pi0242 & ~pi0810;
  assign n13551 = ~n7249 & ~n13550;
  assign n13552 = ~pi0759 & ~n13343;
  assign n13553 = ~n13547 & ~n13552;
  assign n13554 = ~n13546 & n13553;
  assign n13555 = ~n13551 & ~n13554;
  assign n13556 = ~pi0809 & n13555;
  assign n13557 = n13362 & ~n13554;
  assign n13558 = ~n13556 & ~n13557;
  assign n13559 = ~n13348 & n13558;
  assign n13560 = ~n13549 & n13559;
  assign n13561 = ~pi0809 & ~n13357;
  assign n13562 = ~n13550 & ~n13561;
  assign n13563 = ~n7249 & n13562;
  assign n13564 = ~n13554 & ~n13563;
  assign n13565 = n13560 & ~n13564;
  assign n13566 = ~n13371 & n13560;
  assign n13567 = pi0221 & ~pi0808;
  assign n13568 = ~n7135 & ~n13567;
  assign n13569 = ~pi0755 & ~n13568;
  assign n13570 = pi0239 & ~pi0807;
  assign n13571 = ~n7120 & ~n13570;
  assign n13572 = ~pi0806 & ~n13571;
  assign n13573 = ~n13390 & ~n13572;
  assign n13574 = ~pi0755 & ~n13368;
  assign n13575 = ~n7135 & ~n13574;
  assign n13576 = ~n13567 & n13575;
  assign n13577 = ~n13573 & ~n13576;
  assign n13578 = ~n13569 & ~n13577;
  assign n13579 = n13566 & n13578;
  assign n13580 = ~n13565 & ~n13579;
  assign n13581 = ~pi0806 & ~n13380;
  assign n13582 = ~n7120 & ~n13581;
  assign n13583 = ~n13570 & n13582;
  assign n13584 = ~n13554 & ~n13576;
  assign n13585 = ~n13583 & n13584;
  assign n13586 = ~n13563 & n13585;
  assign n13587 = pi0873 & ~n13586;
  assign n13588 = ~n13580 & n13587;
  assign n13589 = ~n6052 & ~n7121;
  assign n13590 = pi0237 & ~pi0804;
  assign n13591 = pi0238 & ~pi0750;
  assign n13592 = ~n13590 & ~n13591;
  assign n13593 = n13589 & n13592;
  assign n13594 = ~pi0257 & pi0859;
  assign n13595 = ~n13593 & ~n13594;
  assign n13596 = ~n13333 & ~n13595;
  assign n13597 = ~n13580 & n13596;
  assign n13598 = pi0237 & n6052;
  assign n13599 = ~pi0750 & n7121;
  assign n13600 = ~n13598 & ~n13599;
  assign n13601 = pi0873 & n13600;
  assign n13602 = n13597 & n13601;
  assign po0852 = n13588 | n13602;
  assign n13604 = pi0744 & n13259;
  assign n13605 = pi0735 & ~n13259;
  assign n13606 = ~n13604 & ~n13605;
  assign po0853 = n13302 | ~n13606;
  assign n13608 = pi0745 & n13259;
  assign n13609 = ~n13278 & n13287;
  assign n13610 = n13278 & ~n13287;
  assign n13611 = ~n13609 & ~n13610;
  assign n13612 = ~n13259 & ~n13611;
  assign n13613 = ~n13608 & ~n13612;
  assign po0854 = n13302 | ~n13613;
  assign n13615 = pi0746 & n13259;
  assign n13616 = n13413 & ~n13455;
  assign n13617 = ~n13413 & n13455;
  assign n13618 = ~n13616 & ~n13617;
  assign n13619 = ~n13259 & ~n13618;
  assign n13620 = ~n13615 & ~n13619;
  assign po0855 = n13302 | ~n13620;
  assign n13622 = pi0747 & n4339;
  assign n13623 = ~pi0048 & ~n4339;
  assign n13624 = ~n13622 & ~n13623;
  assign po0856 = n4458 | ~n13624;
  assign n13626 = pi0748 & ~po1343;
  assign n13627 = ~pi0667 & n6302;
  assign n13628 = ~n13626 & ~n13627;
  assign n13629 = ~pi0398 & po1538;
  assign n13630 = ~pi0497 & n6305;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~pi0580 & n6299;
  assign n13633 = n13631 & ~n13632;
  assign po0857 = ~n13628 | ~n13633;
  assign n13635 = pi0749 & ~po1343;
  assign n13636 = ~pi0704 & n6302;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = ~pi0377 & po1538;
  assign n13639 = ~pi0501 & n6305;
  assign n13640 = ~n13638 & ~n13639;
  assign n13641 = ~pi0581 & n6299;
  assign n13642 = n13640 & ~n13641;
  assign po0858 = ~n13637 | ~n13642;
  assign n13644 = pi0750 & ~po1343;
  assign n13645 = pi1104 & n6302;
  assign n13646 = ~n13644 & ~n13645;
  assign n13647 = pi1280 & po1538;
  assign n13648 = pi1092 & n6305;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = pi1271 & n6299;
  assign n13651 = n13649 & ~n13650;
  assign po0859 = ~n13646 | ~n13651;
  assign n13653 = pi0751 & ~po1343;
  assign n13654 = ~pi0668 & n6302;
  assign n13655 = ~n13653 & ~n13654;
  assign n13656 = ~pi0378 & po1538;
  assign n13657 = ~pi0494 & n6305;
  assign n13658 = ~n13656 & ~n13657;
  assign n13659 = ~pi0578 & n6299;
  assign n13660 = n13658 & ~n13659;
  assign po0860 = ~n13655 | ~n13660;
  assign n13662 = ~pi0752 & ~po1343;
  assign n13663 = ~pi0635 & n6302;
  assign n13664 = ~n13662 & ~n13663;
  assign n13665 = ~pi0318 & po1538;
  assign n13666 = ~pi0366 & n6305;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = ~pi0454 & n6299;
  assign n13669 = n13667 & ~n13668;
  assign po0861 = ~n13664 | ~n13669;
  assign n13671 = n8000 & n8001;
  assign n13672 = pi1760 & n13671;
  assign n13673 = ~pi0417 & n7999;
  assign n13674 = ~pi0440 & n8080;
  assign n13675 = ~n13673 & ~n13674;
  assign n13676 = ~pi1758 & ~pi1759;
  assign n13677 = pi1092 & n13676;
  assign n13678 = pi1758 & ~pi1759;
  assign n13679 = pi1037 & n13678;
  assign n13680 = ~n13677 & ~n13679;
  assign n13681 = n13675 & n13680;
  assign n13682 = n13672 & ~n13681;
  assign n13683 = n8001 & n9427;
  assign n13684 = ~pi1760 & n13683;
  assign n13685 = ~pi0529 & n7999;
  assign n13686 = ~pi0575 & n8080;
  assign n13687 = ~n13685 & ~n13686;
  assign n13688 = pi1271 & n13676;
  assign n13689 = pi1035 & n13678;
  assign n13690 = ~n13688 & ~n13689;
  assign n13691 = n13687 & n13690;
  assign n13692 = n13684 & ~n13691;
  assign n13693 = ~pi0599 & n7999;
  assign n13694 = ~pi0684 & n8080;
  assign n13695 = ~n13693 & ~n13694;
  assign n13696 = pi1104 & n13676;
  assign n13697 = pi1165 & n13678;
  assign n13698 = ~n13696 & ~n13697;
  assign n13699 = n13695 & n13698;
  assign n13700 = pi1760 & n13683;
  assign n13701 = ~n13699 & n13700;
  assign n13702 = ~n13692 & ~n13701;
  assign n13703 = ~pi1760 & n13676;
  assign n13704 = pi1479 & n13703;
  assign n13705 = ~pi1760 & n13678;
  assign n13706 = pi1095 & n13705;
  assign n13707 = ~n13704 & ~n13706;
  assign n13708 = ~pi1760 & n7999;
  assign n13709 = pi1319 & n13708;
  assign n13710 = pi1760 & n13678;
  assign n13711 = pi1684 & n13710;
  assign n13712 = ~pi1760 & n8080;
  assign n13713 = pi1487 & n13712;
  assign n13714 = ~n13711 & ~n13713;
  assign n13715 = pi1760 & n13676;
  assign n13716 = pi0474 & n13715;
  assign n13717 = n13714 & ~n13716;
  assign n13718 = ~n13709 & n13717;
  assign n13719 = n13707 & n13718;
  assign n13720 = ~pi1761 & ~pi1762;
  assign n13721 = n8001 & n13720;
  assign n13722 = ~pi1760 & n13721;
  assign n13723 = ~n13719 & n13722;
  assign n13724 = ~pi1760 & n13671;
  assign n13725 = ~pi0340 & n7999;
  assign n13726 = ~pi0394 & n8080;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = pi1280 & n13676;
  assign n13729 = pi0991 & n13678;
  assign n13730 = ~n13728 & ~n13729;
  assign n13731 = n13727 & n13730;
  assign n13732 = n13724 & ~n13731;
  assign n13733 = pi1760 & n13721;
  assign n13734 = ~n13719 & n13733;
  assign n13735 = ~n13732 & ~n13734;
  assign n13736 = ~n13723 & n13735;
  assign n13737 = n13702 & n13736;
  assign po0862 = n13682 | ~n13737;
  assign n13739 = pi0754 & ~po1343;
  assign n13740 = ~pi0671 & n6302;
  assign n13741 = ~n13739 & ~n13740;
  assign n13742 = ~pi0430 & po1538;
  assign n13743 = ~pi0491 & n6305;
  assign n13744 = ~n13742 & ~n13743;
  assign n13745 = ~pi0573 & n6299;
  assign n13746 = n13744 & ~n13745;
  assign po0863 = ~n13741 | ~n13746;
  assign n13748 = pi0755 & ~po1343;
  assign n13749 = pi1107 & n6302;
  assign n13750 = ~n13748 & ~n13749;
  assign n13751 = pi1272 & po1538;
  assign n13752 = pi1028 & n6305;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = pi1258 & n6299;
  assign n13755 = n13753 & ~n13754;
  assign po0864 = ~n13750 | ~n13755;
  assign n13757 = ~pi0756 & ~po1343;
  assign n13758 = ~pi0609 & n6302;
  assign n13759 = ~n13757 & ~n13758;
  assign n13760 = ~pi0348 & po1538;
  assign n13761 = ~pi0425 & n6305;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = ~pi0531 & n6299;
  assign n13764 = n13762 & ~n13763;
  assign po0865 = ~n13759 | ~n13764;
  assign n13766 = ~pi0757 & ~po1343;
  assign n13767 = ~pi0558 & n6302;
  assign n13768 = ~n13766 & ~n13767;
  assign n13769 = ~pi0324 & po1538;
  assign n13770 = ~pi0371 & n6305;
  assign n13771 = ~n13769 & ~n13770;
  assign n13772 = ~pi0459 & n6299;
  assign n13773 = n13771 & ~n13772;
  assign po0866 = ~n13768 | ~n13773;
  assign n13775 = ~pi0758 & ~po1343;
  assign n13776 = ~pi0636 & n6302;
  assign n13777 = ~n13775 & ~n13776;
  assign n13778 = ~pi0322 & po1538;
  assign n13779 = ~pi0369 & n6305;
  assign n13780 = ~n13778 & ~n13779;
  assign n13781 = ~pi0456 & n6299;
  assign n13782 = n13780 & ~n13781;
  assign po0867 = ~n13777 | ~n13782;
  assign n13784 = pi0759 & ~po1343;
  assign n13785 = pi1110 & n6302;
  assign n13786 = ~n13784 & ~n13785;
  assign n13787 = pi1267 & po1538;
  assign n13788 = pi1029 & n6305;
  assign n13789 = ~n13787 & ~n13788;
  assign n13790 = pi1034 & n6299;
  assign n13791 = n13789 & ~n13790;
  assign po0868 = ~n13786 | ~n13791;
  assign n13793 = pi0760 & ~n6753;
  assign po1782 = ~pi1737 & ~pi1739;
  assign n13795 = pi1674 & po1782;
  assign n13796 = n13793 & ~n13795;
  assign n13797 = ~pi1670 & ~n13796;
  assign n13798 = n6706 & n6712;
  assign n13799 = n6701 & n13798;
  assign n13800 = n6700 & n13799;
  assign n13801 = pi0773 & n13800;
  assign n13802 = ~pi0937 & n13801;
  assign n13803 = ~n13797 & n13802;
  assign n13804 = n6700 & n6702;
  assign n13805 = pi0760 & ~pi1021;
  assign n13806 = n13804 & n13805;
  assign n13807 = n13798 & n13806;
  assign n13808 = n13793 & n13807;
  assign n13809 = ~n13803 & ~n13808;
  assign n13810 = ~n13321 & n13793;
  assign n13811 = ~pi1670 & ~n13810;
  assign n13812 = pi0937 & n6700;
  assign n13813 = ~pi0773 & n13812;
  assign n13814 = n13799 & n13813;
  assign n13815 = ~n13811 & n13814;
  assign n13816 = n13809 & ~n13815;
  assign po1785 = ~pi1747 | pi1757;
  assign po0869 = ~n13816 & ~po1785;
  assign n13819 = ~pi1544 & n13326;
  assign n13820 = pi1345 & n13819;
  assign n13821 = pi0872 & pi1665;
  assign n13822 = pi0761 & ~n13821;
  assign n13823 = pi1673 & n13821;
  assign n13824 = ~n13822 & ~n13823;
  assign po0870 = n13820 & ~n13824;
  assign n13826 = pi0762 & ~po1343;
  assign n13827 = ~pi0542 & n6302;
  assign n13828 = ~n13826 & ~n13827;
  assign n13829 = ~pi0519 & po1538;
  assign n13830 = ~pi0616 & n6305;
  assign n13831 = ~n13829 & ~n13830;
  assign n13832 = ~pi0528 & n6299;
  assign n13833 = n13831 & ~n13832;
  assign po0871 = ~n13828 | ~n13833;
  assign n13835 = ~pi0791 & ~pi0792;
  assign n13836 = ~pi0763 & n13835;
  assign n13837 = pi0763 & ~n13835;
  assign n13838 = ~n13836 & ~n13837;
  assign n13839 = ~pi1665 & n13326;
  assign n13840 = pi1345 & n13839;
  assign po0872 = n13838 & n13840;
  assign n13842 = ~pi0764 & ~n13821;
  assign n13843 = pi1532 & n13821;
  assign n13844 = ~n13842 & ~n13843;
  assign po0873 = n13820 & ~n13844;
  assign n13846 = pi0765 & ~n13821;
  assign n13847 = pi1527 & n13821;
  assign n13848 = ~n13846 & ~n13847;
  assign po0874 = n13820 & ~n13848;
  assign n13850 = ~pi0766 & ~n13821;
  assign n13851 = pi1522 & n13821;
  assign n13852 = ~n13850 & ~n13851;
  assign po0875 = n13820 & ~n13852;
  assign n13854 = pi0767 & ~po1343;
  assign n13855 = pi0992 & n6302;
  assign n13856 = ~n13854 & ~n13855;
  assign n13857 = pi0861 & po1538;
  assign n13858 = pi0938 & n6305;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = pi0967 & n6299;
  assign n13861 = n13859 & ~n13860;
  assign po0876 = ~n13856 | ~n13861;
  assign n13863 = pi0768 & ~po1343;
  assign n13864 = ~pi0608 & n6302;
  assign n13865 = ~n13863 & ~n13864;
  assign n13866 = ~pi0347 & po1538;
  assign n13867 = ~pi0424 & n6305;
  assign n13868 = ~n13866 & ~n13867;
  assign n13869 = ~pi0530 & n6299;
  assign n13870 = n13868 & ~n13869;
  assign po0877 = ~n13865 | ~n13870;
  assign n13872 = pi1060 & ~pi1773;
  assign n13873 = pi1773 & pi1829;
  assign po0878 = n13872 | n13873;
  assign n13875 = pi0770 & ~po1343;
  assign n13876 = ~pi0546 & n6302;
  assign n13877 = ~n13875 & ~n13876;
  assign n13878 = ~pi0342 & po1538;
  assign n13879 = ~pi0419 & n6305;
  assign n13880 = ~n13878 & ~n13879;
  assign n13881 = ~pi0656 & n6299;
  assign n13882 = n13880 & ~n13881;
  assign po0879 = ~n13877 | ~n13882;
  assign n13884 = pi0771 & ~po1343;
  assign n13885 = pi1113 & n6302;
  assign n13886 = ~n13884 & ~n13885;
  assign n13887 = pi1257 & po1538;
  assign n13888 = pi1132 & n6305;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = pi1259 & n6299;
  assign n13891 = n13889 & ~n13890;
  assign po0880 = ~n13886 | ~n13891;
  assign n13893 = pi0772 & ~po1343;
  assign n13894 = ~pi0544 & n6302;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = ~pi0345 & po1538;
  assign n13897 = ~pi0422 & n6305;
  assign n13898 = ~n13896 & ~n13897;
  assign n13899 = ~pi0527 & n6299;
  assign n13900 = n13898 & ~n13899;
  assign po0881 = ~n13895 | ~n13900;
  assign n13902 = pi0773 & ~n6753;
  assign n13903 = ~n6753 & n13321;
  assign n13904 = ~n13902 & ~n13903;
  assign n13905 = n13814 & ~n13904;
  assign n13906 = ~pi1670 & n13905;
  assign n13907 = ~pi0278 & ~pi0773;
  assign n13908 = ~pi1045 & n6712;
  assign n13909 = n6707 & n13908;
  assign n13910 = n6699 & n13909;
  assign n13911 = pi0984 & n13910;
  assign n13912 = ~n13907 & n13911;
  assign n13913 = ~n13906 & ~n13912;
  assign n13914 = n13802 & n13902;
  assign n13915 = ~pi1670 & ~n13795;
  assign n13916 = n13914 & n13915;
  assign n13917 = n13913 & ~n13916;
  assign po0882 = ~po1785 & ~n13917;
  assign n13919 = ~pi0826 & pi0877;
  assign n13920 = ~pi0759 & pi0772;
  assign n13921 = ~pi0810 & pi0825;
  assign n13922 = ~n13920 & ~n13921;
  assign n13923 = pi0772 & pi0825;
  assign n13924 = n13922 & ~n13923;
  assign n13925 = ~n4699 & n13924;
  assign n13926 = ~pi0809 & pi0824;
  assign n13927 = pi0823 & pi0824;
  assign n13928 = ~pi0808 & n13927;
  assign n13929 = pi0823 & n4707;
  assign n13930 = ~n13928 & ~n13929;
  assign n13931 = ~n13926 & n13930;
  assign n13932 = ~n13925 & ~n13931;
  assign n13933 = ~pi0759 & pi0825;
  assign n13934 = ~n13932 & ~n13933;
  assign n13935 = ~pi0810 & n13923;
  assign n13936 = pi0772 & n4699;
  assign n13937 = ~n13935 & ~n13936;
  assign n13938 = n13934 & n13937;
  assign n13939 = ~n13919 & ~n13938;
  assign n13940 = pi0826 & ~pi0877;
  assign n13941 = ~n13939 & ~n13940;
  assign n13942 = ~pi0809 & pi0823;
  assign n13943 = ~pi0808 & pi0824;
  assign n13944 = ~n13942 & ~n13943;
  assign n13945 = ~n13927 & n13944;
  assign n13946 = ~n4707 & n13945;
  assign n13947 = pi0770 & pi0822;
  assign n13948 = ~pi0807 & n13947;
  assign n13949 = pi0770 & n4733;
  assign n13950 = ~n13948 & ~n13949;
  assign n13951 = ~pi0755 & pi0770;
  assign n13952 = ~pi0807 & pi0822;
  assign n13953 = ~n13951 & ~n13952;
  assign n13954 = ~n13947 & n13953;
  assign n13955 = ~n4733 & n13954;
  assign n13956 = pi0750 & ~pi0871;
  assign n13957 = pi0818 & ~n13956;
  assign n13958 = pi0871 & ~n4754;
  assign n13959 = ~n13957 & ~n13958;
  assign n13960 = ~n4757 & n13959;
  assign n13961 = ~pi0806 & pi0819;
  assign n13962 = ~pi0804 & pi0821;
  assign n13963 = ~n13961 & ~n13962;
  assign n13964 = pi0819 & pi0821;
  assign n13965 = n13963 & ~n13964;
  assign n13966 = ~n4737 & n13965;
  assign n13967 = ~n13960 & ~n13966;
  assign n13968 = ~n13955 & n13967;
  assign n13969 = ~pi0804 & n13964;
  assign n13970 = pi0819 & n4737;
  assign n13971 = ~n13969 & ~n13970;
  assign n13972 = ~pi0806 & pi0821;
  assign n13973 = n13971 & ~n13972;
  assign n13974 = ~n13955 & ~n13973;
  assign n13975 = ~pi0755 & pi0822;
  assign n13976 = ~n13974 & ~n13975;
  assign n13977 = ~n13968 & n13976;
  assign n13978 = n13950 & n13977;
  assign n13979 = ~n13919 & ~n13978;
  assign n13980 = ~n13925 & n13979;
  assign n13981 = ~n13946 & n13980;
  assign n13982 = ~pi0762 & ~pi0768;
  assign n13983 = ~n13981 & n13982;
  assign n13984 = ~pi0827 & n13983;
  assign po0885 = n13941 & n13984;
  assign n13986 = pi0777 & n4339;
  assign n13987 = ~pi0050 & ~n4339;
  assign n13988 = ~n13986 & ~n13987;
  assign po0886 = n4458 | ~n13988;
  assign n13990 = pi0778 & n4339;
  assign n13991 = ~pi0060 & ~n4339;
  assign n13992 = ~n13990 & ~n13991;
  assign po0887 = n4458 | ~n13992;
  assign n13994 = pi0779 & n4339;
  assign n13995 = ~pi0052 & ~n4339;
  assign n13996 = ~n13994 & ~n13995;
  assign po0888 = n4458 | ~n13996;
  assign n13998 = pi0780 & ~po1343;
  assign n13999 = ~pi1164 & n6302;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = ~pi1184 & po1538;
  assign n14002 = ~pi1206 & n6305;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = ~pi1225 & n6299;
  assign n14005 = n14003 & ~n14004;
  assign po0889 = ~n14000 | ~n14005;
  assign n14007 = pi1059 & ~pi1773;
  assign n14008 = pi1773 & pi1828;
  assign po0890 = n14007 | n14008;
  assign n14010 = pi1061 & ~pi1773;
  assign n14011 = pi1773 & pi1813;
  assign po0891 = n14010 | n14011;
  assign n14013 = pi0783 & ~n13821;
  assign n14014 = pi1550 & n13821;
  assign n14015 = ~n14013 & ~n14014;
  assign po0892 = n13820 & ~n14015;
  assign n14017 = pi1072 & ~pi1773;
  assign n14018 = pi1773 & pi1814;
  assign po0893 = n14017 | n14018;
  assign n14020 = ~pi0764 & ~pi0790;
  assign n14021 = n13309 & ~n14020;
  assign n14022 = n13326 & ~n14021;
  assign n14023 = ~pi0761 & ~pi0787;
  assign n14024 = ~pi0783 & n14023;
  assign n14025 = ~pi0788 & n14024;
  assign n14026 = n13309 & n14025;
  assign po0894 = n14022 & ~n14026;
  assign n14028 = pi0786 & pi1424;
  assign n14029 = pi1747 & n14028;
  assign n14030 = pi1424 & pi1675;
  assign n14031 = pi1747 & n14030;
  assign n14032 = pi1680 & n14031;
  assign po0895 = n14029 | n14032;
  assign n14034 = pi0787 & ~n13821;
  assign n14035 = pi1705 & n13821;
  assign n14036 = ~n14034 & ~n14035;
  assign po0896 = n13820 & ~n14036;
  assign n14038 = pi0788 & ~n13821;
  assign n14039 = pi1631 & n13821;
  assign n14040 = ~n14038 & ~n14039;
  assign po0897 = n13820 & ~n14040;
  assign n14042 = ~pi0917 & ~n13259;
  assign n14043 = ~pi0789 & ~po1526;
  assign n14044 = ~n14042 & ~n14043;
  assign po0898 = pi1747 & ~n14044;
  assign n14046 = ~pi0790 & ~n13821;
  assign n14047 = pi1546 & n13821;
  assign n14048 = ~n14046 & ~n14047;
  assign po0899 = n13820 & ~n14048;
  assign po0900 = pi0791 & n13840;
  assign n14051 = ~pi0791 & pi0792;
  assign n14052 = pi0791 & ~pi0792;
  assign n14053 = ~n14051 & ~n14052;
  assign po0901 = n13840 & ~n14053;
  assign n14055 = ~pi0793 & n13836;
  assign n14056 = pi0793 & ~n13836;
  assign n14057 = ~n14055 & ~n14056;
  assign po0902 = n13840 & n14057;
  assign n14059 = pi1315 & pi1747;
  assign n14060 = ~pi0794 & ~pi1751;
  assign po0903 = n14059 & ~n14060;
  assign n14062 = pi0795 & ~po1343;
  assign n14063 = ~pi1103 & n6302;
  assign n14064 = ~n14062 & ~n14063;
  assign n14065 = ~pi1120 & po1538;
  assign n14066 = ~pi1084 & n6305;
  assign n14067 = ~n14065 & ~n14066;
  assign n14068 = ~pi1140 & n6299;
  assign n14069 = n14067 & ~n14068;
  assign po0904 = ~n14064 | ~n14069;
  assign n14071 = pi0796 & ~po1343;
  assign n14072 = pi1111 & n6302;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = pi1122 & po1538;
  assign n14075 = pi1131 & n6305;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = pi1143 & n6299;
  assign n14078 = n14076 & ~n14077;
  assign po0905 = ~n14073 | ~n14078;
  assign n14080 = ~pi0797 & ~po1343;
  assign n14081 = pi1051 & n6302;
  assign n14082 = ~n14080 & ~n14081;
  assign n14083 = pi1025 & po1538;
  assign n14084 = ~pi1133 & n6305;
  assign n14085 = ~n14083 & ~n14084;
  assign n14086 = pi1255 & n6299;
  assign n14087 = n14085 & ~n14086;
  assign po0906 = ~n14082 | ~n14087;
  assign n14089 = pi0798 & ~po1343;
  assign n14090 = ~pi1361 & n6302;
  assign n14091 = ~n14089 & ~n14090;
  assign n14092 = ~pi1360 & po1538;
  assign n14093 = ~pi1369 & n6305;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = ~pi1413 & n6299;
  assign n14096 = n14094 & ~n14095;
  assign po0907 = ~n14091 | ~n14096;
  assign n14098 = pi0799 & ~po1343;
  assign n14099 = pi1118 & n6302;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = pi1124 & po1538;
  assign n14102 = ~pi1137 & n6305;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = pi1242 & n6299;
  assign n14105 = n14103 & ~n14104;
  assign po0908 = ~n14100 | ~n14105;
  assign n14107 = pi0800 & ~po1343;
  assign n14108 = pi1074 & n6302;
  assign n14109 = ~n14107 & ~n14108;
  assign n14110 = pi1252 & po1538;
  assign n14111 = ~pi1030 & n6305;
  assign n14112 = ~n14110 & ~n14111;
  assign n14113 = pi1261 & n6299;
  assign n14114 = n14112 & ~n14113;
  assign po0909 = ~n14109 | ~n14114;
  assign n14116 = pi0801 & ~po1343;
  assign n14117 = pi1112 & n6302;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = pi1256 & po1538;
  assign n14120 = pi1080 & n6305;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = pi1144 & n6299;
  assign n14123 = n14121 & ~n14122;
  assign po0910 = ~n14118 | ~n14123;
  assign n14125 = pi0802 & ~po1343;
  assign n14126 = pi0994 & n6302;
  assign n14127 = ~n14125 & ~n14126;
  assign n14128 = pi0863 & po1538;
  assign n14129 = pi0939 & n6305;
  assign n14130 = ~n14128 & ~n14129;
  assign n14131 = pi0969 & n6299;
  assign n14132 = n14130 & ~n14131;
  assign po0911 = ~n14127 | ~n14132;
  assign n14134 = pi0803 & ~po1343;
  assign n14135 = pi1014 & n6302;
  assign n14136 = ~n14134 & ~n14135;
  assign n14137 = pi0876 & po1538;
  assign n14138 = pi0942 & n6305;
  assign n14139 = ~n14137 & ~n14138;
  assign n14140 = pi0973 & n6299;
  assign n14141 = n14139 & ~n14140;
  assign po0912 = ~n14136 | ~n14141;
  assign n14143 = pi0804 & ~po1343;
  assign n14144 = pi1105 & n6302;
  assign n14145 = ~n14143 & ~n14144;
  assign n14146 = pi1022 & po1538;
  assign n14147 = pi1027 & n6305;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = pi1032 & n6299;
  assign n14150 = n14148 & ~n14149;
  assign po0913 = ~n14145 | ~n14150;
  assign n14152 = ~pi0805 & ~po1343;
  assign n14153 = pi0993 & n6302;
  assign n14154 = ~n14152 & ~n14153;
  assign n14155 = pi0862 & po1538;
  assign n14156 = pi0941 & n6305;
  assign n14157 = ~n14155 & ~n14156;
  assign n14158 = pi0968 & n6299;
  assign n14159 = n14157 & ~n14158;
  assign po0914 = ~n14154 | ~n14159;
  assign n14161 = pi0806 & ~po1343;
  assign n14162 = pi1338 & n6302;
  assign n14163 = ~n14161 & ~n14162;
  assign n14164 = pi1277 & po1538;
  assign n14165 = pi1310 & n6305;
  assign n14166 = ~n14164 & ~n14165;
  assign n14167 = pi1342 & n6299;
  assign n14168 = n14166 & ~n14167;
  assign po0915 = ~n14163 | ~n14168;
  assign n14170 = pi0807 & ~po1343;
  assign n14171 = pi1106 & n6302;
  assign n14172 = ~n14170 & ~n14171;
  assign n14173 = pi1023 & po1538;
  assign n14174 = pi1129 & n6305;
  assign n14175 = ~n14173 & ~n14174;
  assign n14176 = pi1141 & n6299;
  assign n14177 = n14175 & ~n14176;
  assign po0916 = ~n14172 | ~n14177;
  assign n14179 = pi0808 & ~po1343;
  assign n14180 = pi1108 & n6302;
  assign n14181 = ~n14179 & ~n14180;
  assign n14182 = pi1121 & po1538;
  assign n14183 = pi1083 & n6305;
  assign n14184 = ~n14182 & ~n14183;
  assign n14185 = pi1033 & n6299;
  assign n14186 = n14184 & ~n14185;
  assign po0917 = ~n14181 | ~n14186;
  assign n14188 = pi0809 & ~po1343;
  assign n14189 = pi1081 & n6302;
  assign n14190 = ~n14188 & ~n14189;
  assign n14191 = pi1274 & po1538;
  assign n14192 = pi1130 & n6305;
  assign n14193 = ~n14191 & ~n14192;
  assign n14194 = pi1142 & n6299;
  assign n14195 = n14193 & ~n14194;
  assign po0918 = ~n14190 | ~n14195;
  assign n14197 = pi0810 & ~po1343;
  assign n14198 = pi1109 & n6302;
  assign n14199 = ~n14197 & ~n14198;
  assign n14200 = pi1270 & po1538;
  assign n14201 = pi1076 & n6305;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = pi1265 & n6299;
  assign n14204 = n14202 & ~n14203;
  assign po0919 = ~n14199 | ~n14204;
  assign n14206 = ~pi0811 & ~po1343;
  assign n14207 = ~pi0593 & n6302;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~pi0337 & po1538;
  assign n14210 = ~pi0612 & n6305;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = ~pi0520 & n6299;
  assign n14213 = n14211 & ~n14212;
  assign po0920 = ~n14208 | ~n14213;
  assign n14215 = ~pi0812 & ~po1343;
  assign n14216 = ~pi0551 & n6302;
  assign n14217 = ~n14215 & ~n14216;
  assign n14218 = ~pi0316 & po1538;
  assign n14219 = ~pi0364 & n6305;
  assign n14220 = ~n14218 & ~n14219;
  assign n14221 = ~pi0451 & n6299;
  assign n14222 = n14220 & ~n14221;
  assign po0921 = ~n14217 | ~n14222;
  assign n14224 = ~pi0813 & ~po1343;
  assign n14225 = ~pi0555 & n6302;
  assign n14226 = ~n14224 & ~n14225;
  assign n14227 = ~pi0319 & po1538;
  assign n14228 = ~pi0367 & n6305;
  assign n14229 = ~n14227 & ~n14228;
  assign n14230 = ~pi0450 & n6299;
  assign n14231 = n14229 & ~n14230;
  assign po0922 = ~n14226 | ~n14231;
  assign n14233 = ~pi0814 & ~po1343;
  assign n14234 = ~pi0601 & n6302;
  assign n14235 = ~n14233 & ~n14234;
  assign n14236 = ~pi0516 & po1538;
  assign n14237 = ~pi0613 & n6305;
  assign n14238 = ~n14236 & ~n14237;
  assign n14239 = ~pi0439 & n6299;
  assign n14240 = n14238 & ~n14239;
  assign po0923 = ~n14235 | ~n14240;
  assign n14242 = ~pi0815 & ~po1343;
  assign n14243 = ~pi0554 & n6302;
  assign n14244 = ~n14242 & ~n14243;
  assign n14245 = ~pi0317 & po1538;
  assign n14246 = ~pi0365 & n6305;
  assign n14247 = ~n14245 & ~n14246;
  assign n14248 = ~pi0453 & n6299;
  assign n14249 = n14247 & ~n14248;
  assign po0924 = ~n14244 | ~n14249;
  assign n14251 = ~pi0816 & ~po1343;
  assign n14252 = ~pi0556 & n6302;
  assign n14253 = ~n14251 & ~n14252;
  assign n14254 = ~pi0320 & po1538;
  assign n14255 = ~pi0368 & n6305;
  assign n14256 = ~n14254 & ~n14255;
  assign n14257 = ~pi0455 & n6299;
  assign n14258 = n14256 & ~n14257;
  assign po0925 = ~n14253 | ~n14258;
  assign n14260 = ~pi0817 & ~po1343;
  assign n14261 = ~pi0595 & n6302;
  assign n14262 = ~n14260 & ~n14261;
  assign n14263 = ~pi0517 & po1538;
  assign n14264 = ~pi0414 & n6305;
  assign n14265 = ~n14263 & ~n14264;
  assign n14266 = ~pi0521 & n6299;
  assign n14267 = n14265 & ~n14266;
  assign po0926 = ~n14262 | ~n14267;
  assign n14269 = pi0818 & ~po1343;
  assign n14270 = ~pi0596 & n6302;
  assign n14271 = ~n14269 & ~n14270;
  assign n14272 = ~pi0518 & po1538;
  assign n14273 = ~pi0614 & n6305;
  assign n14274 = ~n14272 & ~n14273;
  assign n14275 = ~pi0522 & n6299;
  assign n14276 = n14274 & ~n14275;
  assign po0927 = ~n14271 | ~n14276;
  assign n14278 = pi0819 & ~po1343;
  assign n14279 = ~pi0598 & n6302;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = ~pi0339 & po1538;
  assign n14282 = ~pi0416 & n6305;
  assign n14283 = ~n14281 & ~n14282;
  assign n14284 = ~pi0444 & n6299;
  assign n14285 = n14283 & ~n14284;
  assign po0928 = ~n14280 | ~n14285;
  assign n14287 = ~pi0820 & ~po1343;
  assign n14288 = ~pi0599 & n6302;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = ~pi0340 & po1538;
  assign n14291 = ~pi0417 & n6305;
  assign n14292 = ~n14290 & ~n14291;
  assign n14293 = ~pi0529 & n6299;
  assign n14294 = n14292 & ~n14293;
  assign po0929 = ~n14289 | ~n14294;
  assign n14296 = pi0821 & ~po1343;
  assign n14297 = ~pi0600 & n6302;
  assign n14298 = ~n14296 & ~n14297;
  assign n14299 = ~pi0341 & po1538;
  assign n14300 = ~pi0418 & n6305;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = ~pi0524 & n6299;
  assign n14303 = n14301 & ~n14302;
  assign po0930 = ~n14298 | ~n14303;
  assign n14305 = pi0822 & ~po1343;
  assign n14306 = ~pi0604 & n6302;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = ~pi0438 & po1538;
  assign n14309 = ~pi0536 & n6305;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 = ~pi0525 & n6299;
  assign n14312 = n14310 & ~n14311;
  assign po0931 = ~n14307 | ~n14312;
  assign n14314 = pi0823 & ~po1343;
  assign n14315 = ~pi0602 & n6302;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = ~pi0343 & po1538;
  assign n14318 = ~pi0420 & n6305;
  assign n14319 = ~n14317 & ~n14318;
  assign n14320 = ~pi0657 & n6299;
  assign n14321 = n14319 & ~n14320;
  assign po0932 = ~n14316 | ~n14321;
  assign n14323 = pi0824 & ~po1343;
  assign n14324 = ~pi0603 & n6302;
  assign n14325 = ~n14323 & ~n14324;
  assign n14326 = ~pi0344 & po1538;
  assign n14327 = ~pi0421 & n6305;
  assign n14328 = ~n14326 & ~n14327;
  assign n14329 = ~pi0526 & n6299;
  assign n14330 = n14328 & ~n14329;
  assign po0933 = ~n14325 | ~n14330;
  assign n14332 = pi0825 & ~po1343;
  assign n14333 = ~pi0606 & n6302;
  assign n14334 = ~n14332 & ~n14333;
  assign n14335 = ~pi0346 & po1538;
  assign n14336 = ~pi0432 & n6305;
  assign n14337 = ~n14335 & ~n14336;
  assign n14338 = ~pi0629 & n6299;
  assign n14339 = n14337 & ~n14338;
  assign po0934 = ~n14334 | ~n14339;
  assign n14341 = pi0826 & ~po1343;
  assign n14342 = ~pi0605 & n6302;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = ~pi0314 & po1538;
  assign n14345 = ~pi0423 & n6305;
  assign n14346 = ~n14344 & ~n14345;
  assign n14347 = ~pi0658 & n6299;
  assign n14348 = n14346 & ~n14347;
  assign po0935 = ~n14343 | ~n14348;
  assign n14350 = pi0827 & ~po1343;
  assign n14351 = ~pi0515 & n6302;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = ~pi0311 & po1538;
  assign n14354 = ~pi0350 & n6305;
  assign n14355 = ~n14353 & ~n14354;
  assign n14356 = ~pi0427 & n6299;
  assign n14357 = n14355 & ~n14356;
  assign po0936 = ~n14352 | ~n14357;
  assign n14359 = ~pi0828 & ~po1343;
  assign n14360 = ~pi0607 & n6302;
  assign n14361 = ~n14359 & ~n14360;
  assign n14362 = ~pi0435 & po1538;
  assign n14363 = ~pi0534 & n6305;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = ~pi0626 & n6299;
  assign n14366 = n14364 & ~n14365;
  assign po0937 = ~n14361 | ~n14366;
  assign n14368 = ~pi0829 & ~po1343;
  assign n14369 = ~pi0437 & n6302;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = ~pi0312 & po1538;
  assign n14372 = ~pi0351 & n6305;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = ~pi0428 & n6299;
  assign n14375 = n14373 & ~n14374;
  assign po0938 = ~n14370 | ~n14375;
  assign n14377 = ~pi0830 & ~po1343;
  assign n14378 = ~pi0557 & n6302;
  assign n14379 = ~n14377 & ~n14378;
  assign n14380 = ~pi0458 & po1538;
  assign n14381 = ~pi0559 & n6305;
  assign n14382 = ~n14380 & ~n14381;
  assign n14383 = ~pi0632 & n6299;
  assign n14384 = n14382 & ~n14383;
  assign po0939 = ~n14379 | ~n14384;
  assign n14386 = ~pi0831 & ~po1343;
  assign n14387 = ~pi0547 & n6302;
  assign n14388 = ~n14386 & ~n14387;
  assign n14389 = ~pi0447 & po1538;
  assign n14390 = ~pi0548 & n6305;
  assign n14391 = ~n14389 & ~n14390;
  assign n14392 = ~pi0640 & n6299;
  assign n14393 = n14391 & ~n14392;
  assign po0940 = ~n14388 | ~n14393;
  assign n14395 = ~pi0832 & ~po1343;
  assign n14396 = ~pi0550 & n6302;
  assign n14397 = ~n14395 & ~n14396;
  assign n14398 = ~pi0321 & po1538;
  assign n14399 = ~pi0362 & n6305;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = ~pi0449 & n6299;
  assign n14402 = n14400 & ~n14401;
  assign po0941 = ~n14397 | ~n14402;
  assign n14404 = ~pi0833 & ~po1343;
  assign n14405 = ~pi0610 & n6302;
  assign n14406 = ~n14404 & ~n14405;
  assign n14407 = ~pi0349 & po1538;
  assign n14408 = ~pi0356 & n6305;
  assign n14409 = ~n14407 & ~n14408;
  assign n14410 = ~pi0436 & n6299;
  assign n14411 = n14409 & ~n14410;
  assign po0942 = ~n14406 | ~n14411;
  assign n14413 = ~pi0834 & ~po1343;
  assign n14414 = ~pi0611 & n6302;
  assign n14415 = ~n14413 & ~n14414;
  assign n14416 = ~pi0313 & po1538;
  assign n14417 = ~pi0426 & n6305;
  assign n14418 = ~n14416 & ~n14417;
  assign n14419 = ~pi0659 & n6299;
  assign n14420 = n14418 & ~n14419;
  assign po0943 = ~n14415 | ~n14420;
  assign n14422 = ~pi0835 & ~po1343;
  assign n14423 = ~pi0670 & n6302;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = ~pi0389 & po1538;
  assign n14426 = ~pi0487 & n6305;
  assign n14427 = ~n14425 & ~n14426;
  assign n14428 = ~pi0570 & n6299;
  assign n14429 = n14427 & ~n14428;
  assign po0944 = ~n14424 | ~n14429;
  assign n14431 = ~pi0836 & ~po1343;
  assign n14432 = ~pi0638 & n6302;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~pi0325 & po1538;
  assign n14435 = ~pi0372 & n6305;
  assign n14436 = ~n14434 & ~n14435;
  assign n14437 = ~pi0460 & n6299;
  assign n14438 = n14436 & ~n14437;
  assign po0945 = ~n14433 | ~n14438;
  assign n14440 = ~pi0837 & ~po1343;
  assign n14441 = ~pi0680 & n6302;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = ~pi0390 & po1538;
  assign n14444 = ~pi0488 & n6305;
  assign n14445 = ~n14443 & ~n14444;
  assign n14446 = ~pi0571 & n6299;
  assign n14447 = n14445 & ~n14446;
  assign po0946 = ~n14442 | ~n14447;
  assign n14449 = ~pi0838 & ~po1343;
  assign n14450 = ~pi0637 & n6302;
  assign n14451 = ~n14449 & ~n14450;
  assign n14452 = ~pi0323 & po1538;
  assign n14453 = ~pi0370 & n6305;
  assign n14454 = ~n14452 & ~n14453;
  assign n14455 = ~pi0457 & n6299;
  assign n14456 = n14454 & ~n14455;
  assign po0947 = ~n14451 | ~n14456;
  assign n14458 = ~pi0839 & ~po1343;
  assign n14459 = ~pi0639 & n6302;
  assign n14460 = ~n14458 & ~n14459;
  assign n14461 = ~pi0326 & po1538;
  assign n14462 = ~pi0373 & n6305;
  assign n14463 = ~n14461 & ~n14462;
  assign n14464 = ~pi0532 & n6299;
  assign n14465 = n14463 & ~n14464;
  assign po0948 = ~n14460 | ~n14465;
  assign n14467 = ~pi0840 & ~po1343;
  assign n14468 = ~pi0681 & n6302;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = ~pi0391 & po1538;
  assign n14471 = ~pi0489 & n6305;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = ~pi0572 & n6299;
  assign n14474 = n14472 & ~n14473;
  assign po0949 = ~n14469 | ~n14474;
  assign n14476 = pi0841 & ~po1343;
  assign n14477 = ~pi0682 & n6302;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~pi0392 & po1538;
  assign n14480 = ~pi0490 & n6305;
  assign n14481 = ~n14479 & ~n14480;
  assign n14482 = ~pi0543 & n6299;
  assign n14483 = n14481 & ~n14482;
  assign po0950 = ~n14478 | ~n14483;
  assign n14485 = pi0842 & ~po1343;
  assign n14486 = ~pi0683 & n6302;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = ~pi0393 & po1538;
  assign n14489 = ~pi0492 & n6305;
  assign n14490 = ~n14488 & ~n14489;
  assign n14491 = ~pi0574 & n6299;
  assign n14492 = n14490 & ~n14491;
  assign po0951 = ~n14487 | ~n14492;
  assign n14494 = ~pi0843 & ~po1343;
  assign n14495 = ~pi0684 & n6302;
  assign n14496 = ~n14494 & ~n14495;
  assign n14497 = ~pi0394 & po1538;
  assign n14498 = ~pi0440 & n6305;
  assign n14499 = ~n14497 & ~n14498;
  assign n14500 = ~pi0575 & n6299;
  assign n14501 = n14499 & ~n14500;
  assign po0952 = ~n14496 | ~n14501;
  assign n14503 = pi0844 & ~po1343;
  assign n14504 = ~pi0685 & n6302;
  assign n14505 = ~n14503 & ~n14504;
  assign n14506 = ~pi0395 & po1538;
  assign n14507 = ~pi0493 & n6305;
  assign n14508 = ~n14506 & ~n14507;
  assign n14509 = ~pi0538 & n6299;
  assign n14510 = n14508 & ~n14509;
  assign po0953 = ~n14505 | ~n14510;
  assign n14512 = pi0845 & ~po1343;
  assign n14513 = ~pi0686 & n6302;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = ~pi0396 & po1538;
  assign n14516 = ~pi0495 & n6305;
  assign n14517 = ~n14515 & ~n14516;
  assign n14518 = ~pi0576 & n6299;
  assign n14519 = n14517 & ~n14518;
  assign po0954 = ~n14514 | ~n14519;
  assign n14521 = pi0846 & ~po1343;
  assign n14522 = ~pi0687 & n6302;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = ~pi0399 & po1538;
  assign n14525 = ~pi0446 & n6305;
  assign n14526 = ~n14524 & ~n14525;
  assign n14527 = ~pi0577 & n6299;
  assign n14528 = n14526 & ~n14527;
  assign po0955 = ~n14523 | ~n14528;
  assign n14530 = pi0847 & ~po1343;
  assign n14531 = ~pi0688 & n6302;
  assign n14532 = ~n14530 & ~n14531;
  assign n14533 = ~pi0397 & po1538;
  assign n14534 = ~pi0496 & n6305;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~pi0540 & n6299;
  assign n14537 = n14535 & ~n14536;
  assign po0956 = ~n14532 | ~n14537;
  assign n14539 = pi0848 & ~po1343;
  assign n14540 = ~pi0690 & n6302;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = ~pi0401 & po1538;
  assign n14543 = ~pi0498 & n6305;
  assign n14544 = ~n14542 & ~n14543;
  assign n14545 = ~pi0579 & n6299;
  assign n14546 = n14544 & ~n14545;
  assign po0957 = ~n14541 | ~n14546;
  assign n14548 = pi0849 & ~po1343;
  assign n14549 = ~pi0689 & n6302;
  assign n14550 = ~n14548 & ~n14549;
  assign n14551 = ~pi0400 & po1538;
  assign n14552 = ~pi0445 & n6305;
  assign n14553 = ~n14551 & ~n14552;
  assign n14554 = ~pi0539 & n6299;
  assign n14555 = n14553 & ~n14554;
  assign po0958 = ~n14550 | ~n14555;
  assign n14557 = pi0850 & ~po1343;
  assign n14558 = ~pi0651 & n6302;
  assign n14559 = ~n14557 & ~n14558;
  assign n14560 = ~pi0334 & po1538;
  assign n14561 = ~pi0406 & n6305;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = ~pi0504 & n6299;
  assign n14564 = n14562 & ~n14563;
  assign po0959 = ~n14559 | ~n14564;
  assign n14566 = ~pi0851 & ~po1343;
  assign n14567 = ~pi0692 & n6302;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = ~pi0402 & po1538;
  assign n14570 = ~pi0499 & n6305;
  assign n14571 = ~n14569 & ~n14570;
  assign n14572 = ~pi0582 & n6299;
  assign n14573 = n14571 & ~n14572;
  assign po0960 = ~n14568 | ~n14573;
  assign n14575 = pi0852 & ~po1343;
  assign n14576 = ~pi0691 & n6302;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = ~pi0403 & po1538;
  assign n14579 = ~pi0500 & n6305;
  assign n14580 = ~n14578 & ~n14579;
  assign n14581 = ~pi0583 & n6299;
  assign n14582 = n14580 & ~n14581;
  assign po0961 = ~n14577 | ~n14582;
  assign n14584 = ~pi0853 & ~po1343;
  assign n14585 = ~pi0652 & n6302;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = ~pi0335 & po1538;
  assign n14588 = ~pi0407 & n6305;
  assign n14589 = ~n14587 & ~n14588;
  assign n14590 = ~pi0505 & n6299;
  assign n14591 = n14589 & ~n14590;
  assign po0962 = ~n14586 | ~n14591;
  assign n14593 = ~pi0854 & ~po1343;
  assign n14594 = ~pi0641 & n6302;
  assign n14595 = ~n14593 & ~n14594;
  assign n14596 = ~pi0328 & po1538;
  assign n14597 = ~pi0374 & n6305;
  assign n14598 = ~n14596 & ~n14597;
  assign n14599 = ~pi0462 & n6299;
  assign n14600 = n14598 & ~n14599;
  assign po0963 = ~n14595 | ~n14600;
  assign n14602 = ~pi0855 & ~po1343;
  assign n14603 = ~pi0628 & n6302;
  assign n14604 = ~n14602 & ~n14603;
  assign n14605 = ~pi0329 & po1538;
  assign n14606 = ~pi0376 & n6305;
  assign n14607 = ~n14605 & ~n14606;
  assign n14608 = ~pi0463 & n6299;
  assign n14609 = n14607 & ~n14608;
  assign po0964 = ~n14604 | ~n14609;
  assign n14611 = ~pi0856 & ~po1343;
  assign n14612 = ~pi0633 & n6302;
  assign n14613 = ~n14611 & ~n14612;
  assign n14614 = ~pi0327 & po1538;
  assign n14615 = ~pi0357 & n6305;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = ~pi0461 & n6299;
  assign n14618 = n14616 & ~n14617;
  assign po0965 = ~n14613 | ~n14618;
  assign n14620 = ~pi0857 & ~po1343;
  assign n14621 = ~pi0694 & n6302;
  assign n14622 = ~n14620 & ~n14621;
  assign n14623 = ~pi0404 & po1538;
  assign n14624 = ~pi0503 & n6305;
  assign n14625 = ~n14623 & ~n14624;
  assign n14626 = ~pi0584 & n6299;
  assign n14627 = n14625 & ~n14626;
  assign po0966 = ~n14622 | ~n14627;
  assign n14629 = ~pi0858 & ~po1343;
  assign n14630 = ~pi0693 & n6302;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~pi0405 & po1538;
  assign n14633 = ~pi0443 & n6305;
  assign n14634 = ~n14632 & ~n14633;
  assign n14635 = ~pi0585 & n6299;
  assign n14636 = n14634 & ~n14635;
  assign po0967 = ~n14631 | ~n14636;
  assign n14638 = pi0859 & ~po1343;
  assign n14639 = ~pi1237 & n6302;
  assign n14640 = ~n14638 & ~n14639;
  assign n14641 = ~pi1235 & po1538;
  assign n14642 = ~pi1126 & n6305;
  assign n14643 = ~n14641 & ~n14642;
  assign n14644 = ~pi1031 & n6299;
  assign n14645 = n14643 & ~n14644;
  assign po0968 = ~n14640 | ~n14645;
  assign n14647 = pi0860 & ~po1343;
  assign n14648 = ~pi1243 & n6302;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = ~pi1268 & po1538;
  assign n14651 = ~pi1128 & n6305;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = ~pi1273 & n6299;
  assign n14654 = n14652 & ~n14653;
  assign po0969 = ~n14649 | ~n14654;
  assign n14656 = pi1430 & pi1698;
  assign n14657 = pi0064 & n14656;
  assign n14658 = pi0861 & ~n14656;
  assign n14659 = ~n14657 & ~n14658;
  assign po0970 = pi1747 & ~n14659;
  assign n14661 = pi0862 & ~n14656;
  assign n14662 = pi0057 & n14656;
  assign n14663 = ~n14661 & ~n14662;
  assign po0971 = pi1747 & ~n14663;
  assign n14665 = pi1430 & pi1695;
  assign n14666 = pi0056 & n14665;
  assign n14667 = pi0863 & ~n14665;
  assign n14668 = ~n14666 & ~n14667;
  assign po0972 = pi1747 & ~n14668;
  assign n14670 = ~pi0870 & ~po1343;
  assign n14671 = ~pi0553 & n6302;
  assign n14672 = ~n14670 & ~n14671;
  assign n14673 = ~pi0315 & po1538;
  assign n14674 = ~pi0363 & n6305;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = ~pi0452 & n6299;
  assign n14677 = n14675 & ~n14676;
  assign po0979 = ~n14672 | ~n14677;
  assign n14679 = pi0871 & ~po1343;
  assign n14680 = ~pi0597 & n6302;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = ~pi0338 & po1538;
  assign n14683 = ~pi0415 & n6305;
  assign n14684 = ~n14682 & ~n14683;
  assign n14685 = ~pi0523 & n6299;
  assign n14686 = n14684 & ~n14685;
  assign po0980 = ~n14681 | ~n14686;
  assign n14688 = pi0765 & ~n13308;
  assign n14689 = pi0766 & ~n14688;
  assign n14690 = pi0766 & pi0790;
  assign n14691 = n14025 & n14690;
  assign n14692 = n13326 & ~n14691;
  assign po0981 = ~n14689 & n14692;
  assign n14694 = ~pi0873 & ~po1343;
  assign n14695 = pi1114 & n6302;
  assign n14696 = ~n14694 & ~n14695;
  assign n14697 = pi1024 & po1538;
  assign n14698 = ~pi1078 & n6305;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = pi1145 & n6299;
  assign n14701 = n14699 & ~n14700;
  assign po0982 = ~n14696 | ~n14701;
  assign n14703 = pi0876 & ~n14665;
  assign n14704 = pi0049 & n14665;
  assign n14705 = ~n14703 & ~n14704;
  assign po0985 = pi1747 & ~n14705;
  assign n14707 = pi0877 & ~po1343;
  assign n14708 = pi1102 & n6302;
  assign n14709 = ~n14707 & ~n14708;
  assign n14710 = pi1119 & po1538;
  assign n14711 = pi1127 & n6305;
  assign n14712 = ~n14710 & ~n14711;
  assign n14713 = pi1139 & n6299;
  assign n14714 = n14712 & ~n14713;
  assign po0986 = ~n14709 | ~n14714;
  assign n14716 = pi0878 & n4339;
  assign n14717 = ~pi0051 & ~n4339;
  assign n14718 = ~n14716 & ~n14717;
  assign po0987 = n4458 | ~n14718;
  assign n14720 = ~pi0879 & ~po1343;
  assign n14721 = ~pi0624 & n6302;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = ~pi0330 & po1538;
  assign n14724 = ~pi0375 & n6305;
  assign n14725 = ~n14723 & ~n14724;
  assign n14726 = ~pi0464 & n6299;
  assign n14727 = n14725 & ~n14726;
  assign po0988 = ~n14722 | ~n14727;
  assign n14729 = ~pi0880 & ~po1343;
  assign n14730 = ~pi0703 & n6302;
  assign n14731 = ~n14729 & ~n14730;
  assign n14732 = ~pi0360 & po1538;
  assign n14733 = ~pi0502 & n6305;
  assign n14734 = ~n14732 & ~n14733;
  assign n14735 = ~pi0537 & n6299;
  assign n14736 = n14734 & ~n14735;
  assign po0989 = ~n14731 | ~n14736;
  assign n14738 = ~pi0918 & ~n13259;
  assign n14739 = ~pi0881 & n13259;
  assign po0990 = n14738 | n14739;
  assign n14741 = pi1300 & ~pi1773;
  assign n14742 = pi1773 & pi1831;
  assign po0991 = n14741 | n14742;
  assign n14744 = ~pi0612 & n7999;
  assign n14745 = ~pi0487 & n8080;
  assign n14746 = ~n14744 & ~n14745;
  assign n14747 = ~pi1126 & n13676;
  assign n14748 = pi0617 & n13678;
  assign n14749 = ~n14747 & ~n14748;
  assign n14750 = n14746 & n14749;
  assign n14751 = n13672 & ~n14750;
  assign n14752 = ~pi0593 & n7999;
  assign n14753 = ~pi0670 & n8080;
  assign n14754 = ~n14752 & ~n14753;
  assign n14755 = ~pi1237 & n13676;
  assign n14756 = pi0535 & n13678;
  assign n14757 = ~n14755 & ~n14756;
  assign n14758 = n14754 & n14757;
  assign n14759 = n13700 & ~n14758;
  assign n14760 = ~pi0520 & n7999;
  assign n14761 = ~pi0570 & n8080;
  assign n14762 = ~n14760 & ~n14761;
  assign n14763 = ~pi1031 & n13676;
  assign n14764 = pi0592 & n13678;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = n14762 & n14765;
  assign n14767 = n13684 & ~n14766;
  assign n14768 = ~n14759 & ~n14767;
  assign n14769 = pi1038 & n13703;
  assign n14770 = pi1094 & n13705;
  assign n14771 = ~n14769 & ~n14770;
  assign n14772 = pi1291 & n13708;
  assign n14773 = pi1687 & n13710;
  assign n14774 = pi1503 & n13712;
  assign n14775 = ~n14773 & ~n14774;
  assign n14776 = pi0469 & n13715;
  assign n14777 = n14775 & ~n14776;
  assign n14778 = ~n14772 & n14777;
  assign n14779 = n14771 & n14778;
  assign n14780 = n13722 & ~n14779;
  assign n14781 = ~pi0337 & n7999;
  assign n14782 = ~pi0389 & n8080;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = ~pi1235 & n13676;
  assign n14785 = pi0615 & n13678;
  assign n14786 = ~n14784 & ~n14785;
  assign n14787 = n14783 & n14786;
  assign n14788 = n13724 & ~n14787;
  assign n14789 = n13733 & ~n14779;
  assign n14790 = ~n14788 & ~n14789;
  assign n14791 = ~n14780 & n14790;
  assign n14792 = n14768 & n14791;
  assign po0992 = n14751 | ~n14792;
  assign n14794 = ~pi0887 & ~n13259;
  assign n14795 = ~pi0884 & n13259;
  assign po0993 = n14794 | n14795;
  assign n14797 = ~pi0534 & n7999;
  assign n14798 = ~pi0499 & n8080;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = pi1027 & n13676;
  assign n14801 = pi0118 & n13678;
  assign n14802 = ~n14800 & ~n14801;
  assign n14803 = n14799 & n14802;
  assign n14804 = n13672 & ~n14803;
  assign n14805 = ~pi0626 & n7999;
  assign n14806 = ~pi0582 & n8080;
  assign n14807 = ~n14805 & ~n14806;
  assign n14808 = pi1032 & n13676;
  assign n14809 = pi0114 & n13678;
  assign n14810 = ~n14808 & ~n14809;
  assign n14811 = n14807 & n14810;
  assign n14812 = n13684 & ~n14811;
  assign n14813 = ~pi0607 & n7999;
  assign n14814 = ~pi0692 & n8080;
  assign n14815 = ~n14813 & ~n14814;
  assign n14816 = pi1105 & n13676;
  assign n14817 = pi0115 & n13678;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = n14815 & n14818;
  assign n14820 = n13700 & ~n14819;
  assign n14821 = ~n14812 & ~n14820;
  assign n14822 = pi1457 & n13703;
  assign n14823 = pi1096 & n13705;
  assign n14824 = ~n14822 & ~n14823;
  assign n14825 = pi1289 & n13708;
  assign n14826 = pi1682 & n13710;
  assign n14827 = pi1505 & n13712;
  assign n14828 = ~n14826 & ~n14827;
  assign n14829 = pi0433 & n13715;
  assign n14830 = n14828 & ~n14829;
  assign n14831 = ~n14825 & n14830;
  assign n14832 = n14824 & n14831;
  assign n14833 = n13722 & ~n14832;
  assign n14834 = ~pi0435 & n7999;
  assign n14835 = ~pi0402 & n8080;
  assign n14836 = ~n14834 & ~n14835;
  assign n14837 = pi1022 & n13676;
  assign n14838 = pi0116 & n13678;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = n14836 & n14839;
  assign n14841 = n13724 & ~n14840;
  assign n14842 = n13733 & ~n14832;
  assign n14843 = ~n14841 & ~n14842;
  assign n14844 = ~n14833 & n14843;
  assign n14845 = n14821 & n14844;
  assign po0994 = n14804 | ~n14845;
  assign n14847 = ~pi0425 & n7999;
  assign n14848 = ~pi0502 & n8080;
  assign n14849 = ~n14847 & ~n14848;
  assign n14850 = pi1310 & n13676;
  assign n14851 = pi0959 & n13678;
  assign n14852 = ~n14850 & ~n14851;
  assign n14853 = n14849 & n14852;
  assign n14854 = n13672 & ~n14853;
  assign n14855 = ~pi0531 & n7999;
  assign n14856 = ~pi0537 & n8080;
  assign n14857 = ~n14855 & ~n14856;
  assign n14858 = pi1342 & n13676;
  assign n14859 = pi0970 & n13678;
  assign n14860 = ~n14858 & ~n14859;
  assign n14861 = n14857 & n14860;
  assign n14862 = n13684 & ~n14861;
  assign n14863 = ~pi0609 & n7999;
  assign n14864 = ~pi0703 & n8080;
  assign n14865 = ~n14863 & ~n14864;
  assign n14866 = pi1338 & n13676;
  assign n14867 = pi0957 & n13678;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = n14865 & n14868;
  assign n14870 = n13700 & ~n14869;
  assign n14871 = ~n14862 & ~n14870;
  assign n14872 = pi0475 & n13715;
  assign n14873 = pi1069 & n13705;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = pi1320 & n13708;
  assign n14876 = pi1700 & n13710;
  assign n14877 = pi1504 & n13712;
  assign n14878 = ~n14876 & ~n14877;
  assign n14879 = pi1731 & n13703;
  assign n14880 = n14878 & ~n14879;
  assign n14881 = ~n14875 & n14880;
  assign n14882 = n14874 & n14881;
  assign n14883 = n13722 & ~n14882;
  assign n14884 = ~pi0348 & n7999;
  assign n14885 = ~pi0360 & n8080;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = pi1277 & n13676;
  assign n14888 = pi0958 & n13678;
  assign n14889 = ~n14887 & ~n14888;
  assign n14890 = n14886 & n14889;
  assign n14891 = n13724 & ~n14890;
  assign n14892 = n13733 & ~n14882;
  assign n14893 = ~n14891 & ~n14892;
  assign n14894 = ~n14883 & n14893;
  assign n14895 = n14871 & n14894;
  assign po0995 = n14854 | ~n14895;
  assign n14897 = ~pi1740 & ~n13259;
  assign n14898 = ~pi0887 & n13259;
  assign po0996 = n14897 | n14898;
  assign n14900 = pi1301 & ~pi1773;
  assign n14901 = pi1773 & pi1832;
  assign po0997 = n14900 | n14901;
  assign n14903 = ~pi1741 & ~n13259;
  assign n14904 = ~pi0889 & n13259;
  assign po0998 = n14903 | n14904;
  assign n14906 = ~pi1727 & ~n13259;
  assign n14907 = ~pi0890 & n13259;
  assign po0999 = n14906 | n14907;
  assign n14909 = pi0095 & n4173;
  assign n14910 = pi0012 & n14909;
  assign n14911 = pi1510 & n14910;
  assign n14912 = pi1447 & n14911;
  assign n14913 = ~pi0891 & ~n14912;
  assign po1000 = n6201 & ~n14913;
  assign n14915 = pi1480 & n14911;
  assign n14916 = ~pi0892 & ~n14915;
  assign po1001 = n6189 & ~n14916;
  assign n14918 = pi0795 & pi1479;
  assign n14919 = pi0860 & pi1479;
  assign n14920 = n14918 & n14919;
  assign n14921 = pi0799 & n14920;
  assign n14922 = pi0771 & n14921;
  assign n14923 = pi0803 & n14922;
  assign n14924 = ~n4122 & ~n14923;
  assign n14925 = pi0771 & pi0799;
  assign n14926 = n14918 & n14925;
  assign n14927 = ~pi0802 & n14919;
  assign n14928 = n14926 & ~n14927;
  assign n14929 = ~n4122 & ~n14928;
  assign n14930 = n14924 & ~n14929;
  assign n14931 = ~pi0771 & ~pi0802;
  assign n14932 = ~pi0799 & n14931;
  assign n14933 = pi0803 & n14919;
  assign n14934 = ~pi0800 & ~pi0802;
  assign n14935 = ~n14933 & n14934;
  assign n14936 = ~pi0771 & n14918;
  assign n14937 = n14935 & n14936;
  assign n14938 = ~n14932 & ~n14937;
  assign n14939 = ~pi0801 & ~pi0802;
  assign n14940 = ~pi0799 & n14939;
  assign n14941 = n14938 & ~n14940;
  assign n14942 = ~n14930 & ~n14941;
  assign n14943 = ~pi0803 & n14918;
  assign n14944 = n14919 & n14943;
  assign n14945 = n14925 & n14944;
  assign n14946 = ~n14924 & ~n14945;
  assign n14947 = n14924 & n14945;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = n14942 & n14948;
  assign n14950 = ~n14929 & n14946;
  assign n14951 = pi0802 & n4183;
  assign n14952 = n14950 & ~n14951;
  assign n14953 = ~n14949 & ~n14952;
  assign n14954 = pi1494 & n14950;
  assign n14955 = n8887 & n14945;
  assign n14956 = n14924 & n14955;
  assign n14957 = n8887 & ~n14945;
  assign n14958 = ~n14924 & n14957;
  assign n14959 = ~n14956 & ~n14958;
  assign n14960 = n14929 & ~n14959;
  assign n14961 = n14930 & n14957;
  assign n14962 = ~n14960 & ~n14961;
  assign n14963 = ~n14954 & n14962;
  assign po1003 = ~n14953 | ~n14963;
  assign n14965 = pi0549 & ~pi1083;
  assign n14966 = pi0567 & ~pi1130;
  assign n14967 = ~n14965 & ~n14966;
  assign n14968 = ~n7428 & n14967;
  assign n14969 = ~n6354 & n14968;
  assign n14970 = pi0622 & ~pi1129;
  assign n14971 = pi0587 & ~pi1028;
  assign n14972 = ~n14970 & ~n14971;
  assign n14973 = ~n7450 & n14972;
  assign n14974 = ~n6333 & n14973;
  assign n14975 = ~n10187 & ~n14974;
  assign n14976 = ~pi1129 & n6333;
  assign n14977 = pi0587 & n7450;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = ~n14975 & n14978;
  assign n14980 = ~n8790 & n14979;
  assign n14981 = pi1126 & n7421;
  assign n14982 = ~pi1127 & ~pi1130;
  assign n14983 = ~pi1083 & ~pi1310;
  assign n14984 = ~pi1027 & n14983;
  assign n14985 = ~pi1092 & n7450;
  assign n14986 = n14984 & n14985;
  assign n14987 = n14982 & n14986;
  assign n14988 = n14981 & n14987;
  assign n14989 = ~n14980 & ~n14988;
  assign n14990 = pi0483 & ~pi1076;
  assign n14991 = pi0485 & ~pi1029;
  assign n14992 = ~n14990 & ~n14991;
  assign n14993 = ~n7421 & n14992;
  assign n14994 = ~n6345 & n14993;
  assign n14995 = ~n8774 & ~n14994;
  assign n14996 = n14989 & n14995;
  assign n14997 = ~n14969 & n14996;
  assign n14998 = ~pi1083 & n6354;
  assign n14999 = pi0567 & n7428;
  assign n15000 = ~n14998 & ~n14999;
  assign n15001 = ~n8782 & n15000;
  assign n15002 = ~n14994 & ~n15001;
  assign n15003 = ~n8775 & ~n15002;
  assign n15004 = ~pi1076 & n6345;
  assign n15005 = pi0485 & n7421;
  assign n15006 = ~n15004 & ~n15005;
  assign n15007 = n15003 & n15006;
  assign n15008 = ~n8774 & ~n15007;
  assign n15009 = ~pi0468 & ~pi0562;
  assign n15010 = n11019 & n15009;
  assign n15011 = ~n15008 & n15010;
  assign n15012 = ~n14988 & ~n15011;
  assign po1005 = n14997 | n15012;
  assign n15014 = pi0480 & ~pi1121;
  assign n15015 = pi0484 & ~pi1274;
  assign n15016 = ~n15014 & ~n15015;
  assign n15017 = ~n7547 & n15016;
  assign n15018 = ~n6531 & n15017;
  assign n15019 = pi0509 & ~pi1023;
  assign n15020 = pi0508 & ~pi1272;
  assign n15021 = ~n15019 & ~n15020;
  assign n15022 = ~n7569 & n15021;
  assign n15023 = ~n6510 & n15022;
  assign n15024 = ~n9054 & ~n15023;
  assign n15025 = ~pi1023 & n6510;
  assign n15026 = pi0508 & n7569;
  assign n15027 = ~n15025 & ~n15026;
  assign n15028 = ~n15024 & n15027;
  assign n15029 = ~n8726 & n15028;
  assign n15030 = pi1235 & n7540;
  assign n15031 = ~pi1119 & ~pi1274;
  assign n15032 = ~pi1121 & ~pi1277;
  assign n15033 = ~pi1022 & n15032;
  assign n15034 = ~pi1280 & n7569;
  assign n15035 = n15033 & n15034;
  assign n15036 = n15031 & n15035;
  assign n15037 = n15030 & n15036;
  assign n15038 = ~n15029 & ~n15037;
  assign n15039 = pi0386 & ~pi1270;
  assign n15040 = pi0387 & ~pi1267;
  assign n15041 = ~n15039 & ~n15040;
  assign n15042 = ~n7540 & n15041;
  assign n15043 = ~n6522 & n15042;
  assign n15044 = ~n8707 & ~n15043;
  assign n15045 = n15038 & n15044;
  assign n15046 = ~n15018 & n15045;
  assign n15047 = ~pi1121 & n6531;
  assign n15048 = pi0484 & n7547;
  assign n15049 = ~n15047 & ~n15048;
  assign n15050 = ~n8715 & n15049;
  assign n15051 = ~n15043 & ~n15050;
  assign n15052 = ~n8708 & ~n15051;
  assign n15053 = ~pi1270 & n6522;
  assign n15054 = pi0387 & n7540;
  assign n15055 = ~n15053 & ~n15054;
  assign n15056 = n15052 & n15055;
  assign n15057 = ~n8707 & ~n15056;
  assign n15058 = ~pi0381 & ~pi0470;
  assign n15059 = n9915 & n15058;
  assign n15060 = ~n15057 & n15059;
  assign n15061 = ~n15037 & ~n15060;
  assign po1006 = n15046 | n15061;
  assign n15063 = pi0714 & ~pi1108;
  assign n15064 = pi0717 & ~pi1081;
  assign n15065 = ~n15063 & ~n15064;
  assign n15066 = ~n7661 & n15065;
  assign n15067 = ~n6815 & n15066;
  assign n15068 = pi0708 & ~pi1106;
  assign n15069 = pi0719 & ~pi1107;
  assign n15070 = ~n15068 & ~n15069;
  assign n15071 = ~n7683 & n15070;
  assign n15072 = ~n6794 & n15071;
  assign n15073 = ~n12236 & ~n15072;
  assign n15074 = ~pi1106 & n6794;
  assign n15075 = pi0719 & n7683;
  assign n15076 = ~n15074 & ~n15075;
  assign n15077 = ~n15073 & n15076;
  assign n15078 = ~n8508 & n15077;
  assign n15079 = pi1237 & n7654;
  assign n15080 = ~pi1081 & ~pi1102;
  assign n15081 = ~pi1108 & ~pi1338;
  assign n15082 = ~pi1105 & n15081;
  assign n15083 = ~pi1104 & n7683;
  assign n15084 = n15082 & n15083;
  assign n15085 = n15080 & n15084;
  assign n15086 = n15079 & n15085;
  assign n15087 = ~n15078 & ~n15086;
  assign n15088 = pi0675 & ~pi1109;
  assign n15089 = pi0678 & ~pi1110;
  assign n15090 = ~n15088 & ~n15089;
  assign n15091 = ~n7654 & n15090;
  assign n15092 = ~n6806 & n15091;
  assign n15093 = ~n8489 & ~n15092;
  assign n15094 = n15087 & n15093;
  assign n15095 = ~n15067 & n15094;
  assign n15096 = ~pi1108 & n6815;
  assign n15097 = pi0717 & n7661;
  assign n15098 = ~n15096 & ~n15097;
  assign n15099 = ~n8497 & n15098;
  assign n15100 = ~n15092 & ~n15099;
  assign n15101 = ~n8490 & ~n15100;
  assign n15102 = ~pi1109 & n6806;
  assign n15103 = pi0678 & n7654;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = n15101 & n15104;
  assign n15106 = ~n8489 & ~n15105;
  assign n15107 = ~pi0664 & ~pi0665;
  assign n15108 = n12230 & n15107;
  assign n15109 = ~n15106 & n15108;
  assign n15110 = ~n15086 & ~n15109;
  assign po1007 = n15095 | n15110;
  assign n15112 = pi0648 & ~pi1033;
  assign n15113 = pi0650 & ~pi1142;
  assign n15114 = ~n15112 & ~n15113;
  assign n15115 = ~n7604 & n15114;
  assign n15116 = ~n6453 & n15115;
  assign n15117 = pi0654 & ~pi1141;
  assign n15118 = pi0653 & ~pi1258;
  assign n15119 = ~n15117 & ~n15118;
  assign n15120 = ~n7626 & n15119;
  assign n15121 = ~n6432 & n15120;
  assign n15122 = ~n11192 & ~n15121;
  assign n15123 = ~pi1141 & n6432;
  assign n15124 = pi0653 & n7626;
  assign n15125 = ~n15123 & ~n15124;
  assign n15126 = ~n15122 & n15125;
  assign n15127 = ~n8439 & n15126;
  assign n15128 = pi1031 & n7597;
  assign n15129 = ~pi1139 & ~pi1142;
  assign n15130 = ~pi1033 & ~pi1342;
  assign n15131 = ~pi1032 & n15130;
  assign n15132 = ~pi1271 & n7626;
  assign n15133 = n15131 & n15132;
  assign n15134 = n15129 & n15133;
  assign n15135 = n15128 & n15134;
  assign n15136 = ~n15127 & ~n15135;
  assign n15137 = pi0566 & ~pi1265;
  assign n15138 = pi0569 & ~pi1034;
  assign n15139 = ~n15137 & ~n15138;
  assign n15140 = ~n7597 & n15139;
  assign n15141 = ~n6444 & n15140;
  assign n15142 = ~n8420 & ~n15141;
  assign n15143 = n15136 & n15142;
  assign n15144 = ~n15116 & n15143;
  assign n15145 = ~pi1033 & n6453;
  assign n15146 = pi0650 & n7604;
  assign n15147 = ~n15145 & ~n15146;
  assign n15148 = ~n8428 & n15147;
  assign n15149 = ~n15141 & ~n15148;
  assign n15150 = ~n8421 & ~n15149;
  assign n15151 = ~pi1265 & n6444;
  assign n15152 = pi0569 & n7597;
  assign n15153 = ~n15151 & ~n15152;
  assign n15154 = n15150 & n15153;
  assign n15155 = ~n8420 & ~n15154;
  assign n15156 = ~pi0621 & ~pi0645;
  assign n15157 = n11931 & n15156;
  assign n15158 = ~n15155 & n15157;
  assign n15159 = ~n15135 & ~n15158;
  assign po1008 = n15144 | n15159;
  assign n15161 = pi1479 & po1737;
  assign n15162 = pi0966 & n15161;
  assign n15163 = ~pi0995 & ~pi1045;
  assign n15164 = ~pi1050 & n15163;
  assign n15165 = ~pi0954 & n15164;
  assign n15166 = ~pi0773 & ~pi0984;
  assign n15167 = ~pi0937 & n15166;
  assign n15168 = ~pi1021 & n15167;
  assign n15169 = ~pi0966 & ~pi0971;
  assign n15170 = ~pi1019 & n15169;
  assign n15171 = ~pi1046 & n15170;
  assign n15172 = n15168 & n15171;
  assign n15173 = n15165 & n15172;
  assign n15174 = ~pi0916 & ~pi1677;
  assign n15175 = ~pi0966 & n15174;
  assign n15176 = pi0760 & n15175;
  assign n15177 = n15173 & n15176;
  assign n15178 = ~n15162 & ~n15177;
  assign n15179 = pi0262 & n15178;
  assign n15180 = ~pi0916 & n15179;
  assign n15181 = pi1019 & n15180;
  assign n15182 = pi0900 & n15178;
  assign n15183 = ~pi0760 & n15168;
  assign n15184 = ~pi0971 & n6711;
  assign n15185 = n15183 & n15184;
  assign n15186 = ~pi0966 & ~pi0995;
  assign n15187 = ~pi1019 & n15186;
  assign n15188 = pi0916 & pi1019;
  assign n15189 = ~pi0916 & ~pi1019;
  assign n15190 = ~n15188 & ~n15189;
  assign n15191 = pi1677 & n6699;
  assign n15192 = ~pi1045 & n15191;
  assign n15193 = ~n15190 & n15192;
  assign n15194 = n15187 & n15193;
  assign n15195 = n15185 & n15194;
  assign n15196 = n6711 & n15170;
  assign n15197 = pi0954 & ~pi1677;
  assign n15198 = n15183 & n15197;
  assign n15199 = ~pi0760 & ~pi0937;
  assign n15200 = n15166 & n15199;
  assign n15201 = pi1021 & n15200;
  assign n15202 = ~pi0954 & ~pi1677;
  assign n15203 = n15201 & n15202;
  assign n15204 = ~n15198 & ~n15203;
  assign n15205 = ~n15190 & ~n15204;
  assign n15206 = n15164 & n15205;
  assign n15207 = n15196 & n15206;
  assign n15208 = ~n15195 & ~n15207;
  assign n15209 = n15178 & ~n15208;
  assign n15210 = n6740 & ~n6743;
  assign n15211 = n15178 & n15210;
  assign n15212 = pi0916 & ~pi1019;
  assign n15213 = n15211 & n15212;
  assign n15214 = ~n15209 & ~n15213;
  assign n15215 = ~n15182 & n15214;
  assign po1009 = n15181 | ~n15215;
  assign n15217 = pi0901 & pi1747;
  assign n15218 = pi1424 & n15217;
  assign n15219 = ~pi1676 & n6325;
  assign n15220 = ~pi1726 & n15219;
  assign po1010 = n15218 | n15220;
  assign n15222 = pi1286 & ~pi1773;
  assign n15223 = pi1773 & pi1810;
  assign po1011 = n15222 | n15223;
  assign n15225 = pi1459 & n14911;
  assign n15226 = ~pi0903 & ~n15225;
  assign po1012 = n6185 & ~n15226;
  assign n15228 = pi1430 & n14911;
  assign n15229 = ~pi0904 & ~n15228;
  assign po1013 = n6193 & ~n15229;
  assign n15231 = pi1294 & ~pi1773;
  assign n15232 = pi1773 & pi1822;
  assign po1014 = n15231 | n15232;
  assign n15234 = pi1299 & ~pi1773;
  assign n15235 = pi1773 & pi1830;
  assign po1015 = n15234 | n15235;
  assign n15237 = pi1302 & ~pi1773;
  assign n15238 = pi1773 & pi1834;
  assign po1016 = n15237 | n15238;
  assign n15240 = pi1298 & ~pi1773;
  assign n15241 = pi1773 & pi1827;
  assign po1017 = n15240 | n15241;
  assign n15243 = pi1293 & ~pi1773;
  assign n15244 = pi1773 & pi1826;
  assign po1018 = n15243 | n15244;
  assign n15246 = pi1297 & ~pi1773;
  assign n15247 = pi1773 & pi1825;
  assign po1019 = n15246 | n15247;
  assign n15249 = pi1304 & ~pi1773;
  assign n15250 = pi1773 & pi1812;
  assign po1020 = n15249 | n15250;
  assign n15252 = pi1303 & ~pi1773;
  assign n15253 = pi1773 & pi1811;
  assign po1021 = n15252 | n15253;
  assign n15255 = pi1296 & ~pi1773;
  assign n15256 = pi1773 & pi1824;
  assign po1022 = n15255 | n15256;
  assign n15258 = pi1295 & ~pi1773;
  assign n15259 = pi1773 & pi1823;
  assign po1023 = n15258 | n15259;
  assign n15261 = pi0915 & pi1424;
  assign n15262 = pi1747 & n15261;
  assign n15263 = pi1424 & ~pi1675;
  assign n15264 = pi1747 & n15263;
  assign n15265 = ~pi1680 & n15264;
  assign po1024 = n15262 | n15265;
  assign n15267 = pi0916 & ~n6739;
  assign n15268 = n6735 & ~n6743;
  assign n15269 = ~n6738 & n15268;
  assign n15270 = n15267 & n15269;
  assign n15271 = ~pi0276 & ~pi0916;
  assign n15272 = n6705 & n6717;
  assign n15273 = ~pi0971 & n15272;
  assign n15274 = pi0995 & n15273;
  assign n15275 = ~n15271 & n15274;
  assign n15276 = ~pi0916 & ~n6753;
  assign n15277 = n13807 & ~n15276;
  assign n15278 = ~n15275 & ~n15277;
  assign n15279 = ~n15270 & n15278;
  assign n15280 = pi0183 & ~pi0916;
  assign n15281 = n13317 & ~n15280;
  assign n15282 = n15279 & ~n15281;
  assign n15283 = ~pi0760 & pi1021;
  assign n15284 = n13798 & n13804;
  assign n15285 = n15283 & n15284;
  assign n15286 = n15282 & ~n15285;
  assign po1025 = ~po1785 & ~n15286;
  assign n15288 = ~pi0917 & ~po1526;
  assign n15289 = n13259 & ~n15288;
  assign po1026 = pi1747 & ~n15289;
  assign n15291 = ~pi1733 & ~n13259;
  assign n15292 = ~pi0918 & n13259;
  assign po1027 = n15291 | n15292;
  assign n15294 = n13802 & ~n13814;
  assign n15295 = ~pi1670 & n13795;
  assign n15296 = n15294 & n15295;
  assign n15297 = ~n13802 & n13814;
  assign n15298 = ~pi1670 & n13321;
  assign n15299 = n15297 & n15298;
  assign n15300 = ~n15296 & ~n15299;
  assign n15301 = ~pi0919 & n15300;
  assign n15302 = pi0919 & ~pi0963;
  assign n15303 = ~pi0919 & pi0963;
  assign n15304 = ~n15302 & ~n15303;
  assign n15305 = ~n15300 & ~n15304;
  assign n15306 = ~n15301 & ~n15305;
  assign po1028 = ~pi0984 & ~n15306;
  assign n15308 = ~pi1722 & ~n13259;
  assign n15309 = ~pi0920 & n13259;
  assign po1029 = n15308 | n15309;
  assign n15311 = ~pi0921 & n15300;
  assign n15312 = ~pi0919 & ~pi0963;
  assign n15313 = ~pi0921 & ~n15312;
  assign n15314 = pi0921 & n15312;
  assign n15315 = ~n15313 & ~n15314;
  assign n15316 = ~n15300 & ~n15315;
  assign n15317 = ~n15311 & ~n15316;
  assign po1030 = ~pi0984 & ~n15317;
  assign n15319 = ~pi1735 & ~n13259;
  assign n15320 = ~pi0922 & n13259;
  assign po1031 = n15319 | n15320;
  assign n15322 = ~pi1738 & ~n13259;
  assign n15323 = ~pi0923 & n13259;
  assign po1032 = n15322 | n15323;
  assign n15325 = ~pi1725 & ~n13259;
  assign n15326 = ~pi0924 & n13259;
  assign po1033 = n15325 | n15326;
  assign n15328 = ~pi0889 & ~n13259;
  assign n15329 = ~pi0925 & n13259;
  assign po1034 = n15328 | n15329;
  assign n15331 = ~pi0920 & ~n13259;
  assign n15332 = ~pi0926 & n13259;
  assign po1035 = n15331 | n15332;
  assign n15334 = ~pi0890 & ~n13259;
  assign n15335 = ~pi0927 & n13259;
  assign po1036 = n15334 | n15335;
  assign n15337 = ~pi0922 & ~n13259;
  assign n15338 = ~pi0928 & n13259;
  assign po1037 = n15337 | n15338;
  assign n15340 = ~pi0923 & ~n13259;
  assign n15341 = ~pi0929 & n13259;
  assign po1038 = n15340 | n15341;
  assign n15343 = ~pi0924 & ~n13259;
  assign n15344 = ~pi0930 & n13259;
  assign po1039 = n15343 | n15344;
  assign n15346 = ~pi0925 & ~n13259;
  assign n15347 = ~pi0931 & n13259;
  assign po1040 = n15346 | n15347;
  assign n15349 = ~pi0926 & ~n13259;
  assign n15350 = ~pi0932 & n13259;
  assign po1041 = n15349 | n15350;
  assign n15352 = ~pi0927 & ~n13259;
  assign n15353 = ~pi0933 & n13259;
  assign po1042 = n15352 | n15353;
  assign n15355 = ~pi0928 & ~n13259;
  assign n15356 = ~pi0934 & n13259;
  assign po1043 = n15355 | n15356;
  assign n15358 = ~pi0929 & ~n13259;
  assign n15359 = ~pi0935 & n13259;
  assign po1044 = n15358 | n15359;
  assign n15361 = ~pi0930 & ~n13259;
  assign n15362 = ~pi0936 & n13259;
  assign po1045 = n15361 | n15362;
  assign n15364 = pi0937 & ~n6753;
  assign n15365 = n13814 & n15364;
  assign n15366 = ~pi1670 & ~n13321;
  assign n15367 = n15365 & n15366;
  assign n15368 = ~n6753 & n13795;
  assign n15369 = ~n15364 & ~n15368;
  assign n15370 = n13802 & ~n15369;
  assign n15371 = ~pi1670 & n15370;
  assign n15372 = ~n15367 & ~n15371;
  assign po1046 = ~po1785 & ~n15372;
  assign n15374 = pi1447 & pi1698;
  assign n15375 = pi0064 & n15374;
  assign n15376 = pi0938 & ~n15374;
  assign n15377 = ~n15375 & ~n15376;
  assign po1047 = pi1747 & ~n15377;
  assign n15379 = pi1447 & pi1695;
  assign n15380 = pi0056 & n15379;
  assign n15381 = pi0939 & ~n15379;
  assign n15382 = ~n15380 & ~n15381;
  assign po1048 = pi1747 & ~n15382;
  assign n15384 = pi0941 & ~n15374;
  assign n15385 = pi0057 & n15374;
  assign n15386 = ~n15384 & ~n15385;
  assign po1050 = pi1747 & ~n15386;
  assign n15388 = pi0942 & ~n15379;
  assign n15389 = pi0049 & n15379;
  assign n15390 = ~n15388 & ~n15389;
  assign po1051 = pi1747 & ~n15390;
  assign n15392 = ~pi0881 & ~n13259;
  assign n15393 = ~pi0943 & n13259;
  assign po1052 = n15392 | n15393;
  assign n15395 = ~pi0884 & ~n13259;
  assign n15396 = ~pi0944 & n13259;
  assign po1053 = n15395 | n15396;
  assign n15398 = ~pi0715 & pi1269;
  assign n15399 = pi0715 & ~pi1269;
  assign n15400 = ~n15398 & ~n15399;
  assign n15401 = pi0720 & ~pi1158;
  assign n15402 = pi0707 & ~pi1157;
  assign n15403 = ~pi0669 & pi1155;
  assign n15404 = pi0669 & ~pi1155;
  assign n15405 = ~pi0699 & pi1154;
  assign n15406 = ~n15404 & n15405;
  assign n15407 = ~n15403 & ~n15406;
  assign n15408 = ~pi0698 & pi1283;
  assign n15409 = pi0700 & ~pi1331;
  assign n15410 = pi0698 & ~pi1283;
  assign n15411 = ~n15409 & ~n15410;
  assign n15412 = ~n15408 & ~n15411;
  assign n15413 = pi0699 & ~pi1154;
  assign n15414 = ~n15404 & ~n15413;
  assign n15415 = ~n15412 & n15414;
  assign n15416 = n15407 & ~n15415;
  assign n15417 = pi0710 & ~pi1156;
  assign n15418 = ~n15416 & ~n15417;
  assign n15419 = ~n15402 & n15418;
  assign n15420 = ~pi0707 & pi1157;
  assign n15421 = ~pi0710 & pi1156;
  assign n15422 = ~n15402 & n15421;
  assign n15423 = ~n15420 & ~n15422;
  assign n15424 = ~n15419 & n15423;
  assign n15425 = pi0679 & ~pi1275;
  assign n15426 = ~n15424 & ~n15425;
  assign n15427 = ~n15401 & n15426;
  assign n15428 = pi0709 & ~pi1346;
  assign n15429 = pi0663 & ~pi1159;
  assign n15430 = ~n15428 & ~n15429;
  assign n15431 = n15427 & n15430;
  assign n15432 = ~pi0709 & pi1346;
  assign n15433 = ~pi0720 & pi1158;
  assign n15434 = ~pi0679 & pi1275;
  assign n15435 = ~n15401 & n15434;
  assign n15436 = ~n15433 & ~n15435;
  assign n15437 = ~n15428 & ~n15436;
  assign n15438 = ~n15432 & ~n15437;
  assign n15439 = ~n15429 & ~n15438;
  assign n15440 = ~n15431 & ~n15439;
  assign n15441 = ~pi0663 & pi1159;
  assign n15442 = n15440 & ~n15441;
  assign n15443 = n15400 & n15442;
  assign n15444 = ~n15400 & ~n15442;
  assign po1056 = n15443 | n15444;
  assign n15446 = ~pi0481 & pi1177;
  assign n15447 = pi0481 & ~pi1177;
  assign n15448 = ~n15446 & ~n15447;
  assign n15449 = pi0482 & ~pi1089;
  assign n15450 = pi0510 & ~pi1093;
  assign n15451 = ~pi0413 & pi1087;
  assign n15452 = pi0413 & ~pi1087;
  assign n15453 = ~pi0412 & pi1173;
  assign n15454 = ~n15452 & n15453;
  assign n15455 = ~n15451 & ~n15454;
  assign n15456 = ~pi0411 & pi1077;
  assign n15457 = pi0410 & ~pi1241;
  assign n15458 = pi0411 & ~pi1077;
  assign n15459 = ~n15457 & ~n15458;
  assign n15460 = ~n15456 & ~n15459;
  assign n15461 = pi0412 & ~pi1173;
  assign n15462 = ~n15452 & ~n15461;
  assign n15463 = ~n15460 & n15462;
  assign n15464 = n15455 & ~n15463;
  assign n15465 = pi0442 & ~pi1174;
  assign n15466 = ~n15464 & ~n15465;
  assign n15467 = ~n15450 & n15466;
  assign n15468 = ~pi0510 & pi1093;
  assign n15469 = ~pi0442 & pi1174;
  assign n15470 = ~n15450 & n15469;
  assign n15471 = ~n15468 & ~n15470;
  assign n15472 = ~n15467 & n15471;
  assign n15473 = pi0388 & ~pi1175;
  assign n15474 = ~n15472 & ~n15473;
  assign n15475 = ~n15449 & n15474;
  assign n15476 = pi0441 & ~pi1176;
  assign n15477 = pi0384 & ~pi1082;
  assign n15478 = ~n15476 & ~n15477;
  assign n15479 = n15475 & n15478;
  assign n15480 = ~pi0441 & pi1176;
  assign n15481 = ~pi0482 & pi1089;
  assign n15482 = ~pi0388 & pi1175;
  assign n15483 = ~n15449 & n15482;
  assign n15484 = ~n15481 & ~n15483;
  assign n15485 = ~n15476 & ~n15484;
  assign n15486 = ~n15480 & ~n15485;
  assign n15487 = ~n15477 & ~n15486;
  assign n15488 = ~n15479 & ~n15487;
  assign n15489 = ~pi0384 & pi1082;
  assign n15490 = n15488 & ~n15489;
  assign n15491 = n15448 & n15490;
  assign n15492 = ~n15448 & ~n15490;
  assign po1057 = n15491 | n15492;
  assign n15494 = ~pi0564 & pi1201;
  assign n15495 = pi0564 & ~pi1201;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = pi0565 & ~pi1198;
  assign n15498 = pi0588 & ~pi1264;
  assign n15499 = ~pi0514 & pi1195;
  assign n15500 = pi0514 & ~pi1195;
  assign n15501 = ~pi0513 & pi1194;
  assign n15502 = ~n15500 & n15501;
  assign n15503 = ~n15499 & ~n15502;
  assign n15504 = ~pi0512 & pi1276;
  assign n15505 = pi0511 & ~pi1192;
  assign n15506 = pi0512 & ~pi1276;
  assign n15507 = ~n15505 & ~n15506;
  assign n15508 = ~n15504 & ~n15507;
  assign n15509 = pi0513 & ~pi1194;
  assign n15510 = ~n15500 & ~n15509;
  assign n15511 = ~n15508 & n15510;
  assign n15512 = n15503 & ~n15511;
  assign n15513 = pi0541 & ~pi1196;
  assign n15514 = ~n15512 & ~n15513;
  assign n15515 = ~n15498 & n15514;
  assign n15516 = ~pi0588 & pi1264;
  assign n15517 = ~pi0541 & pi1196;
  assign n15518 = ~n15498 & n15517;
  assign n15519 = ~n15516 & ~n15518;
  assign n15520 = ~n15515 & n15519;
  assign n15521 = pi0486 & ~pi1197;
  assign n15522 = ~n15520 & ~n15521;
  assign n15523 = ~n15497 & n15522;
  assign n15524 = pi0560 & ~pi1199;
  assign n15525 = pi0472 & ~pi1249;
  assign n15526 = ~n15524 & ~n15525;
  assign n15527 = n15523 & n15526;
  assign n15528 = ~pi0560 & pi1199;
  assign n15529 = ~pi0565 & pi1198;
  assign n15530 = ~pi0486 & pi1197;
  assign n15531 = ~n15497 & n15530;
  assign n15532 = ~n15529 & ~n15531;
  assign n15533 = ~n15524 & ~n15532;
  assign n15534 = ~n15528 & ~n15533;
  assign n15535 = ~n15525 & ~n15534;
  assign n15536 = ~n15527 & ~n15535;
  assign n15537 = ~pi0472 & pi1249;
  assign n15538 = n15536 & ~n15537;
  assign n15539 = n15496 & n15538;
  assign n15540 = ~n15496 & ~n15538;
  assign po1058 = n15539 | n15540;
  assign n15542 = ~pi0649 & pi1232;
  assign n15543 = pi0649 & ~pi1232;
  assign n15544 = ~n15542 & ~n15543;
  assign n15545 = pi0631 & ~pi1219;
  assign n15546 = pi0655 & ~pi1217;
  assign n15547 = ~pi0591 & pi1216;
  assign n15548 = pi0591 & ~pi1216;
  assign n15549 = ~pi0590 & pi1215;
  assign n15550 = ~n15548 & n15549;
  assign n15551 = ~n15547 & ~n15550;
  assign n15552 = ~pi0589 & pi1214;
  assign n15553 = pi0594 & ~pi1213;
  assign n15554 = pi0589 & ~pi1214;
  assign n15555 = ~n15553 & ~n15554;
  assign n15556 = ~n15552 & ~n15555;
  assign n15557 = pi0590 & ~pi1215;
  assign n15558 = ~n15548 & ~n15557;
  assign n15559 = ~n15556 & n15558;
  assign n15560 = n15551 & ~n15559;
  assign n15561 = pi0627 & ~pi1066;
  assign n15562 = ~n15560 & ~n15561;
  assign n15563 = ~n15546 & n15562;
  assign n15564 = ~pi0655 & pi1217;
  assign n15565 = ~pi0627 & pi1066;
  assign n15566 = ~n15546 & n15565;
  assign n15567 = ~n15564 & ~n15566;
  assign n15568 = ~n15563 & n15567;
  assign n15569 = pi0568 & ~pi1218;
  assign n15570 = ~n15568 & ~n15569;
  assign n15571 = ~n15545 & n15570;
  assign n15572 = pi0642 & ~pi1056;
  assign n15573 = pi0552 & ~pi1057;
  assign n15574 = ~n15572 & ~n15573;
  assign n15575 = n15571 & n15574;
  assign n15576 = ~pi0642 & pi1056;
  assign n15577 = ~pi0631 & pi1219;
  assign n15578 = ~pi0568 & pi1218;
  assign n15579 = ~n15545 & n15578;
  assign n15580 = ~n15577 & ~n15579;
  assign n15581 = ~n15572 & ~n15580;
  assign n15582 = ~n15576 & ~n15581;
  assign n15583 = ~n15573 & ~n15582;
  assign n15584 = ~n15575 & ~n15583;
  assign n15585 = ~pi0552 & pi1057;
  assign n15586 = n15584 & ~n15585;
  assign n15587 = n15544 & n15586;
  assign n15588 = ~n15544 & ~n15586;
  assign po1059 = n15587 | n15588;
  assign n15590 = pi1366 & ~pi1773;
  assign n15591 = pi1773 & pi1836;
  assign po1060 = n15590 | n15591;
  assign n15593 = pi1367 & ~pi1773;
  assign n15594 = pi1773 & pi1837;
  assign po1061 = n15593 | n15594;
  assign n15596 = ~pi1099 & pi1358;
  assign n15597 = pi0257 & pi1099;
  assign po1062 = n15596 | n15597;
  assign n15599 = ~pi0872 & ~pi1683;
  assign n15600 = ~n13795 & ~n15599;
  assign n15601 = pi0954 & n15600;
  assign n15602 = ~n6754 & ~n15601;
  assign n15603 = n6720 & ~n15602;
  assign n15604 = ~n6738 & ~n6739;
  assign n15605 = pi0954 & n15604;
  assign n15606 = ~n6743 & ~n15605;
  assign n15607 = n6735 & ~n15606;
  assign n15608 = pi0954 & ~n13322;
  assign n15609 = ~n6759 & ~n15608;
  assign n15610 = n6709 & ~n15609;
  assign n15611 = ~n15607 & ~n15610;
  assign n15612 = ~pi0277 & pi0954;
  assign n15613 = n6716 & n15612;
  assign n15614 = n15611 & ~n15613;
  assign n15615 = ~n15603 & n15614;
  assign po1063 = ~po1785 & ~n15615;
  assign n15617 = pi1368 & ~pi1773;
  assign n15618 = pi1773 & pi1833;
  assign po1064 = n15617 | n15618;
  assign n15620 = pi1365 & ~pi1773;
  assign n15621 = pi1773 & pi1835;
  assign po1065 = n15620 | n15621;
  assign n15623 = pi0012 & pi0095;
  assign n15624 = ~pi1511 & n15623;
  assign n15625 = ~n4173 & n15624;
  assign n15626 = pi1480 & n15625;
  assign n15627 = ~pi0957 & ~n15626;
  assign po1066 = n6189 & ~n15627;
  assign n15629 = pi1430 & n15625;
  assign n15630 = ~pi0958 & ~n15629;
  assign po1067 = n6193 & ~n15630;
  assign n15632 = pi1447 & n15625;
  assign n15633 = ~pi0959 & ~n15632;
  assign po1068 = n6201 & ~n15633;
  assign po1069 = n13326 & n14021;
  assign n15636 = pi1372 & ~pi1773;
  assign n15637 = pi1773 & pi1817;
  assign po1070 = n15636 | n15637;
  assign n15639 = pi1373 & ~pi1773;
  assign n15640 = pi1773 & pi1815;
  assign po1071 = n15639 | n15640;
  assign n15642 = ~pi0963 & ~n15300;
  assign n15643 = pi0963 & n15300;
  assign n15644 = ~n15642 & ~n15643;
  assign po1072 = ~pi0984 & n15644;
  assign n15646 = pi1392 & ~pi1773;
  assign n15647 = pi1773 & pi1818;
  assign po1073 = n15646 | n15647;
  assign n15649 = ~pi0965 & ~n8082;
  assign po1074 = n6193 & ~n15649;
  assign n15651 = pi0966 & ~po1737;
  assign n15652 = n6730 & n15651;
  assign n15653 = ~pi0277 & ~pi0966;
  assign n15654 = ~pi0984 & n6699;
  assign n15655 = n6706 & n15654;
  assign n15656 = pi1045 & n15655;
  assign n15657 = n6713 & n15656;
  assign n15658 = ~n15653 & n15657;
  assign n15659 = ~n15652 & ~n15658;
  assign n15660 = pi0966 & ~n15599;
  assign n15661 = ~n13795 & ~n15660;
  assign n15662 = n6720 & ~n15661;
  assign n15663 = ~n6754 & n15662;
  assign n15664 = n15659 & ~n15663;
  assign po1075 = ~po1785 & ~n15664;
  assign n15666 = pi1459 & pi1698;
  assign n15667 = pi0064 & n15666;
  assign n15668 = pi0967 & ~n15666;
  assign n15669 = ~n15667 & ~n15668;
  assign po1076 = pi1747 & ~n15669;
  assign n15671 = pi0968 & ~n15666;
  assign n15672 = pi0057 & n15666;
  assign n15673 = ~n15671 & ~n15672;
  assign po1077 = pi1747 & ~n15673;
  assign n15675 = pi1459 & pi1695;
  assign n15676 = pi0056 & n15675;
  assign n15677 = pi0969 & ~n15675;
  assign n15678 = ~n15676 & ~n15677;
  assign po1078 = pi1747 & ~n15678;
  assign n15680 = pi1459 & n15625;
  assign n15681 = ~pi0970 & ~n15680;
  assign po1079 = n6185 & ~n15681;
  assign n15683 = pi0971 & ~n6759;
  assign n15684 = ~n13323 & ~n15683;
  assign n15685 = n6709 & ~n15684;
  assign n15686 = pi0971 & ~n6738;
  assign n15687 = ~n6739 & ~n15686;
  assign n15688 = n6735 & ~n15687;
  assign n15689 = ~n6743 & n15688;
  assign n15690 = ~n15685 & ~n15689;
  assign n15691 = n6720 & ~n13795;
  assign n15692 = ~n15599 & n15691;
  assign n15693 = pi0971 & n15692;
  assign n15694 = ~n6754 & n15693;
  assign n15695 = n15690 & ~n15694;
  assign po1080 = ~po1785 & ~n15695;
  assign n15697 = pi1371 & ~pi1773;
  assign n15698 = pi1773 & pi1816;
  assign po1081 = n15697 | n15698;
  assign n15700 = pi0973 & ~n15675;
  assign n15701 = pi0049 & n15675;
  assign n15702 = ~n15700 & ~n15701;
  assign po1082 = pi1747 & ~n15702;
  assign po1083 = ~pi0789 & ~n13259;
  assign n15705 = pi0954 & ~pi1021;
  assign n15706 = n15200 & n15705;
  assign n15707 = ~pi0937 & n13805;
  assign n15708 = ~pi0954 & ~pi0984;
  assign n15709 = ~pi0773 & n15708;
  assign n15710 = n15707 & n15709;
  assign n15711 = ~n15706 & ~n15710;
  assign n15712 = n15196 & ~n15711;
  assign n15713 = ~pi1677 & n15712;
  assign n15714 = n15164 & n15713;
  assign n15715 = pi0975 & ~n15714;
  assign n15716 = ~n15162 & n15715;
  assign n15717 = ~pi0916 & ~pi0971;
  assign n15718 = ~pi0984 & ~pi1050;
  assign n15719 = ~pi1045 & n15718;
  assign n15720 = ~pi0954 & n15719;
  assign n15721 = ~pi0773 & n15199;
  assign n15722 = ~pi1021 & n15721;
  assign n15723 = n15720 & n15722;
  assign n15724 = n15187 & n15723;
  assign n15725 = n6764 & n15724;
  assign n15726 = n15717 & n15725;
  assign n15727 = pi0966 & ~n15162;
  assign n15728 = pi0975 & n15727;
  assign n15729 = ~n15726 & ~n15728;
  assign n15730 = ~n15716 & n15729;
  assign n15731 = pi0916 & n15210;
  assign n15732 = n15730 & ~n15731;
  assign n15733 = n15171 & n15200;
  assign n15734 = n15165 & n15733;
  assign n15735 = pi1021 & n15174;
  assign n15736 = ~pi0916 & n15735;
  assign n15737 = n15734 & n15736;
  assign po1084 = ~n15732 | n15737;
  assign n15739 = ~n13805 & ~n15283;
  assign n15740 = ~pi0937 & n15164;
  assign n15741 = ~pi0954 & n15740;
  assign n15742 = n15166 & n15741;
  assign n15743 = ~n15739 & n15742;
  assign n15744 = ~pi1046 & n15169;
  assign n15745 = ~pi1019 & n15744;
  assign n15746 = n15174 & n15745;
  assign n15747 = n15743 & n15746;
  assign n15748 = ~pi0966 & n15747;
  assign n15749 = pi0966 & po1737;
  assign n15750 = ~n15748 & ~n15749;
  assign n15751 = pi0976 & n15750;
  assign n15752 = ~pi0995 & n15722;
  assign n15753 = n15174 & n15752;
  assign n15754 = n15171 & n15753;
  assign n15755 = n15719 & n15754;
  assign n15756 = pi0954 & ~pi1019;
  assign n15757 = n15755 & n15756;
  assign n15758 = pi0262 & pi1019;
  assign n15759 = ~n15757 & ~n15758;
  assign po1085 = n15751 | ~n15759;
  assign n15761 = ~pi0977 & pi1543;
  assign po1086 = n6325 & ~n15761;
  assign n15763 = ~n15428 & n15433;
  assign n15764 = ~n15432 & ~n15763;
  assign n15765 = n15420 & ~n15425;
  assign n15766 = ~n15434 & ~n15765;
  assign n15767 = n15403 & ~n15417;
  assign n15768 = ~n15421 & ~n15767;
  assign n15769 = n15408 & ~n15413;
  assign n15770 = ~n15405 & ~n15769;
  assign n15771 = ~n15404 & ~n15417;
  assign n15772 = ~n15770 & n15771;
  assign n15773 = n15768 & ~n15772;
  assign n15774 = ~n15402 & ~n15425;
  assign n15775 = ~n15773 & n15774;
  assign n15776 = n15766 & ~n15775;
  assign n15777 = ~n15401 & ~n15428;
  assign n15778 = ~n15776 & n15777;
  assign n15779 = n15764 & ~n15778;
  assign n15780 = n15441 & ~n15779;
  assign n15781 = ~n15429 & ~n15441;
  assign n15782 = n15774 & n15777;
  assign n15783 = ~n15409 & ~n15413;
  assign n15784 = n15771 & n15783;
  assign n15785 = ~n15410 & n15784;
  assign n15786 = n15782 & n15785;
  assign n15787 = ~n15781 & n15786;
  assign n15788 = ~n15780 & ~n15787;
  assign n15789 = n15779 & n15781;
  assign n15790 = ~n15786 & n15789;
  assign n15791 = n15429 & ~n15779;
  assign n15792 = ~n15790 & ~n15791;
  assign po1087 = ~n15788 | ~n15792;
  assign n15794 = ~n15476 & n15481;
  assign n15795 = ~n15480 & ~n15794;
  assign n15796 = n15468 & ~n15473;
  assign n15797 = ~n15482 & ~n15796;
  assign n15798 = n15451 & ~n15465;
  assign n15799 = ~n15469 & ~n15798;
  assign n15800 = n15456 & ~n15461;
  assign n15801 = ~n15453 & ~n15800;
  assign n15802 = ~n15452 & ~n15465;
  assign n15803 = ~n15801 & n15802;
  assign n15804 = n15799 & ~n15803;
  assign n15805 = ~n15450 & ~n15473;
  assign n15806 = ~n15804 & n15805;
  assign n15807 = n15797 & ~n15806;
  assign n15808 = ~n15449 & ~n15476;
  assign n15809 = ~n15807 & n15808;
  assign n15810 = n15795 & ~n15809;
  assign n15811 = n15477 & ~n15810;
  assign n15812 = ~n15477 & ~n15489;
  assign n15813 = n15805 & n15808;
  assign n15814 = ~n15457 & ~n15461;
  assign n15815 = n15802 & n15814;
  assign n15816 = ~n15458 & n15815;
  assign n15817 = n15813 & n15816;
  assign n15818 = ~n15812 & n15817;
  assign n15819 = ~n15811 & ~n15818;
  assign n15820 = n15810 & n15812;
  assign n15821 = ~n15817 & n15820;
  assign n15822 = n15489 & ~n15810;
  assign n15823 = ~n15821 & ~n15822;
  assign po1088 = ~n15819 | ~n15823;
  assign n15825 = ~n15524 & n15529;
  assign n15826 = ~n15528 & ~n15825;
  assign n15827 = n15516 & ~n15521;
  assign n15828 = ~n15530 & ~n15827;
  assign n15829 = n15499 & ~n15513;
  assign n15830 = ~n15517 & ~n15829;
  assign n15831 = n15504 & ~n15509;
  assign n15832 = ~n15501 & ~n15831;
  assign n15833 = ~n15500 & ~n15513;
  assign n15834 = ~n15832 & n15833;
  assign n15835 = n15830 & ~n15834;
  assign n15836 = ~n15498 & ~n15521;
  assign n15837 = ~n15835 & n15836;
  assign n15838 = n15828 & ~n15837;
  assign n15839 = ~n15497 & ~n15524;
  assign n15840 = ~n15838 & n15839;
  assign n15841 = n15826 & ~n15840;
  assign n15842 = n15537 & ~n15841;
  assign n15843 = ~n15525 & ~n15537;
  assign n15844 = n15836 & n15839;
  assign n15845 = ~n15505 & ~n15509;
  assign n15846 = n15833 & n15845;
  assign n15847 = ~n15506 & n15846;
  assign n15848 = n15844 & n15847;
  assign n15849 = ~n15843 & n15848;
  assign n15850 = ~n15842 & ~n15849;
  assign n15851 = n15841 & n15843;
  assign n15852 = ~n15848 & n15851;
  assign n15853 = n15525 & ~n15841;
  assign n15854 = ~n15852 & ~n15853;
  assign po1089 = ~n15850 | ~n15854;
  assign n15856 = ~n15572 & n15577;
  assign n15857 = ~n15576 & ~n15856;
  assign n15858 = n15564 & ~n15569;
  assign n15859 = ~n15578 & ~n15858;
  assign n15860 = n15547 & ~n15561;
  assign n15861 = ~n15565 & ~n15860;
  assign n15862 = n15552 & ~n15557;
  assign n15863 = ~n15549 & ~n15862;
  assign n15864 = ~n15548 & ~n15561;
  assign n15865 = ~n15863 & n15864;
  assign n15866 = n15861 & ~n15865;
  assign n15867 = ~n15546 & ~n15569;
  assign n15868 = ~n15866 & n15867;
  assign n15869 = n15859 & ~n15868;
  assign n15870 = ~n15545 & ~n15572;
  assign n15871 = ~n15869 & n15870;
  assign n15872 = n15857 & ~n15871;
  assign n15873 = n15573 & ~n15872;
  assign n15874 = ~n15573 & ~n15585;
  assign n15875 = n15867 & n15870;
  assign n15876 = ~n15553 & ~n15557;
  assign n15877 = n15864 & n15876;
  assign n15878 = ~n15554 & n15877;
  assign n15879 = n15875 & n15878;
  assign n15880 = ~n15874 & n15879;
  assign n15881 = ~n15873 & ~n15880;
  assign n15882 = n15872 & n15874;
  assign n15883 = ~n15879 & n15882;
  assign n15884 = n15585 & ~n15872;
  assign n15885 = ~n15883 & ~n15884;
  assign po1090 = ~n15881 | ~n15885;
  assign n15887 = ~n14919 & n14925;
  assign n15888 = ~n14918 & n15887;
  assign n15889 = n4122 & ~n15888;
  assign n15890 = ~n4122 & n15888;
  assign n15891 = ~n15889 & ~n15890;
  assign n15892 = pi0799 & n14918;
  assign n15893 = n14934 & n15892;
  assign n15894 = ~n14919 & n15893;
  assign n15895 = ~pi0800 & n14944;
  assign n15896 = pi0799 & ~n15895;
  assign n15897 = pi0802 & ~n15896;
  assign n15898 = ~n15894 & ~n15897;
  assign n15899 = n15891 & ~n15898;
  assign n15900 = ~pi0771 & n15899;
  assign n15901 = ~pi0800 & ~pi0803;
  assign n15902 = n15892 & n15901;
  assign n15903 = n6070 & ~n14919;
  assign n15904 = ~n15902 & ~n15903;
  assign n15905 = ~pi0801 & ~n15904;
  assign n15906 = ~pi0801 & pi0802;
  assign n15907 = ~pi0799 & n15906;
  assign n15908 = ~n15905 & ~n15907;
  assign n15909 = n15891 & ~n15908;
  assign n15910 = ~n15900 & ~n15909;
  assign n15911 = ~pi1494 & n15889;
  assign n15912 = pi0803 & ~n4183;
  assign n15913 = ~n14951 & ~n15912;
  assign n15914 = n15911 & ~n15913;
  assign n15915 = ~n8883 & n15890;
  assign n15916 = ~n8882 & n15915;
  assign n15917 = ~n15914 & ~n15916;
  assign po1091 = ~n15910 | ~n15917;
  assign n15919 = ~n14930 & n14948;
  assign n15920 = ~pi0771 & pi0802;
  assign n15921 = ~pi0800 & n15920;
  assign n15922 = n15919 & n15921;
  assign n15923 = pi0799 & n15922;
  assign n15924 = n14944 & n15923;
  assign n15925 = n14950 & ~n15912;
  assign n15926 = n14930 & n14955;
  assign n15927 = ~n15925 & ~n15926;
  assign n15928 = ~n15924 & n15927;
  assign po1092 = n14954 | ~n15928;
  assign n15930 = ~pi0277 & ~pi0984;
  assign n15931 = n6716 & ~n15930;
  assign n15932 = ~pi0278 & n13911;
  assign n15933 = pi0984 & n15932;
  assign n15934 = ~n15931 & ~n15933;
  assign po1093 = ~po1785 & ~n15934;
  assign n15936 = n15750 & n15759;
  assign po1094 = pi0985 & n15936;
  assign n15938 = ~pi0986 & pi1548;
  assign po1095 = n6325 & ~n15938;
  assign n15940 = ~pi0987 & pi1523;
  assign po1096 = n6325 & ~n15940;
  assign n15942 = pi1414 & ~pi1773;
  assign n15943 = pi1773 & pi1819;
  assign po1097 = n15942 | n15943;
  assign n15945 = pi1415 & ~pi1773;
  assign n15946 = pi1773 & pi1821;
  assign po1098 = n15945 | n15946;
  assign n15948 = ~pi0990 & ~n8403;
  assign po1099 = n6201 & ~n15948;
  assign n15950 = pi1430 & n5440;
  assign n15951 = ~pi0991 & ~n15950;
  assign po1100 = n6193 & ~n15951;
  assign n15953 = pi1480 & pi1698;
  assign n15954 = pi0992 & ~n15953;
  assign n15955 = pi0064 & n15953;
  assign n15956 = ~n15954 & ~n15955;
  assign po1101 = pi1747 & ~n15956;
  assign n15958 = pi0993 & ~n15953;
  assign n15959 = pi0057 & n15953;
  assign n15960 = ~n15958 & ~n15959;
  assign po1102 = pi1747 & ~n15960;
  assign n15962 = pi1480 & pi1695;
  assign n15963 = pi0994 & ~n15962;
  assign n15964 = pi0056 & n15962;
  assign n15965 = ~n15963 & ~n15964;
  assign po1103 = pi1747 & ~n15965;
  assign n15967 = ~pi0995 & ~po1737;
  assign n15968 = n6730 & ~n15967;
  assign n15969 = ~pi0276 & n15274;
  assign n15970 = pi0995 & n15969;
  assign n15971 = ~n15968 & ~n15970;
  assign po1104 = ~po1785 & ~n15971;
  assign po1105 = ~n4173 & n5094;
  assign n15974 = ~pi0811 & n4173;
  assign n15975 = ~pi0835 & ~n4173;
  assign po1106 = n15974 | n15975;
  assign n15977 = ~pi0820 & n4173;
  assign n15978 = ~pi0843 & ~n4173;
  assign po1107 = n15977 | n15978;
  assign n15980 = ~pi0828 & n4173;
  assign n15981 = ~pi0851 & ~n4173;
  assign po1108 = n15980 | n15981;
  assign n15983 = ~pi0814 & n4173;
  assign n15984 = ~pi0837 & ~n4173;
  assign po1109 = n15983 | n15984;
  assign n15986 = ~pi0815 & n4173;
  assign n15987 = ~pi0838 & ~n4173;
  assign po1110 = n15986 | n15987;
  assign n15989 = ~pi0870 & n4173;
  assign n15990 = ~pi0752 & ~n4173;
  assign po1111 = n15989 | n15990;
  assign n15992 = ~pi0816 & n4173;
  assign n15993 = ~pi0839 & ~n4173;
  assign po1112 = n15992 | n15993;
  assign n15995 = ~pi0817 & n4173;
  assign n15996 = ~pi0840 & ~n4173;
  assign po1113 = n15995 | n15996;
  assign n15998 = ~pi0756 & n4173;
  assign n15999 = ~pi0880 & ~n4173;
  assign po1114 = n15998 | n15999;
  assign n16001 = ~pi0830 & n4173;
  assign n16002 = ~pi0854 & ~n4173;
  assign po1115 = n16001 | n16002;
  assign n16004 = ~pi0831 & n4173;
  assign n16005 = ~pi0855 & ~n4173;
  assign po1116 = n16004 | n16005;
  assign n16007 = ~pi0832 & n4173;
  assign n16008 = ~pi0856 & ~n4173;
  assign po1117 = n16007 | n16008;
  assign n16010 = ~pi0757 & n4173;
  assign n16011 = ~pi0879 & ~n4173;
  assign po1118 = n16010 | n16011;
  assign n16013 = ~pi0833 & n4173;
  assign n16014 = ~pi0857 & ~n4173;
  assign po1119 = n16013 | n16014;
  assign n16016 = ~pi0834 & n4173;
  assign n16017 = ~pi0858 & ~n4173;
  assign po1120 = n16016 | n16017;
  assign n16019 = ~pi0812 & n4173;
  assign n16020 = ~pi0758 & ~n4173;
  assign po1121 = n16019 | n16020;
  assign n16022 = ~pi0813 & n4173;
  assign n16023 = ~pi0836 & ~n4173;
  assign po1122 = n16022 | n16023;
  assign n16025 = pi1014 & ~n15962;
  assign n16026 = pi0049 & n15962;
  assign n16027 = ~n16025 & ~n16026;
  assign po1123 = pi1747 & ~n16027;
  assign n16029 = pi0987 & ~pi1325;
  assign n16030 = ~pi1611 & ~n16029;
  assign n16031 = pi1612 & pi1620;
  assign n16032 = pi1613 & n16031;
  assign n16033 = n16030 & n16032;
  assign n16034 = pi0901 & ~pi1328;
  assign n16035 = pi0915 & ~pi1327;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = n16033 & n16036;
  assign n16038 = pi0136 & ~pi1326;
  assign n16039 = pi0786 & ~pi1288;
  assign n16040 = ~n16038 & ~n16039;
  assign n16041 = pi0977 & ~pi1330;
  assign n16042 = pi0644 & ~pi1324;
  assign n16043 = ~n16041 & ~n16042;
  assign n16044 = pi0986 & ~pi1339;
  assign n16045 = pi0728 & ~pi1329;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = n16043 & n16046;
  assign n16048 = n16040 & n16047;
  assign po1124 = ~n16037 | ~n16048;
  assign n16050 = n14944 & n15891;
  assign n16051 = n14934 & n16050;
  assign n16052 = ~pi0771 & n16051;
  assign n16053 = pi0799 & n16052;
  assign n16054 = ~pi0802 & n14918;
  assign n16055 = ~n14944 & ~n16054;
  assign n16056 = ~pi0800 & ~pi0801;
  assign n16057 = n15891 & n16056;
  assign n16058 = pi0799 & n16057;
  assign n16059 = ~n16055 & n16058;
  assign n16060 = n8885 & n15890;
  assign n16061 = ~n16059 & ~n16060;
  assign po1125 = n16053 | ~n16061;
  assign n16063 = n8879 & n12688;
  assign n16064 = ~pi1738 & n16063;
  assign n16065 = pi1017 & ~n16063;
  assign po1126 = n16064 | n16065;
  assign n16067 = ~pi0076 & n3955;
  assign n16068 = n5575 & n5588;
  assign n16069 = n5580 & n16068;
  assign n16070 = pi0073 & n16069;
  assign n16071 = n16067 & n16070;
  assign n16072 = ~po1655 & ~n16071;
  assign n16073 = pi1018 & n16072;
  assign n16074 = ~n5585 & ~n16073;
  assign po1127 = pi1747 & ~n16074;
  assign n16076 = ~pi0262 & n6726;
  assign n16077 = pi1019 & n16076;
  assign n16078 = ~pi1019 & ~n15599;
  assign n16079 = n6720 & ~n16078;
  assign n16080 = ~n13795 & n16079;
  assign n16081 = ~n6754 & n16080;
  assign n16082 = ~n16077 & ~n16081;
  assign po1128 = ~po1785 & ~n16082;
  assign n16084 = pi0987 & pi1319;
  assign n16085 = ~pi1617 & ~n16084;
  assign n16086 = pi1618 & pi1619;
  assign n16087 = pi1616 & n16086;
  assign n16088 = n16085 & n16087;
  assign n16089 = pi0901 & pi1321;
  assign n16090 = pi0915 & pi1290;
  assign n16091 = ~n16089 & ~n16090;
  assign n16092 = n16088 & n16091;
  assign n16093 = pi0136 & pi1289;
  assign n16094 = pi0786 & pi1320;
  assign n16095 = ~n16093 & ~n16094;
  assign n16096 = pi0977 & ~pi1287;
  assign n16097 = pi0644 & pi1291;
  assign n16098 = ~n16096 & ~n16097;
  assign n16099 = pi0986 & ~pi1323;
  assign n16100 = pi0728 & pi1322;
  assign n16101 = ~n16099 & ~n16100;
  assign n16102 = n16098 & n16101;
  assign n16103 = n16095 & n16102;
  assign po1129 = ~n16092 | ~n16103;
  assign n16105 = ~pi1670 & n6753;
  assign n16106 = pi1021 & n13915;
  assign n16107 = ~n16105 & ~n16106;
  assign n16108 = n13802 & ~n16107;
  assign n16109 = pi1021 & ~n13321;
  assign n16110 = ~pi1670 & n16109;
  assign n16111 = ~n16105 & ~n16110;
  assign n16112 = n13814 & ~n16111;
  assign n16113 = ~n16108 & ~n16112;
  assign po1130 = ~po1785 & ~n16113;
  assign n16115 = n8006 & n13676;
  assign n16116 = pi1776 & n16115;
  assign n16117 = pi1022 & ~n16115;
  assign n16118 = ~n16116 & ~n16117;
  assign po1131 = pi1747 & ~n16118;
  assign n16120 = pi1778 & n16115;
  assign n16121 = pi1023 & ~n16115;
  assign n16122 = ~n16120 & ~n16121;
  assign po1132 = pi1747 & ~n16122;
  assign n16124 = pi1790 & n16115;
  assign n16125 = pi1024 & ~n16115;
  assign n16126 = ~n16124 & ~n16125;
  assign po1133 = pi1747 & ~n16126;
  assign n16128 = pi1791 & n16115;
  assign n16129 = pi1025 & ~n16115;
  assign n16130 = ~n16128 & ~n16129;
  assign po1134 = pi1747 & ~n16130;
  assign n16132 = pi1792 & n16115;
  assign n16133 = pi1026 & ~n16115;
  assign n16134 = ~n16132 & ~n16133;
  assign po1135 = pi1747 & ~n16134;
  assign n16136 = n8355 & n13676;
  assign n16137 = pi1776 & n16136;
  assign n16138 = pi1027 & ~n16136;
  assign n16139 = ~n16137 & ~n16138;
  assign po1136 = pi1747 & ~n16139;
  assign n16141 = pi1779 & n16136;
  assign n16142 = pi1028 & ~n16136;
  assign n16143 = ~n16141 & ~n16142;
  assign po1137 = pi1747 & ~n16143;
  assign n16145 = pi1783 & n16136;
  assign n16146 = pi1029 & ~n16136;
  assign n16147 = ~n16145 & ~n16146;
  assign po1138 = pi1747 & ~n16147;
  assign n16149 = pi1799 & n16136;
  assign n16150 = ~pi1030 & ~n16136;
  assign n16151 = ~n16149 & ~n16150;
  assign po1139 = pi1747 & ~n16151;
  assign n16153 = n9429 & n13676;
  assign n16154 = pi1774 & n16153;
  assign n16155 = ~pi1031 & ~n16153;
  assign n16156 = ~n16154 & ~n16155;
  assign po1140 = pi1747 & ~n16156;
  assign n16158 = pi1776 & n16153;
  assign n16159 = pi1032 & ~n16153;
  assign n16160 = ~n16158 & ~n16159;
  assign po1141 = pi1747 & ~n16160;
  assign n16162 = pi1780 & n16153;
  assign n16163 = pi1033 & ~n16153;
  assign n16164 = ~n16162 & ~n16163;
  assign po1142 = pi1747 & ~n16164;
  assign n16166 = pi1783 & n16153;
  assign n16167 = pi1034 & ~n16153;
  assign n16168 = ~n16166 & ~n16167;
  assign po1143 = pi1747 & ~n16168;
  assign n16170 = pi1459 & n5440;
  assign n16171 = ~pi1035 & ~n16170;
  assign po1144 = n6185 & ~n16171;
  assign n16173 = pi1036 & ~n8356;
  assign n16174 = pi1747 & ~n16173;
  assign po1145 = n9397 | ~n16174;
  assign n16176 = pi1447 & n5440;
  assign n16177 = ~pi1037 & ~n16176;
  assign po1146 = n6201 & ~n16177;
  assign n16179 = ~pi1021 & n15163;
  assign n16180 = n15199 & n16179;
  assign n16181 = n6699 & n16180;
  assign n16182 = n15166 & n16181;
  assign n16183 = n15170 & n16182;
  assign n16184 = ~pi0971 & n6764;
  assign n16185 = n16183 & n16184;
  assign n16186 = pi0971 & n6754;
  assign n16187 = ~n16185 & ~n16186;
  assign n16188 = ~n6723 & ~n6727;
  assign n16189 = n16182 & ~n16188;
  assign n16190 = n15184 & n16189;
  assign n16191 = ~pi1677 & n16190;
  assign po1424 = ~n16187 | n16191;
  assign n16193 = n6696 & n13323;
  assign n16194 = n6733 & n13312;
  assign n16195 = ~n16193 & ~n16194;
  assign n16196 = ~pi1038 & n16195;
  assign po1147 = ~po1424 & ~n16196;
  assign n16198 = ~pi1733 & n16063;
  assign n16199 = pi1039 & ~n16063;
  assign po1148 = n16198 | n16199;
  assign n16201 = ~pi1741 & n16063;
  assign n16202 = pi1040 & ~n16063;
  assign po1149 = n16201 | n16202;
  assign n16204 = ~pi1727 & n16063;
  assign n16205 = pi1041 & ~n16063;
  assign po1150 = n16204 | n16205;
  assign n16207 = ~pi1740 & n16063;
  assign n16208 = pi1042 & ~n16063;
  assign po1151 = n16207 | n16208;
  assign n16210 = ~pi1735 & n16063;
  assign n16211 = pi1043 & ~n16063;
  assign po1152 = n16210 | n16211;
  assign n16213 = ~pi1725 & n16063;
  assign n16214 = pi1044 & ~n16063;
  assign po1153 = n16213 | n16214;
  assign n16216 = ~pi0262 & ~pi1045;
  assign n16217 = n6726 & ~n16216;
  assign n16218 = ~pi0277 & n15657;
  assign n16219 = pi1045 & n16218;
  assign n16220 = ~n16217 & ~n16219;
  assign po1154 = ~po1785 & ~n16220;
  assign n16222 = ~n6739 & ~n6743;
  assign n16223 = pi1046 & n16222;
  assign n16224 = ~n15210 & ~n16223;
  assign n16225 = n6735 & ~n16224;
  assign n16226 = n6709 & ~n6759;
  assign n16227 = pi1046 & n16226;
  assign n16228 = ~n13322 & n16227;
  assign n16229 = ~n16225 & ~n16228;
  assign po1155 = ~po1785 & ~n16229;
  assign po1156 = n4173 & n5094;
  assign n16232 = ~pi1048 & ~n9731;
  assign po1157 = n6185 & ~n16232;
  assign n16234 = ~pi1722 & n16063;
  assign n16235 = pi1049 & ~n16063;
  assign po1158 = n16234 | n16235;
  assign n16237 = pi0183 & n13317;
  assign n16238 = pi1050 & n16237;
  assign n16239 = ~n6765 & ~n16238;
  assign po1159 = ~po1785 & ~n16239;
  assign n16241 = n9549 & n13676;
  assign n16242 = pi1791 & n16241;
  assign n16243 = pi1051 & ~n16241;
  assign n16244 = ~n16242 & ~n16243;
  assign po1160 = pi1747 & ~n16244;
  assign n16246 = ~pi1052 & ~n16241;
  assign n16247 = pi1787 & n16241;
  assign n16248 = ~n16246 & ~n16247;
  assign po1161 = pi1747 & ~n16248;
  assign n16250 = ~pi1053 & ~n8007;
  assign n16251 = pi1747 & ~n16250;
  assign po1162 = n8136 | ~n16251;
  assign n16253 = pi1792 & n16136;
  assign n16254 = pi1054 & ~n16136;
  assign n16255 = ~n16253 & ~n16254;
  assign po1163 = pi1747 & ~n16255;
  assign n16257 = ~pi1055 & ~n8007;
  assign n16258 = pi1747 & ~n16257;
  assign po1164 = n8343 | ~n16258;
  assign n16260 = pi1056 & ~n9430;
  assign n16261 = pi1747 & ~n16260;
  assign po1165 = n12098 | ~n16261;
  assign n16263 = pi1057 & ~n9430;
  assign n16264 = pi1747 & ~n16263;
  assign po1166 = n9431 | ~n16264;
  assign n16266 = n8873 & n8905;
  assign n16267 = ~pi0382 & n16266;
  assign n16268 = ~pi1738 & n16267;
  assign n16269 = pi1058 & ~n16267;
  assign n16270 = ~n16268 & ~n16269;
  assign po1167 = ~pi1747 | ~n16270;
  assign n16272 = pi0273 & n13715;
  assign n16273 = pi0136 & n13712;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = ~pi1329 & n13708;
  assign n16276 = n16274 & ~n16275;
  assign n16277 = n13722 & ~n16276;
  assign n16278 = ~pi1360 & n13676;
  assign n16279 = ~pi0438 & n7999;
  assign n16280 = ~pi0396 & n8080;
  assign n16281 = ~n16279 & ~n16280;
  assign n16282 = ~n16278 & n16281;
  assign n16283 = n13724 & ~n16282;
  assign n16284 = n13733 & ~n16276;
  assign n16285 = ~n16283 & ~n16284;
  assign n16286 = ~pi1369 & n13676;
  assign n16287 = ~pi0536 & n7999;
  assign n16288 = ~pi0495 & n8080;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = ~n16286 & n16289;
  assign n16291 = n13672 & ~n16290;
  assign n16292 = ~pi0525 & n7999;
  assign n16293 = ~pi0576 & n8080;
  assign n16294 = ~n16292 & ~n16293;
  assign n16295 = ~pi1413 & n13676;
  assign n16296 = n16294 & ~n16295;
  assign n16297 = n13684 & ~n16296;
  assign n16298 = ~n16291 & ~n16297;
  assign n16299 = ~pi1361 & n13676;
  assign n16300 = ~pi0604 & n7999;
  assign n16301 = ~pi0686 & n8080;
  assign n16302 = ~n16300 & ~n16301;
  assign n16303 = ~n16299 & n16302;
  assign n16304 = n13700 & ~n16303;
  assign n16305 = n16298 & ~n16304;
  assign n16306 = n16285 & n16305;
  assign po1168 = n16277 | ~n16306;
  assign n16308 = pi0252 & n13715;
  assign n16309 = pi0786 & n13712;
  assign n16310 = ~n16308 & ~n16309;
  assign n16311 = ~pi1339 & n13708;
  assign n16312 = n16310 & ~n16311;
  assign n16313 = n13722 & ~n16312;
  assign n16314 = ~pi1184 & n13676;
  assign n16315 = ~pi0343 & n7999;
  assign n16316 = ~pi0399 & n8080;
  assign n16317 = ~n16315 & ~n16316;
  assign n16318 = ~n16314 & n16317;
  assign n16319 = n13724 & ~n16318;
  assign n16320 = n13733 & ~n16312;
  assign n16321 = ~n16319 & ~n16320;
  assign n16322 = ~pi1206 & n13676;
  assign n16323 = ~pi0420 & n7999;
  assign n16324 = ~pi0446 & n8080;
  assign n16325 = ~n16323 & ~n16324;
  assign n16326 = ~n16322 & n16325;
  assign n16327 = n13672 & ~n16326;
  assign n16328 = ~pi0602 & n7999;
  assign n16329 = ~pi0687 & n8080;
  assign n16330 = ~n16328 & ~n16329;
  assign n16331 = ~pi1164 & n13676;
  assign n16332 = n16330 & ~n16331;
  assign n16333 = n13700 & ~n16332;
  assign n16334 = ~n16327 & ~n16333;
  assign n16335 = ~pi0657 & n7999;
  assign n16336 = ~pi0577 & n8080;
  assign n16337 = ~n16335 & ~n16336;
  assign n16338 = ~pi1225 & n13676;
  assign n16339 = n16337 & ~n16338;
  assign n16340 = n13684 & ~n16339;
  assign n16341 = n16334 & ~n16340;
  assign n16342 = n16321 & n16341;
  assign po1169 = n16313 | ~n16342;
  assign n16344 = pi0467 & n13715;
  assign n16345 = pi1685 & n13710;
  assign n16346 = ~n16344 & ~n16345;
  assign n16347 = ~pi1323 & n13708;
  assign n16348 = n16346 & ~n16347;
  assign n16349 = n13722 & ~n16348;
  assign n16350 = pi1274 & n13676;
  assign n16351 = ~pi0324 & n7999;
  assign n16352 = ~pi0330 & n8080;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = ~n16350 & n16353;
  assign n16355 = n13724 & ~n16354;
  assign n16356 = n13733 & ~n16348;
  assign n16357 = ~n16355 & ~n16356;
  assign n16358 = pi1130 & n13676;
  assign n16359 = ~pi0371 & n7999;
  assign n16360 = ~pi0375 & n8080;
  assign n16361 = ~n16359 & ~n16360;
  assign n16362 = ~n16358 & n16361;
  assign n16363 = n13672 & ~n16362;
  assign n16364 = pi1142 & n13676;
  assign n16365 = ~pi0459 & n7999;
  assign n16366 = ~pi0464 & n8080;
  assign n16367 = ~n16365 & ~n16366;
  assign n16368 = ~n16364 & n16367;
  assign n16369 = n13684 & ~n16368;
  assign n16370 = ~n16363 & ~n16369;
  assign n16371 = pi1081 & n13676;
  assign n16372 = ~pi0558 & n7999;
  assign n16373 = ~pi0624 & n8080;
  assign n16374 = ~n16372 & ~n16373;
  assign n16375 = ~n16371 & n16374;
  assign n16376 = n13700 & ~n16375;
  assign n16377 = n16370 & ~n16376;
  assign n16378 = n16357 & n16377;
  assign po1170 = n16349 | ~n16378;
  assign n16380 = ~pi1062 & ~n9430;
  assign n16381 = pi1747 & ~n16380;
  assign po1171 = n9710 | ~n16381;
  assign n16383 = ~pi1063 & ~n8356;
  assign n16384 = pi1747 & ~n16383;
  assign po1172 = n8592 | ~n16384;
  assign n16386 = ~pi1064 & ~n9430;
  assign n16387 = pi1747 & ~n16386;
  assign po1173 = n10618 | ~n16387;
  assign n16389 = ~pi1065 & ~n8356;
  assign n16390 = pi1747 & ~n16389;
  assign po1174 = n11588 | ~n16390;
  assign n16392 = pi1066 & ~n9430;
  assign n16393 = pi1747 & ~n16392;
  assign po1175 = n12088 | ~n16393;
  assign n16395 = ~pi1067 & ~n8007;
  assign n16396 = pi1747 & ~n16395;
  assign po1176 = n9765 | ~n16396;
  assign n16398 = ~pi1759 & ~pi1760;
  assign n16399 = n8005 & n13721;
  assign n16400 = n16398 & n16399;
  assign n16401 = pi1758 & n16400;
  assign n16402 = pi1779 & n16401;
  assign n16403 = pi1068 & ~n16401;
  assign n16404 = ~n16402 & ~n16403;
  assign po1177 = pi1747 & ~n16404;
  assign n16406 = pi1777 & n16401;
  assign n16407 = pi1069 & ~n16401;
  assign n16408 = ~n16406 & ~n16407;
  assign po1178 = pi1747 & ~n16408;
  assign n16410 = pi1795 & n16241;
  assign n16411 = pi1070 & ~n16241;
  assign n16412 = ~n16410 & ~n16411;
  assign po1179 = pi1747 & ~n16412;
  assign n16414 = ~pi1071 & ~n9430;
  assign n16415 = pi1747 & ~n16414;
  assign po1180 = n10538 | ~n16415;
  assign n16417 = ~pi1287 & n13708;
  assign n16418 = pi0479 & n13715;
  assign n16419 = ~n16417 & ~n16418;
  assign n16420 = n13733 & ~n16419;
  assign n16421 = ~pi0349 & n7999;
  assign n16422 = ~pi0404 & n8080;
  assign n16423 = ~n16421 & ~n16422;
  assign n16424 = pi1270 & n13676;
  assign n16425 = n16423 & ~n16424;
  assign n16426 = n13724 & ~n16425;
  assign n16427 = ~n16420 & ~n16426;
  assign n16428 = n13722 & ~n16419;
  assign n16429 = n16427 & ~n16428;
  assign n16430 = pi1265 & n13676;
  assign n16431 = ~pi0436 & n7999;
  assign n16432 = ~pi0584 & n8080;
  assign n16433 = ~n16431 & ~n16432;
  assign n16434 = ~n16430 & n16433;
  assign n16435 = n13684 & ~n16434;
  assign n16436 = pi1109 & n13676;
  assign n16437 = ~pi0610 & n7999;
  assign n16438 = ~pi0694 & n8080;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = ~n16436 & n16439;
  assign n16441 = n13700 & ~n16440;
  assign n16442 = pi1076 & n13676;
  assign n16443 = ~pi0356 & n7999;
  assign n16444 = ~pi0503 & n8080;
  assign n16445 = ~n16443 & ~n16444;
  assign n16446 = ~n16442 & n16445;
  assign n16447 = n13672 & ~n16446;
  assign n16448 = ~n16441 & ~n16447;
  assign n16449 = ~n16435 & n16448;
  assign po1181 = ~n16429 | ~n16449;
  assign n16451 = ~pi1073 & ~n8007;
  assign n16452 = pi1747 & ~n16451;
  assign po1182 = n8112 | ~n16452;
  assign n16454 = pi1799 & n16241;
  assign n16455 = pi1074 & ~n16241;
  assign n16456 = ~n16454 & ~n16455;
  assign po1183 = pi1747 & ~n16456;
  assign n16458 = ~pi1075 & ~n8007;
  assign n16459 = pi1747 & ~n16458;
  assign po1184 = n8020 | ~n16459;
  assign n16461 = pi1782 & n16136;
  assign n16462 = pi1076 & ~n16136;
  assign n16463 = ~n16461 & ~n16462;
  assign po1185 = pi1747 & ~n16463;
  assign n16465 = pi1077 & ~n8007;
  assign n16466 = pi1747 & ~n16465;
  assign po1186 = n8263 | ~n16466;
  assign n16468 = pi1790 & n16136;
  assign n16469 = ~pi1078 & ~n16136;
  assign n16470 = ~n16468 & ~n16469;
  assign po1187 = pi1747 & ~n16470;
  assign n16472 = ~pi1725 & n16267;
  assign n16473 = pi1079 & ~n16267;
  assign n16474 = ~n16472 & ~n16473;
  assign po1188 = ~pi1747 | ~n16474;
  assign n16476 = pi1080 & ~n16136;
  assign n16477 = pi1800 & n16136;
  assign n16478 = ~n16476 & ~n16477;
  assign po1189 = pi1747 & ~n16478;
  assign n16480 = pi1781 & n16241;
  assign n16481 = pi1081 & ~n16241;
  assign n16482 = ~n16480 & ~n16481;
  assign po1190 = pi1747 & ~n16482;
  assign n16484 = pi1082 & ~n8007;
  assign n16485 = pi1747 & ~n16484;
  assign po1191 = n8008 | ~n16485;
  assign n16487 = pi1780 & n16136;
  assign n16488 = pi1083 & ~n16136;
  assign n16489 = ~n16487 & ~n16488;
  assign po1192 = pi1747 & ~n16489;
  assign n16491 = pi1786 & n16136;
  assign n16492 = ~pi1084 & ~n16136;
  assign n16493 = ~n16491 & ~n16492;
  assign po1193 = pi1747 & ~n16493;
  assign n16495 = ~pi1085 & ~n9430;
  assign n16496 = pi1747 & ~n16495;
  assign po1194 = n9700 | ~n16496;
  assign n16498 = ~pi1086 & ~n9430;
  assign n16499 = pi1747 & ~n16498;
  assign po1195 = n9571 | ~n16499;
  assign n16501 = pi1087 & ~n8007;
  assign n16502 = pi1747 & ~n16501;
  assign po1196 = n9561 | ~n16502;
  assign n16504 = ~pi0138 & pi1088;
  assign n16505 = ~n12119 & ~n16504;
  assign n16506 = n3720 & ~n16505;
  assign n16507 = pi1088 & n8211;
  assign n16508 = n3724 & n16507;
  assign n16509 = ~n16506 & ~n16508;
  assign n16510 = ~pi1088 & ~n7987;
  assign n16511 = n7986 & n7991;
  assign n16512 = ~n16510 & n16511;
  assign n16513 = n16509 & ~n16512;
  assign po1197 = pi1747 & ~n16513;
  assign n16515 = pi1089 & ~n8007;
  assign n16516 = ~n8313 & ~n16515;
  assign po1198 = ~pi1747 | ~n16516;
  assign po1687 = pi1090 & n8211;
  assign n16519 = ~n3714 & n3725;
  assign n16520 = po1687 & ~n16519;
  assign n16521 = ~pi1090 & ~n7972;
  assign n16522 = n7971 & ~n16521;
  assign n16523 = ~n16520 & ~n16522;
  assign po1199 = pi1747 & ~n16523;
  assign n16525 = pi1091 & n8212;
  assign n16526 = pi1091 & ~n7972;
  assign n16527 = ~n7970 & ~n16526;
  assign n16528 = n7968 & ~n16527;
  assign n16529 = ~n16525 & ~n16528;
  assign po1200 = pi1747 & ~n16529;
  assign n16531 = pi1775 & n16136;
  assign n16532 = pi1092 & ~n16136;
  assign n16533 = ~n16531 & ~n16532;
  assign po1201 = pi1747 & ~n16533;
  assign n16535 = pi1093 & ~n8007;
  assign n16536 = pi1747 & ~n16535;
  assign po1202 = n8293 | ~n16536;
  assign n16538 = pi1774 & n16401;
  assign n16539 = pi1094 & ~n16401;
  assign n16540 = ~n16538 & ~n16539;
  assign po1203 = pi1747 & ~n16540;
  assign n16542 = pi1775 & n16401;
  assign n16543 = pi1095 & ~n16401;
  assign n16544 = ~n16542 & ~n16543;
  assign po1204 = pi1747 & ~n16544;
  assign n16546 = pi1776 & n16401;
  assign n16547 = pi1096 & ~n16401;
  assign n16548 = ~n16546 & ~n16547;
  assign po1205 = pi1747 & ~n16548;
  assign n16550 = pi1778 & n16401;
  assign n16551 = pi1097 & ~n16401;
  assign n16552 = ~n16550 & ~n16551;
  assign po1206 = pi1747 & ~n16552;
  assign n16554 = pi1780 & n16401;
  assign n16555 = pi1098 & ~n16401;
  assign n16556 = ~n16554 & ~n16555;
  assign po1207 = pi1747 & ~n16556;
  assign n16558 = pi0112 & n4182;
  assign n16559 = pi0239 & ~pi0806;
  assign n16560 = ~pi0239 & pi0806;
  assign n16561 = ~n16559 & ~n16560;
  assign n16562 = ~pi0238 & ~pi0804;
  assign n16563 = pi0238 & pi0804;
  assign n16564 = ~n16562 & ~n16563;
  assign n16565 = n16561 & ~n16564;
  assign n16566 = pi0237 & ~pi0750;
  assign n16567 = ~pi0237 & pi0750;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = ~n13338 & ~n13594;
  assign n16570 = n16568 & n16569;
  assign n16571 = ~pi0221 & pi0755;
  assign n16572 = pi0221 & ~pi0755;
  assign n16573 = ~n16571 & ~n16572;
  assign n16574 = ~pi0240 & ~pi0807;
  assign n16575 = pi0240 & pi0807;
  assign n16576 = ~n16574 & ~n16575;
  assign n16577 = n16573 & ~n16576;
  assign n16578 = n16570 & n16577;
  assign n16579 = n16565 & n16578;
  assign n16580 = ~n13343 & ~n13348;
  assign n16581 = pi0243 & ~pi0759;
  assign n16582 = ~pi0243 & pi0759;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = n16580 & n16583;
  assign n16585 = ~n13357 & n16584;
  assign n16586 = ~n13362 & n16585;
  assign n16587 = n16579 & n16586;
  assign n16588 = pi0242 & ~pi0809;
  assign n16589 = ~pi0242 & pi0809;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = ~n13368 & ~n13371;
  assign n16592 = n16590 & n16591;
  assign n16593 = n16587 & n16592;
  assign po1208 = n16558 & ~n16593;
  assign n16595 = ~pi1100 & ~n16153;
  assign n16596 = pi1787 & n16153;
  assign n16597 = ~n16595 & ~n16596;
  assign po1209 = pi1747 & ~n16597;
  assign n16599 = pi1784 & n16241;
  assign n16600 = pi1102 & ~n16241;
  assign n16601 = ~n16599 & ~n16600;
  assign po1211 = pi1747 & ~n16601;
  assign n16603 = pi1786 & n16241;
  assign n16604 = ~pi1103 & ~n16241;
  assign n16605 = ~n16603 & ~n16604;
  assign po1212 = pi1747 & ~n16605;
  assign n16607 = pi1775 & n16241;
  assign n16608 = pi1104 & ~n16241;
  assign n16609 = ~n16607 & ~n16608;
  assign po1213 = pi1747 & ~n16609;
  assign n16611 = pi1776 & n16241;
  assign n16612 = pi1105 & ~n16241;
  assign n16613 = ~n16611 & ~n16612;
  assign po1214 = pi1747 & ~n16613;
  assign n16615 = pi1778 & n16241;
  assign n16616 = pi1106 & ~n16241;
  assign n16617 = ~n16615 & ~n16616;
  assign po1215 = pi1747 & ~n16617;
  assign n16619 = pi1779 & n16241;
  assign n16620 = pi1107 & ~n16241;
  assign n16621 = ~n16619 & ~n16620;
  assign po1216 = pi1747 & ~n16621;
  assign n16623 = pi1780 & n16241;
  assign n16624 = pi1108 & ~n16241;
  assign n16625 = ~n16623 & ~n16624;
  assign po1217 = pi1747 & ~n16625;
  assign n16627 = pi1782 & n16241;
  assign n16628 = pi1109 & ~n16241;
  assign n16629 = ~n16627 & ~n16628;
  assign po1218 = pi1747 & ~n16629;
  assign n16631 = pi1783 & n16241;
  assign n16632 = pi1110 & ~n16241;
  assign n16633 = ~n16631 & ~n16632;
  assign po1219 = pi1747 & ~n16633;
  assign n16635 = pi1111 & ~n16241;
  assign n16636 = pi1789 & n16241;
  assign n16637 = ~n16635 & ~n16636;
  assign po1220 = pi1747 & ~n16637;
  assign n16639 = pi1112 & ~n16241;
  assign n16640 = pi1800 & n16241;
  assign n16641 = ~n16639 & ~n16640;
  assign po1221 = pi1747 & ~n16641;
  assign n16643 = pi1113 & ~n16241;
  assign n16644 = pi1801 & n16241;
  assign n16645 = ~n16643 & ~n16644;
  assign po1222 = pi1747 & ~n16645;
  assign n16647 = pi1790 & n16241;
  assign n16648 = pi1114 & ~n16241;
  assign n16649 = ~n16647 & ~n16648;
  assign po1223 = pi1747 & ~n16649;
  assign n16651 = pi1792 & n16241;
  assign n16652 = pi1115 & ~n16241;
  assign n16653 = ~n16651 & ~n16652;
  assign po1224 = pi1747 & ~n16653;
  assign n16655 = pi1793 & n16241;
  assign n16656 = pi1116 & ~n16241;
  assign n16657 = ~n16655 & ~n16656;
  assign po1225 = pi1747 & ~n16657;
  assign n16659 = pi1794 & n16241;
  assign n16660 = pi1117 & ~n16241;
  assign n16661 = ~n16659 & ~n16660;
  assign po1226 = pi1747 & ~n16661;
  assign n16663 = pi1798 & n16241;
  assign n16664 = pi1118 & ~n16241;
  assign n16665 = ~n16663 & ~n16664;
  assign po1227 = pi1747 & ~n16665;
  assign n16667 = pi1784 & n16115;
  assign n16668 = pi1119 & ~n16115;
  assign n16669 = ~n16667 & ~n16668;
  assign po1228 = pi1747 & ~n16669;
  assign n16671 = pi1786 & n16115;
  assign n16672 = ~pi1120 & ~n16115;
  assign n16673 = ~n16671 & ~n16672;
  assign po1229 = pi1747 & ~n16673;
  assign n16675 = pi1780 & n16115;
  assign n16676 = pi1121 & ~n16115;
  assign n16677 = ~n16675 & ~n16676;
  assign po1230 = pi1747 & ~n16677;
  assign n16679 = pi1122 & ~n16115;
  assign n16680 = pi1789 & n16115;
  assign n16681 = ~n16679 & ~n16680;
  assign po1231 = pi1747 & ~n16681;
  assign n16683 = pi1794 & n16115;
  assign n16684 = pi1123 & ~n16115;
  assign n16685 = ~n16683 & ~n16684;
  assign po1232 = pi1747 & ~n16685;
  assign n16687 = pi1798 & n16115;
  assign n16688 = pi1124 & ~n16115;
  assign n16689 = ~n16687 & ~n16688;
  assign po1233 = pi1747 & ~n16689;
  assign n16691 = ~pi1125 & ~n16115;
  assign n16692 = pi1787 & n16115;
  assign n16693 = ~n16691 & ~n16692;
  assign po1234 = pi1747 & ~n16693;
  assign n16695 = pi1774 & n16136;
  assign n16696 = ~pi1126 & ~n16136;
  assign n16697 = ~n16695 & ~n16696;
  assign po1235 = pi1747 & ~n16697;
  assign n16699 = pi1784 & n16136;
  assign n16700 = pi1127 & ~n16136;
  assign n16701 = ~n16699 & ~n16700;
  assign po1236 = pi1747 & ~n16701;
  assign n16703 = pi1785 & n16136;
  assign n16704 = ~pi1128 & ~n16136;
  assign n16705 = ~n16703 & ~n16704;
  assign po1237 = pi1747 & ~n16705;
  assign n16707 = pi1778 & n16136;
  assign n16708 = pi1129 & ~n16136;
  assign n16709 = ~n16707 & ~n16708;
  assign po1238 = pi1747 & ~n16709;
  assign n16711 = pi1781 & n16136;
  assign n16712 = pi1130 & ~n16136;
  assign n16713 = ~n16711 & ~n16712;
  assign po1239 = pi1747 & ~n16713;
  assign n16715 = pi1131 & ~n16136;
  assign n16716 = pi1789 & n16136;
  assign n16717 = ~n16715 & ~n16716;
  assign po1240 = pi1747 & ~n16717;
  assign n16719 = pi1132 & ~n16136;
  assign n16720 = pi1801 & n16136;
  assign n16721 = ~n16719 & ~n16720;
  assign po1241 = pi1747 & ~n16721;
  assign n16723 = pi1791 & n16136;
  assign n16724 = ~pi1133 & ~n16136;
  assign n16725 = ~n16723 & ~n16724;
  assign po1242 = pi1747 & ~n16725;
  assign n16727 = pi1793 & n16136;
  assign n16728 = pi1134 & ~n16136;
  assign n16729 = ~n16727 & ~n16728;
  assign po1243 = pi1747 & ~n16729;
  assign n16731 = pi1794 & n16136;
  assign n16732 = pi1135 & ~n16136;
  assign n16733 = ~n16731 & ~n16732;
  assign po1244 = pi1747 & ~n16733;
  assign n16735 = pi1795 & n16136;
  assign n16736 = pi1136 & ~n16136;
  assign n16737 = ~n16735 & ~n16736;
  assign po1245 = pi1747 & ~n16737;
  assign n16739 = pi1798 & n16136;
  assign n16740 = ~pi1137 & ~n16136;
  assign n16741 = ~n16739 & ~n16740;
  assign po1246 = pi1747 & ~n16741;
  assign n16743 = ~pi1138 & ~n16136;
  assign n16744 = pi1787 & n16136;
  assign n16745 = ~n16743 & ~n16744;
  assign po1247 = pi1747 & ~n16745;
  assign n16747 = pi1784 & n16153;
  assign n16748 = pi1139 & ~n16153;
  assign n16749 = ~n16747 & ~n16748;
  assign po1248 = pi1747 & ~n16749;
  assign n16751 = pi1786 & n16153;
  assign n16752 = ~pi1140 & ~n16153;
  assign n16753 = ~n16751 & ~n16752;
  assign po1249 = pi1747 & ~n16753;
  assign n16755 = pi1778 & n16153;
  assign n16756 = pi1141 & ~n16153;
  assign n16757 = ~n16755 & ~n16756;
  assign po1250 = pi1747 & ~n16757;
  assign n16759 = pi1781 & n16153;
  assign n16760 = pi1142 & ~n16153;
  assign n16761 = ~n16759 & ~n16760;
  assign po1251 = pi1747 & ~n16761;
  assign n16763 = pi1143 & ~n16153;
  assign n16764 = pi1789 & n16153;
  assign n16765 = ~n16763 & ~n16764;
  assign po1252 = pi1747 & ~n16765;
  assign n16767 = pi1144 & ~n16153;
  assign n16768 = pi1800 & n16153;
  assign n16769 = ~n16767 & ~n16768;
  assign po1253 = pi1747 & ~n16769;
  assign n16771 = pi1790 & n16153;
  assign n16772 = pi1145 & ~n16153;
  assign n16773 = ~n16771 & ~n16772;
  assign po1254 = pi1747 & ~n16773;
  assign n16775 = pi1792 & n16153;
  assign n16776 = pi1146 & ~n16153;
  assign n16777 = ~n16775 & ~n16776;
  assign po1255 = pi1747 & ~n16777;
  assign n16779 = pi1795 & n16153;
  assign n16780 = pi1147 & ~n16153;
  assign n16781 = ~n16779 & ~n16780;
  assign po1256 = pi1747 & ~n16781;
  assign n16783 = pi1794 & n16153;
  assign n16784 = pi1148 & ~n16153;
  assign n16785 = ~n16783 & ~n16784;
  assign po1257 = pi1747 & ~n16785;
  assign n16787 = ~pi1149 & ~n9550;
  assign n16788 = pi1747 & ~n16787;
  assign po1258 = n11398 | ~n16788;
  assign n16790 = ~pi1150 & ~n9550;
  assign n16791 = pi1747 & ~n16790;
  assign po1259 = n11478 | ~n16791;
  assign n16793 = ~pi1151 & ~n9550;
  assign n16794 = pi1747 & ~n16793;
  assign po1260 = n10912 | ~n16794;
  assign n16796 = ~pi1152 & ~n9550;
  assign n16797 = pi1747 & ~n16796;
  assign po1261 = n10942 | ~n16797;
  assign n16799 = ~pi1153 & ~n9550;
  assign n16800 = pi1747 & ~n16799;
  assign po1262 = n11418 | ~n16800;
  assign n16802 = pi1154 & ~n9550;
  assign n16803 = pi1747 & ~n16802;
  assign po1263 = n10785 | ~n16803;
  assign n16805 = pi1155 & ~n9550;
  assign n16806 = pi1747 & ~n16805;
  assign po1264 = n11508 | ~n16806;
  assign n16808 = pi1156 & ~n9550;
  assign n16809 = pi1747 & ~n16808;
  assign po1265 = n11488 | ~n16809;
  assign n16811 = pi1157 & ~n9550;
  assign n16812 = pi1747 & ~n16811;
  assign po1266 = n11498 | ~n16812;
  assign n16814 = pi1158 & ~n9550;
  assign n16815 = pi1747 & ~n16814;
  assign po1267 = n11528 | ~n16815;
  assign n16817 = pi1159 & ~n9550;
  assign n16818 = pi1747 & ~n16817;
  assign po1268 = n10478 | ~n16818;
  assign n16820 = pi1160 & ~n9550;
  assign n16821 = pi1747 & ~n16820;
  assign po1269 = n11548 | ~n16821;
  assign n16823 = ~pi1161 & ~n9550;
  assign n16824 = pi1747 & ~n16823;
  assign po1270 = n9551 | ~n16824;
  assign n16826 = ~pi1162 & ~n9550;
  assign n16827 = pi1747 & ~n16826;
  assign po1271 = n10795 | ~n16827;
  assign n16829 = ~pi1163 & ~n9550;
  assign n16830 = pi1747 & ~n16829;
  assign po1272 = n11568 | ~n16830;
  assign n16832 = pi1747 & ~n16241;
  assign n16833 = ~pi1052 & pi1729;
  assign n16834 = n16832 & ~n16833;
  assign n16835 = ~pi1164 & n16834;
  assign n16836 = pi1747 & pi1797;
  assign n16837 = n16241 & n16836;
  assign po1273 = n16835 | n16837;
  assign n16839 = pi1480 & n5440;
  assign n16840 = ~pi1165 & ~n16839;
  assign po1274 = n6189 & ~n16840;
  assign n16842 = ~pi1166 & ~n8007;
  assign n16843 = pi1747 & ~n16842;
  assign po1275 = n8060 | ~n16843;
  assign n16845 = ~pi1167 & ~n8007;
  assign n16846 = pi1747 & ~n16845;
  assign po1276 = n8092 | ~n16846;
  assign n16848 = ~pi1168 & ~n8007;
  assign n16849 = pi1747 & ~n16848;
  assign po1277 = n10488 | ~n16849;
  assign n16851 = ~pi1169 & ~n8007;
  assign n16852 = pi1747 & ~n16851;
  assign po1278 = n8050 | ~n16852;
  assign n16854 = ~pi1170 & ~n8007;
  assign n16855 = pi1747 & ~n16854;
  assign po1279 = n10498 | ~n16855;
  assign n16857 = ~pi1171 & ~n8007;
  assign n16858 = pi1747 & ~n16857;
  assign po1280 = n8233 | ~n16858;
  assign n16860 = ~pi1172 & ~n8007;
  assign n16861 = pi1747 & ~n16860;
  assign po1281 = n8253 | ~n16861;
  assign n16863 = pi1173 & ~n8007;
  assign n16864 = ~n8273 & ~n16863;
  assign po1282 = ~pi1747 | ~n16864;
  assign n16866 = pi1174 & ~n8007;
  assign n16867 = pi1747 & ~n16866;
  assign po1283 = n8283 | ~n16867;
  assign n16869 = pi1175 & ~n8007;
  assign n16870 = pi1747 & ~n16869;
  assign po1284 = n8303 | ~n16870;
  assign n16872 = pi1176 & ~n8007;
  assign n16873 = ~n8040 & ~n16872;
  assign po1285 = ~pi1747 | ~n16873;
  assign n16875 = pi1177 & ~n8007;
  assign n16876 = pi1747 & ~n16875;
  assign po1286 = n10518 | ~n16876;
  assign n16878 = ~pi1178 & ~n8007;
  assign n16879 = ~n9528 & ~n16878;
  assign po1287 = ~pi1747 | ~n16879;
  assign n16881 = pi1179 & ~n8007;
  assign n16882 = pi1747 & ~n16881;
  assign po1288 = n8323 | ~n16882;
  assign n16884 = ~pi1180 & ~n8007;
  assign n16885 = pi1747 & ~n16884;
  assign po1289 = n8333 | ~n16885;
  assign n16887 = ~pi1181 & ~n8007;
  assign n16888 = pi1747 & ~n16887;
  assign po1290 = n9659 | ~n16888;
  assign n16890 = ~pi1182 & ~n8007;
  assign n16891 = pi1747 & ~n16890;
  assign po1291 = n8030 | ~n16891;
  assign n16893 = ~pi1183 & ~n9550;
  assign n16894 = pi1747 & ~n16893;
  assign po1292 = n11578 | ~n16894;
  assign n16896 = pi1747 & ~n16115;
  assign n16897 = ~pi1125 & pi1729;
  assign n16898 = n16896 & ~n16897;
  assign n16899 = ~pi1184 & n16898;
  assign n16900 = n16115 & n16836;
  assign po1293 = n16899 | n16900;
  assign n16902 = ~pi1185 & ~n8356;
  assign n16903 = pi1747 & ~n16902;
  assign po1294 = n8582 | ~n16903;
  assign n16905 = ~pi1186 & ~n8356;
  assign n16906 = pi1747 & ~n16905;
  assign po1295 = n8609 | ~n16906;
  assign n16908 = ~pi1187 & ~n8356;
  assign n16909 = pi1747 & ~n16908;
  assign po1296 = n11598 | ~n16909;
  assign n16911 = ~pi1188 & ~n8356;
  assign n16912 = pi1747 & ~n16911;
  assign po1297 = n8572 | ~n16912;
  assign n16914 = ~pi1189 & ~n8356;
  assign n16915 = pi1747 & ~n16914;
  assign po1298 = n8619 | ~n16915;
  assign n16917 = ~pi1190 & ~n8356;
  assign n16918 = pi1747 & ~n16917;
  assign po1299 = n9297 | ~n16918;
  assign n16920 = ~pi1191 & ~n8356;
  assign n16921 = pi1747 & ~n16920;
  assign po1300 = n9307 | ~n16921;
  assign n16923 = pi1192 & ~n8356;
  assign n16924 = pi1747 & ~n16923;
  assign po1301 = n9317 | ~n16924;
  assign n16926 = ~pi1193 & ~n8356;
  assign n16927 = pi1747 & ~n16926;
  assign po1302 = n9327 | ~n16927;
  assign n16929 = pi1194 & ~n8356;
  assign n16930 = pi1747 & ~n16929;
  assign po1303 = n9347 | ~n16930;
  assign n16932 = pi1195 & ~n8356;
  assign n16933 = pi1747 & ~n16932;
  assign po1304 = n10700 | ~n16933;
  assign n16935 = pi1196 & ~n8356;
  assign n16936 = pi1747 & ~n16935;
  assign po1305 = n9357 | ~n16936;
  assign n16938 = pi1197 & ~n8356;
  assign n16939 = pi1747 & ~n16938;
  assign po1306 = n9377 | ~n16939;
  assign n16941 = pi1198 & ~n8356;
  assign n16942 = pi1747 & ~n16941;
  assign po1307 = n9510 | ~n16942;
  assign n16944 = pi1199 & ~n8356;
  assign n16945 = pi1747 & ~n16944;
  assign po1308 = n9387 | ~n16945;
  assign n16947 = ~pi1200 & ~n8356;
  assign n16948 = pi1747 & ~n16947;
  assign po1309 = n10680 | ~n16948;
  assign n16950 = pi1201 & ~n8356;
  assign n16951 = pi1747 & ~n16950;
  assign po1310 = n11621 | ~n16951;
  assign n16953 = ~pi1202 & ~n8356;
  assign n16954 = pi1747 & ~n16953;
  assign po1311 = n9407 | ~n16954;
  assign n16956 = ~pi1203 & ~n8356;
  assign n16957 = pi1747 & ~n16956;
  assign po1312 = n10972 | ~n16957;
  assign n16959 = ~pi1204 & ~n8356;
  assign n16960 = pi1747 & ~n16959;
  assign po1313 = n10805 | ~n16960;
  assign n16962 = ~pi1205 & ~n8356;
  assign n16963 = pi1747 & ~n16962;
  assign po1314 = n8643 | ~n16963;
  assign n16965 = pi1747 & ~n16136;
  assign n16966 = ~pi1138 & pi1729;
  assign n16967 = n16965 & ~n16966;
  assign n16968 = ~pi1206 & n16967;
  assign n16969 = n16136 & n16836;
  assign po1315 = n16968 | n16969;
  assign n16971 = ~pi1207 & ~n9430;
  assign n16972 = pi1747 & ~n16971;
  assign po1316 = n10528 | ~n16972;
  assign n16974 = ~pi1208 & ~n9430;
  assign n16975 = pi1747 & ~n16974;
  assign po1317 = n9690 | ~n16975;
  assign n16977 = ~pi1209 & ~n9430;
  assign n16978 = pi1747 & ~n16977;
  assign po1318 = n9720 | ~n16978;
  assign n16980 = ~pi1210 & ~n9430;
  assign n16981 = pi1747 & ~n16980;
  assign po1319 = n9741 | ~n16981;
  assign n16983 = ~pi1211 & ~n9430;
  assign n16984 = pi1747 & ~n16983;
  assign po1320 = n10548 | ~n16984;
  assign n16986 = ~pi1212 & ~n9430;
  assign n16987 = pi1747 & ~n16986;
  assign po1321 = n10558 | ~n16987;
  assign n16989 = pi1213 & ~n9430;
  assign n16990 = pi1747 & ~n16989;
  assign po1322 = n9635 | ~n16990;
  assign n16992 = pi1214 & ~n9430;
  assign n16993 = pi1747 & ~n16992;
  assign po1323 = n10568 | ~n16993;
  assign n16995 = pi1215 & ~n9430;
  assign n16996 = pi1747 & ~n16995;
  assign po1324 = n12078 | ~n16996;
  assign n16998 = pi1216 & ~n9430;
  assign n16999 = pi1747 & ~n16998;
  assign po1325 = n10578 | ~n16999;
  assign n17001 = pi1217 & ~n9430;
  assign n17002 = pi1747 & ~n17001;
  assign po1326 = n10588 | ~n17002;
  assign n17004 = pi1218 & ~n9430;
  assign n17005 = pi1747 & ~n17004;
  assign po1327 = n10598 | ~n17005;
  assign n17007 = pi1219 & ~n9430;
  assign n17008 = pi1747 & ~n17007;
  assign po1328 = n11779 | ~n17008;
  assign n17010 = ~pi1220 & ~n9430;
  assign n17011 = pi1747 & ~n17010;
  assign po1329 = n11746 | ~n17011;
  assign n17013 = ~pi1221 & ~n9430;
  assign n17014 = pi1747 & ~n17013;
  assign po1330 = n9441 | ~n17014;
  assign n17016 = ~pi1222 & ~n9430;
  assign n17017 = pi1747 & ~n17016;
  assign po1331 = n11817 | ~n17017;
  assign n17019 = ~pi1223 & ~n9430;
  assign n17020 = pi1747 & ~n17019;
  assign po1332 = n9775 | ~n17020;
  assign n17022 = ~pi1224 & ~n9430;
  assign n17023 = pi1747 & ~n17022;
  assign po1333 = n12108 | ~n17023;
  assign n17025 = pi1747 & ~n16153;
  assign n17026 = ~pi1100 & pi1729;
  assign n17027 = n17025 & ~n17026;
  assign n17028 = ~pi1225 & n17027;
  assign n17029 = n16153 & n16836;
  assign po1334 = n17028 | n17029;
  assign n17031 = pi1445 & ~pi1773;
  assign n17032 = pi1773 & pi1820;
  assign po1335 = n17031 | n17032;
  assign n17034 = ~pi1733 & n16267;
  assign n17035 = pi1227 & ~n16267;
  assign n17036 = ~n17034 & ~n17035;
  assign po1336 = pi1747 & ~n17036;
  assign n17038 = ~pi1741 & n16267;
  assign n17039 = pi1228 & ~n16267;
  assign n17040 = ~n17038 & ~n17039;
  assign po1337 = pi1747 & ~n17040;
  assign n17042 = ~pi1722 & n16267;
  assign n17043 = pi1229 & ~n16267;
  assign n17044 = ~n17042 & ~n17043;
  assign po1338 = pi1747 & ~n17044;
  assign n17046 = ~pi1740 & n16267;
  assign n17047 = pi1230 & ~n16267;
  assign n17048 = ~n17046 & ~n17047;
  assign po1339 = ~pi1747 | ~n17048;
  assign n17050 = ~pi1735 & n16267;
  assign n17051 = pi1231 & ~n16267;
  assign n17052 = ~n17050 & ~n17051;
  assign po1340 = ~pi1747 | ~n17052;
  assign n17054 = pi1232 & ~n9430;
  assign n17055 = pi1747 & ~n17054;
  assign po1341 = n10608 | ~n17055;
  assign po1342 = pi1427 | n8901;
  assign n17058 = pi1774 & n16115;
  assign n17059 = ~pi1235 & ~n16115;
  assign n17060 = ~n17058 & ~n17059;
  assign po1344 = pi1747 & ~n17060;
  assign n17062 = ~pi1727 & n16267;
  assign n17063 = pi1236 & ~n16267;
  assign n17064 = ~n17062 & ~n17063;
  assign po1345 = pi1747 & ~n17064;
  assign n17066 = pi1774 & n16241;
  assign n17067 = ~pi1237 & ~n16241;
  assign n17068 = ~n17066 & ~n17067;
  assign po1346 = pi1747 & ~n17068;
  assign n17070 = ~pi1238 & ~n8356;
  assign n17071 = pi1747 & ~n17070;
  assign po1347 = n8369 | ~n17071;
  assign n17073 = ~pi1239 & ~n8007;
  assign n17074 = pi1747 & ~n17073;
  assign po1348 = n8070 | ~n17074;
  assign n17076 = ~pi1240 & ~n8356;
  assign n17077 = pi1747 & ~n17076;
  assign po1349 = n9417 | ~n17077;
  assign n17079 = pi1241 & ~n8007;
  assign n17080 = pi1747 & ~n17079;
  assign po1350 = n8243 | ~n17080;
  assign n17082 = pi1798 & n16153;
  assign n17083 = pi1242 & ~n16153;
  assign n17084 = ~n17082 & ~n17083;
  assign po1351 = pi1747 & ~n17084;
  assign n17086 = pi1785 & n16241;
  assign n17087 = ~pi1243 & ~n16241;
  assign n17088 = ~n17086 & ~n17087;
  assign po1352 = pi1747 & ~n17088;
  assign n17090 = ~pi1244 & ~n8356;
  assign n17091 = pi1747 & ~n17090;
  assign po1353 = n8562 | ~n17091;
  assign n17093 = ~pi1245 & ~n8356;
  assign n17094 = pi1747 & ~n17093;
  assign po1354 = n8392 | ~n17094;
  assign n17096 = ~pi1246 & ~n8007;
  assign n17097 = pi1747 & ~n17096;
  assign po1355 = n8102 | ~n17097;
  assign n17099 = ~pi1247 & ~n8007;
  assign n17100 = pi1747 & ~n17099;
  assign po1356 = n10508 | ~n17100;
  assign n17102 = ~pi1248 & ~n8356;
  assign n17103 = pi1747 & ~n17102;
  assign po1357 = n11608 | ~n17103;
  assign n17105 = pi1249 & ~n8356;
  assign n17106 = pi1747 & ~n17105;
  assign po1358 = n8357 | ~n17106;
  assign po1360 = pi1418 | po1655;
  assign n17109 = pi1799 & n16115;
  assign n17110 = pi1252 & ~n16115;
  assign n17111 = ~n17109 & ~n17110;
  assign po1361 = pi1747 & ~n17111;
  assign n17113 = pi1793 & n16153;
  assign n17114 = pi1253 & ~n16153;
  assign n17115 = ~n17113 & ~n17114;
  assign po1362 = pi1747 & ~n17115;
  assign n17117 = ~pi1254 & ~n8007;
  assign n17118 = pi1747 & ~n17117;
  assign po1363 = n8223 | ~n17118;
  assign n17120 = pi1791 & n16153;
  assign n17121 = pi1255 & ~n16153;
  assign n17122 = ~n17120 & ~n17121;
  assign po1364 = pi1747 & ~n17122;
  assign n17124 = pi1256 & ~n16115;
  assign n17125 = pi1800 & n16115;
  assign n17126 = ~n17124 & ~n17125;
  assign po1365 = pi1747 & ~n17126;
  assign n17128 = pi1257 & ~n16115;
  assign n17129 = pi1801 & n16115;
  assign n17130 = ~n17128 & ~n17129;
  assign po1366 = pi1747 & ~n17130;
  assign n17132 = pi1779 & n16153;
  assign n17133 = pi1258 & ~n16153;
  assign n17134 = ~n17132 & ~n17133;
  assign po1367 = pi1747 & ~n17134;
  assign n17136 = pi1259 & ~n16153;
  assign n17137 = pi1801 & n16153;
  assign n17138 = ~n17136 & ~n17137;
  assign po1368 = pi1747 & ~n17138;
  assign n17140 = pi1793 & n16115;
  assign n17141 = pi1260 & ~n16115;
  assign n17142 = ~n17140 & ~n17141;
  assign po1369 = pi1747 & ~n17142;
  assign n17144 = pi1799 & n16153;
  assign n17145 = pi1261 & ~n16153;
  assign n17146 = ~n17144 & ~n17145;
  assign po1370 = pi1747 & ~n17146;
  assign n17148 = pi1795 & n16115;
  assign n17149 = pi1262 & ~n16115;
  assign n17150 = ~n17148 & ~n17149;
  assign po1371 = pi1747 & ~n17150;
  assign n17152 = ~pi1263 & ~n9550;
  assign n17153 = pi1747 & ~n17152;
  assign po1372 = n11558 | ~n17153;
  assign n17155 = pi1264 & ~n8356;
  assign n17156 = pi1747 & ~n17155;
  assign po1373 = n9367 | ~n17156;
  assign n17158 = pi1782 & n16153;
  assign n17159 = pi1265 & ~n16153;
  assign n17160 = ~n17158 & ~n17159;
  assign po1374 = pi1747 & ~n17160;
  assign n17162 = pi1266 & ~n9430;
  assign n17163 = pi1747 & ~n17162;
  assign po1375 = n10628 | ~n17163;
  assign n17165 = pi1783 & n16115;
  assign n17166 = pi1267 & ~n16115;
  assign n17167 = ~n17165 & ~n17166;
  assign po1376 = pi1747 & ~n17167;
  assign n17169 = pi1785 & n16115;
  assign n17170 = ~pi1268 & ~n16115;
  assign n17171 = ~n17169 & ~n17170;
  assign po1377 = pi1747 & ~n17171;
  assign n17173 = pi1269 & ~n9550;
  assign n17174 = pi1747 & ~n17173;
  assign po1378 = n10754 | ~n17174;
  assign n17176 = pi1782 & n16115;
  assign n17177 = pi1270 & ~n16115;
  assign n17178 = ~n17176 & ~n17177;
  assign po1379 = pi1747 & ~n17178;
  assign n17180 = pi1775 & n16153;
  assign n17181 = pi1271 & ~n16153;
  assign n17182 = ~n17180 & ~n17181;
  assign po1380 = pi1747 & ~n17182;
  assign n17184 = pi1779 & n16115;
  assign n17185 = pi1272 & ~n16115;
  assign n17186 = ~n17184 & ~n17185;
  assign po1381 = pi1747 & ~n17186;
  assign n17188 = pi1785 & n16153;
  assign n17189 = ~pi1273 & ~n16153;
  assign n17190 = ~n17188 & ~n17189;
  assign po1382 = pi1747 & ~n17190;
  assign n17192 = pi1781 & n16115;
  assign n17193 = pi1274 & ~n16115;
  assign n17194 = ~n17192 & ~n17193;
  assign po1383 = pi1747 & ~n17194;
  assign n17196 = pi1275 & ~n9550;
  assign n17197 = pi1747 & ~n17196;
  assign po1384 = n10771 | ~n17197;
  assign n17199 = pi1276 & ~n8356;
  assign n17200 = pi1747 & ~n17199;
  assign po1385 = n9337 | ~n17200;
  assign n17202 = pi1777 & n16115;
  assign n17203 = pi1277 & ~n16115;
  assign n17204 = ~n17202 & ~n17203;
  assign po1386 = pi1747 & ~n17204;
  assign n17206 = ~pi1278 & ~n9430;
  assign n17207 = pi1747 & ~n17206;
  assign po1387 = n9680 | ~n17207;
  assign n17209 = ~pi1279 & ~n9430;
  assign n17210 = pi1747 & ~n17209;
  assign po1388 = n9538 | ~n17210;
  assign n17212 = pi1775 & n16115;
  assign n17213 = pi1280 & ~n16115;
  assign n17214 = ~n17212 & ~n17213;
  assign po1389 = pi1747 & ~n17214;
  assign n17216 = ~pi1281 & ~n9430;
  assign n17217 = pi1747 & ~n17216;
  assign po1390 = n11875 | ~n17217;
  assign n17219 = ~pi1282 & ~n9430;
  assign n17220 = pi1747 & ~n17219;
  assign po1391 = n10638 | ~n17220;
  assign n17222 = pi1283 & ~n9550;
  assign n17223 = pi1747 & ~n17222;
  assign po1392 = n11468 | ~n17223;
  assign n17225 = ~pi1284 & ~n9550;
  assign n17226 = pi1747 & ~n17225;
  assign po1393 = n11438 | ~n17226;
  assign n17228 = pi1285 & ~po1535;
  assign n17229 = ~pi1738 & po1535;
  assign po1394 = n17228 | n17229;
  assign n17231 = ~pi0559 & n7999;
  assign n17232 = ~pi0374 & n8080;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = pi1129 & n13676;
  assign n17235 = pi0891 & n13678;
  assign n17236 = ~n17234 & ~n17235;
  assign n17237 = n17233 & n17236;
  assign n17238 = n13672 & ~n17237;
  assign n17239 = ~pi0557 & n7999;
  assign n17240 = ~pi0641 & n8080;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = pi1106 & n13676;
  assign n17243 = pi0892 & n13678;
  assign n17244 = ~n17242 & ~n17243;
  assign n17245 = n17241 & n17244;
  assign n17246 = n13700 & ~n17245;
  assign n17247 = ~pi0632 & n7999;
  assign n17248 = ~pi0462 & n8080;
  assign n17249 = ~n17247 & ~n17248;
  assign n17250 = pi1141 & n13676;
  assign n17251 = pi0903 & n13678;
  assign n17252 = ~n17250 & ~n17251;
  assign n17253 = n17249 & n17252;
  assign n17254 = n13684 & ~n17253;
  assign n17255 = ~n17246 & ~n17254;
  assign n17256 = pi1097 & n13705;
  assign n17257 = pi1290 & n13708;
  assign n17258 = ~n17256 & ~n17257;
  assign n17259 = pi1686 & n13710;
  assign n17260 = pi1742 & n13703;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = pi0476 & n13715;
  assign n17263 = n17261 & ~n17262;
  assign n17264 = n17258 & n17263;
  assign n17265 = n13722 & ~n17264;
  assign n17266 = ~pi0458 & n7999;
  assign n17267 = ~pi0328 & n8080;
  assign n17268 = ~n17266 & ~n17267;
  assign n17269 = pi1023 & n13676;
  assign n17270 = pi0904 & n13678;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = n17268 & n17271;
  assign n17273 = n13724 & ~n17272;
  assign n17274 = n13733 & ~n17264;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = ~n17265 & n17275;
  assign n17277 = n17255 & n17276;
  assign po1395 = n17238 | ~n17277;
  assign n17279 = ~pi1760 & ~pi1764;
  assign n17280 = ~pi1763 & n17279;
  assign n17281 = ~pi1762 & n17280;
  assign n17282 = pi1759 & ~pi1761;
  assign n17283 = n17281 & n17282;
  assign n17284 = ~pi1758 & n17283;
  assign n17285 = n8005 & n17284;
  assign n17286 = pi1782 & n17285;
  assign n17287 = ~pi1287 & ~n17285;
  assign n17288 = ~n17286 & ~n17287;
  assign po1396 = pi1747 & ~n17288;
  assign n17290 = pi1793 & n17285;
  assign n17291 = ~pi1288 & ~n17285;
  assign n17292 = ~n17290 & ~n17291;
  assign po1397 = pi1747 & ~n17292;
  assign n17294 = pi1776 & n17285;
  assign n17295 = pi1289 & ~n17285;
  assign n17296 = ~n17294 & ~n17295;
  assign po1398 = pi1747 & ~n17296;
  assign n17298 = pi1778 & n17285;
  assign n17299 = pi1290 & ~n17285;
  assign n17300 = ~n17298 & ~n17299;
  assign po1399 = pi1747 & ~n17300;
  assign n17302 = pi1774 & n17285;
  assign n17303 = pi1291 & ~n17285;
  assign n17304 = ~n17302 & ~n17303;
  assign po1400 = pi1747 & ~n17304;
  assign n17306 = ~pi1292 & ~n9550;
  assign n17307 = pi1747 & ~n17306;
  assign po1401 = n11458 | ~n17307;
  assign n17309 = ~pi0418 & n7999;
  assign n17310 = ~pi0493 & n8080;
  assign n17311 = ~n17309 & ~n17310;
  assign n17312 = pi1135 & n13676;
  assign n17313 = ~pi1391 & n13678;
  assign n17314 = ~n17312 & ~n17313;
  assign n17315 = n17311 & n17314;
  assign n17316 = n13672 & ~n17315;
  assign n17317 = ~pi0524 & n7999;
  assign n17318 = ~pi0538 & n8080;
  assign n17319 = ~n17317 & ~n17318;
  assign n17320 = pi1148 & n13676;
  assign n17321 = ~pi1379 & n13678;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = n17319 & n17322;
  assign n17324 = n13684 & ~n17323;
  assign n17325 = ~pi0600 & n7999;
  assign n17326 = ~pi0685 & n8080;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = pi1117 & n13676;
  assign n17329 = ~pi1351 & n13678;
  assign n17330 = ~n17328 & ~n17329;
  assign n17331 = n17327 & n17330;
  assign n17332 = n13700 & ~n17331;
  assign n17333 = ~n17324 & ~n17332;
  assign n17334 = pi0251 & n13715;
  assign n17335 = pi0644 & n13712;
  assign n17336 = ~n17334 & ~n17335;
  assign n17337 = ~pi1327 & n13708;
  assign n17338 = n17336 & ~n17337;
  assign n17339 = n13722 & ~n17338;
  assign n17340 = ~pi0341 & n7999;
  assign n17341 = ~pi0395 & n8080;
  assign n17342 = ~n17340 & ~n17341;
  assign n17343 = pi1123 & n13676;
  assign n17344 = ~pi1388 & n13678;
  assign n17345 = ~n17343 & ~n17344;
  assign n17346 = n17342 & n17345;
  assign n17347 = n13724 & ~n17346;
  assign n17348 = n13733 & ~n17338;
  assign n17349 = ~n17347 & ~n17348;
  assign n17350 = ~n17339 & n17349;
  assign n17351 = n17333 & n17350;
  assign po1402 = n17316 | ~n17351;
  assign n17353 = ~pi0414 & n7999;
  assign n17354 = ~pi0489 & n8080;
  assign n17355 = ~n17353 & ~n17354;
  assign n17356 = ~pi1078 & n13676;
  assign n17357 = ~pi1394 & n13678;
  assign n17358 = ~n17356 & ~n17357;
  assign n17359 = n17355 & n17358;
  assign n17360 = n13672 & ~n17359;
  assign n17361 = ~pi0521 & n7999;
  assign n17362 = ~pi0572 & n8080;
  assign n17363 = ~n17361 & ~n17362;
  assign n17364 = pi1145 & n13676;
  assign n17365 = ~pi1377 & n13678;
  assign n17366 = ~n17364 & ~n17365;
  assign n17367 = n17363 & n17366;
  assign n17368 = n13684 & ~n17367;
  assign n17369 = ~pi0595 & n7999;
  assign n17370 = ~pi0681 & n8080;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = pi1114 & n13676;
  assign n17373 = ~pi1357 & n13678;
  assign n17374 = ~n17372 & ~n17373;
  assign n17375 = n17371 & n17374;
  assign n17376 = n13700 & ~n17375;
  assign n17377 = ~n17368 & ~n17376;
  assign n17378 = pi0269 & n13715;
  assign n17379 = ~pi1324 & n13708;
  assign n17380 = ~n17378 & ~n17379;
  assign n17381 = n13722 & ~n17380;
  assign n17382 = n13733 & ~n17380;
  assign n17383 = ~pi0517 & n7999;
  assign n17384 = ~pi0391 & n8080;
  assign n17385 = ~n17383 & ~n17384;
  assign n17386 = pi1024 & n13676;
  assign n17387 = ~pi1397 & n13678;
  assign n17388 = ~n17386 & ~n17387;
  assign n17389 = n17385 & n17388;
  assign n17390 = n13724 & ~n17389;
  assign n17391 = ~n17382 & ~n17390;
  assign n17392 = ~n17381 & n17391;
  assign n17393 = n17377 & n17392;
  assign po1403 = n17360 | ~n17393;
  assign n17395 = ~pi0614 & n7999;
  assign n17396 = ~pi0490 & n8080;
  assign n17397 = ~n17395 & ~n17396;
  assign n17398 = ~pi1133 & n13676;
  assign n17399 = ~pi1402 & n13678;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = n17397 & n17400;
  assign n17402 = n13672 & ~n17401;
  assign n17403 = ~pi0522 & n7999;
  assign n17404 = ~pi0543 & n8080;
  assign n17405 = ~n17403 & ~n17404;
  assign n17406 = pi1255 & n13676;
  assign n17407 = ~pi1378 & n13678;
  assign n17408 = ~n17406 & ~n17407;
  assign n17409 = n17405 & n17408;
  assign n17410 = n13684 & ~n17409;
  assign n17411 = pi1051 & n13676;
  assign n17412 = ~pi1355 & n13678;
  assign n17413 = ~n17411 & ~n17412;
  assign n17414 = ~pi0596 & n7999;
  assign n17415 = ~pi0682 & n8080;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = n17413 & n17416;
  assign n17418 = n13700 & ~n17417;
  assign n17419 = ~n17410 & ~n17418;
  assign n17420 = pi0271 & n13715;
  assign n17421 = ~pi1325 & n13708;
  assign n17422 = ~n17420 & ~n17421;
  assign n17423 = n13722 & ~n17422;
  assign n17424 = n13733 & ~n17422;
  assign n17425 = ~pi0518 & n7999;
  assign n17426 = ~pi0392 & n8080;
  assign n17427 = ~n17425 & ~n17426;
  assign n17428 = pi1025 & n13676;
  assign n17429 = ~pi1387 & n13678;
  assign n17430 = ~n17428 & ~n17429;
  assign n17431 = n17427 & n17430;
  assign n17432 = n13724 & ~n17431;
  assign n17433 = ~n17424 & ~n17432;
  assign n17434 = ~n17423 & n17433;
  assign n17435 = n17419 & n17434;
  assign po1404 = n17402 | ~n17435;
  assign n17437 = ~pi0415 & n7999;
  assign n17438 = ~pi0491 & n8080;
  assign n17439 = ~n17437 & ~n17438;
  assign n17440 = pi1054 & n13676;
  assign n17441 = ~pi1408 & n13678;
  assign n17442 = ~n17440 & ~n17441;
  assign n17443 = n17439 & n17442;
  assign n17444 = n13672 & ~n17443;
  assign n17445 = ~pi0597 & n7999;
  assign n17446 = ~pi0671 & n8080;
  assign n17447 = ~n17445 & ~n17446;
  assign n17448 = pi1115 & n13676;
  assign n17449 = ~pi1350 & n13678;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = n17447 & n17450;
  assign n17452 = n13700 & ~n17451;
  assign n17453 = ~pi0523 & n7999;
  assign n17454 = ~pi0573 & n8080;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = pi1146 & n13676;
  assign n17457 = ~pi1405 & n13678;
  assign n17458 = ~n17456 & ~n17457;
  assign n17459 = n17455 & n17458;
  assign n17460 = n13684 & ~n17459;
  assign n17461 = ~n17452 & ~n17460;
  assign n17462 = pi0272 & n13715;
  assign n17463 = ~pi1326 & n13708;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = n13722 & ~n17464;
  assign n17466 = n13733 & ~n17464;
  assign n17467 = ~pi0338 & n7999;
  assign n17468 = ~pi0430 & n8080;
  assign n17469 = ~n17467 & ~n17468;
  assign n17470 = pi1026 & n13676;
  assign n17471 = ~pi1395 & n13678;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = n17469 & n17472;
  assign n17474 = n13724 & ~n17473;
  assign n17475 = ~n17466 & ~n17474;
  assign n17476 = ~n17465 & n17475;
  assign n17477 = n17461 & n17476;
  assign po1405 = n17444 | ~n17477;
  assign n17479 = ~pi0416 & n7999;
  assign n17480 = ~pi0492 & n8080;
  assign n17481 = ~n17479 & ~n17480;
  assign n17482 = pi1134 & n13676;
  assign n17483 = ~pi1411 & n13678;
  assign n17484 = ~n17482 & ~n17483;
  assign n17485 = n17481 & n17484;
  assign n17486 = n13672 & ~n17485;
  assign n17487 = ~pi0598 & n7999;
  assign n17488 = ~pi0683 & n8080;
  assign n17489 = ~n17487 & ~n17488;
  assign n17490 = pi1116 & n13676;
  assign n17491 = ~pi1354 & n13678;
  assign n17492 = ~n17490 & ~n17491;
  assign n17493 = n17489 & n17492;
  assign n17494 = n13700 & ~n17493;
  assign n17495 = ~pi0444 & n7999;
  assign n17496 = ~pi0574 & n8080;
  assign n17497 = ~n17495 & ~n17496;
  assign n17498 = pi1253 & n13676;
  assign n17499 = ~pi1380 & n13678;
  assign n17500 = ~n17498 & ~n17499;
  assign n17501 = n17497 & n17500;
  assign n17502 = n13684 & ~n17501;
  assign n17503 = ~n17494 & ~n17502;
  assign n17504 = pi0270 & n13715;
  assign n17505 = ~pi1288 & n13708;
  assign n17506 = ~n17504 & ~n17505;
  assign n17507 = n13722 & ~n17506;
  assign n17508 = n13733 & ~n17506;
  assign n17509 = ~pi0339 & n7999;
  assign n17510 = ~pi0393 & n8080;
  assign n17511 = ~n17509 & ~n17510;
  assign n17512 = pi1260 & n13676;
  assign n17513 = ~pi1389 & n13678;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = n17511 & n17514;
  assign n17516 = n13724 & ~n17515;
  assign n17517 = ~n17508 & ~n17516;
  assign n17518 = ~n17507 & n17517;
  assign n17519 = n17503 & n17518;
  assign po1406 = n17486 | ~n17519;
  assign n17521 = ~pi0419 & n7999;
  assign n17522 = ~pi0494 & n8080;
  assign n17523 = ~n17521 & ~n17522;
  assign n17524 = pi1136 & n13676;
  assign n17525 = ~pi1412 & n13678;
  assign n17526 = ~n17524 & ~n17525;
  assign n17527 = n17523 & n17526;
  assign n17528 = n13672 & ~n17527;
  assign n17529 = ~pi0546 & n7999;
  assign n17530 = ~pi0668 & n8080;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = pi1070 & n13676;
  assign n17533 = ~pi1347 & n13678;
  assign n17534 = ~n17532 & ~n17533;
  assign n17535 = n17531 & n17534;
  assign n17536 = n13700 & ~n17535;
  assign n17537 = ~pi0656 & n7999;
  assign n17538 = ~pi0578 & n8080;
  assign n17539 = ~n17537 & ~n17538;
  assign n17540 = pi1147 & n13676;
  assign n17541 = ~pi1403 & n13678;
  assign n17542 = ~n17540 & ~n17541;
  assign n17543 = n17539 & n17542;
  assign n17544 = n13684 & ~n17543;
  assign n17545 = ~n17536 & ~n17544;
  assign n17546 = pi0263 & n13715;
  assign n17547 = pi0987 & n13712;
  assign n17548 = ~n17546 & ~n17547;
  assign n17549 = ~pi1328 & n13708;
  assign n17550 = n17548 & ~n17549;
  assign n17551 = n13722 & ~n17550;
  assign n17552 = ~pi0342 & n7999;
  assign n17553 = ~pi0378 & n8080;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = pi1262 & n13676;
  assign n17556 = ~pi1393 & n13678;
  assign n17557 = ~n17555 & ~n17556;
  assign n17558 = n17554 & n17557;
  assign n17559 = n13724 & ~n17558;
  assign n17560 = n13733 & ~n17550;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = ~n17551 & n17561;
  assign n17563 = n17545 & n17562;
  assign po1407 = n17528 | ~n17563;
  assign n17565 = ~pi0421 & n7999;
  assign n17566 = ~pi0496 & n8080;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = ~pi1137 & n13676;
  assign n17569 = ~pi1359 & n13678;
  assign n17570 = ~n17568 & ~n17569;
  assign n17571 = n17567 & n17570;
  assign n17572 = n13672 & ~n17571;
  assign n17573 = ~pi0526 & n7999;
  assign n17574 = ~pi0540 & n8080;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = pi1242 & n13676;
  assign n17577 = ~pi1400 & n13678;
  assign n17578 = ~n17576 & ~n17577;
  assign n17579 = n17575 & n17578;
  assign n17580 = n13684 & ~n17579;
  assign n17581 = ~pi0603 & n7999;
  assign n17582 = ~pi0688 & n8080;
  assign n17583 = ~n17581 & ~n17582;
  assign n17584 = pi1118 & n13676;
  assign n17585 = ~pi1381 & n13678;
  assign n17586 = ~n17584 & ~n17585;
  assign n17587 = n17583 & n17586;
  assign n17588 = n13700 & ~n17587;
  assign n17589 = ~n17580 & ~n17588;
  assign n17590 = pi0253 & n13715;
  assign n17591 = pi0915 & n13712;
  assign n17592 = ~n17590 & ~n17591;
  assign n17593 = ~pi1330 & n13708;
  assign n17594 = n17592 & ~n17593;
  assign n17595 = n13722 & ~n17594;
  assign n17596 = ~pi0344 & n7999;
  assign n17597 = ~pi0397 & n8080;
  assign n17598 = ~n17596 & ~n17597;
  assign n17599 = pi1124 & n13676;
  assign n17600 = ~pi1404 & n13678;
  assign n17601 = ~n17599 & ~n17600;
  assign n17602 = n17598 & n17601;
  assign n17603 = n13724 & ~n17602;
  assign n17604 = n13733 & ~n17594;
  assign n17605 = ~n17603 & ~n17604;
  assign n17606 = ~n17595 & n17605;
  assign n17607 = n17589 & n17606;
  assign po1408 = n17572 | ~n17607;
  assign n17609 = ~pi0422 & n7999;
  assign n17610 = ~pi0497 & n8080;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = ~pi1030 & n13676;
  assign n17613 = ~pi1362 & n13678;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = n17611 & n17614;
  assign n17616 = n13672 & ~n17615;
  assign n17617 = ~pi0527 & n7999;
  assign n17618 = ~pi0580 & n8080;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = pi1261 & n13676;
  assign n17621 = ~pi1374 & n13678;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = n17619 & n17622;
  assign n17624 = n13684 & ~n17623;
  assign n17625 = ~pi0544 & n7999;
  assign n17626 = ~pi0667 & n8080;
  assign n17627 = ~n17625 & ~n17626;
  assign n17628 = pi1074 & n13676;
  assign n17629 = ~pi1363 & n13678;
  assign n17630 = ~n17628 & ~n17629;
  assign n17631 = n17627 & n17630;
  assign n17632 = n13700 & ~n17631;
  assign n17633 = ~n17624 & ~n17632;
  assign n17634 = pi0255 & n13715;
  assign n17635 = pi0901 & n13712;
  assign n17636 = ~n17634 & ~n17635;
  assign n17637 = n13722 & ~n17636;
  assign n17638 = n13733 & ~n17636;
  assign n17639 = ~pi0345 & n7999;
  assign n17640 = ~pi0398 & n8080;
  assign n17641 = ~n17639 & ~n17640;
  assign n17642 = pi1252 & n13676;
  assign n17643 = ~pi1383 & n13678;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = n17641 & n17644;
  assign n17646 = n13724 & ~n17645;
  assign n17647 = ~n17638 & ~n17646;
  assign n17648 = ~n17637 & n17647;
  assign n17649 = n17633 & n17648;
  assign po1409 = n17616 | ~n17649;
  assign n17651 = ~pi0432 & n7999;
  assign n17652 = ~pi0498 & n8080;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = ~pi1390 & n13678;
  assign n17655 = pi1080 & n13676;
  assign n17656 = ~n17654 & ~n17655;
  assign n17657 = n17653 & n17656;
  assign n17658 = n13672 & ~n17657;
  assign n17659 = ~pi0629 & n7999;
  assign n17660 = ~pi0579 & n8080;
  assign n17661 = ~n17659 & ~n17660;
  assign n17662 = ~pi1406 & n13678;
  assign n17663 = pi1144 & n13676;
  assign n17664 = ~n17662 & ~n17663;
  assign n17665 = n17661 & n17664;
  assign n17666 = n13684 & ~n17665;
  assign n17667 = ~pi0606 & n7999;
  assign n17668 = ~pi0690 & n8080;
  assign n17669 = ~n17667 & ~n17668;
  assign n17670 = pi1112 & n13676;
  assign n17671 = ~pi1382 & n13678;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = n17669 & n17672;
  assign n17674 = n13700 & ~n17673;
  assign n17675 = ~n17666 & ~n17674;
  assign n17676 = pi0250 & n13715;
  assign n17677 = pi0728 & n13712;
  assign n17678 = ~n17676 & ~n17677;
  assign n17679 = n13722 & ~n17678;
  assign n17680 = n13733 & ~n17678;
  assign n17681 = ~pi0346 & n7999;
  assign n17682 = ~pi0401 & n8080;
  assign n17683 = ~n17681 & ~n17682;
  assign n17684 = ~pi1384 & n13678;
  assign n17685 = pi1256 & n13676;
  assign n17686 = ~n17684 & ~n17685;
  assign n17687 = n17683 & n17686;
  assign n17688 = n13724 & ~n17687;
  assign n17689 = ~n17680 & ~n17688;
  assign n17690 = ~n17679 & n17689;
  assign n17691 = n17675 & n17690;
  assign po1410 = n17658 | ~n17691;
  assign n17693 = ~pi0350 & n7999;
  assign n17694 = ~pi0406 & n8080;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = ~pi1349 & n13678;
  assign n17697 = pi0939 & n13676;
  assign n17698 = ~n17696 & ~n17697;
  assign n17699 = n17695 & n17698;
  assign n17700 = n13672 & ~n17699;
  assign n17701 = ~pi0515 & n7999;
  assign n17702 = ~pi0651 & n8080;
  assign n17703 = ~n17701 & ~n17702;
  assign n17704 = ~pi1353 & n13678;
  assign n17705 = pi0994 & n13676;
  assign n17706 = ~n17704 & ~n17705;
  assign n17707 = n17703 & n17706;
  assign n17708 = n13700 & ~n17707;
  assign n17709 = ~pi1407 & n13678;
  assign n17710 = pi0969 & n13676;
  assign n17711 = ~n17709 & ~n17710;
  assign n17712 = ~pi0427 & n7999;
  assign n17713 = ~pi0504 & n8080;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = n17711 & n17714;
  assign n17716 = n13684 & ~n17715;
  assign n17717 = ~n17708 & ~n17716;
  assign n17718 = pi0186 & n13715;
  assign n17719 = pi0977 & n13712;
  assign n17720 = ~n17718 & ~n17719;
  assign n17721 = n13722 & ~n17720;
  assign n17722 = n13733 & ~n17720;
  assign n17723 = ~pi0311 & n7999;
  assign n17724 = ~pi0334 & n8080;
  assign n17725 = ~n17723 & ~n17724;
  assign n17726 = ~pi1396 & n13678;
  assign n17727 = pi0863 & n13676;
  assign n17728 = ~n17726 & ~n17727;
  assign n17729 = n17725 & n17728;
  assign n17730 = n13724 & ~n17729;
  assign n17731 = ~n17722 & ~n17730;
  assign n17732 = ~n17721 & n17731;
  assign n17733 = n17717 & n17732;
  assign po1411 = n17700 | ~n17733;
  assign n17735 = ~pi0548 & n7999;
  assign n17736 = ~pi0376 & n8080;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = pi1028 & n13676;
  assign n17739 = pi0131 & n13678;
  assign n17740 = ~n17738 & ~n17739;
  assign n17741 = n17737 & n17740;
  assign n17742 = n13672 & ~n17741;
  assign n17743 = ~pi0640 & n7999;
  assign n17744 = ~pi0463 & n8080;
  assign n17745 = ~n17743 & ~n17744;
  assign n17746 = pi1258 & n13676;
  assign n17747 = pi0128 & n13678;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = n17745 & n17748;
  assign n17750 = n13684 & ~n17749;
  assign n17751 = ~pi0547 & n7999;
  assign n17752 = ~pi0628 & n8080;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = pi1107 & n13676;
  assign n17755 = pi0129 & n13678;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = n17753 & n17756;
  assign n17758 = n13700 & ~n17757;
  assign n17759 = ~n17750 & ~n17758;
  assign n17760 = pi1681 & n13710;
  assign n17761 = pi1068 & n13705;
  assign n17762 = ~n17760 & ~n17761;
  assign n17763 = pi0477 & n13715;
  assign n17764 = pi1321 & n13708;
  assign n17765 = ~n17763 & ~n17764;
  assign n17766 = n17762 & n17765;
  assign n17767 = n13722 & ~n17766;
  assign n17768 = ~pi0447 & n7999;
  assign n17769 = ~pi0329 & n8080;
  assign n17770 = ~n17768 & ~n17769;
  assign n17771 = pi1272 & n13676;
  assign n17772 = pi0130 & n13678;
  assign n17773 = ~n17771 & ~n17772;
  assign n17774 = n17770 & n17773;
  assign n17775 = n13724 & ~n17774;
  assign n17776 = n13733 & ~n17766;
  assign n17777 = ~n17775 & ~n17776;
  assign n17778 = ~n17767 & n17777;
  assign n17779 = n17759 & n17778;
  assign po1412 = n17742 | ~n17779;
  assign n17781 = ~pi0362 & n7999;
  assign n17782 = ~pi0357 & n8080;
  assign n17783 = ~n17781 & ~n17782;
  assign n17784 = pi1083 & n13676;
  assign n17785 = pi0990 & n13678;
  assign n17786 = ~n17784 & ~n17785;
  assign n17787 = n17783 & n17786;
  assign n17788 = n13672 & ~n17787;
  assign n17789 = ~pi0449 & n7999;
  assign n17790 = ~pi0461 & n8080;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = pi1033 & n13676;
  assign n17793 = pi1048 & n13678;
  assign n17794 = ~n17792 & ~n17793;
  assign n17795 = n17791 & n17794;
  assign n17796 = n13684 & ~n17795;
  assign n17797 = ~pi0550 & n7999;
  assign n17798 = ~pi0633 & n8080;
  assign n17799 = ~n17797 & ~n17798;
  assign n17800 = pi1108 & n13676;
  assign n17801 = pi1314 & n13678;
  assign n17802 = ~n17800 & ~n17801;
  assign n17803 = n17799 & n17802;
  assign n17804 = n13700 & ~n17803;
  assign n17805 = ~n17796 & ~n17804;
  assign n17806 = pi1098 & n13705;
  assign n17807 = pi1693 & n13710;
  assign n17808 = ~n17806 & ~n17807;
  assign n17809 = pi0448 & n13715;
  assign n17810 = pi1322 & n13708;
  assign n17811 = ~n17809 & ~n17810;
  assign n17812 = n17808 & n17811;
  assign n17813 = n13722 & ~n17812;
  assign n17814 = ~pi0321 & n7999;
  assign n17815 = ~pi0327 & n8080;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = pi1121 & n13676;
  assign n17818 = pi0965 & n13678;
  assign n17819 = ~n17817 & ~n17818;
  assign n17820 = n17816 & n17819;
  assign n17821 = n13724 & ~n17820;
  assign n17822 = n13733 & ~n17812;
  assign n17823 = ~n17821 & ~n17822;
  assign n17824 = ~n17813 & n17823;
  assign n17825 = n17805 & n17824;
  assign po1413 = n17788 | ~n17825;
  assign n17827 = ~pi1305 & ~n9550;
  assign n17828 = pi1747 & ~n17827;
  assign po1414 = n11428 | ~n17828;
  assign n17830 = ~n15428 & ~n15432;
  assign n17831 = ~n15427 & n15436;
  assign n17832 = n17830 & n17831;
  assign n17833 = ~n17830 & ~n17831;
  assign po1415 = n17832 | n17833;
  assign n17835 = ~n15476 & ~n15480;
  assign n17836 = ~n15475 & n15484;
  assign n17837 = n17835 & n17836;
  assign n17838 = ~n17835 & ~n17836;
  assign po1416 = n17837 | n17838;
  assign n17840 = ~n15524 & ~n15528;
  assign n17841 = ~n15523 & n15532;
  assign n17842 = n17840 & n17841;
  assign n17843 = ~n17840 & ~n17841;
  assign po1417 = n17842 | n17843;
  assign n17845 = ~n15572 & ~n15576;
  assign n17846 = ~n15571 & n15580;
  assign n17847 = n17845 & n17846;
  assign n17848 = ~n17845 & ~n17846;
  assign po1418 = n17847 | n17848;
  assign n17850 = pi1777 & n16136;
  assign n17851 = pi1310 & ~n16136;
  assign n17852 = ~n17850 & ~n17851;
  assign po1419 = pi1747 & ~n17852;
  assign n17854 = ~pi1311 & ~n9550;
  assign n17855 = pi1747 & ~n17854;
  assign po1420 = n10932 | ~n17855;
  assign n17857 = ~pi1312 & ~n9550;
  assign n17858 = pi1747 & ~n17857;
  assign po1421 = n10922 | ~n17858;
  assign n17860 = pi1313 & ~po1535;
  assign n17861 = ~pi1733 & po1535;
  assign po1422 = n17860 | n17861;
  assign n17863 = ~pi1314 & ~n11728;
  assign po1423 = n6189 & ~n17863;
  assign n17865 = ~pi1316 & ~n9550;
  assign n17866 = pi1747 & ~n17865;
  assign po1425 = n10841 | ~n17866;
  assign n17868 = pi1317 & ~po1535;
  assign n17869 = ~pi1741 & po1535;
  assign po1426 = n17868 | n17869;
  assign n17871 = pi1318 & ~po1535;
  assign n17872 = ~pi1722 & po1535;
  assign po1427 = n17871 | n17872;
  assign n17874 = pi1775 & n17285;
  assign n17875 = pi1319 & ~n17285;
  assign n17876 = ~n17874 & ~n17875;
  assign po1428 = pi1747 & ~n17876;
  assign n17878 = pi1777 & n17285;
  assign n17879 = pi1320 & ~n17285;
  assign n17880 = ~n17878 & ~n17879;
  assign po1429 = pi1747 & ~n17880;
  assign n17882 = pi1779 & n17285;
  assign n17883 = pi1321 & ~n17285;
  assign n17884 = ~n17882 & ~n17883;
  assign po1430 = pi1747 & ~n17884;
  assign n17886 = pi1780 & n17285;
  assign n17887 = pi1322 & ~n17285;
  assign n17888 = ~n17886 & ~n17887;
  assign po1431 = pi1747 & ~n17888;
  assign n17890 = pi1781 & n17285;
  assign n17891 = ~pi1323 & ~n17285;
  assign n17892 = ~n17890 & ~n17891;
  assign po1432 = pi1747 & ~n17892;
  assign n17894 = pi1790 & n17285;
  assign n17895 = ~pi1324 & ~n17285;
  assign n17896 = ~n17894 & ~n17895;
  assign po1433 = pi1747 & ~n17896;
  assign n17898 = pi1791 & n17285;
  assign n17899 = ~pi1325 & ~n17285;
  assign n17900 = ~n17898 & ~n17899;
  assign po1434 = pi1747 & ~n17900;
  assign n17902 = pi1792 & n17285;
  assign n17903 = ~pi1326 & ~n17285;
  assign n17904 = ~n17902 & ~n17903;
  assign po1435 = pi1747 & ~n17904;
  assign n17906 = pi1794 & n17285;
  assign n17907 = ~pi1327 & ~n17285;
  assign n17908 = ~n17906 & ~n17907;
  assign po1436 = pi1747 & ~n17908;
  assign n17910 = pi1795 & n17285;
  assign n17911 = ~pi1328 & ~n17285;
  assign n17912 = ~n17910 & ~n17911;
  assign po1437 = pi1747 & ~n17912;
  assign n17914 = pi1796 & n17285;
  assign n17915 = ~pi1329 & ~n17285;
  assign n17916 = ~n17914 & ~n17915;
  assign po1438 = pi1747 & ~n17916;
  assign n17918 = pi1798 & n17285;
  assign n17919 = ~pi1330 & ~n17285;
  assign n17920 = ~n17918 & ~n17919;
  assign po1439 = pi1747 & ~n17920;
  assign n17922 = pi1331 & ~n9550;
  assign n17923 = pi1747 & ~n17922;
  assign po1440 = n11448 | ~n17923;
  assign n17925 = ~pi1332 & ~n9550;
  assign n17926 = pi1747 & ~n17925;
  assign po1441 = n10952 | ~n17926;
  assign n17928 = ~pi1333 & ~n9550;
  assign n17929 = pi1747 & ~n17928;
  assign po1442 = n10962 | ~n17929;
  assign n17931 = pi1334 & ~po1535;
  assign n17932 = ~pi1727 & po1535;
  assign po1443 = n17931 | n17932;
  assign n17934 = pi1335 & ~po1535;
  assign n17935 = ~pi1740 & po1535;
  assign po1444 = n17934 | n17935;
  assign n17937 = pi1336 & ~po1535;
  assign n17938 = ~pi1735 & po1535;
  assign po1445 = n17937 | n17938;
  assign n17940 = pi1337 & ~po1535;
  assign n17941 = ~pi1725 & po1535;
  assign po1446 = n17940 | n17941;
  assign n17943 = pi1777 & n16241;
  assign n17944 = pi1338 & ~n16241;
  assign n17945 = ~n17943 & ~n17944;
  assign po1447 = pi1747 & ~n17945;
  assign n17947 = pi1797 & n17285;
  assign n17948 = ~pi1339 & ~n17285;
  assign n17949 = ~n17947 & ~n17948;
  assign po1448 = pi1747 & ~n17949;
  assign n17951 = ~n15447 & ~n15795;
  assign n17952 = ~n15477 & n17951;
  assign n17953 = ~n15458 & n15814;
  assign n17954 = n15801 & ~n17953;
  assign n17955 = n15802 & n15805;
  assign n17956 = ~n17954 & n17955;
  assign n17957 = ~n15799 & n15805;
  assign n17958 = ~n17956 & ~n17957;
  assign n17959 = n15797 & n17958;
  assign n17960 = ~n15447 & ~n17959;
  assign n17961 = n15808 & n17960;
  assign n17962 = ~n15477 & n17961;
  assign n17963 = ~pi1177 & ~n15489;
  assign n17964 = ~n15446 & n15447;
  assign n17965 = pi0481 & ~n15489;
  assign n17966 = ~n17964 & ~n17965;
  assign n17967 = ~n17963 & n17966;
  assign n17968 = ~n17962 & ~n17967;
  assign n17969 = ~n17952 & n17968;
  assign n17970 = pi0383 & ~pi1179;
  assign n17971 = ~pi0383 & pi1179;
  assign n17972 = ~n17970 & ~n17971;
  assign n17973 = ~n17969 & ~n17972;
  assign n17974 = n17969 & n17972;
  assign po1449 = n17973 | n17974;
  assign n17976 = pi0471 & ~pi1036;
  assign n17977 = ~pi0471 & pi1036;
  assign n17978 = ~n17976 & ~n17977;
  assign n17979 = ~n15506 & n15845;
  assign n17980 = n15832 & ~n17979;
  assign n17981 = n15833 & n15836;
  assign n17982 = ~n17980 & n17981;
  assign n17983 = ~n15830 & n15836;
  assign n17984 = ~n17982 & ~n17983;
  assign n17985 = n15828 & n17984;
  assign n17986 = ~n15495 & ~n17985;
  assign n17987 = n15839 & n17986;
  assign n17988 = ~n15525 & n17987;
  assign n17989 = ~pi1201 & ~n15537;
  assign n17990 = ~n15494 & n15495;
  assign n17991 = ~n17989 & ~n17990;
  assign n17992 = pi0564 & ~n15537;
  assign n17993 = n17991 & ~n17992;
  assign n17994 = ~n15495 & ~n15525;
  assign n17995 = ~n15826 & n17994;
  assign n17996 = ~n17993 & ~n17995;
  assign n17997 = ~n17988 & n17996;
  assign n17998 = ~n17978 & ~n17997;
  assign n17999 = n17978 & n17997;
  assign po1450 = n17998 | n17999;
  assign n18001 = pi1777 & n16153;
  assign n18002 = pi1342 & ~n16153;
  assign n18003 = ~n18001 & ~n18002;
  assign po1451 = pi1747 & ~n18003;
  assign n18005 = ~pi1343 & ~n9550;
  assign n18006 = pi1747 & ~n18005;
  assign po1452 = n10831 | ~n18006;
  assign n18008 = ~pi1344 & ~n9550;
  assign n18009 = pi1747 & ~n18008;
  assign po1453 = n11538 | ~n18009;
  assign n18011 = pi1345 & pi1495;
  assign n18012 = ~pi1479 & po1776;
  assign po1603 = n15161 | n18012;
  assign n18014 = ~pi1345 & ~pi1495;
  assign n18015 = po1603 & ~n18014;
  assign n18016 = ~n18011 & ~n18015;
  assign po1454 = pi1747 & ~n18016;
  assign n18018 = pi1346 & ~n9550;
  assign n18019 = pi1747 & ~n18018;
  assign po1455 = n11518 | ~n18019;
  assign n18021 = n9549 & n13678;
  assign n18022 = ~pi1347 & ~n18021;
  assign n18023 = pi1795 & n18021;
  assign n18024 = ~n18022 & ~n18023;
  assign po1456 = pi1747 & ~n18024;
  assign n18026 = ~pi1348 & ~n18021;
  assign n18027 = pi1801 & n18021;
  assign n18028 = ~n18026 & ~n18027;
  assign po1457 = pi1747 & ~n18028;
  assign n18030 = n8355 & n13678;
  assign n18031 = ~pi1349 & ~n18030;
  assign n18032 = pi1802 & n18030;
  assign n18033 = ~n18031 & ~n18032;
  assign po1458 = pi1747 & ~n18033;
  assign n18035 = ~pi1350 & ~n18021;
  assign n18036 = pi1792 & n18021;
  assign n18037 = ~n18035 & ~n18036;
  assign po1459 = pi1747 & ~n18037;
  assign n18039 = ~pi1351 & ~n18021;
  assign n18040 = pi1794 & n18021;
  assign n18041 = ~n18039 & ~n18040;
  assign po1460 = pi1747 & ~n18041;
  assign n18043 = ~pi1352 & ~n18030;
  assign n18044 = pi1803 & n18030;
  assign n18045 = ~n18043 & ~n18044;
  assign po1461 = pi1747 & ~n18045;
  assign n18047 = ~pi1353 & ~n18021;
  assign n18048 = pi1802 & n18021;
  assign n18049 = ~n18047 & ~n18048;
  assign po1462 = pi1747 & ~n18049;
  assign n18051 = ~pi1354 & ~n18021;
  assign n18052 = pi1793 & n18021;
  assign n18053 = ~n18051 & ~n18052;
  assign po1463 = pi1747 & ~n18053;
  assign n18055 = ~pi1355 & ~n18021;
  assign n18056 = pi1791 & n18021;
  assign n18057 = ~n18055 & ~n18056;
  assign po1464 = pi1747 & ~n18057;
  assign n18059 = ~pi1356 & ~n18021;
  assign n18060 = pi1803 & n18021;
  assign n18061 = ~n18059 & ~n18060;
  assign po1465 = pi1747 & ~n18061;
  assign n18063 = ~pi1357 & ~n18021;
  assign n18064 = pi1790 & n18021;
  assign n18065 = ~n18063 & ~n18064;
  assign po1466 = pi1747 & ~n18065;
  assign n18067 = pi0103 & n5524;
  assign po1467 = n5858 | n18067;
  assign n18069 = ~pi1359 & ~n18030;
  assign n18070 = pi1798 & n18030;
  assign n18071 = ~n18069 & ~n18070;
  assign po1468 = pi1747 & ~n18071;
  assign n18073 = pi1360 & ~n16897;
  assign n18074 = n16896 & ~n18073;
  assign n18075 = pi1747 & pi1796;
  assign n18076 = n16115 & n18075;
  assign po1469 = n18074 | n18076;
  assign n18078 = pi1361 & ~n16833;
  assign n18079 = n16832 & ~n18078;
  assign n18080 = n16241 & n18075;
  assign po1470 = n18079 | n18080;
  assign n18082 = ~pi1362 & ~n18030;
  assign n18083 = pi1799 & n18030;
  assign n18084 = ~n18082 & ~n18083;
  assign po1471 = pi1747 & ~n18084;
  assign n18086 = ~pi1363 & ~n18021;
  assign n18087 = pi1799 & n18021;
  assign n18088 = ~n18086 & ~n18087;
  assign po1472 = pi1747 & ~n18088;
  assign n18090 = ~pi1364 & ~n18030;
  assign n18091 = pi1801 & n18030;
  assign n18092 = ~n18090 & ~n18091;
  assign po1473 = pi1747 & ~n18092;
  assign n18094 = ~pi0542 & n7999;
  assign n18095 = ~pi0704 & n8080;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = ~pi1356 & n13678;
  assign n18098 = pi1014 & n13676;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = n18096 & n18099;
  assign n18101 = n13700 & ~n18100;
  assign n18102 = ~n13722 & ~n13733;
  assign n18103 = n13715 & ~n18102;
  assign n18104 = pi0153 & n18103;
  assign n18105 = ~n18101 & ~n18104;
  assign n18106 = ~pi0616 & n7999;
  assign n18107 = ~pi0501 & n8080;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~pi1352 & n13678;
  assign n18110 = pi0942 & n13676;
  assign n18111 = ~n18109 & ~n18110;
  assign n18112 = n18108 & n18111;
  assign n18113 = n13672 & ~n18112;
  assign n18114 = ~pi0528 & n7999;
  assign n18115 = ~pi0581 & n8080;
  assign n18116 = ~n18114 & ~n18115;
  assign n18117 = pi0973 & n13676;
  assign n18118 = ~pi1376 & n13678;
  assign n18119 = ~n18117 & ~n18118;
  assign n18120 = n18116 & n18119;
  assign n18121 = n13684 & ~n18120;
  assign n18122 = ~n18113 & ~n18121;
  assign n18123 = ~pi0519 & n7999;
  assign n18124 = ~pi0377 & n8080;
  assign n18125 = ~n18123 & ~n18124;
  assign n18126 = ~pi1386 & n13678;
  assign n18127 = pi0876 & n13676;
  assign n18128 = ~n18126 & ~n18127;
  assign n18129 = n18125 & n18128;
  assign n18130 = n13724 & ~n18129;
  assign n18131 = n18122 & ~n18130;
  assign po1474 = ~n18105 | ~n18131;
  assign n18133 = pi0938 & n13676;
  assign n18134 = ~pi0424 & n7999;
  assign n18135 = ~pi0500 & n8080;
  assign n18136 = ~n18134 & ~n18135;
  assign n18137 = ~n18133 & n18136;
  assign n18138 = n13672 & ~n18137;
  assign n18139 = pi0861 & n13676;
  assign n18140 = ~pi0347 & n7999;
  assign n18141 = ~pi0403 & n8080;
  assign n18142 = ~n18140 & ~n18141;
  assign n18143 = ~n18139 & n18142;
  assign n18144 = n13724 & ~n18143;
  assign n18145 = pi0967 & n13676;
  assign n18146 = ~pi0530 & n7999;
  assign n18147 = ~pi0583 & n8080;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = ~n18145 & n18148;
  assign n18150 = n13684 & ~n18149;
  assign n18151 = ~n18144 & ~n18150;
  assign n18152 = pi0992 & n13676;
  assign n18153 = ~pi0608 & n7999;
  assign n18154 = ~pi0691 & n8080;
  assign n18155 = ~n18153 & ~n18154;
  assign n18156 = ~n18152 & n18155;
  assign n18157 = n13700 & ~n18156;
  assign n18158 = pi0195 & n18103;
  assign n18159 = ~n18157 & ~n18158;
  assign n18160 = n18151 & n18159;
  assign po1475 = n18138 | ~n18160;
  assign n18162 = pi0941 & n13676;
  assign n18163 = ~pi0351 & n7999;
  assign n18164 = ~pi0407 & n8080;
  assign n18165 = ~n18163 & ~n18164;
  assign n18166 = ~n18162 & n18165;
  assign n18167 = n13672 & ~n18166;
  assign n18168 = pi0862 & n13676;
  assign n18169 = ~pi0312 & n7999;
  assign n18170 = ~pi0335 & n8080;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = ~n18168 & n18171;
  assign n18173 = n13724 & ~n18172;
  assign n18174 = pi0968 & n13676;
  assign n18175 = ~pi0428 & n7999;
  assign n18176 = ~pi0505 & n8080;
  assign n18177 = ~n18175 & ~n18176;
  assign n18178 = ~n18174 & n18177;
  assign n18179 = n13684 & ~n18178;
  assign n18180 = ~n18173 & ~n18179;
  assign n18181 = pi0993 & n13676;
  assign n18182 = ~pi0437 & n7999;
  assign n18183 = ~pi0652 & n8080;
  assign n18184 = ~n18182 & ~n18183;
  assign n18185 = ~n18181 & n18184;
  assign n18186 = n13700 & ~n18185;
  assign n18187 = pi0185 & n18103;
  assign n18188 = ~n18186 & ~n18187;
  assign n18189 = n18180 & n18188;
  assign po1476 = n18167 | ~n18189;
  assign n18191 = ~pi0658 & n7999;
  assign n18192 = ~pi0539 & n8080;
  assign n18193 = ~n18191 & ~n18192;
  assign n18194 = ~pi1375 & n13678;
  assign n18195 = pi1259 & n13676;
  assign n18196 = ~n18194 & ~n18195;
  assign n18197 = n18193 & n18196;
  assign n18198 = n13684 & ~n18197;
  assign n18199 = ~pi0423 & n7999;
  assign n18200 = ~pi0445 & n8080;
  assign n18201 = ~n18199 & ~n18200;
  assign n18202 = pi1132 & n13676;
  assign n18203 = ~pi1364 & n13678;
  assign n18204 = ~n18202 & ~n18203;
  assign n18205 = n18201 & n18204;
  assign n18206 = n13672 & ~n18205;
  assign n18207 = ~n18198 & ~n18206;
  assign n18208 = ~pi0605 & n7999;
  assign n18209 = ~pi0689 & n8080;
  assign n18210 = ~n18208 & ~n18209;
  assign n18211 = ~pi1348 & n13678;
  assign n18212 = pi1113 & n13676;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n18210 & n18213;
  assign n18215 = n13700 & ~n18214;
  assign n18216 = pi0986 & n13712;
  assign n18217 = ~n18102 & n18216;
  assign n18218 = ~n18215 & ~n18217;
  assign n18219 = ~pi0314 & n7999;
  assign n18220 = ~pi0400 & n8080;
  assign n18221 = ~n18219 & ~n18220;
  assign n18222 = ~pi1385 & n13678;
  assign n18223 = pi1257 & n13676;
  assign n18224 = ~n18222 & ~n18223;
  assign n18225 = n18221 & n18224;
  assign n18226 = n13724 & ~n18225;
  assign n18227 = n18218 & ~n18226;
  assign po1477 = ~n18207 | ~n18227;
  assign n18229 = pi1369 & ~n16966;
  assign n18230 = n16965 & ~n18229;
  assign n18231 = n16136 & n18075;
  assign po1478 = n18230 | n18231;
  assign n18233 = ~n7987 & n16511;
  assign n18234 = pi1370 & n18233;
  assign n18235 = ~pi0138 & pi1370;
  assign n18236 = ~n12119 & ~n18235;
  assign n18237 = n3724 & ~n18236;
  assign n18238 = ~n18234 & ~n18237;
  assign po1479 = pi1747 & ~n18238;
  assign n18240 = pi1139 & n13676;
  assign n18241 = ~pi0451 & n7999;
  assign n18242 = ~pi0456 & n8080;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~n18240 & n18243;
  assign n18245 = n13684 & ~n18244;
  assign n18246 = pi1127 & n13676;
  assign n18247 = ~pi0364 & n7999;
  assign n18248 = ~pi0369 & n8080;
  assign n18249 = ~n18247 & ~n18248;
  assign n18250 = ~n18246 & n18249;
  assign n18251 = n13672 & ~n18250;
  assign n18252 = pi1119 & n13676;
  assign n18253 = ~pi0316 & n7999;
  assign n18254 = ~pi0322 & n8080;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = ~n18252 & n18255;
  assign n18257 = n13724 & ~n18256;
  assign n18258 = ~n18251 & ~n18257;
  assign n18259 = pi1102 & n13676;
  assign n18260 = ~pi0551 & n7999;
  assign n18261 = ~pi0636 & n8080;
  assign n18262 = ~n18260 & ~n18261;
  assign n18263 = ~n18259 & n18262;
  assign n18264 = n13700 & ~n18263;
  assign n18265 = pi0473 & n13715;
  assign n18266 = ~n18102 & n18265;
  assign n18267 = ~n18264 & ~n18266;
  assign n18268 = n18258 & n18267;
  assign po1480 = n18245 | ~n18268;
  assign n18270 = ~pi0450 & n7999;
  assign n18271 = ~pi0460 & n8080;
  assign n18272 = ~n18270 & ~n18271;
  assign n18273 = ~pi1273 & n13676;
  assign n18274 = n18272 & ~n18273;
  assign n18275 = n13684 & ~n18274;
  assign n18276 = ~pi1128 & n13676;
  assign n18277 = ~pi0367 & n7999;
  assign n18278 = ~pi0372 & n8080;
  assign n18279 = ~n18277 & ~n18278;
  assign n18280 = ~n18276 & n18279;
  assign n18281 = n13672 & ~n18280;
  assign n18282 = ~pi0319 & n7999;
  assign n18283 = ~pi0325 & n8080;
  assign n18284 = ~n18282 & ~n18283;
  assign n18285 = ~pi1268 & n13676;
  assign n18286 = n18284 & ~n18285;
  assign n18287 = n13724 & ~n18286;
  assign n18288 = ~n18281 & ~n18287;
  assign n18289 = ~pi1243 & n13676;
  assign n18290 = ~pi0555 & n7999;
  assign n18291 = ~pi0638 & n8080;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~n18289 & n18292;
  assign n18294 = n13700 & ~n18293;
  assign n18295 = ~pi0465 & n13715;
  assign n18296 = ~n18102 & n18295;
  assign n18297 = ~n18294 & ~n18296;
  assign n18298 = n18288 & n18297;
  assign po1481 = n18275 | ~n18298;
  assign n18300 = ~pi0659 & n7999;
  assign n18301 = ~pi0585 & n8080;
  assign n18302 = ~n18300 & ~n18301;
  assign n18303 = pi1034 & n13676;
  assign n18304 = n18302 & ~n18303;
  assign n18305 = n13684 & ~n18304;
  assign n18306 = pi1029 & n13676;
  assign n18307 = ~pi0426 & n7999;
  assign n18308 = ~pi0443 & n8080;
  assign n18309 = ~n18307 & ~n18308;
  assign n18310 = ~n18306 & n18309;
  assign n18311 = n13672 & ~n18310;
  assign n18312 = ~pi0313 & n7999;
  assign n18313 = ~pi0405 & n8080;
  assign n18314 = ~n18312 & ~n18313;
  assign n18315 = pi1267 & n13676;
  assign n18316 = n18314 & ~n18315;
  assign n18317 = n13724 & ~n18316;
  assign n18318 = ~n18311 & ~n18317;
  assign n18319 = pi1110 & n13676;
  assign n18320 = ~pi0611 & n7999;
  assign n18321 = ~pi0693 & n8080;
  assign n18322 = ~n18320 & ~n18321;
  assign n18323 = ~n18319 & n18322;
  assign n18324 = n13700 & ~n18323;
  assign n18325 = pi0478 & n13715;
  assign n18326 = ~n18102 & n18325;
  assign n18327 = ~n18324 & ~n18326;
  assign n18328 = n18318 & n18327;
  assign po1482 = n18305 | ~n18328;
  assign n18330 = n9429 & n13678;
  assign n18331 = ~pi1374 & ~n18330;
  assign n18332 = pi1799 & n18330;
  assign n18333 = ~n18331 & ~n18332;
  assign po1483 = pi1747 & ~n18333;
  assign n18335 = ~pi1375 & ~n18330;
  assign n18336 = pi1801 & n18330;
  assign n18337 = ~n18335 & ~n18336;
  assign po1484 = pi1747 & ~n18337;
  assign n18339 = ~pi1376 & ~n18330;
  assign n18340 = pi1803 & n18330;
  assign n18341 = ~n18339 & ~n18340;
  assign po1485 = pi1747 & ~n18341;
  assign n18343 = ~pi1377 & ~n18330;
  assign n18344 = pi1790 & n18330;
  assign n18345 = ~n18343 & ~n18344;
  assign po1486 = pi1747 & ~n18345;
  assign n18347 = ~pi1378 & ~n18330;
  assign n18348 = pi1791 & n18330;
  assign n18349 = ~n18347 & ~n18348;
  assign po1487 = pi1747 & ~n18349;
  assign n18351 = ~pi1379 & ~n18330;
  assign n18352 = pi1794 & n18330;
  assign n18353 = ~n18351 & ~n18352;
  assign po1488 = pi1747 & ~n18353;
  assign n18355 = ~pi1380 & ~n18330;
  assign n18356 = pi1793 & n18330;
  assign n18357 = ~n18355 & ~n18356;
  assign po1489 = pi1747 & ~n18357;
  assign n18359 = ~pi1381 & ~n18021;
  assign n18360 = pi1798 & n18021;
  assign n18361 = ~n18359 & ~n18360;
  assign po1490 = pi1747 & ~n18361;
  assign n18363 = ~pi1382 & ~n18021;
  assign n18364 = pi1800 & n18021;
  assign n18365 = ~n18363 & ~n18364;
  assign po1491 = pi1747 & ~n18365;
  assign n18367 = n8006 & n13678;
  assign n18368 = ~pi1383 & ~n18367;
  assign n18369 = pi1799 & n18367;
  assign n18370 = ~n18368 & ~n18369;
  assign po1492 = pi1747 & ~n18370;
  assign n18372 = ~pi1384 & ~n18367;
  assign n18373 = pi1800 & n18367;
  assign n18374 = ~n18372 & ~n18373;
  assign po1493 = pi1747 & ~n18374;
  assign n18376 = ~pi1385 & ~n18367;
  assign n18377 = pi1801 & n18367;
  assign n18378 = ~n18376 & ~n18377;
  assign po1494 = pi1747 & ~n18378;
  assign n18380 = ~pi1386 & ~n18367;
  assign n18381 = pi1803 & n18367;
  assign n18382 = ~n18380 & ~n18381;
  assign po1495 = pi1747 & ~n18382;
  assign n18384 = ~pi1387 & ~n18367;
  assign n18385 = pi1791 & n18367;
  assign n18386 = ~n18384 & ~n18385;
  assign po1496 = pi1747 & ~n18386;
  assign n18388 = ~pi1388 & ~n18367;
  assign n18389 = pi1794 & n18367;
  assign n18390 = ~n18388 & ~n18389;
  assign po1497 = pi1747 & ~n18390;
  assign n18392 = ~pi1389 & ~n18367;
  assign n18393 = pi1793 & n18367;
  assign n18394 = ~n18392 & ~n18393;
  assign po1498 = pi1747 & ~n18394;
  assign n18396 = ~pi1390 & ~n18030;
  assign n18397 = pi1800 & n18030;
  assign n18398 = ~n18396 & ~n18397;
  assign po1499 = pi1747 & ~n18398;
  assign n18400 = ~pi1391 & ~n18030;
  assign n18401 = pi1794 & n18030;
  assign n18402 = ~n18400 & ~n18401;
  assign po1500 = pi1747 & ~n18402;
  assign n18404 = ~pi1084 & n13676;
  assign n18405 = ~pi0613 & n7999;
  assign n18406 = ~pi0488 & n8080;
  assign n18407 = ~n18405 & ~n18406;
  assign n18408 = ~n18404 & n18407;
  assign n18409 = n13672 & ~n18408;
  assign n18410 = ~pi1103 & n13676;
  assign n18411 = ~pi0601 & n7999;
  assign n18412 = ~pi0680 & n8080;
  assign n18413 = ~n18411 & ~n18412;
  assign n18414 = ~n18410 & n18413;
  assign n18415 = n13700 & ~n18414;
  assign n18416 = ~pi1120 & n13676;
  assign n18417 = ~pi0516 & n7999;
  assign n18418 = ~pi0390 & n8080;
  assign n18419 = ~n18417 & ~n18418;
  assign n18420 = ~n18416 & n18419;
  assign n18421 = n13724 & ~n18420;
  assign n18422 = ~pi1140 & n13676;
  assign n18423 = ~pi0439 & n7999;
  assign n18424 = ~pi0571 & n8080;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = ~n18422 & n18425;
  assign n18427 = n13684 & ~n18426;
  assign n18428 = ~n18421 & ~n18427;
  assign n18429 = ~n18415 & n18428;
  assign po1501 = n18409 | ~n18429;
  assign n18431 = ~pi1393 & ~n18367;
  assign n18432 = pi1795 & n18367;
  assign n18433 = ~n18431 & ~n18432;
  assign po1502 = pi1747 & ~n18433;
  assign n18435 = ~pi1394 & ~n18030;
  assign n18436 = pi1790 & n18030;
  assign n18437 = ~n18435 & ~n18436;
  assign po1503 = pi1747 & ~n18437;
  assign n18439 = ~pi1395 & ~n18367;
  assign n18440 = pi1792 & n18367;
  assign n18441 = ~n18439 & ~n18440;
  assign po1504 = pi1747 & ~n18441;
  assign n18443 = ~pi1396 & ~n18367;
  assign n18444 = pi1802 & n18367;
  assign n18445 = ~n18443 & ~n18444;
  assign po1505 = pi1747 & ~n18445;
  assign n18447 = ~pi1397 & ~n18367;
  assign n18448 = pi1790 & n18367;
  assign n18449 = ~n18447 & ~n18448;
  assign po1506 = pi1747 & ~n18449;
  assign n18451 = pi0674 & ~pi1160;
  assign n18452 = ~pi0674 & pi1160;
  assign n18453 = ~n18451 & ~n18452;
  assign n18454 = ~n15410 & n15783;
  assign n18455 = n15770 & ~n18454;
  assign n18456 = n15771 & n15774;
  assign n18457 = ~n18455 & n18456;
  assign n18458 = ~n15768 & n15774;
  assign n18459 = ~n18457 & ~n18458;
  assign n18460 = n15766 & n18459;
  assign n18461 = ~n15399 & ~n18460;
  assign n18462 = n15777 & n18461;
  assign n18463 = ~n15429 & n18462;
  assign n18464 = ~pi1269 & ~n15441;
  assign n18465 = ~n15398 & n15399;
  assign n18466 = ~n18464 & ~n18465;
  assign n18467 = pi0715 & ~n15441;
  assign n18468 = n18466 & ~n18467;
  assign n18469 = ~n15399 & ~n15429;
  assign n18470 = ~n15764 & n18469;
  assign n18471 = ~n18468 & ~n18470;
  assign n18472 = ~n18463 & n18471;
  assign n18473 = ~n18453 & ~n18472;
  assign n18474 = n18453 & n18472;
  assign po1507 = n18473 | n18474;
  assign n18476 = pi0563 & ~pi1266;
  assign n18477 = ~pi0563 & pi1266;
  assign n18478 = ~n18476 & ~n18477;
  assign n18479 = ~n15554 & n15876;
  assign n18480 = n15863 & ~n18479;
  assign n18481 = n15864 & n15867;
  assign n18482 = ~n18480 & n18481;
  assign n18483 = ~n15861 & n15867;
  assign n18484 = ~n18482 & ~n18483;
  assign n18485 = n15859 & n18484;
  assign n18486 = ~n15543 & ~n18485;
  assign n18487 = n15870 & n18486;
  assign n18488 = ~n15573 & n18487;
  assign n18489 = ~pi1232 & ~n15585;
  assign n18490 = ~n15542 & n15543;
  assign n18491 = ~n18489 & ~n18490;
  assign n18492 = pi0649 & ~n15585;
  assign n18493 = n18491 & ~n18492;
  assign n18494 = ~n15543 & ~n15573;
  assign n18495 = ~n15857 & n18494;
  assign n18496 = ~n18493 & ~n18495;
  assign n18497 = ~n18488 & n18496;
  assign n18498 = ~n18478 & ~n18497;
  assign n18499 = n18478 & n18497;
  assign po1508 = n18498 | n18499;
  assign n18501 = ~pi1400 & ~n18330;
  assign n18502 = pi1798 & n18330;
  assign n18503 = ~n18501 & ~n18502;
  assign po1509 = pi1747 & ~n18503;
  assign n18505 = pi1747 & n3746;
  assign n18506 = pi1401 & n3742;
  assign n18507 = ~n8004 & ~n18506;
  assign n18508 = ~n11649 & n18507;
  assign po1510 = n18505 & ~n18508;
  assign n18510 = ~pi1402 & ~n18030;
  assign n18511 = pi1791 & n18030;
  assign n18512 = ~n18510 & ~n18511;
  assign po1511 = pi1747 & ~n18512;
  assign n18514 = ~pi1403 & ~n18330;
  assign n18515 = pi1795 & n18330;
  assign n18516 = ~n18514 & ~n18515;
  assign po1512 = pi1747 & ~n18516;
  assign n18518 = ~pi1404 & ~n18367;
  assign n18519 = pi1798 & n18367;
  assign n18520 = ~n18518 & ~n18519;
  assign po1513 = pi1747 & ~n18520;
  assign n18522 = ~pi1405 & ~n18330;
  assign n18523 = pi1792 & n18330;
  assign n18524 = ~n18522 & ~n18523;
  assign po1514 = pi1747 & ~n18524;
  assign n18526 = ~pi1406 & ~n18330;
  assign n18527 = pi1800 & n18330;
  assign n18528 = ~n18526 & ~n18527;
  assign po1515 = pi1747 & ~n18528;
  assign n18530 = ~pi1407 & ~n18330;
  assign n18531 = pi1802 & n18330;
  assign n18532 = ~n18530 & ~n18531;
  assign po1516 = pi1747 & ~n18532;
  assign n18534 = ~pi1408 & ~n18030;
  assign n18535 = pi1792 & n18030;
  assign n18536 = ~n18534 & ~n18535;
  assign po1517 = pi1747 & ~n18536;
  assign n18538 = ~pi1411 & ~n18030;
  assign n18539 = pi1793 & n18030;
  assign n18540 = ~n18538 & ~n18539;
  assign po1519 = pi1747 & ~n18540;
  assign n18542 = ~pi1412 & ~n18030;
  assign n18543 = pi1795 & n18030;
  assign n18544 = ~n18542 & ~n18543;
  assign po1520 = pi1747 & ~n18544;
  assign n18546 = pi1413 & ~n17026;
  assign n18547 = n17025 & ~n18546;
  assign n18548 = n16153 & n18075;
  assign po1521 = n18547 | n18548;
  assign n18550 = ~pi1052 & n13676;
  assign n18551 = ~pi0554 & n7999;
  assign n18552 = ~pi0637 & n8080;
  assign n18553 = ~n18551 & ~n18552;
  assign n18554 = ~n18550 & n18553;
  assign n18555 = n13700 & ~n18554;
  assign n18556 = ~pi0453 & n7999;
  assign n18557 = ~pi0457 & n8080;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = ~pi1100 & n13676;
  assign n18560 = n18558 & ~n18559;
  assign n18561 = n13684 & ~n18560;
  assign n18562 = ~n18555 & ~n18561;
  assign n18563 = ~pi1138 & n13676;
  assign n18564 = ~pi0365 & n7999;
  assign n18565 = ~pi0370 & n8080;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = ~n18563 & n18566;
  assign n18568 = n13672 & ~n18567;
  assign n18569 = ~pi0317 & n7999;
  assign n18570 = ~pi0323 & n8080;
  assign n18571 = ~n18569 & ~n18570;
  assign n18572 = ~pi1125 & n13676;
  assign n18573 = n18571 & ~n18572;
  assign n18574 = n13724 & ~n18573;
  assign n18575 = ~n18568 & ~n18574;
  assign po1522 = ~n18562 | ~n18575;
  assign n18577 = pi1111 & n13676;
  assign n18578 = ~pi0556 & n7999;
  assign n18579 = ~pi0639 & n8080;
  assign n18580 = ~n18578 & ~n18579;
  assign n18581 = ~n18577 & n18580;
  assign n18582 = n13700 & ~n18581;
  assign n18583 = pi1143 & n13676;
  assign n18584 = ~pi0455 & n7999;
  assign n18585 = ~pi0532 & n8080;
  assign n18586 = ~n18584 & ~n18585;
  assign n18587 = ~n18583 & n18586;
  assign n18588 = n13684 & ~n18587;
  assign n18589 = ~n18582 & ~n18588;
  assign n18590 = pi1131 & n13676;
  assign n18591 = ~pi0368 & n7999;
  assign n18592 = ~pi0373 & n8080;
  assign n18593 = ~n18591 & ~n18592;
  assign n18594 = ~n18590 & n18593;
  assign n18595 = n13672 & ~n18594;
  assign n18596 = pi1122 & n13676;
  assign n18597 = ~pi0320 & n7999;
  assign n18598 = ~pi0326 & n8080;
  assign n18599 = ~n18597 & ~n18598;
  assign n18600 = ~n18596 & n18599;
  assign n18601 = n13724 & ~n18600;
  assign n18602 = ~n18595 & ~n18601;
  assign po1523 = ~n18589 | ~n18602;
  assign n18604 = ~pi1463 & ~pi1476;
  assign n18605 = pi1465 & ~pi1479;
  assign n18606 = ~pi1465 & pi1479;
  assign n18607 = ~n18605 & ~n18606;
  assign n18608 = n18604 & n18607;
  assign n18609 = ~pi1466 & n18608;
  assign n18610 = pi1464 & n18609;
  assign n18611 = ~pi1472 & n18610;
  assign n18612 = pi1460 & ~pi1479;
  assign n18613 = ~pi1460 & pi1479;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = n18611 & n18614;
  assign n18616 = pi1478 & ~pi1479;
  assign n18617 = ~pi1478 & pi1479;
  assign n18618 = ~n18616 & ~n18617;
  assign po1524 = n18615 & ~n18618;
  assign n18620 = ~pi1516 & ~pi1519;
  assign n18621 = ~pi1479 & pi1518;
  assign n18622 = pi1479 & ~pi1518;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = n18620 & n18623;
  assign n18625 = ~pi1517 & n18624;
  assign n18626 = pi1508 & n18625;
  assign n18627 = ~pi1506 & n18626;
  assign n18628 = ~pi1479 & pi1502;
  assign n18629 = pi1479 & ~pi1502;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = n18627 & n18630;
  assign n18632 = ~pi1479 & pi1521;
  assign n18633 = pi1479 & ~pi1521;
  assign n18634 = ~n18632 & ~n18633;
  assign po1525 = n18631 & ~n18634;
  assign n18636 = n13710 & n16399;
  assign n18637 = pi1776 & n18636;
  assign n18638 = ~pi1419 & ~n18636;
  assign po1527 = n18637 | n18638;
  assign n18640 = ~n15497 & ~n15529;
  assign n18641 = ~n17985 & ~n18640;
  assign n18642 = n17985 & n18640;
  assign po1528 = n18641 | n18642;
  assign n18644 = ~pi1198 & n12899;
  assign n18645 = ~pi1201 & n18644;
  assign n18646 = ~pi1197 & n12892;
  assign n18647 = pi1192 & pi1276;
  assign n18648 = ~pi1194 & ~n18647;
  assign n18649 = ~pi1195 & n18648;
  assign n18650 = n18646 & n18649;
  assign n18651 = n18645 & n18650;
  assign n18652 = pi1036 & ~n18651;
  assign n18653 = ~pi1036 & n18651;
  assign po1529 = n18652 | n18653;
  assign n18655 = pi1422 & ~pi1692;
  assign n18656 = n3935 & n18655;
  assign n18657 = ~n3925 & ~n18656;
  assign n18658 = pi1422 & n3929;
  assign n18659 = n18657 & ~n18658;
  assign n18660 = ~n3932 & n18659;
  assign po1530 = pi1747 & ~n18660;
  assign n18662 = pi1775 & n18636;
  assign n18663 = ~pi1423 & ~n18636;
  assign po1531 = n18662 | n18663;
  assign n18665 = n3855 & n11649;
  assign n18666 = n17282 & n18665;
  assign n18667 = pi1758 & n18666;
  assign po1532 = n17281 & n18667;
  assign n18669 = pi1774 & n18636;
  assign n18670 = ~pi1425 & ~n18636;
  assign po1533 = n18669 | n18670;
  assign n18672 = pi1777 & n18636;
  assign n18673 = ~pi1426 & ~n18636;
  assign po1534 = n18672 | n18673;
  assign n18675 = ~pi1428 & ~pi1707;
  assign n18676 = ~n18636 & ~n18675;
  assign po1536 = pi1747 & ~n18676;
  assign n18678 = ~n3935 & ~n5071;
  assign n18679 = pi1429 & ~n18678;
  assign n18680 = ~n5072 & ~n18679;
  assign po1537 = pi1747 & ~n18680;
  assign n18682 = ~n15401 & ~n15433;
  assign n18683 = ~n18460 & ~n18682;
  assign n18684 = n18460 & n18682;
  assign po1539 = n18683 | n18684;
  assign n18686 = ~n15449 & ~n15481;
  assign n18687 = ~n17959 & ~n18686;
  assign n18688 = n17959 & n18686;
  assign po1540 = n18687 | n18688;
  assign n18690 = ~n15545 & ~n15577;
  assign n18691 = ~n18485 & ~n18690;
  assign n18692 = n18485 & n18690;
  assign po1541 = n18691 | n18692;
  assign n18694 = ~pi1089 & n12478;
  assign n18695 = ~pi1177 & n18694;
  assign n18696 = ~pi1175 & n12471;
  assign n18697 = pi1077 & pi1241;
  assign n18698 = ~pi1173 & ~n18697;
  assign n18699 = ~pi1087 & n18698;
  assign n18700 = n18696 & n18699;
  assign n18701 = n18695 & n18700;
  assign n18702 = pi1179 & ~n18701;
  assign n18703 = ~pi1179 & n18701;
  assign po1542 = n18702 | n18703;
  assign n18705 = ~pi1089 & ~pi1175;
  assign n18706 = ~pi1174 & n12454;
  assign n18707 = ~pi1176 & n18706;
  assign n18708 = ~n18697 & n18707;
  assign n18709 = ~pi1093 & n18708;
  assign n18710 = n18705 & n18709;
  assign n18711 = pi1082 & ~n18710;
  assign n18712 = ~pi1082 & n18710;
  assign po1543 = n18711 | n18712;
  assign n18714 = ~pi1218 & ~pi1219;
  assign n18715 = ~pi1066 & n12988;
  assign n18716 = ~pi1056 & n18715;
  assign n18717 = pi1213 & pi1214;
  assign n18718 = n18716 & ~n18717;
  assign n18719 = ~pi1217 & n18718;
  assign n18720 = n18714 & n18719;
  assign n18721 = pi1057 & ~n18720;
  assign n18722 = ~pi1057 & n18720;
  assign po1544 = n18721 | n18722;
  assign n18724 = n13678 & n18665;
  assign po1545 = n8354 & n18724;
  assign n18726 = ~pi1175 & n18694;
  assign n18727 = ~pi1093 & n18706;
  assign n18728 = ~n18697 & n18727;
  assign n18729 = n18726 & n18728;
  assign n18730 = pi1177 & ~n18729;
  assign n18731 = ~pi1177 & n18729;
  assign po1546 = n18730 | n18731;
  assign po1547 = n9428 & n18724;
  assign po1548 = n8003 & n18724;
  assign n18735 = ~pi1219 & n13001;
  assign n18736 = ~pi1218 & n18735;
  assign n18737 = ~pi1217 & n18715;
  assign n18738 = ~n18717 & n18737;
  assign n18739 = n18736 & n18738;
  assign n18740 = pi1232 & ~n18739;
  assign n18741 = ~pi1232 & n18739;
  assign po1549 = n18740 | n18741;
  assign n18743 = ~n15425 & ~n15434;
  assign n18744 = n15424 & n18743;
  assign n18745 = ~n15424 & ~n18743;
  assign po1550 = n18744 | n18745;
  assign n18747 = ~n15473 & ~n15482;
  assign n18748 = n15472 & n18747;
  assign n18749 = ~n15472 & ~n18747;
  assign po1551 = n18748 | n18749;
  assign n18751 = ~n15521 & ~n15530;
  assign n18752 = n15520 & n18751;
  assign n18753 = ~n15520 & ~n18751;
  assign po1552 = n18752 | n18753;
  assign n18755 = ~pi0553 & n7999;
  assign n18756 = ~pi0635 & n8080;
  assign n18757 = ~n18755 & ~n18756;
  assign n18758 = n13700 & ~n18757;
  assign n18759 = ~pi0452 & n7999;
  assign n18760 = ~pi0454 & n8080;
  assign n18761 = ~n18759 & ~n18760;
  assign n18762 = n13684 & ~n18761;
  assign n18763 = ~n18758 & ~n18762;
  assign n18764 = ~pi0363 & n7999;
  assign n18765 = ~pi0366 & n8080;
  assign n18766 = ~n18764 & ~n18765;
  assign n18767 = n13672 & ~n18766;
  assign n18768 = ~pi0315 & n7999;
  assign n18769 = ~pi0318 & n8080;
  assign n18770 = ~n18768 & ~n18769;
  assign n18771 = n13724 & ~n18770;
  assign n18772 = ~n18767 & ~n18771;
  assign po1553 = ~n18763 | ~n18772;
  assign n18774 = ~n15569 & ~n15578;
  assign n18775 = n15568 & n18774;
  assign n18776 = ~n15568 & ~n18774;
  assign po1554 = n18775 | n18776;
  assign n18778 = ~pi1158 & n13195;
  assign n18779 = ~pi1269 & n18778;
  assign n18780 = ~pi1275 & n13213;
  assign n18781 = pi1283 & pi1331;
  assign n18782 = ~pi1154 & ~n18781;
  assign n18783 = ~pi1155 & n18782;
  assign n18784 = n18780 & n18783;
  assign n18785 = n18779 & n18784;
  assign n18786 = pi1160 & ~n18785;
  assign n18787 = ~pi1160 & n18785;
  assign po1556 = n18786 | n18787;
  assign n18789 = ~pi1232 & n18735;
  assign n18790 = ~pi1218 & n13019;
  assign n18791 = ~pi1215 & ~n18717;
  assign n18792 = ~pi1216 & n18791;
  assign n18793 = n18790 & n18792;
  assign n18794 = n18789 & n18793;
  assign n18795 = pi1266 & ~n18794;
  assign n18796 = ~pi1266 & n18794;
  assign po1557 = n18795 | n18796;
  assign n18798 = ~n15450 & ~n15468;
  assign n18799 = n15804 & ~n15816;
  assign n18800 = n18798 & n18799;
  assign n18801 = ~n18798 & ~n18799;
  assign po1558 = n18800 | n18801;
  assign n18803 = ~n15402 & ~n15420;
  assign n18804 = n15773 & ~n15785;
  assign n18805 = n18803 & n18804;
  assign n18806 = ~n18803 & ~n18804;
  assign po1559 = n18805 | n18806;
  assign n18808 = ~n15498 & ~n15516;
  assign n18809 = n15835 & ~n15847;
  assign n18810 = n18808 & n18809;
  assign n18811 = ~n18808 & ~n18809;
  assign po1560 = n18810 | n18811;
  assign n18813 = ~n15546 & ~n15564;
  assign n18814 = n15866 & ~n15878;
  assign n18815 = n18813 & n18814;
  assign n18816 = ~n18813 & ~n18814;
  assign po1561 = n18815 | n18816;
  assign n18818 = pi1198 & ~n18650;
  assign n18819 = ~pi1198 & n18650;
  assign po1562 = n18818 | n18819;
  assign n18821 = ~pi1197 & ~pi1198;
  assign n18822 = n12892 & n18821;
  assign n18823 = n18649 & n18822;
  assign n18824 = pi1199 & ~n18823;
  assign n18825 = ~pi1199 & n18823;
  assign po1563 = n18824 | n18825;
  assign n18827 = ~pi1197 & n18644;
  assign n18828 = ~pi1196 & n12875;
  assign n18829 = ~pi1264 & n18828;
  assign n18830 = ~n18647 & n18829;
  assign n18831 = n18827 & n18830;
  assign n18832 = pi1201 & ~n18831;
  assign n18833 = ~pi1201 & n18831;
  assign po1564 = n18832 | n18833;
  assign n18835 = ~pi0183 & pi1050;
  assign n18836 = ~pi1457 & ~n18835;
  assign n18837 = n15184 & n15187;
  assign n18838 = n15723 & n18837;
  assign po1565 = ~n18836 & ~n18838;
  assign n18840 = pi1458 & n5234;
  assign n18841 = ~po1678 & ~n18840;
  assign po1566 = pi1747 & ~n18841;
  assign n18843 = pi1465 & pi1466;
  assign n18844 = pi1464 & n18843;
  assign n18845 = pi1472 & n18844;
  assign n18846 = pi1460 & n18845;
  assign n18847 = ~pi1460 & ~n18845;
  assign n18848 = ~n18846 & ~n18847;
  assign po1568 = pi1626 & n18848;
  assign n18850 = pi1089 & ~n18700;
  assign n18851 = ~pi1089 & n18700;
  assign po1569 = n18850 | n18851;
  assign n18853 = n12471 & n18705;
  assign n18854 = n18699 & n18853;
  assign n18855 = pi1176 & ~n18854;
  assign n18856 = ~pi1176 & n18854;
  assign po1570 = n18855 | n18856;
  assign n18858 = pi1460 & pi1478;
  assign n18859 = pi1472 & n18843;
  assign n18860 = pi1464 & n18859;
  assign n18861 = n18858 & n18860;
  assign n18862 = pi1463 & n18861;
  assign n18863 = ~pi1463 & ~n18861;
  assign n18864 = ~n18862 & ~n18863;
  assign po1571 = pi1626 & n18864;
  assign n18866 = ~pi1464 & ~n18843;
  assign n18867 = ~n18844 & ~n18866;
  assign po1572 = pi1626 & n18867;
  assign n18869 = ~pi1465 & ~pi1466;
  assign n18870 = ~n18843 & ~n18869;
  assign po1573 = pi1626 & n18870;
  assign po1574 = ~pi1466 & pi1626;
  assign n18873 = ~pi1158 & ~pi1275;
  assign n18874 = ~pi1156 & n13182;
  assign n18875 = ~pi1346 & n18874;
  assign n18876 = ~n18781 & n18875;
  assign n18877 = ~pi1157 & n18876;
  assign n18878 = n18873 & n18877;
  assign n18879 = pi1159 & ~n18878;
  assign n18880 = ~pi1159 & n18878;
  assign po1575 = n18879 | n18880;
  assign n18882 = ~pi1199 & n18828;
  assign n18883 = ~n18647 & n18882;
  assign n18884 = ~pi1264 & n18883;
  assign n18885 = n18821 & n18884;
  assign n18886 = pi1249 & ~n18885;
  assign n18887 = ~pi1249 & n18885;
  assign po1576 = n18886 | n18887;
  assign n18889 = ~pi1275 & n18778;
  assign n18890 = ~pi1157 & n18874;
  assign n18891 = ~n18781 & n18890;
  assign n18892 = n18889 & n18891;
  assign n18893 = pi1269 & ~n18892;
  assign n18894 = ~pi1269 & n18892;
  assign po1577 = n18893 | n18894;
  assign n18896 = ~pi0811 & ~pi0820;
  assign n18897 = ~pi0812 & ~pi0813;
  assign n18898 = ~pi0834 & n18897;
  assign n18899 = ~pi0814 & n18898;
  assign n18900 = n18896 & n18899;
  assign n18901 = ~pi0815 & ~pi0870;
  assign n18902 = ~pi0817 & n18901;
  assign n18903 = ~pi0816 & n18902;
  assign n18904 = ~pi0831 & ~pi0832;
  assign n18905 = ~pi0833 & n18904;
  assign n18906 = ~pi0757 & n18905;
  assign n18907 = n18903 & n18906;
  assign n18908 = ~pi0828 & n18907;
  assign n18909 = n18900 & n18908;
  assign n18910 = ~pi0756 & ~pi0830;
  assign po1619 = n18909 & n18910;
  assign po1578 = ~pi0829 | po1619;
  assign n18913 = ~pi0835 & ~pi0843;
  assign n18914 = ~pi0758 & ~pi0836;
  assign n18915 = ~pi0858 & n18914;
  assign n18916 = ~pi0837 & n18915;
  assign n18917 = n18913 & n18916;
  assign n18918 = ~pi0855 & ~pi0856;
  assign n18919 = ~pi0857 & n18918;
  assign n18920 = ~pi0879 & n18919;
  assign n18921 = ~pi0752 & ~pi0838;
  assign n18922 = ~pi0840 & n18921;
  assign n18923 = ~pi0839 & n18922;
  assign n18924 = n18920 & n18923;
  assign n18925 = ~pi0851 & n18924;
  assign n18926 = n18917 & n18925;
  assign n18927 = ~pi0854 & ~pi0880;
  assign po1618 = n18926 & n18927;
  assign po1579 = ~pi0853 | po1618;
  assign n18930 = ~pi1472 & ~n18844;
  assign n18931 = ~n18845 & ~n18930;
  assign po1580 = pi1626 & n18931;
  assign n18933 = n9548 & n13678;
  assign po1581 = n18665 & n18933;
  assign n18935 = pi1175 & ~n18728;
  assign n18936 = ~pi1175 & n18728;
  assign po1582 = n18935 | n18936;
  assign n18938 = pi1218 & ~n18738;
  assign n18939 = ~pi1218 & n18738;
  assign po1583 = n18938 | n18939;
  assign n18941 = pi1463 & n18844;
  assign n18942 = pi1472 & n18941;
  assign n18943 = n18858 & n18942;
  assign n18944 = pi1476 & n18943;
  assign n18945 = ~pi1476 & ~n18943;
  assign n18946 = ~n18944 & ~n18945;
  assign po1584 = pi1626 & n18946;
  assign n18948 = ~pi1173 & n12484;
  assign n18949 = n12478 & n18853;
  assign n18950 = ~pi1087 & n18949;
  assign n18951 = n18948 & n18950;
  assign po1585 = n12525 & ~n18951;
  assign n18953 = pi1460 & n18859;
  assign n18954 = pi1464 & n18953;
  assign n18955 = pi1478 & n18954;
  assign n18956 = ~pi1478 & ~n18954;
  assign n18957 = ~n18955 & ~n18956;
  assign po1586 = pi1626 & n18957;
  assign n18959 = ~pi0760 & ~pi1479;
  assign n18960 = n15187 & n15719;
  assign n18961 = n15721 & n18960;
  assign n18962 = n15184 & n18961;
  assign po1587 = ~n18959 & ~n18962;
  assign n18964 = pi0333 & ~pi1099;
  assign n18965 = pi0221 & pi1099;
  assign po1589 = n18964 | n18965;
  assign n18967 = pi1195 & ~n18648;
  assign po1590 = n18649 | n18967;
  assign n18969 = pi1158 & ~n18784;
  assign n18970 = ~pi1158 & n18784;
  assign po1591 = n18969 | n18970;
  assign n18972 = pi1219 & ~n18793;
  assign n18973 = ~pi1219 & n18793;
  assign po1592 = n18972 | n18973;
  assign n18975 = n13213 & n18873;
  assign n18976 = n18783 & n18975;
  assign n18977 = pi1346 & ~n18976;
  assign n18978 = ~pi1346 & n18976;
  assign po1593 = n18977 | n18978;
  assign n18980 = n13019 & n18714;
  assign n18981 = n18792 & n18980;
  assign n18982 = pi1056 & ~n18981;
  assign n18983 = ~pi1056 & n18981;
  assign po1594 = n18982 | n18983;
  assign po1595 = pi1611 | pi1617;
  assign n18986 = pi1196 & ~n18649;
  assign n18987 = ~pi1196 & n18649;
  assign po1596 = n18986 | n18987;
  assign n18989 = pi1194 & n18647;
  assign po1597 = n18648 | n18989;
  assign n18991 = pi1197 & ~n18830;
  assign n18992 = ~pi1197 & n18830;
  assign po1598 = n18991 | n18992;
  assign n18994 = ~pi1215 & n13007;
  assign n18995 = n13001 & n18980;
  assign n18996 = ~pi1216 & n18995;
  assign n18997 = n18994 & n18996;
  assign po1599 = n13055 & ~n18997;
  assign n18999 = ~pi1194 & n12905;
  assign n19000 = n12899 & n18822;
  assign n19001 = ~pi1195 & n19000;
  assign n19002 = n18999 & n19001;
  assign po1600 = n12946 & ~n19002;
  assign n19004 = pi1493 & ~po1678;
  assign n19005 = n5234 & ~n19004;
  assign po1601 = pi1747 & ~n19005;
  assign n19007 = pi1494 & ~po1676;
  assign n19008 = ~po1678 & n19007;
  assign n19009 = ~po1688 & ~n19008;
  assign po1602 = pi1747 & ~n19009;
  assign n19011 = pi1087 & ~n18698;
  assign po1605 = n18699 | n19011;
  assign n19013 = ~n15417 & ~n15421;
  assign n19014 = n15416 & n19013;
  assign n19015 = ~n15416 & ~n19013;
  assign po1606 = n19014 | n19015;
  assign n19017 = ~n15465 & ~n15469;
  assign n19018 = n15464 & n19017;
  assign n19019 = ~n15464 & ~n19017;
  assign po1607 = n19018 | n19019;
  assign n19021 = ~n15513 & ~n15517;
  assign n19022 = n15512 & n19021;
  assign n19023 = ~n15512 & ~n19021;
  assign po1608 = n19022 | n19023;
  assign n19025 = ~n15561 & ~n15565;
  assign n19026 = n15560 & n19025;
  assign n19027 = ~n15560 & ~n19025;
  assign po1609 = n19026 | n19027;
  assign n19029 = pi1517 & pi1518;
  assign n19030 = pi1508 & n19029;
  assign n19031 = pi1506 & n19030;
  assign n19032 = pi1502 & n19031;
  assign n19033 = ~pi1502 & ~n19031;
  assign n19034 = ~n19032 & ~n19033;
  assign po1610 = ~pi1581 & n19034;
  assign po1611 = ~pi1613 | ~pi1616;
  assign po1612 = ~pi1619 | ~pi1620;
  assign po1613 = ~pi1612 | ~pi1618;
  assign n19039 = ~pi1506 & ~n19030;
  assign n19040 = ~n19031 & ~n19039;
  assign po1614 = ~pi1581 & n19040;
  assign n19042 = pi1174 & ~n18699;
  assign n19043 = ~pi1174 & n18699;
  assign po1615 = n19042 | n19043;
  assign n19045 = ~pi1508 & ~n19029;
  assign n19046 = ~n19030 & ~n19045;
  assign po1616 = ~pi1581 & n19046;
  assign n19048 = pi1173 & n18697;
  assign po1617 = n18698 | n19048;
  assign n19050 = ~n18697 & n18706;
  assign n19051 = pi1093 & ~n19050;
  assign n19052 = ~pi1093 & n19050;
  assign po1620 = n19051 | n19052;
  assign n19054 = ~n18647 & n18828;
  assign n19055 = pi1264 & ~n19054;
  assign n19056 = ~pi1264 & n19054;
  assign po1621 = n19055 | n19056;
  assign n19058 = pi1275 & ~n18891;
  assign n19059 = ~pi1275 & n18891;
  assign po1622 = n19058 | n19059;
  assign n19061 = n18715 & ~n18717;
  assign n19062 = pi1217 & ~n19061;
  assign n19063 = ~pi1217 & n19061;
  assign po1623 = n19062 | n19063;
  assign n19065 = pi1502 & pi1521;
  assign n19066 = pi1506 & n19029;
  assign n19067 = pi1508 & n19066;
  assign n19068 = n19065 & n19067;
  assign n19069 = pi1516 & n19068;
  assign n19070 = ~pi1516 & ~n19068;
  assign n19071 = ~n19069 & ~n19070;
  assign po1624 = ~pi1581 & n19071;
  assign po1625 = ~pi1517 & ~pi1581;
  assign n19074 = ~pi1517 & ~pi1518;
  assign n19075 = ~n19029 & ~n19074;
  assign po1626 = ~pi1581 & n19075;
  assign n19077 = pi1516 & n19030;
  assign n19078 = pi1506 & n19077;
  assign n19079 = n19065 & n19078;
  assign n19080 = pi1519 & n19079;
  assign n19081 = ~pi1519 & ~n19079;
  assign n19082 = ~n19080 & ~n19081;
  assign po1627 = ~pi1581 & n19082;
  assign n19084 = ~pi1154 & n13201;
  assign n19085 = n13195 & n18975;
  assign n19086 = ~pi1155 & n19085;
  assign n19087 = n19084 & n19086;
  assign po1628 = n13249 & ~n19087;
  assign n19089 = pi1502 & n19066;
  assign n19090 = pi1508 & n19089;
  assign n19091 = pi1521 & n19090;
  assign n19092 = ~pi1521 & ~n19090;
  assign n19093 = ~n19091 & ~n19092;
  assign po1629 = ~pi1581 & n19093;
  assign n19095 = pi0788 & n13328;
  assign n19096 = ~pi0764 & pi0783;
  assign n19097 = n19095 & n19096;
  assign n19098 = pi0765 & n19097;
  assign n19099 = ~pi0790 & n19098;
  assign n19100 = ~pi0766 & ~n19099;
  assign n19101 = pi0766 & n19099;
  assign po1630 = n19100 | n19101;
  assign n19103 = ~pi1228 & pi1231;
  assign n19104 = pi1228 & ~pi1231;
  assign n19105 = ~n19103 & ~n19104;
  assign n19106 = ~pi1227 & pi1230;
  assign n19107 = pi1227 & ~pi1230;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = pi1079 & ~pi1236;
  assign n19110 = ~pi1079 & pi1236;
  assign n19111 = ~n19109 & ~n19110;
  assign n19112 = pi1058 & ~pi1229;
  assign n19113 = ~pi1058 & pi1229;
  assign n19114 = ~n19112 & ~n19113;
  assign n19115 = ~n19111 & ~n19114;
  assign n19116 = ~n19108 & n19115;
  assign po1631 = n19105 | ~n19116;
  assign n19118 = pi1155 & ~n18782;
  assign po1632 = n18783 | n19118;
  assign n19120 = pi1216 & ~n18791;
  assign po1633 = n18792 | n19120;
  assign po1634 = n4131 & n15623;
  assign n19123 = n13328 & n14020;
  assign n19124 = pi0783 & n19123;
  assign n19125 = pi0788 & n19124;
  assign n19126 = pi0765 & ~n19125;
  assign n19127 = ~pi0765 & n19125;
  assign po1635 = n19126 | n19127;
  assign n19129 = ~n15403 & ~n15404;
  assign n19130 = n18455 & n19129;
  assign n19131 = ~n18455 & ~n19129;
  assign po1636 = n19130 | n19131;
  assign n19133 = ~n15451 & ~n15452;
  assign n19134 = n17954 & n19133;
  assign n19135 = ~n17954 & ~n19133;
  assign po1637 = n19134 | n19135;
  assign n19137 = ~n15499 & ~n15500;
  assign n19138 = n17980 & n19137;
  assign n19139 = ~n17980 & ~n19137;
  assign po1638 = n19138 | n19139;
  assign n19141 = ~n15547 & ~n15548;
  assign n19142 = n18480 & n19141;
  assign n19143 = ~n18480 & ~n19141;
  assign po1639 = n19142 | n19143;
  assign n19145 = pi0783 & n19095;
  assign n19146 = ~pi0764 & ~n19145;
  assign n19147 = pi0764 & n19145;
  assign po1640 = n19146 | n19147;
  assign n19149 = pi1156 & ~n18783;
  assign n19150 = ~pi1156 & n18783;
  assign po1641 = n19149 | n19150;
  assign n19152 = pi0283 & pi0291;
  assign n19153 = pi0289 & n19152;
  assign n19154 = pi0290 & n19153;
  assign n19155 = ~pi1534 & n19154;
  assign n19156 = n7749 & n19155;
  assign n19157 = ~pi0292 & ~pi0293;
  assign po1642 = n19156 & n19157;
  assign n19159 = pi1066 & ~n18792;
  assign n19160 = ~pi1066 & n18792;
  assign po1643 = n19159 | n19160;
  assign n19162 = pi1215 & n18717;
  assign po1644 = n18791 | n19162;
  assign n19164 = ~n18781 & n18874;
  assign n19165 = pi1157 & ~n19164;
  assign n19166 = ~pi1157 & n19164;
  assign po1645 = n19165 | n19166;
  assign n19168 = n10900 & n12978;
  assign po1646 = n5792 & ~n19168;
  assign n19170 = n12194 & n13172;
  assign po1647 = n5886 & ~n19170;
  assign n19172 = n9006 & n12448;
  assign po1648 = n5806 & ~n19172;
  assign n19174 = n10014 & n12869;
  assign po1649 = n5631 & ~n19174;
  assign n19176 = ~pi0787 & n14020;
  assign n19177 = pi0761 & n19176;
  assign n19178 = ~pi0766 & n19177;
  assign n19179 = pi0765 & n19178;
  assign n19180 = pi0783 & ~pi0788;
  assign po1652 = n19179 & n19180;
  assign n19182 = pi1154 & n18781;
  assign po1653 = n18782 | n19182;
  assign n19184 = pi0787 & n19096;
  assign n19185 = pi0788 & n19184;
  assign n19186 = pi0761 & n19185;
  assign n19187 = ~pi0790 & ~n19186;
  assign n19188 = pi0790 & n19186;
  assign po1654 = n19187 | n19188;
  assign n19190 = pi0783 & ~n19095;
  assign n19191 = ~pi0783 & n19095;
  assign po1658 = n19190 | n19191;
  assign n19193 = pi1551 & pi1694;
  assign n19194 = ~pi1840 & ~n19193;
  assign po1659 = pi1747 & ~n19194;
  assign n19196 = ~n15501 & ~n15509;
  assign n19197 = ~n15508 & ~n19196;
  assign n19198 = n15508 & n19196;
  assign po1660 = n19197 | n19198;
  assign n19200 = ~n15453 & ~n15461;
  assign n19201 = ~n15460 & ~n19200;
  assign n19202 = n15460 & n19200;
  assign po1661 = n19201 | n19202;
  assign n19204 = ~n15405 & ~n15413;
  assign n19205 = ~n15412 & ~n19204;
  assign n19206 = n15412 & n19204;
  assign po1662 = n19205 | n19206;
  assign n19208 = ~n15549 & ~n15557;
  assign n19209 = ~n15556 & ~n19208;
  assign n19210 = n15556 & n19208;
  assign po1663 = n19209 | n19210;
  assign n19212 = pi1556 & pi1689;
  assign n19213 = ~pi1839 & ~n19212;
  assign po1664 = pi1747 & ~n19213;
  assign n19215 = ~n15552 & ~n15554;
  assign n19216 = ~n15553 & ~n19215;
  assign n19217 = n15553 & n19215;
  assign po1665 = n19216 | n19217;
  assign n19219 = ~n15504 & ~n15506;
  assign n19220 = ~n15505 & ~n19219;
  assign n19221 = n15505 & n19219;
  assign po1666 = n19220 | n19221;
  assign n19223 = ~n15456 & ~n15458;
  assign n19224 = ~n15457 & ~n19223;
  assign n19225 = n15457 & n19223;
  assign po1667 = n19224 | n19225;
  assign n19227 = ~n15408 & ~n15410;
  assign n19228 = ~n15409 & ~n19227;
  assign n19229 = n15409 & n19227;
  assign po1668 = n19228 | n19229;
  assign n19231 = pi1561 & pi1691;
  assign n19232 = ~pi1838 & ~n19231;
  assign po1669 = pi1747 & ~n19232;
  assign n19234 = pi1562 & pi1696;
  assign n19235 = ~pi1841 & ~n19234;
  assign po1670 = pi1747 & ~n19235;
  assign n19237 = pi0038 & pi1101;
  assign n19238 = pi1825 & n19237;
  assign n19239 = pi1563 & ~n19237;
  assign po1671 = n19238 | n19239;
  assign n19241 = pi1807 & n19237;
  assign n19242 = pi1564 & ~n19237;
  assign po1672 = n19241 | n19242;
  assign n19244 = pi1077 & ~pi1241;
  assign n19245 = ~pi1077 & pi1241;
  assign po1673 = n19244 | n19245;
  assign n19247 = pi1283 & ~pi1331;
  assign n19248 = ~pi1283 & pi1331;
  assign po1674 = n19247 | n19248;
  assign n19250 = ~pi1213 & pi1214;
  assign n19251 = pi1213 & ~pi1214;
  assign po1675 = n19250 | n19251;
  assign n19253 = ~pi1047 & ~pi1526;
  assign po1677 = ~pi1697 & ~n19253;
  assign po1679 = ~pi1690 & ~n19253;
  assign po1680 = ~pi1679 & ~n19253;
  assign n19257 = pi1837 & n19237;
  assign n19258 = pi1573 & ~n19237;
  assign po1681 = n19257 | n19258;
  assign n19260 = pi1836 & n19237;
  assign n19261 = pi1574 & ~n19237;
  assign po1682 = n19260 | n19261;
  assign n19263 = pi1813 & n19237;
  assign n19264 = pi1575 & ~n19237;
  assign po1683 = n19263 | n19264;
  assign n19266 = pi1830 & n19237;
  assign n19267 = pi1576 & ~n19237;
  assign po1684 = n19266 | n19267;
  assign n19269 = pi1827 & n19237;
  assign n19270 = pi1577 & ~n19237;
  assign po1685 = n19269 | n19270;
  assign n19272 = ~pi0092 & ~pi0108;
  assign po1689 = pi0047 | n19272;
  assign n19274 = pi1583 & ~pi1743;
  assign n19275 = pi0713 & ~n19274;
  assign po1691 = pi1747 & ~n19275;
  assign n19277 = pi1832 & n19237;
  assign n19278 = pi1584 & ~n19237;
  assign po1692 = n19277 | n19278;
  assign n19280 = pi1833 & n19237;
  assign n19281 = pi1585 & ~n19237;
  assign po1693 = n19280 | n19281;
  assign n19283 = pi1809 & n19237;
  assign n19284 = pi1586 & ~n19237;
  assign po1694 = n19283 | n19284;
  assign n19286 = pi1806 & n19237;
  assign n19287 = pi1587 & ~n19237;
  assign po1695 = n19286 | n19287;
  assign n19289 = pi1818 & n19237;
  assign n19290 = pi1588 & ~n19237;
  assign po1696 = n19289 | n19290;
  assign n19292 = pi1808 & n19237;
  assign n19293 = pi1589 & ~n19237;
  assign po1697 = n19292 | n19293;
  assign n19295 = pi1814 & n19237;
  assign n19296 = pi1590 & ~n19237;
  assign po1698 = n19295 | n19296;
  assign n19298 = pi1824 & n19237;
  assign n19299 = pi1591 & ~n19237;
  assign po1699 = n19298 | n19299;
  assign n19301 = pi1834 & n19237;
  assign n19302 = pi1592 & ~n19237;
  assign po1700 = n19301 | n19302;
  assign n19304 = pi1820 & n19237;
  assign n19305 = pi1593 & ~n19237;
  assign po1701 = n19304 | n19305;
  assign po1702 = ~pi1699 & ~n19253;
  assign n19308 = pi1812 & n19237;
  assign n19309 = pi1595 & ~n19237;
  assign po1703 = n19308 | n19309;
  assign n19311 = pi1811 & n19237;
  assign n19312 = pi1596 & ~n19237;
  assign po1704 = n19311 | n19312;
  assign n19314 = pi1815 & n19237;
  assign n19315 = pi1597 & ~n19237;
  assign po1705 = n19314 | n19315;
  assign n19317 = pi1826 & n19237;
  assign n19318 = pi1598 & ~n19237;
  assign po1706 = n19317 | n19318;
  assign n19320 = pi1828 & n19237;
  assign n19321 = pi1599 & ~n19237;
  assign po1707 = n19320 | n19321;
  assign n19323 = pi1821 & n19237;
  assign n19324 = pi1600 & ~n19237;
  assign po1708 = n19323 | n19324;
  assign n19326 = pi1829 & n19237;
  assign n19327 = pi1601 & ~n19237;
  assign po1709 = n19326 | n19327;
  assign n19329 = pi1831 & n19237;
  assign n19330 = pi1602 & ~n19237;
  assign po1710 = n19329 | n19330;
  assign n19332 = pi1823 & n19237;
  assign n19333 = pi1603 & ~n19237;
  assign po1711 = n19332 | n19333;
  assign n19335 = pi1604 & ~pi1728;
  assign n19336 = pi0721 & ~n19335;
  assign po1712 = pi1747 & ~n19336;
  assign n19338 = pi1822 & n19237;
  assign n19339 = pi1605 & ~n19237;
  assign po1713 = n19338 | n19339;
  assign n19341 = pi1810 & n19237;
  assign n19342 = pi1606 & ~n19237;
  assign po1714 = n19341 | n19342;
  assign n19344 = pi1607 & ~pi1734;
  assign n19345 = pi0676 & ~n19344;
  assign po1715 = pi1747 & ~n19345;
  assign n19347 = pi1608 & ~pi1730;
  assign n19348 = pi0711 & ~n19347;
  assign po1716 = pi1747 & ~n19348;
  assign n19350 = pi1835 & n19237;
  assign n19351 = pi1609 & ~n19237;
  assign po1717 = n19350 | n19351;
  assign n19353 = pi1816 & n19237;
  assign n19354 = pi1610 & ~n19237;
  assign po1718 = n19353 | n19354;
  assign n19356 = pi0131 & ~pi1391;
  assign n19357 = pi0891 & ~pi1411;
  assign n19358 = ~n19356 & ~n19357;
  assign n19359 = pi0990 & ~pi1412;
  assign n19360 = pi0959 & ~pi1411;
  assign n19361 = pi0118 & ~pi1408;
  assign n19362 = ~n19360 & ~n19361;
  assign n19363 = pi1037 & ~pi1402;
  assign n19364 = pi0617 & ~pi1394;
  assign n19365 = ~n19363 & ~n19364;
  assign n19366 = n19362 & n19365;
  assign n19367 = ~n19359 & n19366;
  assign po1719 = ~n19358 | ~n19367;
  assign n19369 = pi0128 & ~pi1379;
  assign n19370 = pi0903 & ~pi1380;
  assign n19371 = ~n19369 & ~n19370;
  assign n19372 = pi1048 & ~pi1403;
  assign n19373 = pi1035 & ~pi1378;
  assign n19374 = pi0592 & ~pi1377;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = pi0970 & ~pi1380;
  assign n19377 = pi0114 & ~pi1405;
  assign n19378 = ~n19376 & ~n19377;
  assign n19379 = n19375 & n19378;
  assign n19380 = ~n19372 & n19379;
  assign po1720 = ~n19371 | ~n19380;
  assign n19382 = pi0958 & ~pi1389;
  assign n19383 = pi0116 & ~pi1395;
  assign n19384 = ~n19382 & ~n19383;
  assign n19385 = pi0965 & ~pi1393;
  assign n19386 = pi0991 & ~pi1387;
  assign n19387 = pi0615 & ~pi1397;
  assign n19388 = ~n19386 & ~n19387;
  assign n19389 = pi0130 & ~pi1388;
  assign n19390 = pi0904 & ~pi1389;
  assign n19391 = ~n19389 & ~n19390;
  assign n19392 = n19388 & n19391;
  assign n19393 = ~n19385 & n19392;
  assign po1721 = ~n19384 | ~n19393;
  assign n19395 = pi1817 & n19237;
  assign n19396 = pi1614 & ~n19237;
  assign po1722 = n19395 | n19396;
  assign n19398 = pi1819 & n19237;
  assign n19399 = pi1615 & ~n19237;
  assign po1723 = n19398 | n19399;
  assign n19401 = pi0130 & ~pi1396;
  assign n19402 = pi0965 & ~pi1386;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = pi0904 & ~pi1385;
  assign n19405 = pi0116 & ~pi1384;
  assign n19406 = pi0958 & ~pi1385;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = pi0991 & ~pi1383;
  assign n19409 = pi0615 & ~pi1404;
  assign n19410 = ~n19408 & ~n19409;
  assign n19411 = n19407 & n19410;
  assign n19412 = ~n19404 & n19411;
  assign po1724 = ~n19403 | ~n19412;
  assign n19414 = pi0131 & ~pi1349;
  assign n19415 = pi0990 & ~pi1352;
  assign n19416 = ~n19414 & ~n19415;
  assign n19417 = pi0891 & ~pi1364;
  assign n19418 = pi1037 & ~pi1362;
  assign n19419 = pi0617 & ~pi1359;
  assign n19420 = ~n19418 & ~n19419;
  assign n19421 = pi0118 & ~pi1390;
  assign n19422 = pi0959 & ~pi1364;
  assign n19423 = ~n19421 & ~n19422;
  assign n19424 = n19420 & n19423;
  assign n19425 = ~n19417 & n19424;
  assign po1725 = ~n19416 | ~n19425;
  assign n19427 = pi0128 & ~pi1407;
  assign n19428 = pi1048 & ~pi1376;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = pi0903 & ~pi1375;
  assign n19431 = pi1035 & ~pi1374;
  assign n19432 = pi0592 & ~pi1400;
  assign n19433 = ~n19431 & ~n19432;
  assign n19434 = pi0114 & ~pi1406;
  assign n19435 = pi0970 & ~pi1375;
  assign n19436 = ~n19434 & ~n19435;
  assign n19437 = n19433 & n19436;
  assign n19438 = ~n19430 & n19437;
  assign po1726 = ~n19429 | ~n19438;
  assign n19440 = pi0129 & ~pi1353;
  assign n19441 = pi1314 & ~pi1356;
  assign n19442 = ~n19440 & ~n19441;
  assign n19443 = pi0892 & ~pi1348;
  assign n19444 = pi1165 & ~pi1363;
  assign n19445 = pi0535 & ~pi1381;
  assign n19446 = ~n19444 & ~n19445;
  assign n19447 = pi0115 & ~pi1382;
  assign n19448 = pi0957 & ~pi1348;
  assign n19449 = ~n19447 & ~n19448;
  assign n19450 = n19446 & n19449;
  assign n19451 = ~n19443 & n19450;
  assign po1727 = ~n19442 | ~n19451;
  assign n19453 = pi0129 & ~pi1351;
  assign n19454 = pi0892 & ~pi1354;
  assign n19455 = ~n19453 & ~n19454;
  assign n19456 = pi1314 & ~pi1347;
  assign n19457 = pi1165 & ~pi1355;
  assign n19458 = pi0535 & ~pi1357;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = pi0957 & ~pi1354;
  assign n19461 = pi0115 & ~pi1350;
  assign n19462 = ~n19460 & ~n19461;
  assign n19463 = n19459 & n19462;
  assign n19464 = ~n19456 & n19463;
  assign po1728 = ~n19455 | ~n19464;
  assign n19466 = pi0279 & pi0294;
  assign n19467 = ~pi0295 & n19466;
  assign n19468 = ~pi0296 & n19467;
  assign n19469 = pi0307 & n19468;
  assign n19470 = pi0297 & n19469;
  assign n19471 = ~pi0308 & n19470;
  assign po1729 = pi0298 & n19471;
  assign n19473 = ~pi0700 & pi1331;
  assign po1730 = n15409 | n19473;
  assign n19475 = ~pi0594 & pi1213;
  assign po1731 = n15553 | n19475;
  assign n19477 = ~pi0410 & pi1241;
  assign po1732 = n15457 | n19477;
  assign po1734 = pi1747 & pi1755;
  assign po1735 = pi1747 & pi1756;
  assign po1736 = pi1747 & pi1754;
  assign n19482 = ~pi0511 & pi1192;
  assign po1738 = n15505 | n19482;
  assign n19484 = pi0788 & ~n13328;
  assign n19485 = ~pi0788 & n13328;
  assign po1739 = n19484 | n19485;
  assign n19487 = ~pi0038 & pi1101;
  assign n19488 = pi1808 & n19487;
  assign n19489 = pi1632 & ~n19487;
  assign po1740 = n19488 | n19489;
  assign n19491 = pi1837 & n19487;
  assign n19492 = pi1633 & ~n19487;
  assign po1741 = n19491 | n19492;
  assign n19494 = pi1834 & n19487;
  assign n19495 = pi1634 & ~n19487;
  assign po1742 = n19494 | n19495;
  assign n19497 = pi1812 & n19487;
  assign n19498 = pi1635 & ~n19487;
  assign po1743 = n19497 | n19498;
  assign n19500 = pi1829 & n19487;
  assign n19501 = pi1636 & ~n19487;
  assign po1744 = n19500 | n19501;
  assign n19503 = pi1192 & ~pi1276;
  assign n19504 = ~pi1192 & pi1276;
  assign po1745 = n19503 | n19504;
  assign n19506 = pi1825 & n19487;
  assign n19507 = pi1638 & ~n19487;
  assign po1746 = n19506 | n19507;
  assign n19509 = pi1830 & n19487;
  assign n19510 = pi1639 & ~n19487;
  assign po1747 = n19509 | n19510;
  assign n19512 = pi1824 & n19487;
  assign n19513 = pi1640 & ~n19487;
  assign po1748 = n19512 | n19513;
  assign n19515 = pi1816 & n19487;
  assign n19516 = pi1641 & ~n19487;
  assign po1749 = n19515 | n19516;
  assign n19518 = pi1810 & n19487;
  assign n19519 = pi1642 & ~n19487;
  assign po1750 = n19518 | n19519;
  assign n19521 = pi1836 & n19487;
  assign n19522 = pi1643 & ~n19487;
  assign po1751 = n19521 | n19522;
  assign n19524 = pi1833 & n19487;
  assign n19525 = pi1644 & ~n19487;
  assign po1752 = n19524 | n19525;
  assign n19527 = pi1809 & n19487;
  assign n19528 = pi1645 & ~n19487;
  assign po1753 = n19527 | n19528;
  assign n19530 = pi1811 & n19487;
  assign n19531 = pi1646 & ~n19487;
  assign po1754 = n19530 | n19531;
  assign n19533 = pi1814 & n19487;
  assign n19534 = pi1647 & ~n19487;
  assign po1755 = n19533 | n19534;
  assign n19536 = pi1832 & n19487;
  assign n19537 = pi1648 & ~n19487;
  assign po1756 = n19536 | n19537;
  assign n19539 = pi1820 & n19487;
  assign n19540 = pi1649 & ~n19487;
  assign po1757 = n19539 | n19540;
  assign n19542 = pi1806 & n19487;
  assign n19543 = pi1650 & ~n19487;
  assign po1758 = n19542 | n19543;
  assign n19545 = pi1807 & n19487;
  assign n19546 = pi1651 & ~n19487;
  assign po1759 = n19545 | n19546;
  assign n19548 = pi1835 & n19487;
  assign n19549 = pi1652 & ~n19487;
  assign po1760 = n19548 | n19549;
  assign n19551 = pi1815 & n19487;
  assign n19552 = pi1653 & ~n19487;
  assign po1761 = n19551 | n19552;
  assign n19554 = pi1827 & n19487;
  assign n19555 = pi1654 & ~n19487;
  assign po1762 = n19554 | n19555;
  assign n19557 = pi1826 & n19487;
  assign n19558 = pi1655 & ~n19487;
  assign po1763 = n19557 | n19558;
  assign n19560 = pi1822 & n19487;
  assign n19561 = pi1656 & ~n19487;
  assign po1764 = n19560 | n19561;
  assign n19563 = pi1823 & n19487;
  assign n19564 = pi1657 & ~n19487;
  assign po1765 = n19563 | n19564;
  assign n19566 = pi1813 & n19487;
  assign n19567 = pi1658 & ~n19487;
  assign po1766 = n19566 | n19567;
  assign n19569 = pi1828 & n19487;
  assign n19570 = pi1659 & ~n19487;
  assign po1767 = n19569 | n19570;
  assign n19572 = pi1819 & n19487;
  assign n19573 = pi1660 & ~n19487;
  assign po1768 = n19572 | n19573;
  assign n19575 = pi1831 & n19487;
  assign n19576 = pi1661 & ~n19487;
  assign po1769 = n19575 | n19576;
  assign n19578 = pi1818 & n19487;
  assign n19579 = pi1662 & ~n19487;
  assign po1770 = n19578 | n19579;
  assign n19581 = pi1821 & n19487;
  assign n19582 = pi1663 & ~n19487;
  assign po1771 = n19581 | n19582;
  assign n19584 = pi1817 & n19487;
  assign n19585 = pi1664 & ~n19487;
  assign po1772 = n19584 | n19585;
  assign n19587 = ~pi0763 & ~pi0793;
  assign po1773 = n14051 & n19587;
  assign po1774 = pi0012 & ~pi1099;
  assign po1777 = pi0409 | ~n3716;
  assign n19591 = ~pi0919 & ~pi0921;
  assign po1778 = pi0963 & n19591;
  assign n19593 = ~pi0268 & ~pi0331;
  assign n19594 = pi0274 & n19593;
  assign n19595 = pi0285 & n19594;
  assign po1779 = pi0275 & n19595;
  assign po1780 = ~pi0200 & ~pi1099;
  assign n19598 = ~pi0761 & pi0787;
  assign n19599 = pi0761 & ~pi0787;
  assign po1781 = n19598 | n19599;
  assign po1796 = pi1749 & pi1750;
  assign po0074 = 1'b1;
  assign po0144 = 1'b1;
  assign po0883 = ~pi1000;
  assign po0884 = ~pi1004;
  assign po0973 = ~pi1013;
  assign po0974 = ~pi1002;
  assign po0975 = ~pi1003;
  assign po0976 = ~pi1008;
  assign po0977 = ~pi1009;
  assign po0978 = ~pi1010;
  assign po0984 = ~pi1011;
  assign po1604 = ~pi1626;
  assign po1650 = ~pi1625;
  assign po1657 = ~pi1667;
  assign po1784 = ~pi1726;
  assign po1786 = ~pi1192;
  assign po1804 = ~pi1241;
  assign po1805 = ~pi1213;
  assign po1806 = ~pi1331;
  assign po1807 = ~pi0787;
  assign po1808 = ~pi1426;
  assign po1809 = ~pi1428;
  assign po1810 = ~pi1425;
  assign po1811 = ~pi0944;
  assign po1812 = ~pi1419;
  assign po1813 = ~pi0936;
  assign po1814 = ~pi0943;
  assign po1815 = ~pi0932;
  assign po1816 = ~pi0933;
  assign po1817 = ~pi1423;
  assign po1818 = ~pi0931;
  assign po1819 = ~pi0934;
  assign po1820 = ~pi0935;
  assign po0000 = pi0661;
  assign po0001 = pi0561;
  assign po0002 = pi0666;
  assign po0003 = pi0643;
  assign po0004 = pi0902;
  assign po0005 = pi0912;
  assign po0006 = pi0911;
  assign po0007 = pi0782;
  assign po0008 = pi0784;
  assign po0009 = pi0962;
  assign po0010 = pi0972;
  assign po0011 = pi0961;
  assign po0012 = pi0964;
  assign po0013 = pi0988;
  assign po0014 = pi1226;
  assign po0015 = pi0989;
  assign po0016 = pi0905;
  assign po0017 = pi0914;
  assign po0018 = pi0913;
  assign po0019 = pi0910;
  assign po0020 = pi0909;
  assign po0021 = pi0908;
  assign po0022 = pi0781;
  assign po0023 = pi0769;
  assign po0024 = pi0906;
  assign po0025 = pi0882;
  assign po0026 = pi0888;
  assign po0027 = pi0955;
  assign po0028 = pi0907;
  assign po0029 = pi0956;
  assign po0030 = pi0951;
  assign po0031 = pi0952;
  assign po0064 = pi0256;
  assign po0065 = pi1020;
  assign po0066 = pi1015;
  assign po0067 = pi1701;
  assign po0068 = pi1747;
  assign po0069 = pi0047;
  assign po0070 = pi0975;
  assign po0071 = pi0900;
  assign po0073 = pi1707;
  assign po0076 = pi0085;
  assign po0077 = pi0072;
  assign po0078 = pi0084;
  assign po0079 = pi0087;
  assign po0080 = pi0021;
  assign po0081 = pi0020;
  assign po0082 = pi0002;
  assign po0083 = pi0000;
  assign po0084 = pi0017;
  assign po0085 = pi0026;
  assign po0086 = pi0003;
  assign po0087 = pi0001;
  assign po0088 = pi0985;
  assign po0089 = pi0976;
  assign po0090 = pi1708;
  assign po0091 = pi1715;
  assign po0092 = pi1710;
  assign po0093 = pi1706;
  assign po0109 = pi1752;
  assign po0169 = pi0062;
  assign po0183 = pi1746;
  assign po0333 = pi0267;
  assign po0464 = pi0434;
  assign po0544 = pi0630;
  assign po0848 = pi1012;
  assign po0849 = pi1001;
  assign po0850 = pi1005;
  assign po0851 = pi1006;
  assign po0983 = pi0974;
  assign po1004 = pi0997;
  assign po1049 = pi0999;
  assign po1054 = pi1007;
  assign po1055 = pi0998;
  assign po1359 = pi1410;
  assign po1518 = pi1418;
  assign po1651 = pi1578;
  assign po1656 = pi1627;
  assign po1686 = pi0954;
  assign po1783 = pi1680;
  assign po1787 = pi1730;
  assign po1788 = pi1038;
  assign po1789 = pi1719;
  assign po1790 = pi1723;
  assign po1791 = pi1724;
  assign po1792 = pi1720;
  assign po1793 = pi1736;
  assign po1794 = pi1732;
  assign po1795 = pi1745;
  assign po1797 = pi1734;
  assign po1798 = pi1753;
  assign po1799 = pi1744;
  assign po1800 = pi1743;
  assign po1801 = pi0112;
  assign po1802 = pi1728;
  assign po1803 = pi1721;
  assign po1821 = pi1855;
  assign po1822 = pi1851;
  assign po1823 = pi1853;
  assign po1824 = pi1844;
  assign po1825 = pi1852;
  assign po1826 = pi0794;
  assign po1827 = pi1849;
  assign po1828 = pi1457;
  assign po1829 = pi1845;
  assign po1830 = pi1562;
  assign po1831 = pi1099;
  assign po1832 = pi1556;
  assign po1833 = pi1858;
  assign po1834 = pi1854;
  assign po1835 = pi1842;
  assign po1836 = pi1561;
  assign po1837 = pi1847;
  assign po1838 = pi1857;
  assign po1839 = pi1859;
  assign po1840 = pi1848;
  assign po1841 = pi1846;
  assign po1842 = pi1843;
  assign po1843 = pi1551;
  assign po1844 = pi1856;
  assign po1845 = pi1850;
endmodule


