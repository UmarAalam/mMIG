//Written by the Majority Logic Package Thu Apr 30 21:04:38 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15;
wire one, i0,i1,i2, i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17,i18,i19,i20,i21,i22,i23,i24,i25,i26,i27,i28,i29,i30,
i31, i32, i33, i34, i35, i36, i37, i38,i39, i40,i41, i42,i43,i44, i45, i46, i47, i48, i49,i50,i51, i52, i53, i54, i55, i56, i57, i58, i59
i60, i61, i62, i63, i64,i65,i65,i66,i67,i68,i69,i70,
i71,i72,i73,i74,i78,i79,i80,i81,i82,i83,i84,i85,i86,i87,i88,i89,i90,i91,i92,i93,i94,i95,
i96,i97,i98,i99,i100,i101, i102, i103, i104, i105, i106, i107, i108, i109, i110, i111, i112, i113, i114,
i115, i116, i117, i118, i119, i120, i121, i122, i123, i124, i125,
i126, i127, i128, i129, i130, i131, i131, i132, i133, i134, i135,
i136, i137, i138, i139, i140, i141, i142, i143, i144, i145, i146, i147, i148, i149,i150,
i151, i152, i153, i154, i155, i156, i157, i158, i159,
i160, i161, i162, i163, i164, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155;
assign i0 = ~(pi30 | pi31);
assign w0 = i0;
assign w1 = pi30 & pi31;
assign i1 = ~(pi28 | pi29);
assign i1 = ~(pi28 | pi29);
assign w2 = i1;
assign i2 = ~(pi30 | w2);
assign w3 = i2;
assign i3 = ~(w1 | w3);
assign w4 = i3;
assign w5 = pi30 & ~pi31;
assign w6 = (pi29 & w5) | (pi29 & w1179) | (w5 & w1179);
assign w7 = w1 & w2;
assign i4 = ~(w6 | w7);
assign w8 = i4;
assign w9 = ~w0 & w8;
assign w10 = pi28 & ~w5;
assign i5 = ~(pi26 | pi27);
assign w11 = i5;
assign w12 = ~pi28 & w11;
assign i6 = ~(w10 | w12);
assign w13 = i6;
assign w14 = ~w9 & w13;
assign w15 = w0 & w6;
assign w16 = pi30 & w2;
assign w17 = (pi31 & w2) | (pi31 & w1) | (w2 & w1);
assign w18 = ~w16 & w17;
assign i7 = ~(w15 | w18);
assign w19 = i7;
assign w20 = ~w14 & w19;
assign w21 = ~w14 & w1432;
assign w22 = (~pi26 & w14) | (~pi26 & w1180) | (w14 & w1180);
assign w23 = ~pi27 & w22;
assign w24 = (pi28 & w23) | (pi28 & w1433) | (w23 & w1433);
assign w25 = ~w23 & w1434;
assign i8 = ~(w24 | w25);
assign w26 = i8;
assign i9 = ~(pi24 | pi25);
assign w27 = i9;
assign i10 = ~(pi26 | w27);
assign w28 = i10;
assign w29 = ~w14 & w1181;
assign w30 = (w4 & w29) | (w4 & w1753) | (w29 & w1753);
assign w31 = ~w29 & w1182;
assign w32 = pi27 & ~w22;
assign w33 = ~w23 & ~w32;
assign w34 = ~w31 & ~w33;
assign w35 = (~w30 & w33) | (~w30 & w1754) | (w33 & w1754);
assign w36 = (w1183 & w33) | (w1183 & w1976) | (w33 & w1976);
assign w37 = w26 & ~w36;
assign w38 = w9 & ~w13;
assign w39 = ~w14 & w1617;
assign w40 = (~w15 & w9) | (~w15 & w1618) | (w9 & w1618);
assign w41 = ~w38 & w40;
assign w42 = ~w39 & w41;
assign w43 = (~w34 & w1435) | (~w34 & w1436) | (w1435 & w1436);
assign w44 = ~w37 & w43;
assign w45 = (w27 & w37) | (w27 & w1437) | (w37 & w1437);
assign w46 = ~w37 & w1438;
assign i11 = ~(w45 | w46);
assign w47 = i11;
assign w48 = pi26 & ~w47;
assign w49 = ~pi26 & w47;
assign i12 = ~(w48 | w49);
assign w50 = i12;
assign i13 = ~(w4 | w50);
assign w51 = i13;
assign w52 = w4 & w50;
assign i14 = ~(pi22 | pi23);
assign w53 = i14;
assign i15 = ~(pi24 | w53);
assign w54 = i15;
assign w55 = (w37 & w1439) | (w37 & w1440) | (w1439 & w1440);
assign w56 = ~w20 & w55;
assign w57 = (~w1440 & w1977) | (~w1440 & w1978) | (w1977 & w1978);
assign w58 = (~w37 & w1441) | (~w37 & w1442) | (w1441 & w1442);
assign i16 = ~(w45 | w58);
assign w59 = i16;
assign w60 = ~w57 & w59;
assign i17 = ~(w56 | w60);
assign w61 = i17;
assign i18 = ~(w52 | w61);
assign w62 = i18;
assign i19 = ~(w30 | w31);
assign w63 = i19;
assign w64 = (w63 & w37) | (w63 & w1755) | (w37 & w1755);
assign w65 = w33 & ~w64;
assign w66 = ~w33 & w64;
assign i20 = ~(w65 | w66);
assign w67 = i20;
assign w68 = (~w62 & w1443) | (~w62 & w1444) | (w1443 & w1444);
assign w69 = ~w62 & w1188;
assign w70 = ~w35 & w42;
assign i21 = ~(w26 | w70);
assign w71 = i21;
assign i22 = ~(w37 | w71);
assign w72 = i22;
assign w73 = (~w72 & w62) | (~w72 & w1445) | (w62 & w1445);
assign w74 = ~w68 & w73;
assign w75 = w53 & ~w74;
assign w76 = ~w44 & w74;
assign i23 = ~(w75 | w76);
assign w77 = i23;
assign w78 = pi24 & ~w77;
assign w79 = ~pi24 & w77;
assign i24 = ~(w78 | w79);
assign w80 = i24;
assign w81 = w20 & w80;
assign i25 = ~(pi22 | w74);
assign w82 = i25;
assign w83 = (pi23 & w74) | (pi23 & w1189) | (w74 & w1189);
assign i26 = ~(w75 | w83);
assign w84 = i26;
assign w85 = pi22 & w74;
assign i27 = ~(pi20 | pi21);
assign w86 = i27;
assign i28 = ~(pi22 | w86);
assign w87 = i28;
assign w88 = (~w87 & w37) | (~w87 & w1756) | (w37 & w1756);
assign w89 = ~w37 & w1757;
assign i29 = ~(w88 | w89);
assign w90 = i29;
assign w91 = (w90 & ~w74) | (w90 & w1190) | (~w74 & w1190);
assign w92 = w74 & w1191;
assign i30 = ~(w91 | w92);
assign w93 = i30;
assign w94 = w84 & ~w93;
assign w95 = (w88 & ~w74) | (w88 & w1758) | (~w74 & w1758);
assign i31 = ~(w94 | w95);
assign w96 = i31;
assign i32 = ~(w81 | w96);
assign w97 = i32;
assign w98 = ~w97 & w1192;
assign i33 = ~(w56 | w57);
assign w99 = i33;
assign w100 = (w59 & w74) | (w59 & w1759) | (w74 & w1759);
assign w101 = ~w74 & w1760;
assign i34 = ~(w100 | w101);
assign w102 = i34;
assign w103 = (~w102 & w97) | (~w102 & w1446) | (w97 & w1446);
assign w104 = (~w4 & w97) | (~w4 & w1193) | (w97 & w1193);
assign w105 = (~w97 & w1360) | (~w97 & w1447) | (w1360 & w1447);
assign w106 = ~w103 & w105;
assign w107 = w72 & w2059;
assign i35 = ~(w67 | w107);
assign w108 = i35;
assign i36 = ~(w68 | w69);
assign w109 = i36;
assign w110 = ~w108 & w109;
assign i37 = ~(w51 | w52);
assign w111 = i37;
assign w112 = ~w4 & w74;
assign i38 = ~(w61 | w74);
assign w113 = i38;
assign i39 = ~(w112 | w113);
assign w114 = i39;
assign w115 = w111 & ~w114;
assign w116 = ~w111 & w114;
assign i40 = ~(w115 | w116);
assign w117 = i40;
assign w118 = ~w110 & w117;
assign w119 = ~w106 & w118;
assign w120 = (~w97 & w1448) | (~w97 & w1449) | (w1448 & w1449);
assign w121 = (~w0 & w97) | (~w0 & w1450) | (w97 & w1450);
assign w122 = ~w120 & w121;
assign w123 = ~w110 & w122;
assign i41 = ~(w119 | w123);
assign w124 = i41;
assign w125 = (~w20 & w94) | (~w20 & w1761) | (w94 & w1761);
assign w126 = ~w94 & w1762;
assign i42 = ~(w125 | w126);
assign w127 = i42;
assign w128 = w124 & w1763;
assign i43 = ~(w80 | w124)    //saving #I = 2 
assign w129 = i43 | (~w80 & w1764) | (~w124 & w1764);
assign i44 = ~(w128 | w129);
assign w130 = i44;
assign i45 = ~(w4 | w130);
assign w131 = i45;
assign w132 = w4 & w130;
assign i46 = ~(w82 | w85);
assign w133 = i46;
assign i47 = ~(w124 | w133);
assign w134 = i47;
assign w135 = pi22 & w86;
assign i48 = ~(w87 | w135);
assign w136 = i48;
assign w137 = w124 & w136;
assign i49 = ~(w134 | w137);
assign w138 = i49;
assign w139 = ~w44 & w138;
assign w140 = w44 & ~w138;
assign w141 = (pi21 & ~w124) | (pi21 & w1194) | (~w124 & w1194);
assign w142 = w86 & w124;
assign i50 = ~(w141 | w142);
assign w143 = i50;
assign i51 = ~(pi18 | pi19);
assign w144 = i51;
assign w145 = ~pi20 & w144;
assign w146 = ~w74 & w145;
assign w147 = w74 & ~w145;
assign i52 = ~(w146 | w147);
assign w148 = i52;
assign i53 = ~(w148 | w124);
assign w149 = (i53) | (~w148 & w1195) | (~w124 & w1195);
assign w150 = w124 & w1196;
assign i54 = ~(w146 | w124);
assign w151 = (i54) | (~w146 & w1765) | (~w124 & w1765);
assign w152 = (w151 & ~w143) | (w151 & w1766) | (~w143 & w1766);
assign w153 = ~w20 & w2060;
assign w154 = (w84 & ~w124) | (w84 & w1767) | (~w124 & w1767);
assign w155 = w124 & w1768;
assign i55 = ~(w154 | w155);
assign w156 = i55;
assign w157 = w20 & ~w156;
assign w158 = (~w1197 & w1769) | (~w1197 & w1770) | (w1769 & w1770);
assign i56 = ~(w20 | w156);
assign w159 = i56;
assign w160 = (w1197 & w1771) | (w1197 & w1772) | (w1771 & w1772);
assign i57 = ~(w158 | w160);
assign w161 = i57;
assign i58 = ~(w132 | w161);
assign w162 = (i58) | (~w132 & w1198) | (~w161 & w1198);
assign w163 = (~w0 & w1199) | (~w0 & w162) | (w1199 & w162);
assign i58 = ~(w98 | w104);
assign w164 = i58;
assign w165 = (w102 & ~w124) | (w102 & w1773) | (~w124 & w1773);
assign w166 = w124 & w1774;
assign i59 = ~(w165 | w166);
assign w167 = i59;
assign w168 = (~w1452 & w1775) | (~w1452 & w1776) | (w1775 & w1776);
assign w169 = ~w162 & w1200;
assign i60 = ~(w106 | w122);
assign w170 = i60;
assign w171 = w110 & w117;
assign w172 = w170 & w171;
assign i61 = ~(w117 | w170);
assign w173 = i61;
assign i62 = ~(w172 | w173);
assign w174 = i62;
assign w175 = (w174 & w1201) | (w174 & w162) | (w1201 & w162);
assign w176 = ~w168 & w175;
assign i63 = ~(pi14 | pi15);
assign w177 = i63;
assign i64 = ~(w139 | w140);
assign w178 = i64;
assign w179 = ~w44 & w176;
assign i65 = ~(w152 | w176);
assign w180 = i65;
assign i66 = ~(w179 | w180);
assign w181 = i66;
assign w182 = w178 & ~w181;
assign w183 = ~w178 & w181;
assign i67 = ~(w182 | w183);
assign w184 = i67;
assign w185 = ~w20 & w184;
assign w186 = w20 & ~w184;
assign i68 = ~(w185 | w186);
assign w187 = i68;
assign i69 = ~(w149 | w150);
assign w188 = i69;
assign w189 = (w1777 & w2079) | (w1777 & w1453) | (w2079 & w1453);
assign w190 = (~w1453 & w2080) | (~w1453 & w2081) | (w2080 & w2081);
assign i70 = ~(w189 | w190);
assign w191 = i70;
assign w192 = (w144 & w168) | (w144 & w1202) | (w168 & w1202);
assign w193 = ~w168 & w1203;
assign i71 = ~(w192 | w193);
assign w194 = i71;
assign w195 = pi20 & w194;
assign i72 = ~(pi20 | w194);
assign w196 = i72;
assign i73 = ~(w195 | w196);
assign w197 = i73;
assign w198 = ~w74 & w197;
assign w199 = w74 & ~w197;
assign w200 = (~pi18 & w168) | (~pi18 & w1204) | (w168 & w1204);
assign w201 = (~w168 & w2149) | (~w168 & w2150) | (w2149 & w2150);
assign i74 = ~(w192 | w201);
assign w202 = i74;
assign w203 = ~w168 & w1205;
assign i75 = ~(pi16 | pi17);
assign w204 = i75;
assign i76 = ~(pi18 | w204);
assign w205 = i76;
assign w206 = w124 & ~w205;
assign w207 = ~w124 & w205;
assign i77 = ~(w206 | w207);
assign w208 = i77;
assign w209 = (w208 & w168) | (w208 & w1979) | (w168 & w1979);
assign w210 = ~w168 & w1980;
assign i78 = ~(w209 | w210);
assign w211 = i78;
assign w212 = w202 & ~w211;
assign w213 = ~w203 & w206;
assign i79 = ~(w212 | w213);
assign w214 = i79;
assign i80 = ~(w199 | w214);
assign w215 = i80;
assign w216 = w44 & w191;
assign w217 = (w216 & w215) | (w216 & w1206) | (w215 & w1206);
assign w218 = ~w44 & w191;
assign w219 = ~w215 & w1207;
assign i81 = ~(w217 | w219);
assign w220 = i81;
assign w221 = (~w44 & w215) | (~w44 & w1208) | (w215 & w1208);
assign w222 = w220 & ~w221;
assign i82 = ~(w161 | w176);
assign w223 = i82;
assign w224 = ~w139 & w2061;
assign i83 = ~(w153 | w224);
assign w225 = i83;
assign w226 = (w156 & w176) | (w156 & w1779) | (w176 & w1779);
assign i84 = ~(w223 | w226);
assign w227 = i84;
assign w228 = w220 & w1209;
assign w229 = (w4 & w228) | (w4 & w1210) | (w228 & w1210);
assign w230 = (~w228 & w1454) | (~w228 & w1455) | (w1454 & w1455);
assign w231 = ~w228 & w1211;
assign w232 = (w0 & w228) | (w0 & w1456) | (w228 & w1456);
assign w233 = ~w230 & w232;
assign i85 = ~(w4 | w161);
assign w234 = (i85) | (~w4 & w1780) | (~w161 & w1780);
assign w235 = w161 & w1781;
assign i86 = ~(w234 | w235);
assign w236 = i86;
assign w237 = ~w176 & w1782;
assign w238 = (~w130 & w176) | (~w130 & w1783) | (w176 & w1783);
assign i87 = ~(w237 | w238);
assign w239 = i87;
assign i88 = ~(w163 | w169);
assign w240 = i87;
assign w241 = (w167 & ~w240) | (w167 & w1784) | (~w240 & w1784);
assign w242 = ~w167 & w240;
assign i88 = ~(w241 | w242);
assign w243 = i88;
assign i89 = ~(w239 | w243);
assign w244 = i89;
assign w245 = ~w233 & w244;
assign w246 = (~w227 & w228) | (~w227 & w1212) | (w228 & w1212);
assign w247 = (~w228 & w1213) | (~w228 & w1214) | (w1213 & w1214);
assign w248 = ~w246 & w247;
assign i90 = ~(w243 | w248);
assign w249 = i90;
assign i91 = ~(w245 | w249);
assign w250 = i91;
assign w251 = ~w222 & w250;
assign i92 = ~(w20 | w250);
assign w252 = i92;
assign i93 = ~(w251 | w252);
assign w253 = i93;
assign w254 = w187 & ~w253;
assign w255 = ~w187 & w253;
assign i94 = ~(w254 | w255);
assign w256 = i94;
assign w257 = w4 & ~w256;
assign w258 = ~w4 & w256;
assign w259 = ~w220 & w250;
assign w260 = ~w215 & w1785;
assign i95 = ~(w221 | w260);
assign w261 = i95;
assign i96 = ~(w191 | w250);
assign w262 = (i96) | (~w191 & w1786) | (~w250 & w1786);
assign i97 = ~(w259 | w262);
assign w263 = i97;
assign i98 = ~(w198 | w199);
assign w264 = i98;
assign w265 = ~w214 & w250;
assign i99 = ~(w74 | w250);
assign w266 = i99;
assign i100 = ~(w265 | w266);
assign w267 = i100;
assign w268 = w264 & ~w267;
assign w269 = ~w264 & w267;
assign i101 = ~(w268 | w269);
assign w270 = i101;
assign w271 = w44 & ~w270;
assign w272 = ~w44 & w270;
assign w273 = w250 & w1787;
assign w274 = (w202 & ~w250) | (w202 & w1788) | (~w250 & w1788);

assign i102 = ~(w273 | w274);
assign w275 = i102;
assign i103 = ~(w200 | w203);
assign w276 = i103;
assign i104 = ~(w250 | w276);
assign w277 = i104;
assign w278 = pi18 & w204;
assign i105 = ~(w205 | w278);
assign w279 = i105;
assign w280 = w250 & w279;
assign i106 = ~(w277 | w280);
assign w281 = i106;
assign w282 = w124 & w281;
assign i107 = ~(w124 | w281);
assign w283 = i107;
assign w284 = ~w245 & w1215;
assign w285 = pi17 & ~w284;
assign w286 = ~w245 & w1216;
assign i108 = ~(w285 | w286);
assign w287 = i108;
assign w288 = ~pi16 & w177;
assign w289 = ~w176 & w288;
assign w290 = w176 & ~w288;
assign i109 = ~(w289 | w290);
assign w291 = i109;
assign i110 = ~(w291 | w1217);
assign w292 = (i110) | (~w291 & w1457) | (~w1217 & w1457);
assign w293 = w287 & ~w292;
assign w294 = w1217 & w1458;
assign i111 = ~(w289 | w294);
assign w295 = i111;
assign w296 = ~w293 & w295;
assign w297 = (~w282 & w296) | (~w282 & w1218) | (w296 & w1218);
assign w298 = w74 & ~w275;
assign w299 = ~w297 & w298;
assign i112 = ~(w74 | w275);
assign w300 = i112;
assign w301 = w297 & w300;
assign i113 = ~(w299 | w301);
assign w302 = i113;
assign i114 = ~(w74 | w297);
assign w303 = i114;
assign w304 = w302 & ~w303;
assign w305 = w302 & w1219;
assign w306 = w20 & w263;
assign w307 = ~w305 & w1220;
assign w308 = ~w20 & w263;
assign w309 = (w308 & w305) | (w308 & w1221) | (w305 & w1221);
assign i115 = ~(w307 | w309);
assign w310 = i115;
assign w311 = ~w305 & w1222;
assign w312 = w310 & ~w311;
assign w313 = (w1224 & ~w310) | (w1224 & w1459) | (~w310 & w1459);
assign i116 = ~(w229 | w231);
assign w314 = i116;
assign w315 = (w227 & ~w250) | (w227 & w1789) | (~w250 & w1789);
assign w316 = w250 & w1790;
assign i117 = ~(w315 | w316);
assign w317 = i117;
assign w318 = (w310 & w1619) | (w310 & w1620) | (w1619 & w1620);
assign w319 = (w310 & w1791) | (w310 & w1792) | (w1791 & w1792);
assign i118 = ~(w233 | w248);
assign w320 = i118;
assign w321 = w239 & ~w320;
assign w322 = ~w239 & w243;
assign w323 = w320 & w322;
assign i119 = ~(w321 | w323);
assign w324 = i119;
assign w325 = (~w310 & w2082) | (~w310 & w2083) | (w2082 & w2083);
assign w326 = ~w318 & w325;
assign w327 = (w177 & w318) | (w177 & w1228) | (w318 & w1228);
assign w328 = ~w318 & w1229;
assign i120 = ~(w327 | w328);
assign w329 = i120;
assign w330 = pi16 & w329;
assign i121 = ~(pi16 | w329);
assign w331 = i121;
assign i122 = ~(w330 | w331);
assign w332 = i122;
assign w333 = ~w176 & w332;
assign w334 = w176 & ~w332;
assign i123 = ~(w333 | w334);
assign w335 = i123;
assign w336 = (~pi14 & w318) | (~pi14 & w1230) | (w318 & w1230);
assign w337 = pi15 & ~w336;
assign i124 = ~(w327 | w337);
assign w338 = i124;
assign w339 = ~w318 & w1231;
assign i125 = ~(pi12 | pi13);
assign w340 = i125;
assign i126 = ~(pi14 | w340);
assign w341 = i126;
assign w342 = w250 & ~w341;
assign w343 = ~w250 & w341;
assign i127 = ~(w342 | w343);
assign w344 = i127;
assign w345 = ~w339 & w344;
assign w346 = w250 & w339;
assign i128 = ~(w345 | w346);
assign w347 = i128;
assign w348 = w338 & ~w347;
assign w349 = ~w339 & w342;
assign i129 = ~(w348 | w349);
assign w350 = i129;
assign i130 = ~(w310 | w326);
assign w351 = i130;
assign w352 = (w20 & w305) | (w20 & w1793) | (w305 & w1793);
assign i131 = ~(w311 | w352);
assign w353 = i131;
assign w354 = (~w263 & w326) | (~w263 & w1794) | (w326 & w1794);

assign w355 = ~w351 & ~w354;
assign w356 = ~w271 & ~w272;
assign w357 = ~w44 & w326;
assign w358 = ~w304 & ~w326;
assign w359 = ~w357 & ~w358;
assign w360 = w356 & ~w359;
assign w361 = ~w356 & w359;
assign w362 = ~w360 & ~w361;
assign w363 = w20 & ~w362;
assign w364 = ~w20 & w362;
assign w365 = ~w282 & ~w283;
assign w366 = ~w124 & w326;
assign w367 = w296 & ~w326;
assign w368 = ~w366 & ~w367;
assign w369 = w365 & ~w368;
assign w370 = ~w365 & w368;
assign w371 = ~w369 & ~w370;
assign w372 = ~w74 & ~w371;
assign w373 = w74 & w371;
assign w374 = ~w292 & ~w294;
assign w375 = (w1460 & w1621) | (w1460 & w1622) | (w1621 & w1622);
assign w376 = (~w1460 & w1623) | (~w1460 & w1624) | (w1623 & w1624);
assign w377 = ~w375 & ~w376;
assign w378 = ~w334 & ~w350;
assign w379 = ~w124 & w377;
assign w380 = (w379 & w378) | (w379 & w1232) | (w378 & w1232);
assign w381 = w124 & w377;
assign w382 = ~w378 & w1233;
assign w383 = ~w380 & ~w382;
assign w384 = (w124 & w378) | (w124 & w1234) | (w378 & w1234);
assign w385 = w383 & ~w384;
assign w386 = (~w373 & ~w383) | (~w373 & w1235) | (~w383 & w1235);
assign w387 = ~w302 & ~w326;
assign w388 = w74 & w297;
assign w389 = ~w303 & ~w388;
assign w390 = (w275 & w326) | (w275 & w1795) | (w326 & w1795);
assign w391 = ~w387 & ~w390;
assign w392 = w44 & w391;
assign w393 = (w392 & w386) | (w392 & w1236) | (w386 & w1236);
assign w394 = ~w44 & w391;
assign w395 = ~w386 & w1237;
assign w396 = ~w393 & ~w395;
assign w397 = (~w44 & w386) | (~w44 & w1238) | (w386 & w1238);
assign w398 = w396 & ~w397;
assign w399 = w4 & w355;
assign w400 = (w1239 & ~w396) | (w1239 & w1461) | (~w396 & w1461);
assign w401 = ~w4 & w355;
assign w402 = (w396 & w1462) | (w396 & w1463) | (w1462 & w1463);
assign w403 = ~w400 & ~w402;
assign w404 = (w1241 & ~w396) | (w1241 & w1464) | (~w396 & w1464);
assign w405 = (w396 & w1625) | (w396 & w1626) | (w1625 & w1626);
assign w406 = w403 & w405;
assign w407 = ~w313 & ~w319;
assign w408 = (~w317 & ~w407) | (~w317 & w1796) | (~w407 & w1796);
assign w409 = w317 & w407;
assign w410 = ~w408 & ~w409;
assign w411 = ~w257 & ~w258;
assign w412 = ~w4 & w326;
assign w413 = ~w312 & ~w326;
assign w414 = ~w412 & ~w413;
assign w415 = w411 & ~w414;
assign w416 = ~w411 & w414;
assign w417 = ~w415 & ~w416;
assign w418 = ~w410 & w417;
assign w419 = (w418 & ~w403) | (w418 & w1627) | (~w403 & w1627);
assign w420 = (w396 & w1628) | (w396 & w1629) | (w1628 & w1629);
assign w421 = (w396 & w1465) | (w396 & w1466) | (w1465 & w1466);
assign w422 = (~w396 & w1630) | (~w396 & w1631) | (w1630 & w1631);
assign w423 = ~w420 & w422;
assign w424 = ~w410 & w423;
assign w425 = ~w419 & ~w424;
assign w426 = ~w350 & w425;
assign w427 = ~w176 & ~w425;
assign w428 = ~w426 & ~w427;
assign w429 = w335 & ~w428;
assign w430 = ~w335 & w428;
assign w431 = ~w429 & ~w430;
assign w432 = w425 & w1797;
assign w433 = (w338 & ~w425) | (w338 & w1798) | (~w425 & w1798);
assign w434 = ~w432 & ~w433;
assign w435 = ~w336 & ~w339;
assign w436 = ~w425 & ~w435;
assign w437 = pi14 & w340;
assign w438 = ~w341 & ~w437;
assign w439 = w425 & w438;
assign w440 = ~w436 & ~w439;
assign w441 = w250 & w440;
assign w442 = ~w250 & ~w440;
assign w443 = ~w318 & ~w319;
assign w444 = ~pi10 & ~pi11;
assign w445 = pi12 & w444;
assign w446 = ~w406 & ~w423;
assign w447 = ~w406 & w1799;
assign w448 = pi12 & w410;
assign w449 = (~w444 & w410) | (~w444 & w1800) | (w410 & w1800);
assign w450 = ~w448 & w449;
assign w451 = (w446 & w1711) | (w446 & w1712) | (w1711 & w1712);
assign w452 = (~w446 & w2084) | (~w446 & w2085) | (w2084 & w2085);
assign w453 = ~pi12 & w425;
assign w454 = (pi13 & ~w425) | (pi13 & w1244) | (~w425 & w1244);
assign w455 = w340 & w425;
assign w456 = (w443 & ~w425) | (w443 & w1245) | (~w425 & w1245);
assign w457 = ~w454 & w456;
assign w458 = w451 & ~w457;
assign w459 = (~w443 & ~w425) | (~w443 & w1246) | (~w425 & w1246);
assign w460 = ~w454 & w459;
assign w461 = ~w451 & ~w460;
assign w462 = ~w458 & ~w461;
assign w463 = ~w452 & ~w462;
assign w464 = (~w442 & w462) | (~w442 & w1247) | (w462 & w1247);
assign w465 = ~w464 & w1248;
assign w466 = (~w434 & w464) | (~w434 & w1468) | (w464 & w1468);
assign w467 = (~w176 & w464) | (~w176 & w1249) | (w464 & w1249);
assign w468 = (~w464 & w1469) | (~w464 & w1470) | (w1469 & w1470);
assign w469 = ~w466 & w468;
assign w470 = (w124 & w466) | (w124 & w1250) | (w466 & w1250);
assign w471 = ~w403 & w425;
assign w472 = ~w404 & ~w421;
assign w473 = (~w355 & ~w425) | (~w355 & w1801) | (~w425 & w1801);
assign w474 = ~w471 & ~w473;
assign w475 = ~w363 & ~w364;
assign w476 = ~w398 & w425;
assign w477 = ~w20 & ~w425;
assign w478 = ~w476 & ~w477;
assign w479 = w475 & ~w478;
assign w480 = ~w475 & w478;
assign w481 = ~w479 & ~w480;
assign w482 = w4 & ~w481;
assign w483 = ~w4 & w481;
assign w484 = ~w396 & w425;
assign w485 = ~w386 & w1802;
assign w486 = ~w397 & ~w485;
assign w487 = (~w391 & ~w425) | (~w391 & w1803) | (~w425 & w1803);
assign w488 = ~w484 & ~w487;
assign w489 = ~w372 & ~w373;
assign w490 = ~w385 & w425;
assign w491 = ~w74 & ~w425;
assign w492 = ~w490 & ~w491;
assign w493 = w489 & ~w492;
assign w494 = ~w489 & w492;
assign w495 = ~w493 & ~w494;
assign w496 = w44 & ~w495;
assign w497 = ~w44 & w495;
assign w498 = w431 & ~w469;
assign w499 = ~w383 & w425;
assign w500 = ~w378 & w1804;
assign w501 = ~w384 & ~w500;
assign w502 = (~w377 & ~w425) | (~w377 & w1805) | (~w425 & w1805);
assign w503 = ~w499 & ~w502;
assign w504 = w74 & w503;
assign w505 = (w504 & w498) | (w504 & w1251) | (w498 & w1251);
assign w506 = ~w74 & w503;
assign w507 = ~w498 & w1252;
assign w508 = ~w505 & ~w507;
assign w509 = (~w74 & w498) | (~w74 & w1253) | (w498 & w1253);
assign w510 = w508 & ~w509;
assign w511 = (~w496 & ~w508) | (~w496 & w1806) | (~w508 & w1806);
assign w512 = w20 & w488;
assign w513 = (w1255 & ~w508) | (w1255 & w1634) | (~w508 & w1634);
assign w514 = ~w20 & w488;
assign w515 = (w508 & w1635) | (w508 & w1636) | (w1635 & w1636);
assign w516 = ~w513 & ~w515;
assign w517 = (w1257 & ~w508) | (w1257 & w1807) | (~w508 & w1807);
assign w518 = w516 & ~w517;
assign w519 = (w1259 & ~w516) | (w1259 & w1471) | (~w516 & w1471);
assign w520 = (w516 & w1713) | (w516 & w1714) | (w1713 & w1714);
assign w521 = (w516 & w1808) | (w516 & w1809) | (w1808 & w1809);
assign w522 = w417 & ~w446;
assign w523 = ~w418 & ~w447;
assign w524 = ~w522 & w523;
assign w525 = (~w516 & w1472) | (~w516 & w1473) | (w1472 & w1473);
assign w526 = ~w520 & w525;
assign w527 = ~w469 & ~w470;
assign w528 = (w431 & w526) | (w431 & w1810) | (w526 & w1810);
assign w529 = ~w526 & w1811;
assign w530 = ~w528 & ~w529;
assign w531 = ~w74 & ~w530;
assign w532 = w74 & w530;
assign w533 = ~w531 & ~w532;
assign w534 = ~w441 & ~w442;
assign w535 = ~w520 & w1637;
assign w536 = (w463 & w520) | (w463 & w1638) | (w520 & w1638);
assign w537 = (w534 & w535) | (w534 & w2086) | (w535 & w2086);
assign w538 = ~w535 & w2087;
assign w539 = ~w537 & ~w538;
assign w540 = ~w176 & ~w539;
assign w541 = w176 & w539;
assign w542 = w462 & ~w526;
assign w543 = ~w454 & ~w455;
assign w544 = ~w443 & w451;
assign w545 = ~w452 & ~w544;
assign w546 = (~w1474 & w2088) | (~w1474 & w2089) | (w2088 & w2089);
assign w547 = ~w542 & ~w546;
assign w548 = pi12 & ~w425;
assign w549 = ~w453 & ~w548;
assign w550 = (w446 & w1812) | (w446 & w1813) | (w1812 & w1813);
assign w551 = w444 & w2062;
assign w552 = ~w550 & ~w551;
assign w553 = (w552 & w520) | (w552 & w1475) | (w520 & w1475);
assign w554 = w549 & w553;
assign w555 = ~w549 & ~w553;
assign w556 = ~w554 & ~w555;
assign w557 = w326 & ~w556;
assign w558 = ~w326 & w556;
assign w559 = (~pi10 & w520) | (~pi10 & w1263) | (w520 & w1263);
assign w560 = pi11 & ~w559;
assign w561 = (w444 & w520) | (w444 & w1476) | (w520 & w1476);
assign w562 = ~w560 & ~w561;
assign w563 = ~w520 & w1264;
assign w564 = ~pi08 & ~pi09;
assign w565 = ~pi10 & ~w564;
assign w566 = w425 & ~w565;
assign w567 = ~w425 & w565;
assign w568 = ~w566 & ~w567;
assign w569 = ~w563 & ~w568;
assign w570 = ~w425 & w563;
assign w571 = ~w569 & ~w570;
assign w572 = w562 & w571;
assign w573 = ~w563 & w566;
assign w574 = ~w572 & ~w573;
assign w575 = ~w558 & w574;
assign w576 = (~w557 & ~w574) | (~w557 & w1814) | (~w574 & w1814);
assign w577 = ~w250 & w547;
assign w578 = ~w575 & w1265;
assign w579 = w250 & w547;
assign w580 = (w579 & w575) | (w579 & w1266) | (w575 & w1266);
assign w581 = ~w578 & ~w580;
assign w582 = (w1267 & ~w574) | (w1267 & w1477) | (~w574 & w1477);
assign w583 = w581 & ~w582;
assign w584 = (w581 & w1815) | (w581 & w1816) | (w1815 & w1816);
assign w585 = ~w465 & ~w467;
assign w586 = ~w526 & w1817;
assign w587 = (~w434 & w526) | (~w434 & w1818) | (w526 & w1818);
assign w588 = ~w586 & ~w587;
assign w589 = w124 & ~w588;
assign w590 = (w581 & w1478) | (w581 & w1479) | (w1478 & w1479);
assign w591 = ~w124 & ~w588;
assign w592 = (~w581 & w1480) | (~w581 & w1481) | (w1480 & w1481);
assign w593 = ~w590 & ~w592;
assign w594 = (w124 & w1271) | (w124 & w2063) | (w1271 & w2063);
assign w595 = w593 & ~w594;
assign w596 = ~w516 & ~w526;
assign w597 = w20 & ~w511;
assign w598 = ~w517 & ~w597;
assign w599 = (~w488 & w526) | (~w488 & w1819) | (w526 & w1819);
assign w600 = ~w596 & ~w599;
assign w601 = ~w496 & ~w497;
assign w602 = ~w44 & w526;
assign w603 = ~w510 & ~w526;
assign w604 = ~w602 & ~w603;
assign w605 = w601 & ~w604;
assign w606 = ~w601 & w604;
assign w607 = ~w605 & ~w606;
assign w608 = w20 & ~w607;
assign w609 = ~w20 & w607;
assign w610 = ~w508 & ~w526;
assign w611 = ~w498 & w1820;
assign w612 = ~w509 & ~w611;
assign w613 = (~w503 & w526) | (~w503 & w1821) | (w526 & w1821);
assign w614 = ~w610 & ~w613;
assign w615 = (w593 & w1822) | (w593 & w1823) | (w1822 & w1823);
assign w616 = w44 & w614;
assign w617 = (~w593 & w1725) | (~w593 & w1726) | (w1725 & w1726);
assign w618 = ~w44 & w614;
assign w619 = (w593 & w1727) | (w593 & w1728) | (w1727 & w1728);
assign w620 = ~w617 & ~w619;
assign w621 = (~w44 & w1275) | (~w44 & w2064) | (w1275 & w2064);
assign w622 = w620 & ~w621;
assign w623 = (w620 & w1482) | (w620 & w1483) | (w1482 & w1483);
assign w624 = (~w620 & w1639) | (~w620 & w1640) | (w1639 & w1640);
assign w625 = (w1277 & ~w620) | (w1277 & w1484) | (~w620 & w1484);
assign w626 = (w620 & w1641) | (w620 & w1642) | (w1641 & w1642);
assign w627 = ~w624 & w626;
assign w628 = ~w519 & ~w521;
assign w629 = (w474 & ~w628) | (w474 & w1824) | (~w628 & w1824);
assign w630 = ~w474 & w628;
assign w631 = ~w629 & ~w630;
assign w632 = ~w482 & ~w483;
assign w633 = ~w4 & w526;
assign w634 = ~w518 & ~w526;
assign w635 = ~w633 & ~w634;
assign w636 = w632 & ~w635;
assign w637 = ~w632 & w635;
assign w638 = ~w636 & ~w637;
assign w639 = ~w631 & w638;
assign w640 = ~w627 & w639;
assign w641 = (w620 & w1485) | (w620 & w1486) | (w1485 & w1486);
assign w642 = (~w620 & w1487) | (~w620 & w1488) | (w1487 & w1488);
assign w643 = ~w641 & w642;
assign w644 = ~w631 & w643;
assign w645 = ~w640 & ~w644;
assign w646 = ~w595 & w645;
assign w647 = ~w74 & ~w645;
assign w648 = ~w646 & ~w647;
assign w649 = w533 & ~w648;
assign w650 = ~w533 & w648;
assign w651 = ~w649 & ~w650;
assign w652 = w44 & ~w651;
assign w653 = ~w44 & w651;
assign w654 = ~w652 & ~w653;
assign w655 = ~w608 & ~w609;
assign w656 = ~w622 & w645;
assign w657 = ~w20 & ~w645;
assign w658 = ~w656 & ~w657;
assign w659 = w655 & ~w658;
assign w660 = ~w655 & w658;
assign w661 = ~w659 & ~w660;
assign w662 = w4 & ~w661;
assign w663 = ~w4 & w661;
assign w664 = ~w620 & w645;
assign w665 = w44 & w615;
assign w666 = ~w621 & ~w665;
assign w667 = (~w614 & ~w645) | (~w614 & w1825) | (~w645 & w1825);
assign w668 = ~w664 & ~w667;
assign w669 = ~w593 & w645;
assign w670 = ~w124 & w584;
assign w671 = ~w594 & ~w670;
assign w672 = (w588 & ~w645) | (w588 & w1826) | (~w645 & w1826);
assign w673 = ~w669 & ~w672;
assign w674 = ~w540 & ~w541;
assign w675 = ~w583 & w645;
assign w676 = ~w176 & ~w645;
assign w677 = ~w675 & ~w676;
assign w678 = w674 & ~w677;
assign w679 = ~w674 & w677;
assign w680 = ~w678 & ~w679;
assign w681 = ~w124 & ~w680;
assign w682 = w124 & w680;
assign w683 = ~w581 & w645;
assign w684 = ~w250 & ~w576;
assign w685 = ~w582 & ~w684;
assign w686 = (~w547 & ~w645) | (~w547 & w1827) | (~w645 & w1827);
assign w687 = ~w683 & ~w686;
assign w688 = ~w557 & ~w558;
assign w689 = ~w574 & w645;
assign w690 = ~w326 & ~w645;
assign w691 = ~w689 & ~w690;
assign w692 = w688 & ~w691;
assign w693 = ~w688 & w691;
assign w694 = ~w692 & ~w693;
assign w695 = ~w250 & ~w694;
assign w696 = w250 & w694;
assign w697 = w645 & w1715;
assign w698 = (w562 & ~w645) | (w562 & w1716) | (~w645 & w1716);
assign w699 = ~w697 & ~w698;
assign w700 = ~w559 & ~w563;
assign w701 = (~w700 & w640) | (~w700 & w1489) | (w640 & w1489);
assign w702 = pi10 & w564;
assign w703 = ~w565 & ~w702;
assign w704 = ~w640 & w1490;
assign w705 = ~w701 & w1643;
assign w706 = (~w425 & w701) | (~w425 & w1644) | (w701 & w1644);
assign w707 = (pi09 & w640) | (pi09 & w1491) | (w640 & w1491);
assign w708 = ~w640 & w1280;
assign w709 = ~w707 & ~w708;
assign w710 = ~w640 & w1281;
assign w711 = ~pi06 & ~pi07;
assign w712 = ~pi08 & w711;
assign w713 = ~w526 & w712;
assign w714 = w526 & ~w712;
assign w715 = ~w713 & ~w714;
assign w716 = ~w710 & ~w715;
assign w717 = w709 & ~w716;
assign w718 = ~w526 & w710;
assign w719 = (~w713 & ~w710) | (~w713 & w1492) | (~w710 & w1492);
assign w720 = ~w717 & w719;
assign w721 = (~w705 & w720) | (~w705 & w1282) | (w720 & w1282);
assign w722 = w326 & ~w699;
assign w723 = ~w721 & w722;
assign w724 = ~w326 & ~w699;
assign w725 = w721 & w724;
assign w726 = ~w723 & ~w725;
assign w727 = ~w326 & ~w721;
assign w728 = w726 & ~w727;
assign w729 = w726 & w1283;
assign w730 = w176 & w687;
assign w731 = ~w729 & w1284;
assign w732 = ~w176 & w687;
assign w733 = (w732 & w729) | (w732 & w1285) | (w729 & w1285);
assign w734 = ~w731 & ~w733;
assign w735 = ~w729 & w1286;
assign w736 = w734 & ~w735;
assign w737 = (~w681 & ~w734) | (~w681 & w1828) | (~w734 & w1828);
assign w738 = ~w74 & w673;
assign w739 = (w734 & w1493) | (w734 & w1494) | (w1493 & w1494);
assign w740 = w74 & w673;
assign w741 = (w1289 & ~w734) | (w1289 & w1495) | (~w734 & w1495);
assign w742 = ~w739 & ~w741;
assign w743 = (w1290 & ~w734) | (w1290 & w1829) | (~w734 & w1829);
assign w744 = w742 & ~w743;
assign w745 = (~w652 & ~w742) | (~w652 & w1830) | (~w742 & w1830);
assign w746 = w20 & w668;
assign w747 = (w1292 & ~w742) | (w1292 & w1645) | (~w742 & w1645);
assign w748 = ~w20 & w668;
assign w749 = (w742 & w1646) | (w742 & w1647) | (w1646 & w1647);
assign w750 = ~w747 & ~w749;
assign w751 = (w1294 & ~w742) | (w1294 & w1831) | (~w742 & w1831);
assign w752 = w750 & ~w751;
assign w753 = (w1296 & ~w750) | (w1296 & w1496) | (~w750 & w1496);
assign w754 = ~w623 & ~w625;
assign w755 = (w600 & ~w645) | (w600 & w1832) | (~w645 & w1832);
assign w756 = w645 & w1833;
assign w757 = ~w755 & ~w756;
assign w758 = (w750 & w2040) | (w750 & w2041) | (w2040 & w2041);
assign w759 = (w750 & w1834) | (w750 & w1835) | (w1834 & w1835);
assign w760 = ~w627 & ~w643;
assign w761 = w631 & w638;
assign w762 = w760 & w761;
assign w763 = ~w638 & ~w760;
assign w764 = ~w762 & ~w763;
assign w765 = (~w750 & w1497) | (~w750 & w1498) | (w1497 & w1498);
assign w766 = ~w758 & w765;
assign w767 = ~w758 & w1836;
assign w768 = (~w744 & w758) | (~w744 & w1837) | (w758 & w1837);
assign w769 = ~w767 & ~w768;
assign w770 = w654 & ~w769;
assign w771 = ~w654 & w769;
assign w772 = ~w770 & ~w771;
assign w773 = ~w20 & w772;
assign w774 = w20 & ~w772;
assign w775 = ~w773 & ~w774;
assign w776 = (~w742 & w758) | (~w742 & w1838) | (w758 & w1838);
assign w777 = w74 & ~w737;
assign w778 = ~w743 & ~w777;
assign w779 = (w778 & w758) | (w778 & w1839) | (w758 & w1839);
assign w780 = ~w673 & ~w779;
assign w781 = ~w776 & ~w780;
assign w782 = ~w681 & ~w682;
assign w783 = ~w758 & w1840;
assign w784 = (w736 & w758) | (w736 & w1841) | (w758 & w1841);
assign w785 = ~w783 & ~w784;
assign w786 = w782 & ~w785;
assign w787 = ~w782 & w785;
assign w788 = ~w786 & ~w787;
assign w789 = ~w74 & ~w788;
assign w790 = w74 & w788;
assign w791 = (~w734 & w758) | (~w734 & w1842) | (w758 & w1842);
assign w792 = (w176 & w729) | (w176 & w1843) | (w729 & w1843);
assign w793 = ~w735 & ~w792;
assign w794 = (w793 & w758) | (w793 & w1844) | (w758 & w1844);
assign w795 = ~w687 & ~w794;
assign w796 = ~w791 & ~w795;
assign w797 = ~w695 & ~w696;
assign w798 = ~w758 & w1845;
assign w799 = (w728 & w758) | (w728 & w1846) | (w758 & w1846);
assign w800 = ~w798 & ~w799;
assign w801 = w797 & ~w800;
assign w802 = ~w797 & w800;
assign w803 = ~w801 & ~w802;
assign w804 = ~w176 & ~w803;
assign w805 = w176 & w803;
assign w806 = ~w705 & ~w706;
assign w807 = ~w758 & w1847;
assign w808 = (w720 & w758) | (w720 & w1848) | (w758 & w1848);
assign w809 = ~w807 & ~w808;
assign w810 = w806 & ~w809;
assign w811 = ~w806 & w809;
assign w812 = ~w810 & ~w811;
assign w813 = ~w326 & ~w812;
assign w814 = w326 & w812;
assign w815 = ~w716 & ~w718;
assign w816 = (w2042 & w2090) | (w2042 & w1499) | (w2090 & w1499);
assign w817 = (~w1499 & w2091) | (~w1499 & w2092) | (w2091 & w2092);
assign w818 = ~w816 & ~w817;
assign w819 = (w711 & w758) | (w711 & w1300) | (w758 & w1300);
assign w820 = ~w758 & w1301;
assign w821 = ~w819 & ~w820;
assign w822 = pi08 & w821;
assign w823 = ~pi08 & ~w821;
assign w824 = ~w822 & ~w823;
assign w825 = ~w526 & w824;
assign w826 = w526 & ~w824;
assign w827 = (~pi06 & w758) | (~pi06 & w1302) | (w758 & w1302);
assign w828 = (~w758 & w1648) | (~w758 & w1649) | (w1648 & w1649);
assign w829 = ~w819 & ~w828;
assign w830 = ~w758 & w1303;
assign w831 = ~pi04 & ~pi05;
assign w832 = ~pi06 & ~w831;
assign w833 = w645 & ~w832;
assign w834 = ~w645 & w832;
assign w835 = ~w833 & ~w834;
assign w836 = (w835 & w758) | (w835 & w1650) | (w758 & w1650);
assign w837 = ~w758 & w1651;
assign w838 = ~w836 & ~w837;
assign w839 = (w833 & w758) | (w833 & w1849) | (w758 & w1849);
assign w840 = (~w839 & ~w829) | (~w839 & w2151) | (~w829 & w2151);
assign w841 = ~w826 & ~w840;
assign w842 = ~w425 & w818;
assign w843 = (w842 & w841) | (w842 & w1304) | (w841 & w1304);
assign w844 = w425 & w818;
assign w845 = ~w841 & w1305;
assign w846 = ~w843 & ~w845;
assign w847 = (w425 & w841) | (w425 & w1306) | (w841 & w1306);
assign w848 = w846 & ~w847;
assign w849 = (~w814 & ~w846) | (~w814 & w1307) | (~w846 & w1307);
assign w850 = (~w726 & w758) | (~w726 & w1850) | (w758 & w1850);
assign w851 = w326 & w721;
assign w852 = ~w727 & ~w851;
assign w853 = (w852 & w758) | (w852 & w1851) | (w758 & w1851);
assign w854 = w699 & ~w853;
assign w855 = ~w850 & ~w854;
assign w856 = ~w854 & w1852;
assign w857 = (~w846 & w1981) | (~w846 & w1982) | (w1981 & w1982);
assign w858 = ~w854 & w1853;
assign w859 = (w846 & w1983) | (w846 & w1984) | (w1983 & w1984);
assign w860 = ~w857 & ~w859;
assign w861 = (w250 & w849) | (w250 & w1310) | (w849 & w1310);
assign w862 = (w860 & w1854) | (w860 & w1855) | (w1854 & w1855);
assign w863 = ~w795 & w1856;
assign w864 = (~w860 & w1500) | (~w860 & w1501) | (w1500 & w1501);
assign w865 = ~w795 & w1857;
assign w866 = (w860 & w1502) | (w860 & w1503) | (w1502 & w1503);
assign w867 = ~w864 & ~w866;
assign w868 = (w124 & w1314) | (w124 & w2065) | (w1314 & w2065);
assign w869 = (w867 & w1858) | (w867 & w1859) | (w1858 & w1859);
assign w870 = ~w780 & w1860;
assign w871 = (w867 & w1652) | (w867 & w1653) | (w1652 & w1653);
assign w872 = ~w780 & w1861;
assign w873 = (~w867 & w1654) | (~w867 & w1655) | (w1654 & w1655);
assign w874 = ~w871 & ~w873;
assign w875 = (~w44 & w1318) | (~w44 & w2066) | (w1318 & w2066);
assign w876 = w874 & ~w875;
assign w877 = (~w750 & w758) | (~w750 & w1862) | (w758 & w1862);
assign w878 = w20 & ~w745;
assign w879 = ~w751 & ~w878;
assign w880 = (w879 & w758) | (w879 & w1863) | (w758 & w1863);
assign w881 = ~w668 & ~w880;
assign w882 = ~w877 & ~w881;
assign w883 = (w874 & w1504) | (w874 & w1505) | (w1504 & w1505);
assign w884 = (~w874 & w1729) | (~w874 & w1730) | (w1729 & w1730);
assign w885 = (w1320 & ~w874) | (w1320 & w1506) | (~w874 & w1506);
assign w886 = (w874 & w1731) | (w874 & w1732) | (w1731 & w1732);
assign w887 = ~w884 & w886;
assign w888 = ~w753 & ~w759;
assign w889 = (~w757 & ~w888) | (~w757 & w1864) | (~w888 & w1864);
assign w890 = w757 & w888;
assign w891 = ~w889 & ~w890;
assign w892 = ~w662 & ~w663;
assign w893 = ~w758 & w1865;
assign w894 = (~w752 & w758) | (~w752 & w1866) | (w758 & w1866);
assign w895 = ~w893 & ~w894;
assign w896 = w892 & ~w895;
assign w897 = ~w892 & w895;
assign w898 = ~w896 & ~w897;
assign w899 = ~w891 & w898;
assign w900 = ~w887 & w899;
assign w901 = (w874 & w1507) | (w874 & w1508) | (w1507 & w1508);
assign w902 = (~w874 & w1509) | (~w874 & w1510) | (w1509 & w1510);
assign w903 = ~w901 & w902;
assign w904 = ~w891 & w903;
assign w905 = ~w900 & ~w904;
assign w906 = ~w876 & w905;
assign w907 = ~w20 & ~w905;
assign w908 = ~w906 & ~w907;
assign w909 = w775 & ~w908;
assign w910 = ~w775 & w908;
assign w911 = ~w909 & ~w910;
assign w912 = ~w4 & w911;
assign w913 = w4 & ~w911;
assign w914 = ~w912 & ~w913;
assign w915 = (~w74 & ~w867) | (~w74 & w1867) | (~w867 & w1867);
assign w916 = w867 & w1868;
assign w917 = ~w915 & ~w916;
assign w918 = w905 & w1869;
assign w919 = (~w788 & ~w905) | (~w788 & w1870) | (~w905 & w1870);
assign w920 = ~w918 & ~w919;
assign w921 = ~w44 & ~w920;
assign w922 = w44 & w920;
assign w923 = (~w176 & ~w860) | (~w176 & w1871) | (~w860 & w1871);
assign w924 = w860 & w1872;
assign w925 = ~w923 & ~w924;
assign w926 = w905 & w1873;
assign w927 = (~w803 & ~w905) | (~w803 & w1874) | (~w905 & w1874);
assign w928 = ~w926 & ~w927;
assign w929 = w124 & ~w928;
assign w930 = ~w124 & w928;
assign w931 = ~w860 & w905;
assign w932 = ~w849 & w1875;
assign w933 = ~w861 & ~w932;
assign w934 = (~w855 & ~w905) | (~w855 & w1876) | (~w905 & w1876);
assign w935 = ~w931 & ~w934;
assign w936 = ~w813 & ~w814;
assign w937 = ~w848 & w905;
assign w938 = ~w326 & ~w905;
assign w939 = ~w937 & ~w938;
assign w940 = w936 & ~w939;
assign w941 = ~w936 & w939;
assign w942 = ~w940 & ~w941;
assign w943 = ~w250 & ~w942;
assign w944 = w250 & w942;
assign w945 = ~w846 & w905;
assign w946 = ~w841 & w1877;
assign w947 = ~w847 & ~w946;
assign w948 = (~w818 & ~w905) | (~w818 & w1878) | (~w905 & w1878);
assign w949 = ~w945 & ~w948;
assign w950 = ~w825 & ~w826;
assign w951 = ~w900 & w1656;
assign w952 = (~w526 & w900) | (~w526 & w1657) | (w900 & w1657);
assign w953 = ~w951 & ~w952;
assign w954 = w950 & ~w953;
assign w955 = ~w950 & w953;
assign w956 = ~w954 & ~w955;
assign w957 = ~w425 & ~w956;
assign w958 = w425 & w956;
assign w959 = w1658 & w1733;
assign w960 = (w829 & ~w1658) | (w829 & w1734) | (~w1658 & w1734);
assign w961 = ~w959 & ~w960;
assign w962 = ~w827 & ~w830;
assign w963 = (~w962 & w900) | (~w962 & w1511) | (w900 & w1511);
assign w964 = pi06 & w831;
assign w965 = ~w832 & ~w964;
assign w966 = ~w900 & w1512;
assign w967 = ~w963 & ~w966;
assign w968 = w645 & w967;
assign w969 = ~w645 & ~w967;
assign w970 = (pi05 & w900) | (pi05 & w1513) | (w900 & w1513);
assign w971 = ~w900 & w1323;
assign w972 = ~w970 & ~w971;
assign w973 = ~w900 & w1324;
assign w974 = ~pi02 & ~pi03;
assign w975 = ~pi04 & w974;
assign w976 = (w975 & w758) | (w975 & w1879) | (w758 & w1879);
assign w977 = ~w758 & w1880;
assign w978 = ~w976 & ~w977;
assign w979 = (~w978 & w900) | (~w978 & w1659) | (w900 & w1659);
assign w980 = w972 & ~w979;
assign w981 = ~w766 & w973;
assign w982 = (~w976 & ~w973) | (~w976 & w1514) | (~w973 & w1514);
assign w983 = ~w980 & w982;
assign w984 = (~w968 & w983) | (~w968 & w1325) | (w983 & w1325);
assign w985 = w526 & ~w961;
assign w986 = ~w984 & w985;
assign w987 = ~w526 & ~w961;
assign w988 = w984 & w987;
assign w989 = ~w986 & ~w988;
assign w990 = ~w526 & ~w984;
assign w991 = w989 & ~w990;
assign w992 = w989 & w1326;
assign w993 = w326 & w949;
assign w994 = ~w992 & w1327;
assign w995 = ~w326 & w949;
assign w996 = (w995 & w992) | (w995 & w1328) | (w992 & w1328);
assign w997 = ~w994 & ~w996;
assign w998 = ~w992 & w1329;
assign w999 = w997 & ~w998;
assign w1000 = (~w943 & ~w997) | (~w943 & w1881) | (~w997 & w1881);
assign w1001 = w176 & w935;
assign w1002 = (w1331 & ~w997) | (w1331 & w1515) | (~w997 & w1515);
assign w1003 = ~w176 & w935;
assign w1004 = (w997 & w1516) | (w997 & w1517) | (w1516 & w1517);
assign w1005 = ~w1002 & ~w1004;
assign w1006 = (w1333 & ~w997) | (w1333 & w1882) | (~w997 & w1882);
assign w1007 = w1005 & ~w1006;
assign w1008 = (w1005 & w1883) | (w1005 & w1884) | (w1883 & w1884);
assign w1009 = ~w867 & w905;
assign w1010 = ~w124 & w862;
assign w1011 = ~w868 & ~w1010;
assign w1012 = (~w796 & ~w905) | (~w796 & w1885) | (~w905 & w1885);
assign w1013 = ~w1009 & ~w1012;
assign w1014 = w74 & w1013;
assign w1015 = (~w1005 & w1660) | (~w1005 & w1661) | (w1660 & w1661);
assign w1016 = ~w74 & w1013;
assign w1017 = (w1005 & w1662) | (w1005 & w1663) | (w1662 & w1663);
assign w1018 = ~w1015 & ~w1017;
assign w1019 = (~w74 & w1337) | (~w74 & w2067) | (w1337 & w2067);
assign w1020 = w1018 & ~w1019;
assign w1021 = (w1018 & w1886) | (w1018 & w1887) | (w1886 & w1887);
assign w1022 = ~w874 & w905;
assign w1023 = w44 & w869;
assign w1024 = ~w875 & ~w1023;
assign w1025 = (~w781 & ~w905) | (~w781 & w1888) | (~w905 & w1888);
assign w1026 = ~w1022 & ~w1025;
assign w1027 = ~w20 & w1026;
assign w1028 = (w1018 & w1518) | (w1018 & w1519) | (w1518 & w1519);
assign w1029 = w20 & w1026;
assign w1030 = (~w1018 & w1520) | (~w1018 & w1521) | (w1520 & w1521);
assign w1031 = ~w1028 & ~w1030;
assign w1032 = (~w20 & w1341) | (~w20 & w2068) | (w1341 & w2068);
assign w1033 = w1031 & ~w1032;
assign w1034 = (~w913 & ~w1031) | (~w913 & w1889) | (~w1031 & w1889);
assign w1035 = (w1343 & ~w1031) | (w1343 & w1890) | (~w1031 & w1890);
assign w1036 = ~w883 & ~w885;
assign w1037 = (w882 & ~w905) | (w882 & w1891) | (~w905 & w1891);
assign w1038 = w905 & w1892;
assign w1039 = ~w1037 & ~w1038;
assign w1040 = (w1031 & w1664) | (w1031 & w1665) | (w1664 & w1665);
assign w1041 = (w1031 & w1893) | (w1031 & w1894) | (w1893 & w1894);
assign w1042 = ~w887 & ~w903;
assign w1043 = ~w898 & w1042;
assign w1044 = (~w899 & w1042) | (~w899 & w1895) | (w1042 & w1895);
assign w1045 = ~w1043 & w1044;
assign w1046 = (~w1031 & w1666) | (~w1031 & w1667) | (w1666 & w1667);
assign w1047 = ~w1040 & w1046;
assign w1048 = ~w4 & w1047;
assign w1049 = ~w1033 & ~w1047;
assign w1050 = ~w1048 & ~w1049;
assign w1051 = w914 & ~w1050;
assign w1052 = ~w914 & w1050;
assign w1053 = ~w1051 & ~w1052;
assign w1054 = ~w0 & w1053;
assign w1055 = ~w943 & ~w944;
assign w1056 = ~w250 & w1047;
assign w1057 = w999 & ~w1047;
assign w1058 = ~w1056 & ~w1057;
assign w1059 = w1055 & ~w1058;
assign w1060 = ~w1055 & w1058;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = w176 & w1061;
assign w1063 = ~w997 & ~w1047;
assign w1064 = (w326 & w992) | (w326 & w1896) | (w992 & w1896);
assign w1065 = ~w998 & ~w1064;
assign w1066 = (~w949 & w1047) | (~w949 & w1897) | (w1047 & w1897);
assign w1067 = ~w1063 & ~w1066;
assign w1068 = w250 & w1067;
assign w1069 = ~w957 & ~w958;
assign w1070 = ~w425 & w1047;
assign w1071 = w991 & ~w1047;
assign w1072 = ~w1070 & ~w1071;
assign w1073 = w1069 & ~w1072;
assign w1074 = ~w1069 & w1072;
assign w1075 = ~w1073 & ~w1074;
assign w1076 = ~w326 & ~w1075;
assign w1077 = (~w974 & w1040) | (~w974 & w1347) | (w1040 & w1347);
assign w1078 = ~w1040 & w1348;
assign w1079 = ~w1077 & ~w1078;
assign w1080 = pi04 & ~w1079;
assign w1081 = ~pi04 & w1079;
assign w1082 = ~w1080 & ~w1081;
assign w1083 = ~w766 & w1082;
assign w1084 = ~pi00 & ~pi01;
assign w1085 = ~pi02 & w1084;
assign w1086 = w905 & w1085;
assign w1087 = (w1523 & w2093) | (w1523 & w1349) | (w2093 & w1349);
assign w1088 = ~w905 & ~w1085;
assign w1089 = pi03 & w1047;
assign w1090 = (~w1349 & w2094) | (~w1349 & w2095) | (w2094 & w2095);
assign w1091 = ~w1089 & w1090;
assign w1092 = ~w1086 & ~w1087;
assign w1093 = ~w1091 & w1092;
assign w1094 = ~w1083 & w1093;
assign w1095 = ~w979 & ~w981;
assign w1096 = (w1524 & w2096) | (w1524 & w1350) | (w2096 & w1350);
assign w1097 = (~w1350 & w2097) | (~w1350 & w2098) | (w2097 & w2098);
assign w1098 = ~w1096 & ~w1097;
assign w1099 = ~w645 & ~w1098;
assign w1100 = w766 & ~w1082;
assign w1101 = ~w1099 & ~w1100;
assign w1102 = ~w1094 & w1101;
assign w1103 = ~w989 & ~w1047;
assign w1104 = w526 & w984;
assign w1105 = ~w990 & ~w1104;
assign w1106 = (~w1351 & w1668) | (~w1351 & w1669) | (w1668 & w1669);
assign w1107 = ~w1103 & ~w1106;
assign w1108 = w425 & w1107;
assign w1109 = ~w968 & ~w969;
assign w1110 = ~w1040 & w1352;
assign w1111 = (w983 & w1040) | (w983 & w1353) | (w1040 & w1353);
assign w1112 = ~w1110 & ~w1111;
assign w1113 = w1109 & ~w1112;
assign w1114 = ~w1109 & w1112;
assign w1115 = ~w1113 & ~w1114;
assign w1116 = ~w526 & ~w1115;
assign w1117 = w645 & w1098;
assign w1118 = ~w1108 & ~w1117;
assign w1119 = ~w1116 & w1118;
assign w1120 = ~w1102 & w1119;
assign w1121 = (~w425 & w1103) | (~w425 & w2025) | (w1103 & w2025);
assign w1122 = (w1103 & w2026) | (w1103 & w2027) | (w2026 & w2027);
assign w1123 = (~w1121 & ~w1115) | (~w1121 & w1526) | (~w1115 & w1526);
assign w1124 = ~w250 & ~w1067;
assign w1125 = (w1120 & w1985) | (w1120 & w1986) | (w1985 & w1986);
assign w1126 = ~w929 & ~w930;
assign w1127 = ~w124 & w1047;
assign w1128 = w1007 & ~w1047;
assign w1129 = ~w1127 & ~w1128;
assign w1130 = w1126 & ~w1129;
assign w1131 = ~w1126 & w1129;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = ~w176 & ~w1061;
assign w1134 = ~w1005 & ~w1047;
assign w1135 = w176 & ~w1000;
assign w1136 = ~w1006 & ~w1135;
assign w1137 = (~w935 & w1047) | (~w935 & w1899) | (w1047 & w1899);
assign w1138 = ~w1134 & ~w1137;
assign w1139 = w124 & w1138;
assign w1140 = (~w1139 & w1132) | (~w1139 & w1900) | (w1132 & w1900);
assign w1141 = ~w1133 & w1140;
assign w1142 = ~w1018 & ~w1047;
assign w1143 = w74 & w1008;
assign w1144 = ~w1019 & ~w1143;
assign w1145 = (~w1013 & w1047) | (~w1013 & w1901) | (w1047 & w1901);
assign w1146 = ~w1142 & ~w1145;
assign w1147 = w44 & ~w1146;
assign w1148 = ~w124 & ~w1138;
assign w1149 = (w1148 & w1132) | (w1148 & w1902) | (w1132 & w1902);
assign w1150 = (~w1147 & ~w1132) | (~w1147 & w1987) | (~w1132 & w1987);
assign w1151 = ~w1149 & w1150;
assign w1152 = ~w44 & w1146;
assign w1153 = ~w921 & ~w922;
assign w1154 = ~w44 & w1047;
assign w1155 = ~w1020 & ~w1047;
assign w1156 = ~w1154 & ~w1155;
assign w1157 = w1153 & ~w1156;
assign w1158 = ~w1153 & w1156;
assign w1159 = ~w1157 & ~w1158;
assign w1160 = ~w20 & w1159;
assign w1161 = ~w1031 & ~w1047;
assign w1162 = w20 & w1021;
assign w1163 = ~w1032 & ~w1162;
assign w1164 = (~w1026 & w1047) | (~w1026 & w1903) | (w1047 & w1903);
assign w1165 = ~w1161 & ~w1164;
assign w1166 = ~w4 & w1165;
assign w1167 = ~w1152 & ~w1166;
assign w1168 = ~w1160 & w1167;
assign w1169 = w4 & ~w1165;
assign w1170 = w20 & ~w1159;
assign w1171 = (~w1169 & ~w1170) | (~w1169 & w1670) | (~w1170 & w1670);
assign w1172 = (~w1527 & w1988) | (~w1527 & w1989) | (w1988 & w1989);
assign w1173 = ~w1034 & w1039;
assign w1174 = (~w1039 & w1035) | (~w1039 & w1905) | (w1035 & w1905);
assign w1175 = ~w1040 & ~w1041;
assign w1176 = ~w1174 & w1175;
assign w1177 = (w1053 & w1906) | (w1053 & w1907) | (w1906 & w1907);
assign w1178 = ~w1172 & w1177;
assign w1179 = pi28 & pi29;
assign w1180 = ~w19 & ~pi26;
assign w1181 = w19 & pi26;
assign w1182 = ~w28 & ~w4;
assign w1183 = (~w29 & w1908) | (~w29 & w1909) | (w1908 & w1909);
assign w1184 = (w1360 & w29) | (w1360 & w1529) | (w29 & w1529);
assign w1185 = w53 & ~pi24;
assign w1186 = pi24 & pi25;
assign w1187 = ~w50 & w1213;
assign w1188 = (w0 & w50) | (w0 & w1360) | (w50 & w1360);
assign w1189 = pi22 & pi23;
assign w1190 = ~pi22 & w90;
assign w1191 = (pi22 & w37) | (pi22 & w1910) | (w37 & w1910);
assign w1192 = (w4 & w80) | (w4 & w1361) | (w80 & w1361);
assign w1193 = ~w80 & w1362;
assign w1194 = pi20 & pi21;
assign w1195 = ~pi20 & ~w148;
assign w1196 = pi20 & ~w74;
assign w1197 = w140 & ~w139;
assign w1198 = (~w1197 & w2099) | (~w1197 & w2100) | (w2099 & w2100);
assign w1199 = w131 & ~w0;
assign w1200 = (w0 & w130) | (w0 & w1360) | (w130 & w1360);
assign w1201 = w174 & ~w1200;
assign w1202 = (w161 & w1911) | (w161 & w1912) | (w1911 & w1912);
assign w1203 = (~w161 & w1913) | (~w161 & w1914) | (w1913 & w1914);
assign w1204 = (w161 & w1915) | (w161 & w1916) | (w1915 & w1916);
assign w1205 = (~w161 & w1917) | (~w161 & w1918) | (w1917 & w1918);
assign w1206 = w198 & w216;
assign w1207 = ~w198 & w218;
assign w1208 = w197 & w1372;
assign w1209 = ~w221 & ~w185;
assign w1210 = ~w184 & w1361;
assign w1211 = (~w4 & w184) | (~w4 & w1362) | (w184 & w1362);
assign w1212 = ~w227 & ~w1211;
assign w1213 = (~w0 & w3) | (~w0 & w1919) | (w3 & w1919);
assign w1214 = (~w0 & w184) | (~w0 & w1583) | (w184 & w1583);
assign w1215 = (~pi16 & ~w248) | (~pi16 & w1373) | (~w248 & w1373);
assign w1216 = (w204 & ~w248) | (w204 & w1530) | (~w248 & w1530);
assign w1217 = (pi16 & ~w248) | (pi16 & w1920) | (~w248 & w1920);
assign w1218 = w283 & ~w282;
assign w1219 = ~w303 & ~w272;
assign w1220 = (w306 & w270) | (w306 & w1921) | (w270 & w1921);
assign w1221 = ~w270 & w1922;
assign w1222 = (~w20 & w270) | (~w20 & w1671) | (w270 & w1671);
assign w1223 = (~w258 & w305) | (~w258 & w1374) | (w305 & w1374);
assign w1224 = (~w0 & w256) | (~w0 & w1923) | (w256 & w1923);
assign w1225 = ~w256 & w1360;
assign w1226 = w324 & ~w0;
assign w1227 = (w324 & w256) | (w324 & w1924) | (w256 & w1924);
assign w1228 = (w310 & w1531) | (w310 & w1532) | (w1531 & w1532);
assign w1229 = (~w310 & w1533) | (~w310 & w1534) | (w1533 & w1534);
assign w1230 = (w310 & w1535) | (w310 & w1536) | (w1535 & w1536);
assign w1231 = (~w310 & w1537) | (~w310 & w1538) | (w1537 & w1538);
assign w1232 = w333 & w379;
assign w1233 = ~w333 & w381;
assign w1234 = w332 & w1383;
assign w1235 = w384 & ~w373;
assign w1236 = ~w371 & w1925;
assign w1237 = (w394 & w371) | (w394 & w1926) | (w371 & w1926);
assign w1238 = ~w371 & w1372;
assign w1239 = (w399 & w362) | (w399 & w1927) | (w362 & w1927);
assign w1240 = ~w362 & w1928;
assign w1241 = (~w4 & w362) | (~w4 & w1362) | (w362 & w1362);
assign w1242 = ~w362 & w1361;
assign w1243 = (w417 & ~w403) | (w417 & w1672) | (~w403 & w1672);
assign w1244 = pi12 & pi13;
assign w1245 = ~w340 & w443;
assign w1246 = ~w340 & ~w443;
assign w1247 = (w452 & w440) | (w452 & w1929) | (w440 & w1929);
assign w1248 = (w176 & ~w440) | (w176 & w1539) | (~w440 & w1539);
assign w1249 = w440 & w1540;
assign w1250 = (w462 & w1930) | (w462 & w1931) | (w1930 & w1931);
assign w1251 = (w466 & w1387) | (w466 & w1388) | (w1387 & w1388);
assign w1252 = (~w466 & w1389) | (~w466 & w1390) | (w1389 & w1390);
assign w1253 = (w466 & w1391) | (w466 & w1392) | (w1391 & w1392);
assign w1254 = (~w498 & w1393) | (~w498 & w1394) | (w1393 & w1394);
assign w1255 = (w512 & w495) | (w512 & w1932) | (w495 & w1932);
assign w1256 = ~w495 & w1933;
assign w1257 = (~w20 & w495) | (~w20 & w1671) | (w495 & w1671);
assign w1258 = (w508 & w1673) | (w508 & w1674) | (w1673 & w1674);
assign w1259 = (~w0 & w481) | (~w0 & w1923) | (w481 & w1923);
assign w1260 = ~w481 & w1360;
assign w1261 = ~w524 & ~w0;
assign w1262 = (~w524 & w481) | (~w524 & w1934) | (w481 & w1934);
assign w1263 = (w516 & w1541) | (w516 & w1542) | (w1541 & w1542);
assign w1264 = (~w516 & w1543) | (~w516 & w1544) | (w1543 & w1544);
assign w1265 = ~w557 & w577;
assign w1266 = w557 & w579;
assign w1267 = (w250 & w556) | (w250 & w1400) | (w556 & w1400);
assign w1268 = w582 & ~w541;
assign w1269 = ~w540 & w589;
assign w1270 = w540 & w591;
assign w1271 = ~w539 & w1383;
assign w1272 = (~w581 & w1675) | (~w581 & w1676) | (w1675 & w1676);
assign w1273 = w531 & w616;
assign w1274 = ~w531 & w618;
assign w1275 = ~w530 & w1372;
assign w1276 = ~w607 & w1361;
assign w1277 = (~w4 & w607) | (~w4 & w1362) | (w607 & w1362);
assign w1278 = ~w600 & ~w1277;
assign w1279 = (~w0 & w607) | (~w0 & w1583) | (w607 & w1583);
assign w1280 = (w564 & ~w643) | (w564 & w1545) | (~w643 & w1545);
assign w1281 = (pi08 & ~w643) | (pi08 & w1546) | (~w643 & w1546);
assign w1282 = w706 & ~w705;
assign w1283 = ~w727 & ~w696;
assign w1284 = (w730 & w694) | (w730 & w1935) | (w694 & w1935);
assign w1285 = ~w694 & w1936;
assign w1286 = (~w176 & w694) | (~w176 & w1540) | (w694 & w1540);
assign w1287 = (~w682 & w729) | (~w682 & w1406) | (w729 & w1406);
assign w1288 = ~w680 & w1937;
assign w1289 = (w740 & w680) | (w740 & w1938) | (w680 & w1938);
assign w1290 = (~w74 & w680) | (~w74 & w1391) | (w680 & w1391);
assign w1291 = (w734 & w1547) | (w734 & w1548) | (w1547 & w1548);
assign w1292 = (w746 & w651) | (w746 & w1939) | (w651 & w1939);
assign w1293 = ~w651 & w1940;
assign w1294 = (~w20 & w651) | (~w20 & w1671) | (w651 & w1671);
assign w1295 = (w742 & w1549) | (w742 & w1550) | (w1549 & w1550);
assign w1296 = (~w0 & w661) | (~w0 & w1923) | (w661 & w1923);
assign w1297 = ~w661 & w1360;
assign w1298 = w764 & ~w0;
assign w1299 = (w764 & w661) | (w764 & w1941) | (w661 & w1941);
assign w1300 = (w750 & w1551) | (w750 & w1552) | (w1551 & w1552);
assign w1301 = (~w750 & w1553) | (~w750 & w1554) | (w1553 & w1554);
assign w1302 = (w750 & w1555) | (w750 & w1556) | (w1555 & w1556);
assign w1303 = (~w750 & w1557) | (~w750 & w1558) | (w1557 & w1558);
assign w1304 = w825 & w842;
assign w1305 = ~w825 & w844;
assign w1306 = w824 & w1413;
assign w1307 = (w841 & w1942) | (w841 & w1943) | (w1942 & w1943);
assign w1308 = ~w812 & w1944;
assign w1309 = (w858 & w812) | (w858 & w1945) | (w812 & w1945);
assign w1310 = ~w812 & w1400;
assign w1311 = (w1415 & w1414) | (w1415 & w849) | (w1414 & w849);
assign w1312 = ~w803 & w1946;
assign w1313 = (w865 & w803) | (w865 & w1947) | (w803 & w1947);
assign w1314 = ~w803 & w1383;
assign w1315 = (~w860 & w1559) | (~w860 & w1560) | (w1559 & w1560);
assign w1316 = (w870 & w788) | (w870 & w1948) | (w788 & w1948);
assign w1317 = ~w788 & w1949;
assign w1318 = ~w788 & w1372;
assign w1319 = ~w772 & w1361;
assign w1320 = (~w4 & w772) | (~w4 & w1362) | (w772 & w1362);
assign w1321 = ~w882 & ~w1320;
assign w1322 = (~w0 & w772) | (~w0 & w1583) | (w772 & w1583);
assign w1323 = (w831 & ~w903) | (w831 & w1563) | (~w903 & w1563);
assign w1324 = (pi04 & ~w903) | (pi04 & w1564) | (~w903 & w1564);
assign w1325 = w969 & ~w968;
assign w1326 = ~w990 & ~w958;
assign w1327 = ~w957 & w993;
assign w1328 = w957 & w995;
assign w1329 = (~w326 & w956) | (~w326 & w1565) | (w956 & w1565);
assign w1330 = (~w944 & w992) | (~w944 & w1421) | (w992 & w1421);
assign w1331 = (w1001 & w942) | (w1001 & w1950) | (w942 & w1950);
assign w1332 = ~w942 & w1951;
assign w1333 = (~w176 & w942) | (~w176 & w1540) | (w942 & w1540);
assign w1334 = (w1422 & ~w997) | (w1422 & w1566) | (~w997 & w1566);
assign w1335 = w929 & w1014;
assign w1336 = ~w929 & w1016;
assign w1337 = ~w928 & w1391;
assign w1338 = (~w1005 & w1567) | (~w1005 & w1568) | (w1567 & w1568);
assign w1339 = ~w921 & w1027;
assign w1340 = w921 & w1029;
assign w1341 = ~w920 & w1671;
assign w1342 = (w1018 & w1569) | (w1018 & w1570) | (w1569 & w1570);
assign w1343 = (~w0 & w911) | (~w0 & w1923) | (w911 & w1923);
assign w1344 = ~w911 & w1360;
assign w1345 = ~w1045 & ~w0;
assign w1346 = (~w1045 & w911) | (~w1045 & w1952) | (w911 & w1952);
assign w1347 = (w1031 & w1571) | (w1031 & w1572) | (w1571 & w1572);
assign w1348 = (~w1031 & w1573) | (~w1031 & w1574) | (w1573 & w1574);
assign w1349 = ~w1046 & ~pi03;
assign w1350 = ~w1046 & w1095;
assign w1351 = (w1031 & w1953) | (w1031 & w1954) | (w1953 & w1954);
assign w1352 = (~w1031 & w2101) | (~w1031 & w2102) | (w2101 & w2102);
assign w1353 = (w1031 & w1677) | (w1031 & w1678) | (w1677 & w1678);
assign w1354 = ~w1123 & ~w1076;
assign w1355 = (w1075 & w2028) | (w1075 & w2029) | (w2028 & w2029);
assign w1356 = w1140 & w1431;
assign w1357 = w1151 & ~w1141;
assign w1358 = w1151 & ~w1356;
assign w1359 = ~w1168 & w1171;
assign w1360 = ~w3 & w1955;
assign w1361 = ~w14 & w1956;
assign w1362 = (~w4 & w14) | (~w4 & w1957) | (w14 & w1957);
assign w1363 = (~w20 & ~w130) | (~w20 & w1362) | (~w130 & w1362);
assign w1364 = w144 & ~w174;
assign w1365 = w144 & ~w1201;
assign w1366 = w124 & w174;
assign w1367 = w124 & w1201;
assign w1368 = ~pi18 & ~w174;
assign w1369 = ~pi18 & ~w1201;
assign w1370 = pi18 & w174;
assign w1371 = pi18 & w1201;
assign w1372 = ~w74 & ~w44;
assign w1373 = w243 & ~pi16;
assign w1374 = ~w1222 & ~w258;
assign w1375 = (w177 & ~w324) | (w177 & w1958) | (~w324 & w1958);
assign w1376 = w177 & ~w1227;
assign w1377 = w324 & w1959;
assign w1378 = (w256 & w1960) | (w256 & w1961) | (w1960 & w1961);
assign w1379 = (~pi14 & ~w324) | (~pi14 & w1962) | (~w324 & w1962);
assign w1380 = ~pi14 & ~w1227;
assign w1381 = w324 & w1963;
assign w1382 = (w256 & w1964) | (w256 & w1965) | (w1964 & w1965);
assign w1383 = (w124 & w168) | (w124 & w1966) | (w168 & w1966);
assign w1384 = (w44 & ~w362) | (w44 & w1967) | (~w362 & w1967);
assign w1385 = ~w364 & ~w1238;
assign w1386 = w440 & w1679;
assign w1387 = w503 & w1968;
assign w1388 = (w464 & w1577) | (w464 & w1578) | (w1577 & w1578);
assign w1389 = w503 & w1969;
assign w1390 = (~w464 & w2103) | (~w464 & w2104) | (w2103 & w2104);
assign w1391 = ~w74 & w124;
assign w1392 = (w464 & w1579) | (w464 & w1580) | (w1579 & w1580);
assign w1393 = (w74 & ~w495) | (w74 & w1970) | (~w495 & w1970);
assign w1394 = ~w497 & ~w1253;
assign w1395 = ~w1257 & ~w483;
assign w1396 = (~pi10 & w524) | (~pi10 & w1971) | (w524 & w1971);
assign w1397 = ~pi10 & ~w1262;
assign w1398 = ~w524 & w1972;
assign w1399 = (w481 & w1973) | (w481 & w1974) | (w1973 & w1974);
assign w1400 = ~w326 & w250;
assign w1401 = (w124 & ~w530) | (w124 & w1391) | (~w530 & w1391);
assign w1402 = ~w532 & w1271;
assign w1403 = (w44 & ~w607) | (w44 & w1967) | (~w607 & w1967);
assign w1404 = (~w1275 & ~w607) | (~w1275 & w1975) | (~w607 & w1975);
assign w1405 = w631 & ~pi08;
assign w1406 = ~w1286 & ~w682;
assign w1407 = ~w1290 & ~w653;
assign w1408 = ~w1294 & ~w663;
assign w1409 = w645 & w1298;
assign w1410 = w645 & w1299;
assign w1411 = pi06 & w1298;
assign w1412 = pi06 & w1299;
assign w1413 = ~w526 & w425;
assign w1414 = (w250 & ~w803) | (w250 & w1540) | (~w803 & w1540);
assign w1415 = ~w805 & w1310;
assign w1416 = (w124 & ~w788) | (w124 & w1391) | (~w788 & w1391);
assign w1417 = ~w790 & w1314;
assign w1418 = ~w773 & w44;
assign w1419 = ~w773 & ~w1318;
assign w1420 = w891 & ~pi04;
assign w1421 = ~w1329 & ~w944;
assign w1422 = w1333 & ~w930;
assign w1423 = ~w922 & ~w74;
assign w1424 = ~w922 & w1337;
assign w1425 = ~w912 & w20;
assign w1426 = ~w912 & ~w1341;
assign w1427 = ~w974 & ~w1345;
assign w1428 = ~w974 & ~w1346;
assign w1429 = ~w905 & w1345;
assign w1430 = ~w905 & w1346;
assign w1431 = ~w1133 & w1062;
assign w1432 = w19 & ~w4;
assign w1433 = w21 & pi28;
assign w1434 = ~w21 & ~pi28;
assign w1435 = ~w42 & ~w0;
assign w1436 = ~w42 & ~w1184;
assign w1437 = (w34 & w1680) | (w34 & w1681) | (w1680 & w1681);
assign w1438 = (~w34 & w1682) | (~w34 & w1683) | (w1682 & w1683);
assign w1439 = w1185 | ~w54;
assign w1440 = (~w54 & w1185) | (~w54 & ~w43) | (w1185 & ~w43);
assign w1441 = w1186 & pi25;
assign w1442 = (~w34 & w2105) | (~w34 & w2106) | (w2105 & w2106);
assign w1443 = w67 & w0;
assign w1444 = w67 & ~w1187;
assign w1445 = (~w50 & w2107) | (~w50 & w2108) | (w2107 & w2108);
assign w1446 = (~w80 & w2109) | (~w80 & w2110) | (w2109 & w2110);
assign w1447 = (w0 & w80) | (w0 & w1581) | (w80 & w1581);
assign w1448 = w102 & w4;
assign w1449 = (w102 & w80) | (w102 & w1582) | (w80 & w1582);
assign w1450 = (~w80 & w1213) | (~w80 & w1583) | (w1213 & w1583);
assign w1451 = (~w0 & w1199) | (~w0 & ~w132) | (w1199 & ~w132);
assign w1452 = (~w0 & w1199) | (~w0 & w1198) | (w1199 & w1198);
assign w1453 = ~w175 & w188;
assign w1454 = w227 & ~w4;
assign w1455 = w227 & ~w1210;
assign w1456 = ~w1211 & w0;
assign w1457 = w245 & ~w291;
assign w1458 = ~w245 & ~w176;
assign w1459 = w1224 & ~w1223;
assign w1460 = ~w325 & w374;
assign w1461 = (w386 & w1586) | (w386 & w1587) | (w1586 & w1587);
assign w1462 = w1240 & w401;
assign w1463 = (~w386 & w2111) | (~w386 & w2112) | (w2111 & w2112);
assign w1464 = (w386 & w1588) | (w386 & w1589) | (w1588 & w1589);
assign w1465 = w1242 & w4;
assign w1466 = (w4 & w1242) | (w4 & w2069) | (w1242 & w2069);
assign w1467 = w450 & ~w445;
assign w1468 = ~w1248 & ~w434;
assign w1469 = ~w124 & w176;
assign w1470 = ~w124 & ~w1249;
assign w1471 = (~w508 & w1684) | (~w508 & w1685) | (w1684 & w1685);
assign w1472 = w1262 | w1261;
assign w1473 = (~w508 & w1686) | (~w508 & w1687) | (w1686 & w1687);
assign w1474 = ~w525 & w545;
assign w1475 = (w516 & w1596) | (w516 & w1597) | (w1596 & w1597);
assign w1476 = (w516 & w1717) | (w516 & w1718) | (w1717 & w1718);
assign w1477 = w558 & w1267;
assign w1478 = w1269 & w541;
assign w1479 = w1269 & ~w1268;
assign w1480 = (w591 & w1270) | (w591 & ~w541) | (w1270 & ~w541);
assign w1481 = (w591 & w1270) | (w591 & w1268) | (w1270 & w1268);
assign w1482 = w1276 & w4;
assign w1483 = (w593 & w1688) | (w593 & w1689) | (w1688 & w1689);
assign w1484 = (~w593 & w1690) | (~w593 & w1691) | (w1690 & w1691);
assign w1485 = w1278 & ~w600;
assign w1486 = (w593 & w1735) | (w593 & w1736) | (w1735 & w1736);
assign w1487 = w1279 | w1213;
assign w1488 = (~w593 & w2113) | (~w593 & w2114) | (w2113 & w2114);
assign w1489 = w643 & w1692;
assign w1490 = (w703 & ~w643) | (w703 & w1604) | (~w643 & w1604);
assign w1491 = (w643 & w1605) | (w643 & w1606) | (w1605 & w1606);
assign w1492 = w526 & ~w713;
assign w1493 = w1288 & w738;
assign w1494 = (w729 & w1607) | (w729 & w1608) | (w1607 & w1608);
assign w1495 = (~w729 & w2115) | (~w729 & w2116) | (w2115 & w2116);
assign w1496 = (~w742 & w2030) | (~w742 & w2031) | (w2030 & w2031);
assign w1497 = w1299 | w1298;
assign w1498 = (~w742 & w2032) | (~w742 & w2033) | (w2032 & w2033);
assign w1499 = ~w765 & w815;
assign w1500 = (w863 & w1312) | (w863 & ~w805) | (w1312 & ~w805);
assign w1501 = (~w846 & w2117) | (~w846 & w2118) | (w2117 & w2118);
assign w1502 = w1313 & w805;
assign w1503 = (w846 & w1990) | (w846 & w1991) | (w1990 & w1991);
assign w1504 = w1319 & w4;
assign w1505 = (w867 & w1719) | (w867 & w1720) | (w1719 & w1720);
assign w1506 = (~w867 & w1721) | (~w867 & w1722) | (w1721 & w1722);
assign w1507 = w1321 & ~w882;
assign w1508 = (w867 & w1737) | (w867 & w1738) | (w1737 & w1738);
assign w1509 = w1322 | w1213;
assign w1510 = (~w867 & w2152) | (~w867 & w2153) | (w2152 & w2153);
assign w1511 = w903 & w1611;
assign w1512 = (w965 & ~w903) | (w965 & w1612) | (~w903 & w1612);
assign w1513 = (w903 & w1613) | (w903 & w1614) | (w1613 & w1614);
assign w1514 = w766 & ~w976;
assign w1515 = (~w992 & w2119) | (~w992 & w2120) | (w2119 & w2120);
assign w1516 = w1332 & w1003;
assign w1517 = (w992 & w1615) | (w992 & w1616) | (w1615 & w1616);
assign w1518 = w1339 & w922;
assign w1519 = (w1005 & w2034) | (w1005 & w2035) | (w2034 & w2035);
assign w1520 = (w1029 & w1340) | (w1029 & ~w922) | (w1340 & ~w922);
assign w1521 = (~w1005 & w2154) | (~w1005 & w2155) | (w2154 & w2155);
assign w1522 = ~w1343 & w1039;
assign w1523 = pi02 & w1040;
assign w1524 = w972 & w1040;
assign w1525 = ~w425 & w526;
assign w1526 = ~w1122 & ~w1121;
assign w1527 = (w1171 & w1359) | (w1171 & w1358) | (w1359 & w1358);
assign w1528 = (w1171 & w1359) | (w1171 & w1357) | (w1359 & w1357);
assign w1529 = w28 & w1360;
assign w1530 = w243 & w204;
assign w1531 = w1376 & w1375;
assign w1532 = (w305 & w1992) | (w305 & w1993) | (w1992 & w1993);
assign w1533 = w1378 | w1377;
assign w1534 = (~w305 & w2121) | (~w305 & w2122) | (w2121 & w2122);
assign w1535 = w1380 & w1379;
assign w1536 = (w305 & w1994) | (w305 & w1995) | (w1994 & w1995);
assign w1537 = w1382 | w1381;
assign w1538 = (~w305 & w2123) | (~w305 & w2124) | (w2123 & w2124);
assign w1539 = ~w250 & w176;
assign w1540 = w250 & ~w176;
assign w1541 = w1397 & w1396;
assign w1542 = (w1396 & w1397) | (w1396 & w1258) | (w1397 & w1258);
assign w1543 = w1399 | w1398;
assign w1544 = (w1398 & w1399) | (w1398 & ~w1258) | (w1399 & ~w1258);
assign w1545 = w631 & w564;
assign w1546 = w631 & pi08;
assign w1547 = w1407 & ~w653;
assign w1548 = (w729 & w1996) | (w729 & w1997) | (w1996 & w1997);
assign w1549 = w1408 & ~w663;
assign w1550 = (w734 & w1998) | (w734 & w1999) | (w1998 & w1999);
assign w1551 = w711 & ~w1497;
assign w1552 = (w742 & w2043) | (w742 & w2044) | (w2043 & w2044);
assign w1553 = w645 & w1497;
assign w1554 = (~w742 & w2125) | (~w742 & w2126) | (w2125 & w2126);
assign w1555 = ~pi06 & ~w1497;
assign w1556 = (w742 & w2045) | (w742 & w2046) | (w2045 & w2046);
assign w1557 = pi06 & w1497;
assign w1558 = (~w742 & w2127) | (~w742 & w2128) | (w2127 & w2128);
assign w1559 = (w1416 & w1417) | (w1416 & ~w805) | (w1417 & ~w805);
assign w1560 = (~w846 & w2129) | (~w846 & w2130) | (w2129 & w2130);
assign w1561 = ~w773 & w2070;
assign w1562 = (w860 & w1695) | (w860 & w1696) | (w1695 & w1696);
assign w1563 = w891 & w831;
assign w1564 = w891 & pi04;
assign w1565 = w425 & ~w326;
assign w1566 = (~w992 & w2131) | (~w992 & w2132) | (w2131 & w2132);
assign w1567 = ~w922 & w2071;
assign w1568 = (~w997 & w2000) | (~w997 & w2001) | (w2000 & w2001);
assign w1569 = ~w912 & w2072;
assign w1570 = (w1005 & w2002) | (w1005 & w2003) | (w2002 & w2003);
assign w1571 = ~w974 & ~w1666;
assign w1572 = (w1018 & w2004) | (w1018 & w2005) | (w2004 & w2005);
assign w1573 = ~w905 & w1666;
assign w1574 = (~w1018 & w2006) | (~w1018 & w2007) | (w2006 & w2007);
assign w1575 = ~w645 & w1345;
assign w1576 = ~w645 & w1346;
assign w1577 = w504 & w1383;
assign w1578 = w504 & w1386;
assign w1579 = ~w74 & w1383;
assign w1580 = ~w74 & w1386;
assign w1581 = ~w1362 & w0;
assign w1582 = ~w1362 & w102;
assign w1583 = ~w0 & ~w1361;
assign w1584 = w1224 & w258;
assign w1585 = w1224 & ~w1374;
assign w1586 = w1239 & ~w1384;
assign w1587 = w1239 & ~w1385;
assign w1588 = w1241 & ~w1384;
assign w1589 = w1241 & ~w1385;
assign w1590 = (w4 & w1242) | (w4 & w1384) | (w1242 & w1384);
assign w1591 = (w4 & w1242) | (w4 & w1385) | (w1242 & w1385);
assign w1592 = w1259 & w483;
assign w1593 = w1259 & ~w1395;
assign w1594 = (w1261 & w1262) | (w1261 & w483) | (w1262 & w483);
assign w1595 = (w1261 & w1262) | (w1261 & ~w1395) | (w1262 & ~w1395);
assign w1596 = w552 & ~w1472;
assign w1597 = w552 & ~w1473;
assign w1598 = (w4 & w1276) | (w4 & w1404) | (w1276 & w1404);
assign w1599 = (w4 & w1276) | (w4 & w1403) | (w1276 & w1403);
assign w1600 = w1277 & ~w1404;
assign w1601 = w1277 & ~w1403;
assign w1602 = (w1213 & w1279) | (w1213 & ~w1404) | (w1279 & ~w1404);
assign w1603 = (w1213 & w1279) | (w1213 & ~w1403) | (w1279 & ~w1403);
assign w1604 = w631 & w703;
assign w1605 = pi09 & pi08;
assign w1606 = pi09 & ~w1405;
assign w1607 = (w738 & w1288) | (w738 & ~w682) | (w1288 & ~w682);
assign w1608 = (w738 & w1288) | (w738 & w1406) | (w1288 & w1406);
assign w1609 = (w863 & w1312) | (w863 & w1414) | (w1312 & w1414);
assign w1610 = (w863 & w1312) | (w863 & w1415) | (w1312 & w1415);
assign w1611 = ~w891 & ~w962;
assign w1612 = w891 & w965;
assign w1613 = pi05 & pi04;
assign w1614 = pi05 & ~w1420;
assign w1615 = (w1003 & w1332) | (w1003 & ~w944) | (w1332 & ~w944);
assign w1616 = (w1003 & w1332) | (w1003 & w1421) | (w1332 & w1421);
assign w1617 = w19 & w8;
assign w1618 = ~w13 & ~w15;
assign w1619 = w317 & ~w1224;
assign w1620 = (w305 & w1697) | (w305 & w1698) | (w1697 & w1698);
assign w1621 = w287 & w374;
assign w1622 = w287 & w318;
assign w1623 = ~w287 & ~w374;
assign w1624 = ~w287 & ~w318;
assign w1625 = w0 & ~w1241;
assign w1626 = (~w386 & w1699) | (~w386 & w1700) | (w1699 & w1700);
assign w1627 = (~w396 & w1701) | (~w396 & w1702) | (w1701 & w1702);
assign w1628 = ~w355 & ~w1241;
assign w1629 = (~w386 & w1703) | (~w386 & w1704) | (w1703 & w1704);
assign w1630 = ~w0 & ~w1465;
assign w1631 = (w386 & w1705) | (w386 & w1706) | (w1705 & w1706);
assign w1632 = w443 & w445;
assign w1633 = w443 & ~w1467;
assign w1634 = ~w1254 & w1255;
assign w1635 = w1256 & w514;
assign w1636 = (w514 & w1256) | (w514 & w1254) | (w1256 & w1254);
assign w1637 = ~w250 & w525;
assign w1638 = (w516 & w1723) | (w516 & w1724) | (w1723 & w1724);
assign w1639 = w600 & ~w1482;
assign w1640 = w600 & ~w1483;
assign w1641 = w0 & ~w1277;
assign w1642 = w0 & ~w1484;
assign w1643 = ~w704 & w425;
assign w1644 = w704 & ~w425;
assign w1645 = (~w734 & w2133) | (~w734 & w2134) | (w2133 & w2134);
assign w1646 = w1293 & w748;
assign w1647 = (w734 & w2008) | (w734 & w2009) | (w2008 & w2009);
assign w1648 = pi07 & pi06;
assign w1649 = pi07 & ~w1302;
assign w1650 = (w750 & w2047) | (w750 & w2048) | (w2047 & w2048);
assign w1651 = (~w750 & w2049) | (~w750 & w2050) | (w2049 & w2050);
assign w1652 = w1316 & w790;
assign w1653 = (w860 & w1707) | (w860 & w1708) | (w1707 & w1708);
assign w1654 = (w872 & w1317) | (w872 & ~w790) | (w1317 & ~w790);
assign w1655 = (~w860 & w1709) | (~w860 & w1710) | (w1709 & w1710);
assign w1656 = (~w840 & ~w903) | (~w840 & w1739) | (~w903 & w1739);
assign w1657 = w903 & w1740;
assign w1658 = ~w904 & ~w838;
assign w1659 = (w903 & w1741) | (w903 & w1742) | (w1741 & w1742);
assign w1660 = (w1014 & w1335) | (w1014 & ~w930) | (w1335 & ~w930);
assign w1661 = (~w997 & w2010) | (~w997 & w2011) | (w2010 & w2011);
assign w1662 = w1336 & w930;
assign w1663 = (w997 & w2012) | (w997 & w2013) | (w2012 & w2013);
assign w1664 = w1522 & w1039;
assign w1665 = (w1018 & w2014) | (w1018 & w2015) | (w2014 & w2015);
assign w1666 = w1346 | w1345;
assign w1667 = (~w1018 & w2016) | (~w1018 & w2017) | (w2016 & w2017);
assign w1668 = w961 & ~w1105;
assign w1669 = (~w1031 & w2018) | (~w1031 & w2019) | (w2018 & w2019);
assign w1670 = w1166 & ~w1169;
assign w1671 = ~w44 & ~w20;
assign w1672 = ~w405 & w417;
assign w1673 = w1395 & ~w483;
assign w1674 = (~w483 & w1395) | (~w483 & w1254) | (w1395 & w1254);
assign w1675 = (w1401 & w1402) | (w1401 & ~w541) | (w1402 & ~w541);
assign w1676 = (w1401 & w1402) | (w1401 & w1268) | (w1402 & w1268);
assign w1677 = w983 & ~w1666;
assign w1678 = (w1342 & w2135) | (w1342 & w2136) | (w2135 & w2136);
assign w1679 = w1540 & w124;
assign w1680 = w27 & ~w1436;
assign w1681 = (w27 & w42) | (w27 & w2020) | (w42 & w2020);
assign w1682 = ~w20 & w1436;
assign w1683 = ~w42 & w2021;
assign w1684 = w1259 & ~w1673;
assign w1685 = (w1592 & w1593) | (w1592 & ~w1254) | (w1593 & ~w1254);
assign w1686 = (w1261 & w1262) | (w1261 & ~w1673) | (w1262 & ~w1673);
assign w1687 = (w1595 & w1594) | (w1595 & ~w1254) | (w1594 & ~w1254);
assign w1688 = (w4 & w1276) | (w4 & w2073) | (w1276 & w2073);
assign w1689 = (w1599 & w1598) | (w1599 & ~w1272) | (w1598 & ~w1272);
assign w1690 = w1277 & ~w2073;
assign w1691 = (w1601 & w1600) | (w1601 & w1272) | (w1600 & w1272);
assign w1692 = ~w631 & ~w700;
assign w1693 = (w1416 & w1417) | (w1416 & w1414) | (w1417 & w1414);
assign w1694 = (w1416 & w1417) | (w1416 & w1415) | (w1417 & w1415);
assign w1695 = ~w773 & w2074;
assign w1696 = (w1418 & w1419) | (w1418 & ~w1560) | (w1419 & ~w1560);
assign w1697 = w317 & ~w1585;
assign w1698 = w317 & ~w1584;
assign w1699 = w0 & ~w1589;
assign w1700 = w0 & ~w1588;
assign w1701 = w418 & ~w1625;
assign w1702 = w418 & ~w1626;
assign w1703 = ~w355 & ~w1589;
assign w1704 = ~w355 & ~w1588;
assign w1705 = ~w0 & ~w1591;
assign w1706 = ~w0 & ~w1590;
assign w1707 = w1316 & ~w1559;
assign w1708 = w1316 & ~w1560;
assign w1709 = (w872 & w1317) | (w872 & w1559) | (w1317 & w1559);
assign w1710 = (w872 & w1317) | (w872 & w1560) | (w1317 & w1560);
assign w1711 = (~w445 & w1467) | (~w445 & ~w1243) | (w1467 & ~w1243);
assign w1712 = (~w445 & w1467) | (~w445 & w406) | (w1467 & w406);
assign w1713 = ~w474 & ~w1259;
assign w1714 = ~w474 & ~w1471;
assign w1715 = w571 & ~w562;
assign w1716 = ~w571 & w562;
assign w1717 = w444 & ~w1472;
assign w1718 = w444 & ~w1473;
assign w1719 = (w4 & w1319) | (w4 & w1561) | (w1319 & w1561);
assign w1720 = (w860 & w1745) | (w860 & w1746) | (w1745 & w1746);
assign w1721 = w1320 & ~w1561;
assign w1722 = (~w860 & w1747) | (~w860 & w1748) | (w1747 & w1748);
assign w1723 = w463 & ~w1472;
assign w1724 = w463 & ~w1473;
assign w1725 = (w616 & w1273) | (w616 & ~w532) | (w1273 & ~w532);
assign w1726 = (w616 & w1273) | (w616 & w1272) | (w1273 & w1272);
assign w1727 = w1274 & w532;
assign w1728 = w1274 & ~w1272;
assign w1729 = w882 & ~w1504;
assign w1730 = (~w867 & w1749) | (~w867 & w1750) | (w1749 & w1750);
assign w1731 = w0 & ~w1320;
assign w1732 = (w867 & w1751) | (w867 & w1752) | (w1751 & w1752);
assign w1733 = ~w900 & ~w829;
assign w1734 = w900 & w829;
assign w1735 = (~w600 & w1278) | (~w600 & w2073) | (w1278 & w2073);
assign w1736 = (~w1272 & w2137) | (~w1272 & w2138) | (w2137 & w2138);
assign w1737 = (~w882 & w1321) | (~w882 & w1561) | (w1321 & w1561);
assign w1738 = (~w882 & w1321) | (~w882 & w1562) | (w1321 & w1562);
assign w1739 = w891 & ~w840;
assign w1740 = ~w891 & ~w526;
assign w1741 = ~w978 & ~pi04;
assign w1742 = ~w978 & ~w1564;
assign w1743 = (~w1694 & w1418) | (~w1694 & w1419) | (w1418 & w1419);
assign w1744 = (~w1693 & w1418) | (~w1693 & w1419) | (w1418 & w1419);
assign w1745 = (w4 & w1319) | (w4 & w1695) | (w1319 & w1695);
assign w1746 = (~w849 & w2139) | (~w849 & w2140) | (w2139 & w2140);
assign w1747 = w1320 & ~w1695;
assign w1748 = (w849 & w2022) | (w849 & w2023) | (w2022 & w2023);
assign w1749 = w882 & ~w1719;
assign w1750 = w882 & ~w1720;
assign w1751 = w0 & ~w1721;
assign w1752 = w0 & ~w1722;
assign w1753 = w28 & w4;
assign w1754 = w31 & ~w30;
assign w1755 = ~w43 & w63;
assign w1756 = ~w43 & ~w87;
assign w1757 = w43 & w87;
assign w1758 = ~pi22 & w88;
assign w1759 = ~w99 & w59;
assign w1760 = w99 & ~w59;
assign w1761 = w95 & ~w20;
assign w1762 = ~w95 & w20;
assign w1763 = w127 & w80;
assign w1764 = ~w127 & ~w80;
assign w1765 = ~w1196 & ~w146;
assign w1766 = w149 & w151;
assign w1767 = w93 & w84;
assign w1768 = ~w93 & ~w84;
assign w1769 = w157 & w139;
assign w1770 = w157 & ~w152;
assign w1771 = w159 & ~w139;
assign w1772 = w159 & w152;
assign w1773 = ~w164 & w102;
assign w1774 = w164 & ~w102;
assign w1775 = ~w167 & ~w1451;
assign w1776 = ~w167 & w161;
assign w1777 = w143 & w168;
assign w1778 = w20 & w152;
assign w1779 = ~w225 & w156;
assign w1780 = w153 & ~w4;
assign w1781 = ~w153 & w4;
assign w1782 = w236 & w130;
assign w1783 = ~w236 & ~w130;
assign w1784 = w174 & w167;
assign w1785 = ~w198 & w44;
assign w1786 = ~w261 & ~w191;
assign w1787 = ~w211 & ~w202;
assign w1788 = w211 & w202;
assign w1789 = ~w314 & w227;
assign w1790 = w314 & ~w227;
assign w1791 = w1225 & w0;
assign w1792 = (w0 & w1225) | (w0 & w1223) | (w1225 & w1223);
assign w1793 = w271 & w20;
assign w1794 = ~w353 & ~w263;
assign w1795 = ~w389 & w275;
assign w1796 = w324 & ~w317;
assign w1797 = ~w347 & ~w338;
assign w1798 = w347 & w338;
assign w1799 = ~w423 & ~w417;
assign w1800 = pi12 & ~w444;
assign w1801 = ~w472 & ~w355;
assign w1802 = ~w372 & w44;
assign w1803 = ~w486 & ~w391;
assign w1804 = ~w333 & ~w124;
assign w1805 = ~w501 & ~w377;
assign w1806 = ~w1254 & ~w496;
assign w1807 = ~w1254 & w1257;
assign w1808 = w1260 & w0;
assign w1809 = (w0 & w1260) | (w0 & w1258) | (w1260 & w1258);
assign w1810 = ~w527 & w431;
assign w1811 = w527 & ~w431;
assign w1812 = ~w444 & ~w1243;
assign w1813 = ~w444 & w406;
assign w1814 = w558 & ~w557;
assign w1815 = ~w540 & w541;
assign w1816 = ~w540 & ~w1268;
assign w1817 = w585 & w434;
assign w1818 = ~w585 & ~w434;
assign w1819 = ~w598 & ~w488;
assign w1820 = ~w470 & w74;
assign w1821 = ~w612 & ~w503;
assign w1822 = ~w531 & w532;
assign w1823 = ~w531 & ~w1272;
assign w1824 = ~w524 & w474;
assign w1825 = ~w666 & ~w614;
assign w1826 = ~w671 & w588;
assign w1827 = ~w685 & ~w547;
assign w1828 = ~w1287 & ~w681;
assign w1829 = ~w1287 & w1290;
assign w1830 = ~w1291 & ~w652;
assign w1831 = ~w1291 & w1294;
assign w1832 = ~w754 & w600;
assign w1833 = w754 & ~w600;
assign w1834 = w1297 & w0;
assign w1835 = (w0 & w1297) | (w0 & w1295) | (w1297 & w1295);
assign w1836 = w765 & ~w44;
assign w1837 = ~w765 & ~w744;
assign w1838 = ~w765 & ~w742;
assign w1839 = ~w765 & w778;
assign w1840 = (~w750 & w2051) | (~w750 & w2052) | (w2051 & w2052);
assign w1841 = (w750 & w2053) | (w750 & w2054) | (w2053 & w2054);
assign w1842 = ~w765 & ~w734;
assign w1843 = w695 & w176;
assign w1844 = ~w765 & w793;
assign w1845 = (~w750 & w2055) | (~w750 & w2056) | (w2055 & w2056);
assign w1846 = (w750 & w2057) | (w750 & w2058) | (w2057 & w2058);
assign w1847 = (~w750 & w2036) | (~w750 & w2037) | (w2036 & w2037);
assign w1848 = (w750 & w2038) | (w750 & w2039) | (w2038 & w2039);
assign w1849 = ~w1303 & w833;
assign w1850 = ~w765 & ~w726;
assign w1851 = ~w765 & w852;
assign w1852 = ~w850 & ~w250;
assign w1853 = ~w850 & w250;
assign w1854 = ~w804 & w805;
assign w1855 = ~w804 & ~w1311;
assign w1856 = ~w791 & ~w124;
assign w1857 = ~w791 & w124;
assign w1858 = ~w789 & w790;
assign w1859 = ~w789 & ~w1315;
assign w1860 = ~w776 & ~w44;
assign w1861 = ~w776 & w44;
assign w1862 = ~w765 & ~w750;
assign w1863 = ~w765 & w879;
assign w1864 = w764 & ~w757;
assign w1865 = w765 & ~w4;
assign w1866 = ~w765 & ~w752;
assign w1867 = w868 & ~w74;
assign w1868 = ~w868 & w74;
assign w1869 = w917 & w788;
assign w1870 = ~w917 & ~w788;
assign w1871 = w861 & ~w176;
assign w1872 = ~w861 & w176;
assign w1873 = w925 & w803;
assign w1874 = ~w925 & ~w803;
assign w1875 = ~w813 & ~w250;
assign w1876 = ~w933 & ~w855;
assign w1877 = ~w825 & ~w425;
assign w1878 = ~w947 & ~w818;
assign w1879 = ~w765 & w975;
assign w1880 = w765 & ~w975;
assign w1881 = ~w1330 & ~w943;
assign w1882 = ~w1330 & w1333;
assign w1883 = ~w929 & w930;
assign w1884 = ~w929 & ~w1334;
assign w1885 = ~w1011 & ~w796;
assign w1886 = ~w921 & w922;
assign w1887 = ~w921 & ~w1338;
assign w1888 = ~w1024 & ~w781;
assign w1889 = ~w1342 & ~w913;
assign w1890 = ~w1342 & w1343;
assign w1891 = ~w1036 & w882;
assign w1892 = w1036 & ~w882;
assign w1893 = w1344 & w0;
assign w1894 = (w0 & w1344) | (w0 & w1342) | (w1344 & w1342);
assign w1895 = ~w898 & ~w899;
assign w1896 = w957 & w326;
assign w1897 = ~w1065 & ~w949;
assign w1898 = (~w326 & w1067) | (~w326 & w1400) | (w1067 & w1400);
assign w1899 = ~w1136 & ~w935;
assign w1900 = (w74 & ~w1138) | (w74 & w2024) | (~w1138 & w2024);
assign w1901 = ~w1144 & ~w1013;
assign w1902 = ~w1138 & w2024;
assign w1903 = ~w1163 & ~w1026;
assign w1904 = w1173 & w0;
assign w1905 = ~w1045 & ~w1039;
assign w1906 = ~w1176 & ~w0;
assign w1907 = ~w1176 & ~w1904;
assign w1908 = w1213 & ~w0;
assign w1909 = (~w0 & w1213) | (~w0 & ~w28) | (w1213 & ~w28);
assign w1910 = ~w43 & pi22;
assign w1911 = w144 & w2075;
assign w1912 = (w1364 & w1365) | (w1364 & ~w1198) | (w1365 & ~w1198);
assign w1913 = w124 & ~w2075;
assign w1914 = (w1366 & w1367) | (w1366 & w1198) | (w1367 & w1198);
assign w1915 = ~pi18 & w2075;
assign w1916 = (w1368 & w1369) | (w1368 & ~w1198) | (w1369 & ~w1198);
assign w1917 = pi18 & ~w2075;
assign w1918 = (w1370 & w1371) | (w1370 & w1198) | (w1371 & w1198);
assign w1919 = w1 & ~w0;
assign w1920 = w243 & pi16;
assign w1921 = ~w44 & w306;
assign w1922 = w44 & w308;
assign w1923 = ~w4 & ~w0;
assign w1924 = ~w1360 & w324;
assign w1925 = ~w74 & w392;
assign w1926 = w74 & w394;
assign w1927 = ~w20 & w399;
assign w1928 = w20 & w401;
assign w1929 = w250 & w452;
assign w1930 = (w1383 & w1386) | (w1383 & w1247) | (w1386 & w1247);
assign w1931 = (w1383 & w1386) | (w1383 & ~w442) | (w1386 & ~w442);
assign w1932 = ~w44 & w512;
assign w1933 = w44 & w514;
assign w1934 = ~w1360 & ~w524;
assign w1935 = w250 & w730;
assign w1936 = ~w250 & w732;
assign w1937 = ~w124 & w738;
assign w1938 = w124 & w740;
assign w1939 = ~w44 & w746;
assign w1940 = w44 & w748;
assign w1941 = ~w1360 & w764;
assign w1942 = (w425 & ~w812) | (w425 & w1565) | (~w812 & w1565);
assign w1943 = ~w814 & w1306;
assign w1944 = ~w326 & w856;
assign w1945 = w326 & w858;
assign w1946 = ~w176 & w863;
assign w1947 = w176 & w865;
assign w1948 = w74 & w870;
assign w1949 = ~w74 & w872;
assign w1950 = w250 & w1001;
assign w1951 = ~w250 & w1003;
assign w1952 = ~w1360 & ~w1045;
assign w1953 = w1105 & ~w1666;
assign w1954 = (w1342 & w2141) | (w1342 & w2142) | (w2141 & w2142);
assign w1955 = ~w1 & w0;
assign w1956 = w19 & w4;
assign w1957 = ~w19 & ~w4;
assign w1958 = w0 & w177;
assign w1959 = ~w0 & w250;
assign w1960 = w250 & w324;
assign w1961 = w250 & w1924;
assign w1962 = w0 & ~pi14;
assign w1963 = ~w0 & pi14;
assign w1964 = pi14 & w324;
assign w1965 = pi14 & w1924;
assign w1966 = ~w175 & w124;
assign w1967 = w20 & w44;
assign w1968 = w74 & w124;
assign w1969 = ~w74 & ~w124;
assign w1970 = w44 & w74;
assign w1971 = w0 & ~pi10;
assign w1972 = ~w0 & pi10;
assign w1973 = pi10 & ~w524;
assign w1974 = pi10 & w1934;
assign w1975 = w20 & ~w1275;
assign w1976 = w31 & w1183;
assign w1977 = w20 & ~w1439;
assign w1978 = w20 & ~w37;
assign w1979 = ~w1205 & w208;
assign w1980 = w1205 & w124;
assign w1981 = (w856 & w1308) | (w856 & ~w814) | (w1308 & ~w814);
assign w1982 = (w856 & w1308) | (w856 & w1307) | (w1308 & w1307);
assign w1983 = w1309 & w814;
assign w1984 = w1309 & ~w1307;
assign w1985 = (~w1068 & w1355) | (~w1068 & ~w1076) | (w1355 & ~w1076);
assign w1986 = (~w1068 & w1355) | (~w1068 & w1354) | (w1355 & w1354);
assign w1987 = (~w74 & w1146) | (~w74 & w1372) | (w1146 & w1372);
assign w1988 = ~w1054 & ~w1528;
assign w1989 = ~w1054 & w1125;
assign w1990 = w1313 & w2076;
assign w1991 = (~w1307 & w2143) | (~w1307 & w2144) | (w2143 & w2144);
assign w1992 = (w1375 & w1376) | (w1375 & ~w258) | (w1376 & ~w258);
assign w1993 = (w1375 & w1376) | (w1375 & w1374) | (w1376 & w1374);
assign w1994 = (w1379 & w1380) | (w1379 & ~w258) | (w1380 & ~w258);
assign w1995 = (w1379 & w1380) | (w1379 & w1374) | (w1380 & w1374);
assign w1996 = (~w653 & w1407) | (~w653 & ~w682) | (w1407 & ~w682);
assign w1997 = (~w653 & w1407) | (~w653 & w1406) | (w1407 & w1406);
assign w1998 = (~w663 & w1408) | (~w663 & w1547) | (w1408 & w1547);
assign w1999 = (~w663 & w1408) | (~w663 & w1548) | (w1408 & w1548);
assign w2000 = ~w922 & w2077;
assign w2001 = (w1423 & w1424) | (w1423 & w1566) | (w1424 & w1566);
assign w2002 = ~w912 & w2078;
assign w2003 = (w1426 & w1425) | (w1426 & ~w1568) | (w1425 & ~w1568);
assign w2004 = ~w974 & ~w2016;
assign w2005 = (w1427 & w1428) | (w1427 & w1570) | (w1428 & w1570);
assign w2006 = ~w905 & w2016;
assign w2007 = (w1429 & w1430) | (w1429 & ~w1570) | (w1430 & ~w1570);
assign w2008 = (w748 & w1293) | (w748 & w1547) | (w1293 & w1547);
assign w2009 = (w748 & w1293) | (w748 & w1548) | (w1293 & w1548);
assign w2010 = (w1014 & w1335) | (w1014 & w1422) | (w1335 & w1422);
assign w2011 = (w1014 & w1335) | (w1014 & w1566) | (w1335 & w1566);
assign w2012 = w1336 & ~w1422;
assign w2013 = w1336 & ~w1566;
assign w2014 = (w1039 & w1522) | (w1039 & w1569) | (w1522 & w1569);
assign w2015 = (w1039 & w1522) | (w1039 & w1570) | (w1522 & w1570);
assign w2016 = (w1345 & w1346) | (w1345 & ~w1569) | (w1346 & ~w1569);
assign w2017 = (w1345 & w1346) | (w1345 & ~w1570) | (w1346 & ~w1570);
assign w2018 = w961 & ~w1664;
assign w2019 = w961 & ~w1665;
assign w2020 = w0 & w27;
assign w2021 = ~w0 & ~w20;
assign w2022 = w1320 & ~w1744;
assign w2023 = w1320 & ~w1743;
assign w2024 = ~w124 & w74;
assign w2025 = w1106 & ~w425;
assign w2026 = w1525 | w526;
assign w2027 = (w526 & w1525) | (w526 & w1106) | (w1525 & w1106);
assign w2028 = ~w1068 & ~w1898;
assign w2029 = ~w1068 & w1124;
assign w2030 = w1296 & ~w1549;
assign w2031 = w1296 & ~w1550;
assign w2032 = (w1298 & w1299) | (w1298 & ~w1549) | (w1299 & ~w1549);
assign w2033 = (w1298 & w1299) | (w1298 & ~w1550) | (w1299 & ~w1550);
assign w2034 = w1339 & ~w1567;
assign w2035 = w1339 & ~w1568;
assign w2036 = ~w425 & w1497;
assign w2037 = ~w425 & w1498;
assign w2038 = w720 & ~w1497;
assign w2039 = w720 & ~w1498;
assign w2040 = w757 & ~w1296;
assign w2041 = w757 & ~w1496;
assign w2042 = w709 & w758;
assign w2043 = w711 & ~w2032;
assign w2044 = (w1550 & w2145) | (w1550 & w2146) | (w2145 & w2146);
assign w2045 = ~pi06 & ~w2032;
assign w2046 = (w1550 & w2147) | (w1550 & w2148) | (w2147 & w2148);
assign w2047 = w835 & ~w1557;
assign w2048 = w835 & ~w1558;
assign w2049 = w645 & w1557;
assign w2050 = w645 & w1558;
assign w2051 = ~w124 & w1497;
assign w2052 = ~w124 & w1498;
assign w2053 = w736 & ~w1497;
assign w2054 = w736 & ~w1498;
assign w2055 = ~w250 & w1497;
assign w2056 = ~w250 & w1498;
assign w2057 = w728 & ~w1497;
assign w2058 = w728 & ~w1498;
assign w2059 = (w0 & ~w1187) | (w0 & ~w62) | (~w1187 & ~w62);
assign w2060 = (w139 & ~w152) | (w139 & ~w1197) | (~w152 & ~w1197);
assign w2061 = (w140 & w20) | (w140 & w1778) | (w20 & w1778);
assign w2062 = (w1243 & ~w406) | (w1243 & ~w446) | (~w406 & ~w446);
assign w2063 = (~w541 & w1268) | (~w541 & ~w581) | (w1268 & ~w581);
assign w2064 = (~w532 & w1272) | (~w532 & ~w593) | (w1272 & ~w593);
assign w2065 = (~w805 & w1311) | (~w805 & ~w860) | (w1311 & ~w860);
assign w2066 = (~w790 & w1315) | (~w790 & ~w867) | (w1315 & ~w867);
assign w2067 = (~w930 & w1334) | (~w930 & ~w1005) | (w1334 & ~w1005);
assign w2068 = (~w922 & w1338) | (~w922 & ~w1018) | (w1338 & ~w1018);
assign w2069 = (w1384 & w1385) | (w1384 & ~w386) | (w1385 & ~w386);
assign w2070 = (w44 & ~w1318) | (w44 & w790) | (~w1318 & w790);
assign w2071 = (~w74 & w1337) | (~w74 & ~w930) | (w1337 & ~w930);
assign w2072 = (~w1341 & w20) | (~w1341 & w922) | (w20 & w922);
assign w2073 = (w1403 & w1404) | (w1403 & w532) | (w1404 & w532);
assign w2074 = (w44 & ~w1318) | (w44 & ~w1559) | (~w1318 & ~w1559);
assign w2075 = (~w174 & ~w1201) | (~w174 & w132) | (~w1201 & w132);
assign w2076 = (~w1415 & ~w1414) | (~w1415 & w814) | (~w1414 & w814);
assign w2077 = (~w74 & w1337) | (~w74 & w1422) | (w1337 & w1422);
assign w2078 = (~w1341 & w20) | (~w1341 & ~w1567) | (w20 & ~w1567);
assign w2079 = w188 & w143;
assign w2080 = ~w143 & ~w188;
assign w2081 = ~w143 & ~w168;
assign w2082 = w1227 | w1226;
assign w2083 = (w1226 & w1227) | (w1226 & ~w1223) | (w1227 & ~w1223);
assign w2084 = (w1632 & w1633) | (w1632 & w1243) | (w1633 & w1243);
assign w2085 = (w1632 & w1633) | (w1632 & ~w406) | (w1633 & ~w406);
assign w2086 = w536 & w534;
assign w2087 = ~w536 & ~w534;
assign w2088 = ~w543 & ~w545;
assign w2089 = ~w543 & ~w520;
assign w2090 = w815 & w709;
assign w2091 = ~w709 & ~w815;
assign w2092 = ~w709 & ~w758;
assign w2093 = ~pi03 & pi02;
assign w2094 = ~w1088 & pi03;
assign w2095 = ~w1088 & ~w1040;
assign w2096 = w1095 & w972;
assign w2097 = ~w972 & ~w1095;
assign w2098 = ~w972 & ~w1040;
assign w2099 = w1363 & w139;
assign w2100 = w1363 & ~w152;
assign w2101 = w1576 | w1575;
assign w2102 = (w1575 & w1576) | (w1575 & ~w1342) | (w1576 & ~w1342);
assign w2103 = w506 & ~w1383;
assign w2104 = w506 & ~w1386;
assign w2105 = (pi25 & w1186) | (pi25 & w1436) | (w1186 & w1436);
assign w2106 = (pi25 & w1186) | (pi25 & w1435) | (w1186 & w1435);
assign w2107 = ~w72 & ~w0;
assign w2108 = ~w72 & ~w1360;
assign w2109 = ~w102 & ~w4;
assign w2110 = ~w102 & ~w1361;
assign w2111 = (w401 & w1240) | (w401 & w1384) | (w1240 & w1384);
assign w2112 = (w401 & w1240) | (w401 & w1385) | (w1240 & w1385);
assign w2113 = (w1603 & w1602) | (w1603 & ~w532) | (w1602 & ~w532);
assign w2114 = (w1603 & w1602) | (w1603 & w1272) | (w1602 & w1272);
assign w2115 = w1289 & w682;
assign w2116 = w1289 & ~w1406;
assign w2117 = (w1610 & w1609) | (w1610 & ~w814) | (w1609 & ~w814);
assign w2118 = (w1610 & w1609) | (w1610 & w1307) | (w1609 & w1307);
assign w2119 = w1331 & w944;
assign w2120 = w1331 & ~w1421;
assign w2121 = (w1377 & w1378) | (w1377 & w258) | (w1378 & w258);
assign w2122 = (w1377 & w1378) | (w1377 & ~w1374) | (w1378 & ~w1374);
assign w2123 = (w1381 & w1382) | (w1381 & w258) | (w1382 & w258);
assign w2124 = (w1381 & w1382) | (w1381 & ~w1374) | (w1382 & ~w1374);
assign w2125 = (w1409 & w1410) | (w1409 & ~w1549) | (w1410 & ~w1549);
assign w2126 = (w1409 & w1410) | (w1409 & ~w1550) | (w1410 & ~w1550);
assign w2127 = (w1411 & w1412) | (w1411 & ~w1549) | (w1412 & ~w1549);
assign w2128 = (w1411 & w1412) | (w1411 & ~w1550) | (w1412 & ~w1550);
assign w2129 = (w1694 & w1693) | (w1694 & ~w814) | (w1693 & ~w814);
assign w2130 = (w1694 & w1693) | (w1694 & w1307) | (w1693 & w1307);
assign w2131 = w1422 & w944;
assign w2132 = w1422 & ~w1421;
assign w2133 = w1292 & ~w1547;
assign w2134 = w1292 & ~w1548;
assign w2135 = w983 & ~w1345;
assign w2136 = w983 & ~w1346;
assign w2137 = (~w600 & w1278) | (~w600 & w1403) | (w1278 & w1403);
assign w2138 = (~w600 & w1278) | (~w600 & w1404) | (w1278 & w1404);
assign w2139 = (w4 & w1319) | (w4 & w1744) | (w1319 & w1744);
assign w2140 = (w4 & w1319) | (w4 & w1743) | (w1319 & w1743);
assign w2141 = w1105 & ~w1345;
assign w2142 = w1105 & ~w1346;
assign w2143 = w1313 & ~w1414;
assign w2144 = w1313 & ~w1415;
assign w2145 = w711 & ~w1298;
assign w2146 = w711 & ~w1299;
assign w2147 = ~pi06 & ~w1298;
assign w2148 = ~pi06 & ~w1299;
assign w2149 = pi19 & pi18;
assign w2150 = pi19 & ~w1204;
assign w2151 = w838 & ~w839;
assign w2152 = (w1213 & w1322) | (w1213 & ~w1561) | (w1322 & ~w1561);
assign w2153 = (w1213 & w1322) | (w1213 & ~w1562) | (w1322 & ~w1562);
assign w2154 = (w1029 & w1340) | (w1029 & w1567) | (w1340 & w1567);
assign w2155 = (w1029 & w1340) | (w1029 & w1568) | (w1340 & w1568);
assign one = 1;
assign po00 = ~w1178;// level 164
assign po01 = ~w1047;// level 153
assign po02 = w905;// level 136
assign po03 = ~w766;// level 119
assign po04 = w645;// level 104
assign po05 = ~w526;// level 89
assign po06 = w425;// level 75
assign po07 = ~w326;// level 61
assign po08 = w250;// level 49
assign po09 = ~w176;// level 37
assign po10 = w124;// level 28
assign po11 = ~w74;// level 18
assign po12 = ~w44;// level 11
assign po13 = ~w20;// level 6
assign po14 = ~w4;// level 3
assign po15 = ~w0;// level 1
endmodule
