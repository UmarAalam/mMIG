// Benchmark "diffeq1" written by ABC on Wed Apr 29 17:21:40 2015

module diffeq1 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288;
  wire n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n834, n835,
    n836, n837, n839, n840, n842, n843, n845, n846, n848, n849, n851, n852,
    n854, n855, n857, n858, n860, n861, n863, n864, n866, n867, n869, n870,
    n872, n873, n875, n876, n878, n879, n881, n882, n884, n885, n887, n888,
    n890, n891, n893, n894, n896, n897, n899, n900, n902, n903, n905, n906,
    n908, n909, n911, n912, n914, n915, n917, n918, n920, n921, n923, n924,
    n926, n927, n929, n930, n932, n933, n935, n936, n938, n939, n941, n942,
    n944, n945, n947, n948, n950, n951, n953, n954, n956, n957, n959, n960,
    n962, n963, n965, n966, n968, n969, n971, n972, n974, n975, n977, n978,
    n980, n981, n983, n984, n986, n987, n989, n990, n992, n993, n995, n996,
    n998, n999, n1001, n1002, n1004, n1005, n1006, n1007, n1009, n1010,
    n1012, n1013, n1015, n1016, n1018, n1019, n1021, n1022, n1024, n1025,
    n1027, n1028, n1030, n1031, n1033, n1034, n1036, n1037, n1039, n1040,
    n1042, n1043, n1045, n1046, n1048, n1049, n1051, n1052, n1054, n1055,
    n1057, n1058, n1060, n1061, n1063, n1064, n1066, n1067, n1069, n1070,
    n1072, n1073, n1075, n1076, n1078, n1079, n1081, n1082, n1084, n1085,
    n1087, n1088, n1090, n1091, n1093, n1094, n1096, n1097, n1099, n1100,
    n1102, n1103, n1105, n1106, n1108, n1109, n1111, n1112, n1114, n1115,
    n1117, n1118, n1120, n1121, n1123, n1124, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
    n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
    n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
    n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
    n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
    n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
    n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
    n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
    n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
    n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
    n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
    n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
    n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
    n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
    n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
    n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
    n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
    n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
    n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
    n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
    n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
    n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
    n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
    n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
    n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
    n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
    n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
    n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
    n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
    n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
    n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
    n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
    n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
    n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
    n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
    n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
    n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
    n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
    n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
    n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
    n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
    n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
    n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
    n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
    n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
    n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
    n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
    n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
    n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
    n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
    n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
    n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
    n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
    n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
    n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
    n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
    n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
    n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
    n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
    n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
    n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
    n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
    n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
    n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
    n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
    n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
    n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
    n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
    n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
    n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
    n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
    n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
    n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
    n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
    n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
    n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
    n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
    n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
    n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
    n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
    n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
    n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
    n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
    n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
    n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
    n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
    n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
    n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
    n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
    n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
    n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
    n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
    n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
    n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
    n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
    n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
    n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
    n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
    n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
    n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
    n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
    n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
    n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
    n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
    n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
    n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
    n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
    n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
    n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
    n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
    n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
    n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
    n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
    n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
    n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
    n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
    n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
    n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
    n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
    n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
    n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
    n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
    n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
    n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
    n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
    n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
    n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
    n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
    n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
    n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
    n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
    n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
    n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
    n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
    n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
    n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
    n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
    n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
    n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
    n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
    n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
    n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
    n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
    n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
    n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
    n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
    n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
    n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
    n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
    n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
    n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
    n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
    n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
    n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
    n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
    n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
    n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
    n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
    n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
    n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
    n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
    n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
    n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
    n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
    n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
    n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
    n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
    n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
    n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
    n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
    n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
    n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
    n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
    n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
    n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
    n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
    n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
    n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
    n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
    n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
    n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
    n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
    n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
    n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
    n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
    n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
    n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
    n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
    n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
    n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
    n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
    n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
    n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
    n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
    n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
    n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
    n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
    n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
    n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
    n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
    n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
    n11951, n11952, n11953, n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
    n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
    n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
    n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
    n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
    n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
    n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
    n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
    n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
    n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
    n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
    n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
    n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
    n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
    n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
    n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
    n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
    n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
    n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
    n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
    n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
    n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
    n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
    n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
    n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
    n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
    n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
    n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
    n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
    n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
    n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
    n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
    n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
    n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
    n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
    n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13207, n13208, n13209, n13210, n13211, n13212,
    n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
    n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
    n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
    n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
    n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
    n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
    n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
    n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
    n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
    n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
    n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
    n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
    n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
    n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
    n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
    n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
    n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
    n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
    n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
    n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
    n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
    n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
    n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
    n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
    n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
    n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
    n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
    n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
    n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
    n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
    n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
    n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
    n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
    n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
    n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
    n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
    n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
    n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
    n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
    n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
    n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
    n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
    n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
    n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
    n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
    n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
    n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
    n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
    n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
    n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
    n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
    n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
    n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
    n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
    n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
    n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
    n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
    n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
    n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
    n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
    n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
    n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
    n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
    n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
    n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
    n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
    n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
    n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
    n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
    n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
    n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
    n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
    n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
    n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
    n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
    n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
    n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
    n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
    n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
    n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
    n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
    n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
    n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
    n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
    n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
    n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
    n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
    n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
    n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
    n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
    n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
    n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
    n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
    n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
    n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
    n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
    n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
    n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
    n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
    n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
    n14536, n14537, n14538, n14539, n14540, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
    n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
    n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
    n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
    n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
    n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
    n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
    n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
    n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
    n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
    n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
    n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
    n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
    n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
    n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
    n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
    n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
    n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
    n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
    n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
    n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
    n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
    n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
    n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
    n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
    n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
    n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
    n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
    n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
    n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
    n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
    n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
    n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
    n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
    n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
    n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
    n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
    n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
    n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
    n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
    n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
    n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
    n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
    n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
    n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
    n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
    n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
    n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
    n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
    n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
    n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
    n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
    n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
    n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
    n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
    n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
    n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
    n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
    n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
    n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
    n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
    n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
    n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
    n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
    n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
    n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
    n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
    n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
    n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
    n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
    n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
    n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
    n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
    n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
    n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
    n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
    n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
    n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
    n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
    n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
    n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
    n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
    n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
    n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
    n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
    n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
    n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
    n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
    n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
    n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
    n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
    n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
    n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
    n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
    n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
    n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
    n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
    n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
    n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
    n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
    n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
    n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
    n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
    n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
    n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
    n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
    n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
    n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
    n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
    n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
    n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
    n17400, n17401, n17402, n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
    n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
    n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
    n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
    n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
    n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
    n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
    n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
    n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
    n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
    n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
    n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
    n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
    n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
    n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
    n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
    n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
    n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
    n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
    n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
    n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
    n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
    n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
    n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
    n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
    n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
    n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
    n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
    n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
    n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
    n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
    n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
    n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
    n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
    n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
    n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
    n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
    n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
    n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
    n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
    n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
    n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
    n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
    n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
    n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
    n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
    n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
    n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
    n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
    n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
    n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
    n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
    n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
    n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
    n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
    n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
    n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
    n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
    n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
    n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
    n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
    n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
    n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
    n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
    n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
    n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
    n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
    n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
    n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
    n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
    n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
    n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
    n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
    n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
    n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
    n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
    n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
    n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
    n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
    n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
    n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
    n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
    n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
    n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
    n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
    n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
    n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
    n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
    n18400, n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
    n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
    n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
    n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
    n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
    n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
    n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
    n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
    n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
    n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
    n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
    n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
    n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
    n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
    n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542, n18543,
    n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
    n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
    n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
    n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
    n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
    n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
    n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
    n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
    n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
    n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
    n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
    n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
    n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687,
    n18688, n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
    n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
    n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
    n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
    n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
    n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
    n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
    n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759,
    n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
    n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
    n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
    n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
    n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
    n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
    n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
    n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831,
    n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
    n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
    n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
    n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
    n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
    n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
    n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966, n18967,
    n18968, n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
    n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
    n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
    n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
    n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
    n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
    n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
    n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038, n19039,
    n19040, n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
    n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
    n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
    n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
    n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
    n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
    n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110, n19111,
    n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
    n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
    n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
    n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
    n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
    n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
    n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182, n19183,
    n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
    n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
    n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
    n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
    n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
    n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
    n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255,
    n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
    n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
    n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
    n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
    n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
    n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
    n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326, n19327,
    n19328, n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
    n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
    n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
    n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
    n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
    n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
    n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
    n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
    n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
    n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
    n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
    n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
    n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
    n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
    n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
    n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
    n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
    n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
    n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
    n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831,
    n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
    n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
    n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
    n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
    n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
    n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
    n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
    n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903,
    n19904, n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912,
    n19913, n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
    n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
    n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
    n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
    n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
    n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
    n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974, n19975,
    n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984,
    n19985, n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
    n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
    n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
    n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046, n20047,
    n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
    n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
    n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
    n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
    n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
    n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
    n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119,
    n20120, n20121, n20122, n20123, n20124, n20125, n20126, n20127, n20128,
    n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
    n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
    n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
    n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
    n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
    n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
    n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200,
    n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
    n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
    n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
    n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262, n20263,
    n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272,
    n20273, n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
    n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
    n20291, n20292, n20293, n20294, n20295, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
    n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327,
    n20328, n20329, n20330, n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
    n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
    n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
    n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399,
    n20400, n20401, n20402, n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
    n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
    n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
    n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470, n20471,
    n20472, n20473, n20474, n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
    n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
    n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
    n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543,
    n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
    n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
    n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
    n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614, n20615,
    n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
    n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
    n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
    n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686, n20687,
    n20688, n20689, n20690, n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
    n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
    n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
    n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
    n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
    n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
    n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
    n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
    n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
    n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
    n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
    n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
    n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
    n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
    n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
    n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
    n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
    n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
    n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
    n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
    n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
    n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119,
    n21120, n21121, n21122, n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
    n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
    n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
    n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191,
    n21192, n21193, n21194, n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
    n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
    n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
    n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263,
    n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
    n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
    n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
    n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335,
    n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
    n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
    n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
    n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406, n21407,
    n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
    n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
    n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478, n21479,
    n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
    n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
    n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
    n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550, n21551,
    n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
    n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
    n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766, n21767,
    n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
    n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
    n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
    n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838, n21839,
    n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
    n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
    n21876, n21877, n21878, n21879, n21880, n21882, n21883, n21884, n21885,
    n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
    n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902, n21903,
    n21904, n21905, n21906, n21907, n21908, n21909, n21910, n21911, n21912,
    n21913, n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
    n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
    n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
    n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947, n21948,
    n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
    n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
    n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975,
    n21976, n21977, n21978, n21979, n21980, n21981, n21982, n21983, n21984,
    n21985, n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
    n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
    n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
    n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019, n22020,
    n22021, n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
    n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
    n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046, n22047,
    n22048, n22049, n22050, n22051, n22052, n22053, n22054, n22055, n22056,
    n22057, n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
    n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
    n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
    n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091, n22092,
    n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
    n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
    n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118, n22119,
    n22120, n22121, n22122, n22123, n22124, n22125, n22126, n22127, n22128,
    n22129, n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
    n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
    n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
    n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163, n22164,
    n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
    n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
    n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191,
    n22192, n22193, n22194, n22195, n22196, n22197, n22198, n22199, n22200,
    n22201, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
    n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
    n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
    n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
    n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263,
    n22264, n22265, n22266, n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
    n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
    n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
    n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
    n22309, n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
    n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
    n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334, n22335,
    n22336, n22337, n22338, n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
    n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
    n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
    n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
    n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
    n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452,
    n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461,
    n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470,
    n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479,
    n22480, n22481, n22482, n22483, n22484, n22485, n22486, n22487, n22488,
    n22489, n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
    n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
    n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
    n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524,
    n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533,
    n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542,
    n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551,
    n22552, n22553, n22554, n22555, n22556, n22557, n22558, n22559, n22560,
    n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
    n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
    n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
    n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595, n22596,
    n22597, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
    n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
    n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622, n22623,
    n22624, n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632,
    n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
    n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
    n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
    n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668,
    n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
    n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
    n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695,
    n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703, n22704,
    n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
    n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
    n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
    n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740,
    n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
    n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
    n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
    n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776,
    n22777, n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
    n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
    n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
    n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812,
    n22813, n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
    n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
    n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
    n22840, n22841, n22842, n22843, n22844, n22845, n22846, n22847, n22848,
    n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
    n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
    n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
    n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
    n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
    n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901, n22902,
    n22903, n22904, n22905, n22906, n22907, n22908, n22909, n22910, n22911,
    n22912, n22913, n22914, n22915, n22916, n22917, n22918, n22919, n22920,
    n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
    n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
    n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
    n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956,
    n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
    n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974,
    n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983,
    n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992,
    n22993, n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
    n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
    n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028,
    n23029, n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
    n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045, n23046,
    n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055,
    n23056, n23057, n23058, n23059, n23060, n23061, n23062, n23063, n23064,
    n23065, n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
    n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
    n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
    n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100,
    n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109,
    n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
    n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126, n23127,
    n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136,
    n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
    n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
    n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
    n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171, n23172,
    n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181,
    n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
    n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199,
    n23200, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208,
    n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
    n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
    n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
    n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243, n23244,
    n23245, n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
    n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
    n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270, n23271,
    n23272, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280,
    n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
    n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
    n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
    n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316,
    n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
    n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
    n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342, n23343,
    n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352,
    n23353, n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
    n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
    n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
    n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388,
    n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
    n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
    n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414, n23415,
    n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424,
    n23425, n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
    n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
    n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
    n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460,
    n23461, n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
    n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
    n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486, n23487,
    n23488, n23489, n23490, n23491, n23492, n23493, n23494, n23495, n23496,
    n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
    n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
    n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
    n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531, n23532,
    n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
    n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568,
    n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
    n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596,
    n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
    n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
    n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622, n23623,
    n23624, n23625, n23626, n23627, n23628, n23629, n23630, n23631, n23632,
    n23633, n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
    n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
    n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
    n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667, n23668,
    n23669, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
    n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
    n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694, n23695,
    n23696, n23697, n23698, n23699, n23700, n23701, n23702, n23703, n23704,
    n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
    n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
    n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
    n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740,
    n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
    n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
    n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767,
    n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23775, n23776,
    n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
    n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
    n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
    n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812,
    n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
    n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
    n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839,
    n23840, n23841, n23842, n23843, n23844, n23845, n23846, n23847, n23848,
    n23849, n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
    n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
    n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
    n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911,
    n23912, n23913, n23914, n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
    n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
    n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
    n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983,
    n23984, n23985, n23986, n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
    n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
    n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
    n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052, n24053, n24054, n24055,
    n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
    n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
    n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
    n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127,
    n24128, n24129, n24130, n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
    n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
    n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
    n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196, n24197, n24198, n24199,
    n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
    n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
    n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244,
    n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
    n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277, n24278, n24279, n24280,
    n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316,
    n24317, n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
    n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349, n24350, n24351, n24352,
    n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
    n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388,
    n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
    n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
    n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415,
    n24416, n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424,
    n24425, n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
    n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
    n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
    n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460,
    n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
    n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
    n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486, n24487,
    n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496,
    n24497, n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
    n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
    n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
    n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532,
    n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
    n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
    n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558, n24559,
    n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568,
    n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
    n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
    n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
    n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603, n24604,
    n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
    n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621, n24622,
    n24623, n24624, n24625, n24626, n24627, n24628, n24629, n24630, n24631,
    n24632, n24633, n24634, n24635, n24636, n24637, n24638, n24639, n24640,
    n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
    n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
    n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
    n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676,
    n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
    n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694,
    n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703,
    n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
    n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
    n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
    n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766,
    n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774, n24775,
    n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
    n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
    n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
    n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820,
    n24821, n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
    n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838,
    n24839, n24840, n24841, n24842, n24843, n24844, n24845, n24846, n24847,
    n24848, n24849, n24850, n24851, n24852, n24853, n24854, n24855, n24856,
    n24857, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
    n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
    n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
    n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891, n24892,
    n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
    n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910,
    n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919,
    n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928,
    n24929, n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
    n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
    n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
    n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964,
    n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
    n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982,
    n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991,
    n24992, n24993, n24994, n24995, n24996, n24997, n24998, n24999, n25000,
    n25001, n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
    n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
    n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
    n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035, n25036,
    n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
    n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054,
    n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25062, n25063,
    n25064, n25065, n25066, n25067, n25068, n25069, n25070, n25071, n25072,
    n25073, n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
    n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108,
    n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125, n25126,
    n25127, n25128, n25129, n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144,
    n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
    n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180,
    n25181, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198,
    n25199, n25200, n25201, n25202, n25203, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213, n25214, n25215, n25216,
    n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
    n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252,
    n25253, n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270,
    n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288,
    n25289, n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
    n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324,
    n25325, n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341, n25342,
    n25343, n25344, n25345, n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
    n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
    n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415,
    n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
    n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
    n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
    n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487,
    n25488, n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496,
    n25497, n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
    n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
    n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
    n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532,
    n25533, n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
    n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550,
    n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559,
    n25560, n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568,
    n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
    n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
    n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604,
    n25605, n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613,
    n25614, n25615, n25616, n25617, n25618, n25619, n25620, n25621, n25622,
    n25623, n25624, n25625, n25626, n25627, n25628, n25629, n25630, n25631,
    n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640,
    n25641, n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
    n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
    n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
    n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685,
    n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703,
    n25704, n25705, n25706, n25707, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
    n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
    n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
    n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772, n25773, n25774, n25775,
    n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
    n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
    n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
    n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844, n25845, n25846, n25847,
    n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
    n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
    n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
    n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919,
    n25920, n25921, n25922, n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
    n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
    n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25972, n25973,
    n25974, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988, n25989, n25990, n25991,
    n25992, n25993, n25994, n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
    n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
    n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045,
    n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063,
    n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
    n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
    n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
    n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135,
    n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
    n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
    n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
    n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207,
    n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
    n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
    n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
    n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
    n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
    n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
    n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351,
    n26352, n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360,
    n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
    n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
    n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
    n26406, n26407, n26408, n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423,
    n26424, n26425, n26426, n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
    n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
    n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
    n26478, n26479, n26480, n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492, n26493, n26494, n26495,
    n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
    n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
    n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
    n26550, n26551, n26552, n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564, n26565, n26566, n26567,
    n26568, n26569, n26570, n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
    n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
    n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
    n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639,
    n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
    n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
    n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
    n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708, n26709, n26710, n26711,
    n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
    n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
    n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765,
    n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780, n26781, n26782, n26783,
    n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
    n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
    n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
    n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855,
    n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
    n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
    n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
    n26910, n26911, n26912, n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924, n26925, n26926, n26927,
    n26928, n26929, n26930, n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
    n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
    n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
    n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999,
    n27000, n27001, n27002, n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
    n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
    n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
    n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071,
    n27072, n27073, n27074, n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
    n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
    n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
    n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
    n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
    n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180,
    n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
    n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198,
    n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207,
    n27208, n27209, n27210, n27211, n27212, n27213, n27214, n27215, n27216,
    n27217, n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
    n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
    n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
    n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251, n27252,
    n27253, n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
    n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269, n27270,
    n27271, n27272, n27273, n27274, n27275, n27276, n27277, n27278, n27279,
    n27280, n27281, n27282, n27283, n27284, n27285, n27286, n27287, n27288,
    n27289, n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
    n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
    n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
    n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323, n27324,
    n27325, n27326, n27327, n27328, n27329, n27330, n27331, n27332, n27333,
    n27334, n27335, n27336, n27337, n27338, n27339, n27340, n27341, n27342,
    n27343, n27344, n27345, n27346, n27347, n27348, n27349, n27350, n27351,
    n27352, n27353, n27354, n27355, n27356, n27357, n27358, n27359, n27360,
    n27361, n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
    n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
    n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
    n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395, n27396,
    n27397, n27398, n27399, n27400, n27401, n27402, n27403, n27404, n27405,
    n27406, n27407, n27408, n27409, n27410, n27411, n27412, n27413, n27414,
    n27415, n27416, n27417, n27418, n27419, n27420, n27421, n27422, n27423,
    n27424, n27425, n27426, n27427, n27428, n27429, n27430, n27431, n27432,
    n27433, n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
    n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
    n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
    n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467, n27468,
    n27469, n27470, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
    n27478, n27479, n27480, n27481, n27482, n27483, n27484, n27485, n27486,
    n27487, n27488, n27489, n27490, n27491, n27492, n27493, n27494, n27495,
    n27496, n27497, n27498, n27499, n27500, n27501, n27502, n27503, n27504,
    n27505, n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
    n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
    n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
    n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539, n27540,
    n27541, n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
    n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557, n27558,
    n27559, n27560, n27561, n27562, n27563, n27564, n27565, n27566, n27567,
    n27568, n27569, n27570, n27571, n27572, n27573, n27574, n27575, n27576,
    n27577, n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
    n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
    n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
    n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611, n27612,
    n27613, n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
    n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629, n27630,
    n27631, n27632, n27633, n27634, n27635, n27636, n27637, n27638, n27639,
    n27640, n27641, n27642, n27643, n27644, n27645, n27646, n27647, n27648,
    n27649, n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
    n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
    n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
    n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683, n27684,
    n27685, n27686, n27687, n27688, n27689, n27690, n27691, n27692, n27693,
    n27694, n27695, n27696, n27697, n27698, n27699, n27700, n27701, n27702,
    n27703, n27704, n27705, n27706, n27707, n27708, n27709, n27710, n27711,
    n27712, n27713, n27714, n27715, n27716, n27717, n27718, n27719, n27720,
    n27721, n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
    n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
    n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
    n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755, n27756,
    n27757, n27758, n27759, n27760, n27761, n27762, n27763, n27764, n27765,
    n27766, n27767, n27768, n27769, n27770, n27771, n27772, n27773, n27774,
    n27775, n27776, n27777, n27778, n27779, n27780, n27781, n27782, n27783,
    n27784, n27785, n27786, n27787, n27788, n27789, n27790, n27791, n27792,
    n27793, n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
    n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
    n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
    n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827, n27828,
    n27829, n27830, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
    n27838, n27839, n27840, n27841, n27842, n27843, n27844, n27845, n27846,
    n27847, n27848, n27849, n27850, n27851, n27852, n27853, n27854, n27855,
    n27856, n27857, n27858, n27859, n27860, n27861, n27862, n27863, n27864,
    n27865, n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
    n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
    n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
    n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899, n27900,
    n27901, n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
    n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917, n27918,
    n27919, n27920, n27921, n27922, n27923, n27924, n27925, n27926, n27927,
    n27928, n27929, n27930, n27931, n27932, n27933, n27934, n27935, n27936,
    n27937, n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
    n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
    n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
    n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971, n27972,
    n27973, n27974, n27975, n27976, n27977, n27978, n27979, n27980, n27981,
    n27982, n27983, n27984, n27985, n27986, n27987, n27988, n27989, n27990,
    n27991, n27992, n27993, n27994, n27995, n27996, n27997, n27998, n27999,
    n28000, n28001, n28002, n28003, n28004, n28005, n28006, n28007, n28008,
    n28009, n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
    n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
    n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
    n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043, n28044,
    n28045, n28046, n28047, n28048, n28049, n28050, n28051, n28052, n28053,
    n28054, n28055, n28056, n28057, n28058, n28059, n28060, n28061, n28062,
    n28063, n28064, n28065, n28066, n28067, n28068, n28069, n28070, n28071,
    n28072, n28073, n28074, n28075, n28076, n28077, n28078, n28079, n28080,
    n28081, n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
    n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
    n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
    n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115, n28116,
    n28117, n28118, n28119, n28120, n28121, n28122, n28123, n28124, n28125,
    n28126, n28127, n28128, n28129, n28130, n28131, n28132, n28133, n28134,
    n28135, n28136, n28137, n28138, n28139, n28140, n28141, n28142, n28143,
    n28144, n28145, n28146, n28147, n28148, n28149, n28150, n28151, n28152,
    n28153, n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
    n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
    n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
    n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187, n28188,
    n28189, n28190, n28191, n28192, n28193, n28194, n28195, n28196, n28197,
    n28198, n28199, n28200, n28201, n28202, n28203, n28204, n28205, n28206,
    n28207, n28208, n28209, n28210, n28211, n28212, n28213, n28214, n28215,
    n28216, n28217, n28218, n28219, n28220, n28221, n28222, n28223, n28224,
    n28225, n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
    n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
    n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
    n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259, n28260,
    n28261, n28262, n28263, n28264, n28265, n28266, n28267, n28268, n28269,
    n28270, n28271, n28272, n28273, n28274, n28275, n28276, n28277, n28278,
    n28279, n28280, n28281, n28282, n28283, n28284, n28285, n28286, n28287,
    n28288, n28289, n28290, n28291, n28292, n28293, n28294, n28295, n28296,
    n28297, n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
    n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
    n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
    n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331, n28332,
    n28333, n28334, n28335, n28336, n28337, n28338, n28339, n28340, n28341,
    n28342, n28343, n28344, n28345, n28346, n28347, n28348, n28349, n28350,
    n28351, n28352, n28353, n28354, n28355, n28356, n28357, n28358, n28359,
    n28360, n28361, n28362, n28363, n28364, n28365, n28366, n28367, n28368,
    n28369, n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
    n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
    n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
    n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403, n28404,
    n28405, n28406, n28407, n28408, n28409, n28410, n28411, n28412, n28413,
    n28414, n28415, n28416, n28417, n28418, n28419, n28420, n28421, n28422,
    n28423, n28424, n28425, n28426, n28427, n28428, n28429, n28430, n28431,
    n28432, n28433, n28434, n28435, n28436, n28437, n28438, n28439, n28440,
    n28441, n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
    n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
    n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
    n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475, n28476,
    n28477, n28478, n28479, n28480, n28481, n28482, n28483, n28484, n28485,
    n28486, n28487, n28488, n28489, n28490, n28491, n28492, n28493, n28494,
    n28495, n28496, n28497, n28498, n28499, n28500, n28501, n28502, n28503,
    n28504, n28505, n28506, n28507, n28508, n28509, n28510, n28511, n28512,
    n28513, n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
    n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
    n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
    n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547, n28548,
    n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556, n28557,
    n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565, n28566,
    n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574, n28575,
    n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583, n28584,
    n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
    n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
    n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
    n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619, n28620,
    n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628, n28629,
    n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637, n28638,
    n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646, n28647,
    n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655, n28656,
    n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
    n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
    n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
    n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691, n28692,
    n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700, n28701,
    n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709, n28710,
    n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718, n28719,
    n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727, n28728,
    n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
    n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
    n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
    n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763, n28764,
    n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772, n28773,
    n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781, n28782,
    n28783, n28784, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
    n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
    n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
    n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
    n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
    n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
    n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845,
    n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
    n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
    n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
    n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
    n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
    n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
    n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
    n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
    n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
    n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
    n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
    n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
    n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
    n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
    n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
    n29035, n29036, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
    n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
    n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
    n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
    n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
    n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
    n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287,
    n29288, n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
    n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
    n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341,
    n29342, n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359,
    n29360, n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
    n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
    n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413,
    n29414, n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431,
    n29432, n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
    n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
    n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485,
    n29486, n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503,
    n29504, n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
    n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
    n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554, n29555, n29556, n29557,
    n29558, n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574, n29575,
    n29576, n29577, n29578, n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
    n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
    n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626, n29627, n29628, n29629,
    n29630, n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646, n29647,
    n29648, n29649, n29650, n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
    n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
    n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698, n29699, n29700, n29701,
    n29702, n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718, n29719,
    n29720, n29721, n29722, n29723, n29724, n29725, n29726, n29727, n29728,
    n29729, n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
    n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
    n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
    n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763, n29764,
    n29765, n29766, n29767, n29768, n29769, n29770, n29771, n29772, n29773,
    n29774, n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
    n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790, n29791,
    n29792, n29793, n29794, n29795, n29796, n29797, n29798, n29799, n29800,
    n29801, n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
    n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
    n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
    n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835, n29836,
    n29837, n29838, n29839, n29840, n29841, n29842, n29843, n29844, n29845,
    n29846, n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
    n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862, n29863,
    n29864, n29865, n29866, n29867, n29868, n29869, n29870, n29871, n29872,
    n29873, n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
    n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
    n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
    n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907, n29908,
    n29909, n29910, n29911, n29912, n29913, n29914, n29915, n29916, n29917,
    n29918, n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
    n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934, n29935,
    n29936, n29937, n29938, n29939, n29940, n29941, n29942, n29943, n29944,
    n29945, n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
    n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
    n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
    n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979, n29980,
    n29981, n29982, n29983, n29984, n29985, n29986, n29987, n29988, n29989,
    n29990, n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
    n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006, n30007,
    n30008, n30009, n30010, n30011, n30012, n30013, n30014, n30015, n30016,
    n30017, n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
    n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
    n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
    n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051, n30052,
    n30053, n30054, n30055, n30056, n30057, n30058, n30059, n30060, n30061,
    n30062, n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
    n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078, n30079,
    n30080, n30081, n30082, n30083, n30084, n30085, n30086, n30087, n30088,
    n30089, n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
    n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
    n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
    n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123, n30124,
    n30125, n30126, n30127, n30128, n30129, n30130, n30131, n30132, n30133,
    n30134, n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
    n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150, n30151,
    n30152, n30153, n30154, n30155, n30156, n30157, n30158, n30159, n30160,
    n30161, n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
    n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
    n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
    n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195, n30196,
    n30197, n30198, n30199, n30200, n30201, n30202, n30203, n30204, n30205,
    n30206, n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
    n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222, n30223,
    n30224, n30225, n30226, n30227, n30228, n30229, n30230, n30231, n30232,
    n30233, n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
    n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
    n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
    n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267, n30268,
    n30269, n30270, n30271, n30272, n30273, n30274, n30275, n30276, n30277,
    n30278, n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
    n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294, n30295,
    n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30303, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
    n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
    n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339, n30340,
    n30341, n30342, n30343, n30344, n30345, n30346, n30347, n30348, n30349,
    n30350, n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
    n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366, n30367,
    n30368, n30369, n30370, n30371, n30372, n30373, n30374, n30375, n30376,
    n30377, n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
    n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
    n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
    n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411, n30412,
    n30413, n30414, n30415, n30416, n30417, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
    n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438, n30439,
    n30440, n30441, n30442, n30443, n30444, n30445, n30446, n30447, n30448,
    n30449, n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
    n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
    n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511,
    n30512, n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520,
    n30521, n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
    n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
    n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
    n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555, n30556,
    n30557, n30558, n30559, n30560, n30561, n30562, n30563, n30564, n30565,
    n30566, n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
    n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582, n30583,
    n30584, n30585, n30586, n30587, n30588, n30589, n30590, n30591, n30592,
    n30593, n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
    n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
    n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
    n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628,
    n30629, n30630, n30631, n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643, n30644, n30645, n30646,
    n30647, n30648, n30649, n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661, n30662, n30663, n30664,
    n30665, n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
    n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
    n30701, n30702, n30703, n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715, n30716, n30717, n30718,
    n30719, n30720, n30721, n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733, n30734, n30735, n30736,
    n30737, n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
    n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771, n30772,
    n30773, n30774, n30775, n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787, n30788, n30789, n30790,
    n30791, n30792, n30793, n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808,
    n30809, n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
    n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843, n30844,
    n30845, n30846, n30847, n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859, n30860, n30861, n30862,
    n30863, n30864, n30865, n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877, n30878, n30879, n30880,
    n30881, n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
    n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915, n30916,
    n30917, n30918, n30919, n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931, n30932, n30933, n30934,
    n30935, n30936, n30937, n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949, n30950, n30951, n30952,
    n30953, n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
    n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987, n30988,
    n30989, n30990, n30991, n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31004, n31005, n31006, n31007,
    n31008, n31009, n31010, n31011, n31012, n31013, n31014, n31015, n31016,
    n31017, n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
    n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
    n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
    n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052,
    n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061,
    n31062, n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070,
    n31071, n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079,
    n31080, n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088,
    n31089, n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
    n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106,
    n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
    n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124,
    n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133,
    n31134, n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142,
    n31143, n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151,
    n31152, n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160,
    n31161, n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
    n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178,
    n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
    n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196,
    n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205,
    n31206, n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214,
    n31215, n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223,
    n31224, n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232,
    n31233, n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
    n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
    n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
    n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
    n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277,
    n31278, n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286,
    n31287, n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295,
    n31296, n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304,
    n31305, n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
    n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
    n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
    n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340,
    n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349,
    n31350, n31351, n31352, n31353, n31354, n31355, n31356, n31357, n31358,
    n31359, n31360, n31361, n31362, n31363, n31364, n31365, n31366, n31367,
    n31368, n31369, n31370, n31371, n31372, n31373, n31374, n31375, n31376,
    n31377, n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
    n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394,
    n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
    n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
    n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420, n31421,
    n31422, n31423, n31424, n31425, n31426, n31427, n31428, n31429, n31430,
    n31431, n31432, n31433, n31434, n31435, n31436, n31437, n31438, n31439,
    n31440, n31441, n31442, n31443, n31444, n31445, n31446, n31447, n31448,
    n31449, n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
    n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466,
    n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
    n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484,
    n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492, n31493,
    n31494, n31495, n31496, n31497, n31498, n31499, n31500, n31501, n31502,
    n31503, n31504, n31505, n31506, n31507, n31508, n31509, n31510, n31511,
    n31512, n31513, n31514, n31515, n31516, n31517, n31518, n31519, n31520,
    n31521, n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
    n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
    n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
    n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
    n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564, n31565,
    n31566, n31567, n31568, n31569, n31570, n31571, n31572, n31573, n31574,
    n31575, n31576, n31577, n31578, n31579, n31580, n31581, n31582, n31583,
    n31584, n31585, n31586, n31587, n31588, n31589, n31590, n31591, n31592,
    n31593, n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
    n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
    n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
    n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636, n31637,
    n31638, n31639, n31640, n31641, n31642, n31643, n31644, n31645, n31646,
    n31647, n31648, n31649, n31650, n31651, n31652, n31653, n31654, n31655,
    n31656, n31657, n31658, n31659, n31660, n31661, n31662, n31663, n31664,
    n31665, n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
    n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
    n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
    n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
    n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709,
    n31710, n31711, n31712, n31713, n31714, n31715, n31716, n31717, n31718,
    n31719, n31720, n31721, n31722, n31723, n31724, n31725, n31726, n31727,
    n31728, n31729, n31730, n31731, n31732, n31733, n31734, n31735, n31736,
    n31737, n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
    n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
    n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
    n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781,
    n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
    n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
    n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
    n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
    n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
    n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
    n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
    n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853,
    n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
    n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31871,
    n31872, n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880,
    n31881, n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
    n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898,
    n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
    n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
    n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924, n31925,
    n31926, n31927, n31928, n31929, n31930, n31931, n31932, n31933, n31934,
    n31935, n31936, n31937, n31938, n31939, n31940, n31941, n31942, n31943,
    n31944, n31945, n31946, n31947, n31948, n31949, n31950, n31951, n31952,
    n31953, n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
    n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
    n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
    n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
    n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996, n31997,
    n31998, n31999, n32000, n32001, n32002, n32003, n32004, n32005, n32006,
    n32007, n32008, n32009, n32010, n32011, n32012, n32013, n32014, n32015,
    n32016, n32017, n32018, n32019, n32020, n32021, n32022, n32023, n32024,
    n32025, n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
    n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
    n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
    n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
    n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068, n32069,
    n32070, n32071, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
    n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086, n32087,
    n32088, n32089, n32090, n32091, n32092, n32093, n32094, n32095, n32096,
    n32097, n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
    n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
    n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
    n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132,
    n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140, n32141,
    n32142, n32143, n32144, n32145, n32146, n32147, n32148, n32149, n32150,
    n32151, n32152, n32153, n32154, n32155, n32156, n32157, n32158, n32159,
    n32160, n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168,
    n32169, n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
    n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
    n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
    n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204,
    n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212, n32213,
    n32214, n32215, n32216, n32217, n32218, n32219, n32220, n32221, n32222,
    n32223, n32224, n32225, n32226, n32227, n32228, n32229, n32230, n32231,
    n32232, n32233, n32234, n32235, n32236, n32237, n32238, n32239, n32240,
    n32241, n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
    n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
    n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
    n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
    n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285,
    n32286, n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294,
    n32295, n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303,
    n32304, n32305, n32306, n32307, n32308, n32309, n32310, n32311, n32312,
    n32313, n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
    n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
    n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
    n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348,
    n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356, n32357,
    n32358, n32359, n32360, n32361, n32362, n32363, n32364, n32365, n32366,
    n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374, n32375,
    n32376, n32377, n32378, n32379, n32380, n32381, n32382, n32383, n32384,
    n32385, n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
    n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
    n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428, n32429,
    n32430, n32431, n32432, n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444, n32445, n32446, n32447,
    n32448, n32449, n32450, n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
    n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500, n32501,
    n32502, n32503, n32504, n32505, n32506, n32507, n32508, n32509, n32510,
    n32511, n32512, n32513, n32514, n32515, n32516, n32517, n32518, n32519,
    n32520, n32521, n32522, n32523, n32524, n32525, n32526, n32527, n32528,
    n32529, n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
    n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
    n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
    n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
    n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572, n32573,
    n32574, n32575, n32576, n32577, n32578, n32579, n32580, n32581, n32582,
    n32583, n32584, n32585, n32586, n32587, n32588, n32589, n32590, n32591,
    n32592, n32593, n32594, n32595, n32596, n32597, n32598, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
    n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
    n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
    n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
    n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
    n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653, n32654,
    n32655, n32656, n32657, n32658, n32659, n32660, n32661, n32662, n32663,
    n32664, n32665, n32666, n32667, n32668, n32669, n32670, n32671, n32672,
    n32673, n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
    n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
    n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
    n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
    n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716, n32717,
    n32718, n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
    n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734, n32735,
    n32736, n32737, n32738, n32739, n32740, n32741, n32742, n32743, n32744,
    n32745, n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
    n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
    n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
    n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780,
    n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788, n32789,
    n32790, n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
    n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806, n32807,
    n32808, n32809, n32810, n32811, n32812, n32813, n32814, n32815, n32816,
    n32817, n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
    n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
    n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
    n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852,
    n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860, n32861,
    n32862, n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
    n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878, n32879,
    n32880, n32881, n32882, n32883, n32884, n32885, n32886, n32887, n32888,
    n32889, n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
    n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
    n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
    n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924,
    n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932, n32933,
    n32934, n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
    n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950, n32951,
    n32952, n32953, n32954, n32955, n32956, n32957, n32958, n32959, n32960,
    n32961, n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
    n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
    n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
    n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
    n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004, n33005,
    n33006, n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
    n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
    n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
    n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
    n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
    n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068, n33069,
    n33070, n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
    n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087,
    n33088, n33089, n33090, n33091, n33092, n33093, n33094, n33095, n33096,
    n33097, n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
    n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
    n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
    n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132,
    n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140, n33141,
    n33142, n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
    n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33159, n33160,
    n33161, n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
    n33170, n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
    n33180, n33181, n33182, n33183, n33185, n33186, n33187, n33188, n33189,
    n33190, n33191, n33192, n33193, n33194, n33195, n33196, n33198, n33199,
    n33200, n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208,
    n33209, n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33224, n33225, n33226, n33227, n33228,
    n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33237, n33238,
    n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
    n33258, n33259, n33260, n33261, n33263, n33264, n33265, n33266, n33267,
    n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33276, n33277,
    n33278, n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
    n33287, n33289, n33290, n33291, n33292, n33293, n33294, n33295, n33296,
    n33297, n33298, n33299, n33300, n33302, n33303, n33304, n33305, n33306,
    n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33315, n33316,
    n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324, n33325,
    n33326, n33328, n33329, n33330, n33331, n33332, n33333, n33334, n33335,
    n33336, n33337, n33338, n33339, n33341, n33342, n33343, n33344, n33345,
    n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33354, n33355,
    n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
    n33365, n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
    n33375, n33376, n33377, n33378, n33380, n33381, n33382, n33383, n33384,
    n33385, n33386, n33387, n33388, n33389, n33390, n33391, n33393, n33394,
    n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
    n33404, n33406, n33407, n33408, n33409, n33410, n33411, n33412, n33413,
    n33414, n33415, n33416, n33417, n33419, n33420, n33421, n33422, n33423,
    n33424, n33425, n33426, n33427, n33428, n33429, n33430, n33432, n33433,
    n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
    n33443, n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33458, n33459, n33460, n33461, n33462,
    n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33471, n33472,
    n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
    n33482, n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
    n33492, n33493, n33494, n33495, n33497, n33498, n33499, n33500, n33501,
    n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33510, n33511,
    n33512, n33513, n33514, n33515, n33516, n33517, n33518, n33519, n33520,
    n33521, n33522, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
    n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
    n33540, n33541, n33543, n33544, n33545, n33546, n33547, n33548, n33549,
    n33550, n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
    n33560, n33561, n33562, n33563, n33564, n33565, n33566, n33568, n33569,
    n33570, n33571, n33572, n33573, n33574, n33575, n33577, n33578, n33579,
    n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588,
    n33589, n33590, n33591, n33592, n33593, n33595, n33596, n33597, n33598,
    n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606, n33607,
    n33608, n33609, n33610, n33611, n33612, n33613, n33614, n33616, n33617,
    n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626,
    n33627, n33628, n33629, n33630, n33631, n33632, n33634, n33635, n33636,
    n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644, n33645,
    n33646, n33647, n33648, n33649, n33650, n33651, n33652, n33654, n33655,
    n33656, n33657, n33658, n33659, n33660, n33661, n33662, n33663, n33664,
    n33665, n33666, n33667, n33668, n33669, n33670, n33672, n33673, n33674,
    n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
    n33684, n33685, n33686, n33687, n33688, n33689, n33691, n33692, n33693,
    n33694, n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
    n33703, n33704, n33705, n33706, n33707, n33708, n33710, n33711, n33712,
    n33713, n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
    n33722, n33723, n33724, n33725, n33726, n33728, n33729, n33730, n33731,
    n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
    n33741, n33742, n33743, n33744, n33745, n33747, n33748, n33749, n33750,
    n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758, n33759,
    n33760, n33761, n33762, n33763, n33764, n33765, n33767, n33768, n33769,
    n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
    n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33787, n33788,
    n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796, n33797,
    n33798, n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33807,
    n33808, n33809, n33810, n33811, n33812, n33813, n33814, n33815, n33816,
    n33817, n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
    n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
    n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
    n33845, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
    n33864, n33865, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
    n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33887, n33888, n33889, n33890, n33891, n33892,
    n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900, n33901,
    n33902, n33903, n33904, n33905, n33907, n33908, n33909, n33910, n33911,
    n33912, n33913, n33914, n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33927, n33928, n33929, n33930,
    n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
    n33940, n33941, n33942, n33943, n33944, n33945, n33947, n33948, n33949,
    n33950, n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
    n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33967, n33968,
    n33969, n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
    n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33987,
    n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
    n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004, n34005,
    n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015,
    n34016, n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024,
    n34025, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
    n34044, n34045, n34047, n34048, n34049, n34050, n34051, n34052, n34053,
    n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
    n34063, n34064, n34065, n34067, n34068, n34069, n34070, n34071, n34072,
    n34073, n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
    n34082, n34083, n34084, n34085, n34087, n34088, n34089, n34090, n34091,
    n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
    n34101, n34102, n34103, n34104, n34105, n34107, n34108, n34109, n34110,
    n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118, n34119,
    n34120, n34121, n34122, n34123, n34124, n34125, n34127, n34128, n34129,
    n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
    n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34147, n34148,
    n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156, n34157,
    n34158, n34159, n34160, n34161, n34162, n34163, n34165, n34166, n34167,
    n34168, n34169, n34170, n34171, n34172, n34173, n34174, n34175, n34176,
    n34177, n34178;
  assign n644 = pi127 & ~pi353;
  assign n645 = ~pi127 & pi353;
  assign n646 = pi126 & pi352;
  assign n647 = ~pi126 & ~pi352;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n645 & ~n648;
  assign n650 = ~pi351 & n649;
  assign n651 = pi125 & n650;
  assign n652 = ~n644 & ~n651;
  assign n653 = pi125 & ~pi351;
  assign n654 = ~n644 & ~n653;
  assign n655 = ~pi125 & pi351;
  assign n656 = ~pi124 & pi350;
  assign n657 = ~n655 & ~n656;
  assign n658 = n654 & n657;
  assign n659 = n649 & n658;
  assign n660 = ~pi123 & pi349;
  assign n661 = pi122 & ~pi348;
  assign n662 = ~pi122 & pi348;
  assign n663 = ~pi347 & ~n662;
  assign n664 = pi121 & n663;
  assign n665 = ~n661 & ~n664;
  assign n666 = ~n660 & ~n665;
  assign n667 = pi124 & ~pi350;
  assign n668 = pi123 & ~pi349;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n666 & n669;
  assign n671 = n659 & ~n670;
  assign n672 = ~n660 & ~n668;
  assign n673 = ~n667 & n672;
  assign n674 = pi122 & pi348;
  assign n675 = ~pi122 & ~pi348;
  assign n676 = ~n674 & ~n675;
  assign n677 = pi121 & pi347;
  assign n678 = ~pi121 & ~pi347;
  assign n679 = ~n677 & ~n678;
  assign n680 = ~n676 & ~n679;
  assign n681 = n673 & n680;
  assign n682 = n659 & n681;
  assign n683 = pi120 & ~pi346;
  assign n684 = ~pi120 & pi346;
  assign n685 = pi119 & ~pi345;
  assign n686 = ~pi119 & pi345;
  assign n687 = ~pi344 & ~n686;
  assign n688 = pi118 & n687;
  assign n689 = ~n685 & ~n688;
  assign n690 = ~n684 & ~n689;
  assign n691 = ~n683 & ~n690;
  assign n692 = n682 & ~n691;
  assign n693 = ~n671 & ~n692;
  assign n694 = n652 & n693;
  assign n695 = ~pi117 & pi343;
  assign n696 = ~n684 & ~n695;
  assign n697 = ~n683 & n696;
  assign n698 = pi119 & pi345;
  assign n699 = ~pi119 & ~pi345;
  assign n700 = ~n698 & ~n699;
  assign n701 = pi118 & pi344;
  assign n702 = ~pi118 & ~pi344;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n700 & ~n703;
  assign n705 = n697 & n704;
  assign n706 = n682 & n705;
  assign n707 = pi117 & ~pi343;
  assign n708 = pi116 & ~pi342;
  assign n709 = ~n707 & ~n708;
  assign n710 = n706 & ~n709;
  assign n711 = n694 & ~n710;
  assign n712 = pi116 & pi342;
  assign n713 = ~pi116 & ~pi342;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n707 & ~n714;
  assign n716 = n706 & n715;
  assign n717 = ~pi115 & pi341;
  assign n718 = ~pi340 & ~n717;
  assign n719 = pi114 & n718;
  assign n720 = pi115 & ~pi341;
  assign n721 = ~n719 & ~n720;
  assign n722 = n716 & ~n721;
  assign n723 = n711 & ~n722;
  assign n724 = pi115 & pi341;
  assign n725 = ~pi115 & ~pi341;
  assign n726 = ~n724 & ~n725;
  assign n727 = pi114 & pi340;
  assign n728 = ~pi114 & ~pi340;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n726 & ~n729;
  assign n731 = n716 & n730;
  assign n732 = ~pi113 & pi339;
  assign n733 = ~pi338 & ~n732;
  assign n734 = pi112 & n733;
  assign n735 = pi113 & ~pi339;
  assign n736 = ~n734 & ~n735;
  assign n737 = n731 & ~n736;
  assign n738 = n723 & ~n737;
  assign n739 = pi113 & pi339;
  assign n740 = ~pi113 & ~pi339;
  assign n741 = ~n739 & ~n740;
  assign n742 = pi112 & pi338;
  assign n743 = ~pi112 & ~pi338;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n741 & ~n744;
  assign n746 = n731 & n745;
  assign n747 = ~pi111 & pi337;
  assign n748 = ~pi336 & ~n747;
  assign n749 = pi110 & n748;
  assign n750 = pi111 & ~pi337;
  assign n751 = ~n749 & ~n750;
  assign n752 = n746 & ~n751;
  assign n753 = n738 & ~n752;
  assign n754 = pi111 & pi337;
  assign n755 = ~pi111 & ~pi337;
  assign n756 = ~n754 & ~n755;
  assign n757 = pi110 & pi336;
  assign n758 = ~pi110 & ~pi336;
  assign n759 = ~n757 & ~n758;
  assign n760 = ~n756 & ~n759;
  assign n761 = n746 & n760;
  assign n762 = ~pi109 & pi335;
  assign n763 = ~pi334 & ~n762;
  assign n764 = pi108 & n763;
  assign n765 = pi109 & ~pi335;
  assign n766 = ~n764 & ~n765;
  assign n767 = n761 & ~n766;
  assign n768 = n753 & ~n767;
  assign n769 = pi109 & pi335;
  assign n770 = ~pi109 & ~pi335;
  assign n771 = ~n769 & ~n770;
  assign n772 = pi108 & pi334;
  assign n773 = ~pi108 & ~pi334;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n771 & ~n774;
  assign n776 = n761 & n775;
  assign n777 = pi107 & ~pi333;
  assign n778 = ~pi107 & pi333;
  assign n779 = ~pi332 & ~n778;
  assign n780 = pi106 & n779;
  assign n781 = ~n777 & ~n780;
  assign n782 = ~n777 & ~n778;
  assign n783 = pi106 & ~pi332;
  assign n784 = ~pi106 & pi332;
  assign n785 = ~pi105 & pi331;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~n783 & n786;
  assign n788 = n782 & n787;
  assign n789 = pi105 & ~pi331;
  assign n790 = pi104 & ~pi330;
  assign n791 = ~n789 & ~n790;
  assign n792 = pi102 & ~pi328;
  assign n793 = ~pi102 & pi328;
  assign n794 = ~pi100 & pi326;
  assign n795 = pi100 & ~pi326;
  assign n796 = pi098 & ~pi324;
  assign n797 = ~pi098 & pi324;
  assign n798 = pi097 & ~pi323;
  assign n799 = ~pi097 & pi323;
  assign n800 = ~pi322 & ~n799;
  assign n801 = pi096 & n800;
  assign n802 = ~n798 & ~n801;
  assign n803 = ~n797 & ~n802;
  assign n804 = ~n796 & ~n803;
  assign n805 = pi325 & n804;
  assign n806 = ~pi325 & ~n804;
  assign n807 = ~pi099 & ~n806;
  assign n808 = ~n805 & ~n807;
  assign n809 = ~n795 & ~n808;
  assign n810 = ~n794 & ~n809;
  assign n811 = pi327 & ~n810;
  assign n812 = pi101 & ~n811;
  assign n813 = ~pi327 & n810;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n793 & ~n814;
  assign n816 = ~n792 & ~n815;
  assign n817 = ~pi329 & ~n816;
  assign n818 = ~pi103 & ~n817;
  assign n819 = pi329 & n816;
  assign n820 = ~pi104 & pi330;
  assign n821 = n791 & ~n820;
  assign n822 = ~n819 & n821;
  assign n823 = ~n818 & n822;
  assign n824 = n791 & ~n823;
  assign n825 = n788 & ~n824;
  assign n826 = n781 & ~n825;
  assign n827 = n776 & ~n826;
  assign n828 = n768 & ~n827;
  assign n829 = ~pi352 & ~n645;
  assign n830 = pi126 & n829;
  assign n831 = n828 & ~n830;
  assign n832 = pi161 & n831;
  assign po096 = ~pi160 & ~n832;
  assign n834 = ~pi160 & pi161;
  assign n835 = n831 & n834;
  assign n836 = pi258 & n835;
  assign n837 = pi162 & ~n835;
  assign po097 = n836 | n837;
  assign n839 = pi259 & n835;
  assign n840 = pi163 & ~n835;
  assign po098 = n839 | n840;
  assign n842 = pi268 & n835;
  assign n843 = pi164 & ~n835;
  assign po099 = n842 | n843;
  assign n845 = pi269 & n835;
  assign n846 = pi165 & ~n835;
  assign po100 = n845 | n846;
  assign n848 = pi270 & n835;
  assign n849 = pi166 & ~n835;
  assign po101 = n848 | n849;
  assign n851 = pi271 & n835;
  assign n852 = pi167 & ~n835;
  assign po102 = n851 | n852;
  assign n854 = pi272 & n835;
  assign n855 = pi168 & ~n835;
  assign po103 = n854 | n855;
  assign n857 = pi273 & n835;
  assign n858 = pi169 & ~n835;
  assign po104 = n857 | n858;
  assign n860 = pi274 & n835;
  assign n861 = pi170 & ~n835;
  assign po105 = n860 | n861;
  assign n863 = pi275 & n835;
  assign n864 = pi171 & ~n835;
  assign po106 = n863 | n864;
  assign n866 = pi276 & n835;
  assign n867 = pi172 & ~n835;
  assign po107 = n866 | n867;
  assign n869 = pi277 & n835;
  assign n870 = pi173 & ~n835;
  assign po108 = n869 | n870;
  assign n872 = pi260 & n835;
  assign n873 = pi174 & ~n835;
  assign po109 = n872 | n873;
  assign n875 = pi278 & n835;
  assign n876 = pi175 & ~n835;
  assign po110 = n875 | n876;
  assign n878 = pi279 & n835;
  assign n879 = pi176 & ~n835;
  assign po111 = n878 | n879;
  assign n881 = pi280 & n835;
  assign n882 = pi177 & ~n835;
  assign po112 = n881 | n882;
  assign n884 = pi281 & n835;
  assign n885 = pi178 & ~n835;
  assign po113 = n884 | n885;
  assign n887 = pi282 & n835;
  assign n888 = pi179 & ~n835;
  assign po114 = n887 | n888;
  assign n890 = pi283 & n835;
  assign n891 = pi180 & ~n835;
  assign po115 = n890 | n891;
  assign n893 = pi284 & n835;
  assign n894 = pi181 & ~n835;
  assign po116 = n893 | n894;
  assign n896 = pi285 & n835;
  assign n897 = pi182 & ~n835;
  assign po117 = n896 | n897;
  assign n899 = pi286 & n835;
  assign n900 = pi183 & ~n835;
  assign po118 = n899 | n900;
  assign n902 = pi287 & n835;
  assign n903 = pi184 & ~n835;
  assign po119 = n902 | n903;
  assign n905 = pi261 & n835;
  assign n906 = pi185 & ~n835;
  assign po120 = n905 | n906;
  assign n908 = pi288 & n835;
  assign n909 = pi186 & ~n835;
  assign po121 = n908 | n909;
  assign n911 = pi289 & n835;
  assign n912 = pi187 & ~n835;
  assign po122 = n911 | n912;
  assign n914 = pi262 & n835;
  assign n915 = pi188 & ~n835;
  assign po123 = n914 | n915;
  assign n917 = pi263 & n835;
  assign n918 = pi189 & ~n835;
  assign po124 = n917 | n918;
  assign n920 = pi264 & n835;
  assign n921 = pi190 & ~n835;
  assign po125 = n920 | n921;
  assign n923 = pi265 & n835;
  assign n924 = pi191 & ~n835;
  assign po126 = n923 | n924;
  assign n926 = pi266 & n835;
  assign n927 = pi192 & ~n835;
  assign po127 = n926 | n927;
  assign n929 = pi267 & n835;
  assign n930 = pi193 & ~n835;
  assign po128 = n929 | n930;
  assign n932 = pi322 & n835;
  assign n933 = pi194 & ~n835;
  assign po129 = n932 | n933;
  assign n935 = pi323 & n835;
  assign n936 = pi195 & ~n835;
  assign po130 = n935 | n936;
  assign n938 = pi332 & n835;
  assign n939 = pi196 & ~n835;
  assign po131 = n938 | n939;
  assign n941 = pi333 & n835;
  assign n942 = pi197 & ~n835;
  assign po132 = n941 | n942;
  assign n944 = pi334 & n835;
  assign n945 = pi198 & ~n835;
  assign po133 = n944 | n945;
  assign n947 = pi335 & n835;
  assign n948 = pi199 & ~n835;
  assign po134 = n947 | n948;
  assign n950 = pi336 & n835;
  assign n951 = pi200 & ~n835;
  assign po135 = n950 | n951;
  assign n953 = pi337 & n835;
  assign n954 = pi201 & ~n835;
  assign po136 = n953 | n954;
  assign n956 = pi338 & n835;
  assign n957 = pi202 & ~n835;
  assign po137 = n956 | n957;
  assign n959 = pi339 & n835;
  assign n960 = pi203 & ~n835;
  assign po138 = n959 | n960;
  assign n962 = pi340 & n835;
  assign n963 = pi204 & ~n835;
  assign po139 = n962 | n963;
  assign n965 = pi341 & n835;
  assign n966 = pi205 & ~n835;
  assign po140 = n965 | n966;
  assign n968 = pi324 & n835;
  assign n969 = pi206 & ~n835;
  assign po141 = n968 | n969;
  assign n971 = pi342 & n835;
  assign n972 = pi207 & ~n835;
  assign po142 = n971 | n972;
  assign n974 = pi343 & n835;
  assign n975 = pi208 & ~n835;
  assign po143 = n974 | n975;
  assign n977 = pi344 & n835;
  assign n978 = pi209 & ~n835;
  assign po144 = n977 | n978;
  assign n980 = pi345 & n835;
  assign n981 = pi210 & ~n835;
  assign po145 = n980 | n981;
  assign n983 = pi346 & n835;
  assign n984 = pi211 & ~n835;
  assign po146 = n983 | n984;
  assign n986 = pi347 & n835;
  assign n987 = pi212 & ~n835;
  assign po147 = n986 | n987;
  assign n989 = pi348 & n835;
  assign n990 = pi213 & ~n835;
  assign po148 = n989 | n990;
  assign n992 = pi349 & n835;
  assign n993 = pi214 & ~n835;
  assign po149 = n992 | n993;
  assign n995 = pi350 & n835;
  assign n996 = pi215 & ~n835;
  assign po150 = n995 | n996;
  assign n998 = pi351 & n835;
  assign n999 = pi216 & ~n835;
  assign po151 = n998 | n999;
  assign n1001 = pi325 & n835;
  assign n1002 = pi217 & ~n835;
  assign po152 = n1001 | n1002;
  assign n1004 = ~pi160 & n832;
  assign n1005 = pi218 & ~n1004;
  assign n1006 = pi352 & n828;
  assign n1007 = n834 & n1006;
  assign po153 = n1005 | n1007;
  assign n1009 = pi353 & n835;
  assign n1010 = pi219 & ~n835;
  assign po154 = n1009 | n1010;
  assign n1012 = pi326 & n835;
  assign n1013 = pi220 & ~n835;
  assign po155 = n1012 | n1013;
  assign n1015 = pi327 & n835;
  assign n1016 = pi221 & ~n835;
  assign po156 = n1015 | n1016;
  assign n1018 = pi328 & n835;
  assign n1019 = pi222 & ~n835;
  assign po157 = n1018 | n1019;
  assign n1021 = pi329 & n835;
  assign n1022 = pi223 & ~n835;
  assign po158 = n1021 | n1022;
  assign n1024 = pi330 & n835;
  assign n1025 = pi224 & ~n835;
  assign po159 = n1024 | n1025;
  assign n1027 = pi331 & n835;
  assign n1028 = pi225 & ~n835;
  assign po160 = n1027 | n1028;
  assign n1030 = pi321 & n835;
  assign n1031 = pi226 & ~n835;
  assign po161 = n1030 | n1031;
  assign n1033 = pi320 & n835;
  assign n1034 = pi227 & ~n835;
  assign po162 = n1033 | n1034;
  assign n1036 = pi311 & n835;
  assign n1037 = pi228 & ~n835;
  assign po163 = n1036 | n1037;
  assign n1039 = pi310 & n835;
  assign n1040 = pi229 & ~n835;
  assign po164 = n1039 | n1040;
  assign n1042 = pi309 & n835;
  assign n1043 = pi230 & ~n835;
  assign po165 = n1042 | n1043;
  assign n1045 = pi308 & n835;
  assign n1046 = pi231 & ~n835;
  assign po166 = n1045 | n1046;
  assign n1048 = pi307 & n835;
  assign n1049 = pi232 & ~n835;
  assign po167 = n1048 | n1049;
  assign n1051 = pi306 & n835;
  assign n1052 = pi233 & ~n835;
  assign po168 = n1051 | n1052;
  assign n1054 = pi305 & n835;
  assign n1055 = pi234 & ~n835;
  assign po169 = n1054 | n1055;
  assign n1057 = pi304 & n835;
  assign n1058 = pi235 & ~n835;
  assign po170 = n1057 | n1058;
  assign n1060 = pi303 & n835;
  assign n1061 = pi236 & ~n835;
  assign po171 = n1060 | n1061;
  assign n1063 = pi302 & n835;
  assign n1064 = pi237 & ~n835;
  assign po172 = n1063 | n1064;
  assign n1066 = pi319 & n835;
  assign n1067 = pi238 & ~n835;
  assign po173 = n1066 | n1067;
  assign n1069 = pi301 & n835;
  assign n1070 = pi239 & ~n835;
  assign po174 = n1069 | n1070;
  assign n1072 = pi300 & n835;
  assign n1073 = pi240 & ~n835;
  assign po175 = n1072 | n1073;
  assign n1075 = pi299 & n835;
  assign n1076 = pi241 & ~n835;
  assign po176 = n1075 | n1076;
  assign n1078 = pi298 & n835;
  assign n1079 = pi242 & ~n835;
  assign po177 = n1078 | n1079;
  assign n1081 = pi297 & n835;
  assign n1082 = pi243 & ~n835;
  assign po178 = n1081 | n1082;
  assign n1084 = pi296 & n835;
  assign n1085 = pi244 & ~n835;
  assign po179 = n1084 | n1085;
  assign n1087 = pi295 & n835;
  assign n1088 = pi245 & ~n835;
  assign po180 = n1087 | n1088;
  assign n1090 = pi294 & n835;
  assign n1091 = pi246 & ~n835;
  assign po181 = n1090 | n1091;
  assign n1093 = pi293 & n835;
  assign n1094 = pi247 & ~n835;
  assign po182 = n1093 | n1094;
  assign n1096 = pi292 & n835;
  assign n1097 = pi248 & ~n835;
  assign po183 = n1096 | n1097;
  assign n1099 = pi318 & n835;
  assign n1100 = pi249 & ~n835;
  assign po184 = n1099 | n1100;
  assign n1102 = pi291 & n835;
  assign n1103 = pi250 & ~n835;
  assign po185 = n1102 | n1103;
  assign n1105 = pi290 & n835;
  assign n1106 = pi251 & ~n835;
  assign po186 = n1105 | n1106;
  assign n1108 = pi317 & n835;
  assign n1109 = pi252 & ~n835;
  assign po187 = n1108 | n1109;
  assign n1111 = pi316 & n835;
  assign n1112 = pi253 & ~n835;
  assign po188 = n1111 | n1112;
  assign n1114 = pi315 & n835;
  assign n1115 = pi254 & ~n835;
  assign po189 = n1114 | n1115;
  assign n1117 = pi314 & n835;
  assign n1118 = pi255 & ~n835;
  assign po190 = n1117 | n1118;
  assign n1120 = pi313 & n835;
  assign n1121 = pi256 & ~n835;
  assign po191 = n1120 | n1121;
  assign n1123 = pi312 & n835;
  assign n1124 = pi257 & ~n835;
  assign po192 = n1123 | n1124;
  assign n1126 = pi064 & ~pi161;
  assign n1127 = pi258 & n831;
  assign n1128 = pi258 & pi322;
  assign n1129 = pi128 & ~pi258;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = pi321 & ~n1130;
  assign n1132 = ~pi321 & ~pi322;
  assign n1133 = pi128 & ~n1132;
  assign n1134 = pi258 & ~n1133;
  assign n1135 = ~n1131 & ~n1134;
  assign n1136 = ~n831 & ~n1135;
  assign n1137 = ~n1127 & ~n1136;
  assign n1138 = pi161 & ~n1137;
  assign n1139 = ~n1126 & ~n1138;
  assign po193 = ~pi160 & ~n1139;
  assign n1141 = pi065 & ~pi161;
  assign n1142 = pi259 & n831;
  assign n1143 = pi258 & ~pi322;
  assign n1144 = pi321 & ~n1143;
  assign n1145 = pi128 & n1144;
  assign n1146 = ~pi258 & pi259;
  assign n1147 = pi258 & ~pi259;
  assign n1148 = ~pi129 & n1147;
  assign n1149 = ~n1146 & ~n1148;
  assign n1150 = pi128 & ~n1149;
  assign n1151 = pi128 & ~pi259;
  assign n1152 = pi258 & ~n1151;
  assign n1153 = pi129 & n1152;
  assign n1154 = ~n1150 & ~n1153;
  assign n1155 = pi322 & ~n1154;
  assign n1156 = pi128 & pi258;
  assign n1157 = pi323 & n1156;
  assign n1158 = ~pi259 & ~n1157;
  assign n1159 = pi259 & pi323;
  assign n1160 = n1156 & n1159;
  assign n1161 = ~n1158 & ~n1160;
  assign n1162 = ~n1155 & ~n1161;
  assign n1163 = pi259 & ~n1157;
  assign n1164 = ~pi259 & pi323;
  assign n1165 = n1156 & n1164;
  assign n1166 = ~n1163 & ~n1165;
  assign n1167 = ~n1154 & ~n1166;
  assign n1168 = pi322 & n1167;
  assign n1169 = ~n1162 & ~n1168;
  assign n1170 = ~n1145 & ~n1169;
  assign n1171 = n1145 & n1169;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = pi129 & pi321;
  assign n1174 = ~pi128 & ~n1173;
  assign n1175 = pi128 & pi129;
  assign n1176 = pi321 & ~n1175;
  assign n1177 = ~pi320 & ~n1176;
  assign n1178 = pi320 & pi321;
  assign n1179 = ~pi129 & n1178;
  assign n1180 = ~n1177 & ~n1179;
  assign n1181 = ~n1174 & n1180;
  assign n1182 = ~n1172 & ~n1181;
  assign n1183 = ~n1145 & n1169;
  assign n1184 = n1145 & ~n1169;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = pi320 & ~pi321;
  assign n1187 = ~pi320 & pi321;
  assign n1188 = ~pi129 & n1187;
  assign n1189 = ~n1186 & ~n1188;
  assign n1190 = pi128 & ~n1189;
  assign n1191 = pi128 & ~pi320;
  assign n1192 = pi321 & ~n1191;
  assign n1193 = pi129 & n1192;
  assign n1194 = ~n1190 & ~n1193;
  assign n1195 = ~n1185 & ~n1194;
  assign n1196 = ~n1182 & ~n1195;
  assign n1197 = ~n831 & n1196;
  assign n1198 = ~n1142 & ~n1197;
  assign n1199 = pi161 & ~n1198;
  assign n1200 = ~n1141 & ~n1199;
  assign po194 = ~pi160 & ~n1200;
  assign n1202 = pi260 & n831;
  assign n1203 = pi130 & pi321;
  assign n1204 = ~pi128 & n1203;
  assign n1205 = pi128 & ~pi319;
  assign n1206 = n1186 & n1205;
  assign n1207 = ~n1204 & ~n1206;
  assign n1208 = ~pi129 & ~n1207;
  assign n1209 = pi130 & ~pi319;
  assign n1210 = ~pi130 & pi319;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = pi128 & ~n1211;
  assign n1213 = pi130 & pi320;
  assign n1214 = ~pi130 & ~pi320;
  assign n1215 = pi129 & n1214;
  assign n1216 = ~n1213 & ~n1215;
  assign n1217 = ~pi128 & ~n1216;
  assign n1218 = ~n1212 & ~n1217;
  assign n1219 = pi321 & ~n1218;
  assign n1220 = pi320 & ~n1205;
  assign n1221 = pi129 & n1220;
  assign n1222 = pi319 & ~pi320;
  assign n1223 = pi128 & n1222;
  assign n1224 = ~n1221 & ~n1223;
  assign n1225 = ~pi321 & ~n1224;
  assign n1226 = ~n1219 & ~n1225;
  assign n1227 = ~n1208 & n1226;
  assign n1228 = pi323 & ~n1154;
  assign n1229 = pi324 & n1156;
  assign n1230 = ~pi322 & n1229;
  assign n1231 = pi259 & ~pi260;
  assign n1232 = n1129 & n1231;
  assign n1233 = pi130 & pi258;
  assign n1234 = ~pi128 & n1233;
  assign n1235 = ~n1232 & ~n1234;
  assign n1236 = ~pi129 & ~n1235;
  assign n1237 = pi130 & pi259;
  assign n1238 = ~pi130 & ~pi259;
  assign n1239 = pi129 & n1238;
  assign n1240 = ~n1237 & ~n1239;
  assign n1241 = ~pi128 & ~n1240;
  assign n1242 = pi130 & ~pi260;
  assign n1243 = ~pi130 & pi260;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = pi128 & ~n1244;
  assign n1246 = ~n1241 & ~n1245;
  assign n1247 = pi258 & ~n1246;
  assign n1248 = pi128 & ~pi260;
  assign n1249 = pi259 & ~n1248;
  assign n1250 = pi129 & n1249;
  assign n1251 = ~pi259 & pi260;
  assign n1252 = pi128 & n1251;
  assign n1253 = ~n1250 & ~n1252;
  assign n1254 = ~pi258 & ~n1253;
  assign n1255 = ~n1247 & ~n1254;
  assign n1256 = ~n1236 & n1255;
  assign n1257 = ~n1156 & ~n1256;
  assign n1258 = pi322 & n1257;
  assign n1259 = ~n1230 & ~n1258;
  assign n1260 = ~n1228 & ~n1259;
  assign n1261 = pi324 & n1256;
  assign n1262 = ~pi324 & ~n1256;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n1156 & ~n1263;
  assign n1265 = pi322 & n1264;
  assign n1266 = ~pi322 & ~n1229;
  assign n1267 = ~n1156 & n1256;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~n1154 & ~n1268;
  assign n1270 = pi323 & n1269;
  assign n1271 = ~n1265 & ~n1270;
  assign n1272 = ~n1260 & n1271;
  assign n1273 = n1227 & n1272;
  assign n1274 = ~n1227 & ~n1272;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = pi258 & ~n1155;
  assign n1277 = pi128 & n1276;
  assign n1278 = pi323 & n1277;
  assign n1279 = ~n1154 & ~n1157;
  assign n1280 = pi322 & n1279;
  assign n1281 = ~n1278 & ~n1280;
  assign n1282 = ~pi259 & ~n1281;
  assign n1283 = pi260 & n1282;
  assign n1284 = ~pi260 & ~n1282;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n1275 & ~n1285;
  assign n1287 = ~n1227 & n1272;
  assign n1288 = n1227 & ~n1272;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~pi260 & n1282;
  assign n1291 = pi260 & ~n1282;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = ~n1289 & ~n1292;
  assign n1294 = ~n1286 & ~n1293;
  assign n1295 = ~n1183 & ~n1194;
  assign n1296 = ~n1184 & ~n1295;
  assign n1297 = n1294 & n1296;
  assign n1298 = ~n1294 & ~n1296;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = ~n831 & ~n1299;
  assign n1301 = ~n1202 & ~n1300;
  assign n1302 = pi161 & ~n1301;
  assign n1303 = pi066 & ~pi161;
  assign n1304 = ~n1302 & ~n1303;
  assign po195 = ~pi160 & ~n1304;
  assign n1306 = pi261 & n831;
  assign n1307 = pi129 & pi319;
  assign n1308 = ~pi128 & ~n1307;
  assign n1309 = pi319 & ~n1175;
  assign n1310 = ~pi318 & ~n1309;
  assign n1311 = pi318 & pi319;
  assign n1312 = ~pi129 & n1311;
  assign n1313 = ~n1310 & ~n1312;
  assign n1314 = ~n1308 & n1313;
  assign n1315 = ~pi129 & n1186;
  assign n1316 = ~n1203 & ~n1315;
  assign n1317 = pi319 & ~n1316;
  assign n1318 = pi128 & n1317;
  assign n1319 = pi129 & ~pi130;
  assign n1320 = ~pi320 & ~n1319;
  assign n1321 = pi128 & ~n1320;
  assign n1322 = pi130 & ~pi320;
  assign n1323 = ~pi129 & n1322;
  assign n1324 = ~n1321 & ~n1323;
  assign n1325 = ~pi131 & ~n1324;
  assign n1326 = ~pi128 & ~n1322;
  assign n1327 = pi129 & pi130;
  assign n1328 = ~pi129 & ~pi130;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = ~pi320 & ~n1329;
  assign n1331 = ~n1326 & ~n1330;
  assign n1332 = pi131 & ~n1331;
  assign n1333 = ~n1325 & ~n1332;
  assign n1334 = pi321 & ~n1333;
  assign n1335 = ~pi128 & pi129;
  assign n1336 = pi130 & ~n1335;
  assign n1337 = ~pi128 & n1319;
  assign n1338 = ~n1336 & ~n1337;
  assign n1339 = ~pi321 & ~n1338;
  assign n1340 = pi320 & n1339;
  assign n1341 = ~n1334 & ~n1340;
  assign n1342 = ~n1318 & ~n1341;
  assign n1343 = n1318 & n1341;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1314 & ~n1344;
  assign n1346 = ~n1318 & n1341;
  assign n1347 = n1318 & ~n1341;
  assign n1348 = ~n1346 & ~n1347;
  assign n1349 = pi318 & ~pi319;
  assign n1350 = ~pi318 & pi319;
  assign n1351 = ~pi129 & n1350;
  assign n1352 = ~n1349 & ~n1351;
  assign n1353 = pi128 & ~n1352;
  assign n1354 = pi128 & ~pi318;
  assign n1355 = pi319 & ~n1354;
  assign n1356 = pi129 & n1355;
  assign n1357 = ~n1353 & ~n1356;
  assign n1358 = ~n1348 & ~n1357;
  assign n1359 = ~n1345 & ~n1358;
  assign n1360 = ~n1272 & n1282;
  assign n1361 = n1272 & ~n1282;
  assign n1362 = ~pi260 & ~n1361;
  assign n1363 = ~n1360 & ~n1362;
  assign n1364 = pi322 & ~n1256;
  assign n1365 = ~pi322 & n1228;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = n1156 & ~n1366;
  assign n1368 = pi324 & n1367;
  assign n1369 = ~n1154 & ~n1267;
  assign n1370 = pi323 & n1369;
  assign n1371 = pi322 & n1370;
  assign n1372 = ~n1368 & n1371;
  assign n1373 = n1368 & ~n1371;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = pi323 & ~n1256;
  assign n1376 = pi260 & pi261;
  assign n1377 = ~pi260 & ~pi261;
  assign n1378 = n1156 & n1377;
  assign n1379 = ~n1376 & ~n1378;
  assign n1380 = pi259 & ~n1379;
  assign n1381 = ~pi259 & ~pi261;
  assign n1382 = pi128 & ~n1381;
  assign n1383 = pi260 & ~n1382;
  assign n1384 = ~n1380 & ~n1383;
  assign n1385 = pi129 & ~n1384;
  assign n1386 = pi258 & pi259;
  assign n1387 = ~pi260 & ~n1386;
  assign n1388 = pi129 & ~n1387;
  assign n1389 = pi261 & ~n1388;
  assign n1390 = pi128 & n1389;
  assign n1391 = ~n1385 & ~n1390;
  assign n1392 = ~pi129 & n1233;
  assign n1393 = pi129 & n1146;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~pi128 & ~n1394;
  assign n1396 = pi258 & n1231;
  assign n1397 = ~n1251 & ~n1396;
  assign n1398 = ~n1329 & ~n1397;
  assign n1399 = ~pi259 & ~pi260;
  assign n1400 = pi259 & pi260;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = pi258 & ~n1401;
  assign n1403 = ~pi130 & n1402;
  assign n1404 = pi129 & n1403;
  assign n1405 = ~pi258 & n1251;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1398 & n1406;
  assign n1408 = pi128 & ~n1407;
  assign n1409 = pi130 & n1402;
  assign n1410 = ~pi129 & n1409;
  assign n1411 = ~n1408 & ~n1410;
  assign n1412 = ~n1395 & n1411;
  assign n1413 = ~n1391 & n1412;
  assign n1414 = n1391 & ~n1412;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = pi129 & pi259;
  assign n1417 = ~pi128 & n1416;
  assign n1418 = pi128 & pi260;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = pi258 & ~n1419;
  assign n1421 = pi130 & n1420;
  assign n1422 = ~n1237 & ~n1421;
  assign n1423 = n1237 & n1421;
  assign n1424 = ~n1422 & ~n1423;
  assign n1425 = pi258 & ~n1424;
  assign n1426 = pi131 & n1425;
  assign n1427 = pi131 & pi258;
  assign n1428 = ~n1237 & n1421;
  assign n1429 = n1237 & ~n1421;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = ~n1427 & ~n1430;
  assign n1432 = ~n1426 & ~n1431;
  assign n1433 = ~n1415 & ~n1432;
  assign n1434 = ~n1391 & ~n1412;
  assign n1435 = n1391 & n1412;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = pi258 & ~n1430;
  assign n1438 = pi131 & n1437;
  assign n1439 = ~n1424 & ~n1427;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1436 & ~n1440;
  assign n1442 = ~n1433 & ~n1441;
  assign n1443 = pi322 & n1442;
  assign n1444 = ~n1375 & ~n1443;
  assign n1445 = pi322 & pi323;
  assign n1446 = ~n1256 & n1442;
  assign n1447 = n1445 & n1446;
  assign n1448 = ~n1444 & ~n1447;
  assign n1449 = ~n1374 & ~n1448;
  assign n1450 = n1368 & n1371;
  assign n1451 = ~n1368 & ~n1371;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~n1375 & n1442;
  assign n1454 = pi322 & n1453;
  assign n1455 = ~n1256 & ~n1443;
  assign n1456 = pi323 & n1455;
  assign n1457 = ~n1454 & ~n1456;
  assign n1458 = ~n1452 & ~n1457;
  assign n1459 = ~n1449 & ~n1458;
  assign n1460 = pi324 & ~n1154;
  assign n1461 = n1459 & ~n1460;
  assign n1462 = ~n1154 & ~n1459;
  assign n1463 = pi324 & n1462;
  assign n1464 = ~n1461 & ~n1463;
  assign n1465 = pi325 & n1156;
  assign n1466 = n1464 & ~n1465;
  assign n1467 = pi325 & ~n1464;
  assign n1468 = n1156 & n1467;
  assign n1469 = ~n1466 & ~n1468;
  assign n1470 = ~n1363 & ~n1469;
  assign n1471 = n1363 & n1469;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = pi261 & ~n1472;
  assign n1474 = ~n1363 & n1469;
  assign n1475 = n1363 & ~n1469;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~pi261 & ~n1476;
  assign n1478 = ~n1473 & ~n1477;
  assign n1479 = n1227 & n1296;
  assign n1480 = ~n1227 & ~n1296;
  assign n1481 = ~n1360 & ~n1361;
  assign n1482 = pi260 & ~n1481;
  assign n1483 = ~n1272 & ~n1282;
  assign n1484 = n1272 & n1282;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = ~pi260 & ~n1485;
  assign n1487 = ~n1482 & ~n1486;
  assign n1488 = ~n1480 & ~n1487;
  assign n1489 = ~n1479 & ~n1488;
  assign n1490 = n1478 & ~n1489;
  assign n1491 = ~n1478 & n1489;
  assign n1492 = ~n1490 & ~n1491;
  assign n1493 = ~n1359 & ~n1492;
  assign n1494 = n1478 & n1489;
  assign n1495 = ~n1478 & ~n1489;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = n1359 & ~n1496;
  assign n1498 = ~n1493 & ~n1497;
  assign n1499 = ~n831 & ~n1498;
  assign n1500 = ~n1306 & ~n1499;
  assign n1501 = pi161 & ~n1500;
  assign n1502 = pi067 & ~pi161;
  assign n1503 = ~n1501 & ~n1502;
  assign po196 = ~pi160 & ~n1503;
  assign n1505 = pi262 & n831;
  assign n1506 = ~pi129 & pi319;
  assign n1507 = ~n1344 & ~n1506;
  assign n1508 = pi319 & ~n1348;
  assign n1509 = ~pi129 & n1508;
  assign n1510 = ~n1507 & ~n1509;
  assign n1511 = pi318 & ~n1510;
  assign n1512 = pi128 & n1511;
  assign n1513 = ~pi130 & ~n1335;
  assign n1514 = ~pi128 & n1327;
  assign n1515 = ~n1513 & ~n1514;
  assign n1516 = pi131 & ~pi132;
  assign n1517 = pi128 & n1516;
  assign n1518 = ~pi131 & pi132;
  assign n1519 = pi130 & n1518;
  assign n1520 = ~n1517 & ~n1519;
  assign n1521 = pi129 & ~n1520;
  assign n1522 = ~pi131 & ~pi132;
  assign n1523 = pi131 & pi132;
  assign n1524 = ~pi130 & n1523;
  assign n1525 = ~n1522 & ~n1524;
  assign n1526 = ~pi129 & ~n1525;
  assign n1527 = ~pi128 & n1523;
  assign n1528 = ~n1522 & ~n1527;
  assign n1529 = ~pi130 & ~n1528;
  assign n1530 = pi130 & n1516;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = ~n1526 & n1531;
  assign n1533 = ~n1521 & n1532;
  assign n1534 = pi321 & n1533;
  assign n1535 = pi131 & ~n1319;
  assign n1536 = pi128 & n1535;
  assign n1537 = pi130 & ~pi131;
  assign n1538 = ~pi129 & n1537;
  assign n1539 = ~n1337 & ~n1538;
  assign n1540 = ~n1536 & n1539;
  assign n1541 = pi321 & ~n1540;
  assign n1542 = pi320 & n1541;
  assign n1543 = ~pi130 & pi131;
  assign n1544 = pi128 & n1543;
  assign n1545 = ~n1537 & ~n1544;
  assign n1546 = pi129 & ~n1545;
  assign n1547 = ~pi130 & ~pi131;
  assign n1548 = pi130 & pi131;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~pi129 & ~n1549;
  assign n1551 = ~pi128 & n1547;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = ~n1546 & n1552;
  assign n1554 = pi320 & n1553;
  assign n1555 = n1542 & ~n1554;
  assign n1556 = ~n1542 & n1553;
  assign n1557 = pi320 & n1556;
  assign n1558 = ~n1555 & ~n1557;
  assign n1559 = ~n1534 & ~n1558;
  assign n1560 = ~n1542 & ~n1554;
  assign n1561 = n1542 & n1553;
  assign n1562 = pi320 & n1561;
  assign n1563 = ~n1560 & ~n1562;
  assign n1564 = n1533 & ~n1563;
  assign n1565 = pi321 & n1564;
  assign n1566 = ~n1559 & ~n1565;
  assign n1567 = pi128 & ~pi129;
  assign n1568 = ~n1335 & ~n1567;
  assign n1569 = ~n1346 & ~n1568;
  assign n1570 = pi319 & n1569;
  assign n1571 = ~n1347 & ~n1570;
  assign n1572 = n1566 & ~n1571;
  assign n1573 = ~n1566 & n1571;
  assign n1574 = ~n1572 & ~n1573;
  assign n1575 = n1515 & ~n1574;
  assign n1576 = pi319 & n1575;
  assign n1577 = pi319 & n1515;
  assign n1578 = ~n1566 & ~n1571;
  assign n1579 = n1566 & n1571;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n1577 & ~n1580;
  assign n1582 = ~n1576 & ~n1581;
  assign n1583 = ~pi318 & n1582;
  assign n1584 = pi129 & n1582;
  assign n1585 = pi318 & ~n1582;
  assign n1586 = ~pi129 & n1585;
  assign n1587 = ~n1584 & ~n1586;
  assign n1588 = pi128 & ~n1587;
  assign n1589 = ~n1583 & ~n1588;
  assign n1590 = ~n1512 & ~n1589;
  assign n1591 = ~pi129 & n1582;
  assign n1592 = pi129 & n1585;
  assign n1593 = ~n1591 & ~n1592;
  assign n1594 = ~pi128 & ~n1593;
  assign n1595 = pi129 & ~n1582;
  assign n1596 = ~n1591 & ~n1595;
  assign n1597 = n1512 & ~n1596;
  assign n1598 = ~n1594 & ~n1597;
  assign n1599 = ~n1590 & n1598;
  assign n1600 = pi128 & pi317;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = pi317 & n1599;
  assign n1603 = pi128 & n1602;
  assign n1604 = ~n1601 & ~n1603;
  assign n1605 = ~pi261 & ~n1471;
  assign n1606 = ~n1470 & ~n1605;
  assign n1607 = pi324 & ~n1256;
  assign n1608 = ~n1256 & n1371;
  assign n1609 = pi323 & n1608;
  assign n1610 = ~n1371 & ~n1375;
  assign n1611 = n1442 & ~n1610;
  assign n1612 = pi322 & n1611;
  assign n1613 = ~n1609 & ~n1612;
  assign n1614 = ~n1607 & ~n1613;
  assign n1615 = n1607 & n1613;
  assign n1616 = ~n1614 & ~n1615;
  assign n1617 = pi323 & n1442;
  assign n1618 = ~n1391 & ~n1421;
  assign n1619 = n1391 & n1421;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~n1147 & ~n1237;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = ~n1391 & n1421;
  assign n1624 = n1391 & ~n1421;
  assign n1625 = ~n1623 & ~n1624;
  assign n1626 = ~pi130 & ~n1625;
  assign n1627 = pi258 & ~n1626;
  assign n1628 = pi259 & ~n1627;
  assign n1629 = ~n1622 & ~n1628;
  assign n1630 = pi131 & ~n1629;
  assign n1631 = pi258 & pi261;
  assign n1632 = ~pi260 & ~n1631;
  assign n1633 = pi259 & ~n1632;
  assign n1634 = ~n1376 & ~n1633;
  assign n1635 = pi129 & ~n1634;
  assign n1636 = pi128 & n1635;
  assign n1637 = pi129 & pi261;
  assign n1638 = pi262 & ~n1637;
  assign n1639 = pi128 & n1638;
  assign n1640 = pi128 & pi262;
  assign n1641 = pi261 & ~n1640;
  assign n1642 = pi129 & n1641;
  assign n1643 = ~n1639 & ~n1642;
  assign n1644 = ~n1636 & n1643;
  assign n1645 = n1636 & ~n1643;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = pi130 & pi260;
  assign n1648 = n1237 & ~n1391;
  assign n1649 = ~n1237 & n1391;
  assign n1650 = n1421 & ~n1649;
  assign n1651 = ~n1648 & ~n1650;
  assign n1652 = n1647 & ~n1651;
  assign n1653 = ~n1421 & ~n1648;
  assign n1654 = ~n1649 & ~n1653;
  assign n1655 = ~n1647 & ~n1654;
  assign n1656 = ~n1652 & ~n1655;
  assign n1657 = ~n1646 & ~n1656;
  assign n1658 = ~n1636 & ~n1643;
  assign n1659 = n1636 & n1643;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n1647 & ~n1651;
  assign n1662 = n1647 & ~n1654;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~n1660 & ~n1663;
  assign n1665 = ~n1657 & ~n1664;
  assign n1666 = ~n1630 & ~n1665;
  assign n1667 = n1630 & n1665;
  assign n1668 = ~n1666 & ~n1667;
  assign n1669 = n1237 & n1427;
  assign n1670 = ~n1237 & ~n1427;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = ~n1620 & ~n1671;
  assign n1673 = pi258 & ~n1237;
  assign n1674 = pi131 & n1673;
  assign n1675 = pi259 & ~n1427;
  assign n1676 = pi130 & n1675;
  assign n1677 = ~n1674 & ~n1676;
  assign n1678 = ~n1625 & ~n1677;
  assign n1679 = ~n1672 & ~n1678;
  assign n1680 = ~pi258 & pi260;
  assign n1681 = pi128 & n1680;
  assign n1682 = ~n1234 & ~n1681;
  assign n1683 = ~n1416 & ~n1682;
  assign n1684 = pi258 & ~n1244;
  assign n1685 = pi128 & n1684;
  assign n1686 = ~pi258 & ~pi260;
  assign n1687 = ~pi128 & ~n1233;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = pi259 & ~n1688;
  assign n1690 = pi129 & n1689;
  assign n1691 = ~n1685 & ~n1690;
  assign n1692 = ~n1683 & n1691;
  assign n1693 = pi129 & pi258;
  assign n1694 = pi259 & ~n1693;
  assign n1695 = pi128 & n1694;
  assign n1696 = pi128 & pi259;
  assign n1697 = pi258 & ~n1696;
  assign n1698 = pi129 & n1697;
  assign n1699 = ~n1695 & ~n1698;
  assign n1700 = n1156 & ~n1699;
  assign n1701 = n1692 & ~n1700;
  assign n1702 = pi132 & pi258;
  assign n1703 = ~n1701 & ~n1702;
  assign n1704 = n1701 & n1702;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1679 & ~n1705;
  assign n1707 = n1701 & ~n1702;
  assign n1708 = ~n1692 & ~n1699;
  assign n1709 = ~n1701 & n1702;
  assign n1710 = n1708 & n1709;
  assign n1711 = ~n1707 & ~n1710;
  assign n1712 = n1679 & ~n1711;
  assign n1713 = n1703 & ~n1708;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1706 & n1714;
  assign n1716 = ~n1668 & ~n1715;
  assign n1717 = ~n1630 & n1665;
  assign n1718 = n1630 & ~n1665;
  assign n1719 = ~n1717 & ~n1718;
  assign n1720 = ~n1707 & ~n1709;
  assign n1721 = ~n1679 & ~n1720;
  assign n1722 = ~n1708 & n1709;
  assign n1723 = n1703 & n1708;
  assign n1724 = ~n1704 & ~n1723;
  assign n1725 = n1679 & ~n1724;
  assign n1726 = ~n1722 & ~n1725;
  assign n1727 = ~n1721 & n1726;
  assign n1728 = ~n1719 & ~n1727;
  assign n1729 = ~n1716 & ~n1728;
  assign n1730 = pi322 & n1729;
  assign n1731 = ~n1617 & ~n1730;
  assign n1732 = n1442 & n1729;
  assign n1733 = n1445 & n1732;
  assign n1734 = ~n1731 & ~n1733;
  assign n1735 = ~n1616 & ~n1734;
  assign n1736 = ~n1607 & n1613;
  assign n1737 = n1607 & ~n1613;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = ~n1617 & n1729;
  assign n1740 = pi322 & n1739;
  assign n1741 = n1442 & ~n1730;
  assign n1742 = pi323 & n1741;
  assign n1743 = ~n1740 & ~n1742;
  assign n1744 = ~n1738 & ~n1743;
  assign n1745 = ~n1735 & ~n1744;
  assign n1746 = n1371 & n1442;
  assign n1747 = pi322 & n1746;
  assign n1748 = ~n1371 & ~n1443;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1375 & ~n1749;
  assign n1751 = n1371 & ~n1443;
  assign n1752 = ~n1371 & n1442;
  assign n1753 = pi322 & n1752;
  assign n1754 = ~n1751 & ~n1753;
  assign n1755 = ~n1256 & ~n1754;
  assign n1756 = pi323 & n1755;
  assign n1757 = ~n1750 & ~n1756;
  assign n1758 = n1368 & n1757;
  assign n1759 = ~n1368 & ~n1757;
  assign n1760 = ~n1154 & ~n1759;
  assign n1761 = pi324 & n1760;
  assign n1762 = ~n1758 & ~n1761;
  assign n1763 = n1745 & ~n1762;
  assign n1764 = ~n1745 & n1762;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~pi324 & ~n1154;
  assign n1767 = pi258 & ~n1766;
  assign n1768 = pi128 & n1767;
  assign n1769 = ~n1459 & n1768;
  assign n1770 = ~pi324 & n1459;
  assign n1771 = n1156 & ~n1770;
  assign n1772 = ~n1154 & ~n1771;
  assign n1773 = ~n1769 & ~n1772;
  assign n1774 = pi325 & ~n1773;
  assign n1775 = pi326 & n1156;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = pi326 & n1774;
  assign n1778 = n1156 & n1777;
  assign n1779 = ~n1776 & ~n1778;
  assign n1780 = ~n1765 & ~n1779;
  assign n1781 = ~n1745 & ~n1762;
  assign n1782 = n1745 & n1762;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = n1774 & ~n1775;
  assign n1785 = pi326 & ~n1774;
  assign n1786 = n1156 & n1785;
  assign n1787 = ~n1784 & ~n1786;
  assign n1788 = ~n1783 & ~n1787;
  assign n1789 = ~n1780 & ~n1788;
  assign n1790 = ~n1606 & ~n1789;
  assign n1791 = n1606 & n1789;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = pi262 & ~n1792;
  assign n1794 = ~n1606 & n1789;
  assign n1795 = n1606 & ~n1789;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = ~pi262 & ~n1796;
  assign n1798 = ~n1793 & ~n1797;
  assign n1799 = n1359 & ~n1494;
  assign n1800 = ~n1495 & ~n1799;
  assign n1801 = n1798 & ~n1800;
  assign n1802 = ~n1798 & n1800;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = ~n1604 & ~n1803;
  assign n1805 = n1798 & n1800;
  assign n1806 = ~n1798 & ~n1800;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = n1604 & ~n1807;
  assign n1809 = ~n1804 & ~n1808;
  assign n1810 = ~n831 & ~n1809;
  assign n1811 = ~n1505 & ~n1810;
  assign n1812 = pi161 & ~n1811;
  assign n1813 = pi068 & ~pi161;
  assign n1814 = ~n1812 & ~n1813;
  assign po197 = ~pi160 & ~n1814;
  assign n1816 = pi263 & n831;
  assign n1817 = ~pi132 & pi133;
  assign n1818 = pi128 & pi131;
  assign n1819 = n1817 & n1818;
  assign n1820 = pi132 & ~pi133;
  assign n1821 = pi130 & n1820;
  assign n1822 = ~n1819 & ~n1821;
  assign n1823 = pi129 & ~n1822;
  assign n1824 = pi132 & pi133;
  assign n1825 = ~pi131 & n1824;
  assign n1826 = ~pi132 & ~pi133;
  assign n1827 = ~pi130 & n1826;
  assign n1828 = ~n1825 & ~n1827;
  assign n1829 = ~pi129 & ~n1828;
  assign n1830 = ~pi128 & n1826;
  assign n1831 = ~n1825 & ~n1830;
  assign n1832 = ~pi130 & ~n1831;
  assign n1833 = pi130 & n1817;
  assign n1834 = ~n1820 & ~n1833;
  assign n1835 = pi131 & ~n1834;
  assign n1836 = ~pi131 & n1826;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1832 & n1837;
  assign n1839 = ~n1829 & n1838;
  assign n1840 = ~n1823 & n1839;
  assign n1841 = n1533 & n1542;
  assign n1842 = ~pi320 & ~n1841;
  assign n1843 = ~n1533 & ~n1553;
  assign n1844 = pi320 & n1841;
  assign n1845 = ~n1556 & ~n1844;
  assign n1846 = ~n1843 & n1845;
  assign n1847 = ~n1842 & n1846;
  assign n1848 = n1840 & ~n1847;
  assign n1849 = n1542 & ~n1840;
  assign n1850 = ~pi320 & n1533;
  assign n1851 = n1849 & n1850;
  assign n1852 = ~n1848 & ~n1851;
  assign n1853 = pi321 & ~n1852;
  assign n1854 = ~n1542 & ~n1840;
  assign n1855 = ~n1553 & n1854;
  assign n1856 = ~pi321 & ~n1561;
  assign n1857 = ~n1855 & ~n1856;
  assign n1858 = n1533 & ~n1857;
  assign n1859 = pi321 & n1840;
  assign n1860 = n1542 & ~n1859;
  assign n1861 = ~n1533 & n1860;
  assign n1862 = n1553 & n1861;
  assign n1863 = ~n1858 & ~n1862;
  assign n1864 = pi320 & ~n1863;
  assign n1865 = ~n1853 & ~n1864;
  assign n1866 = n1515 & ~n1579;
  assign n1867 = pi319 & n1866;
  assign n1868 = ~n1578 & ~n1867;
  assign n1869 = ~n1865 & ~n1868;
  assign n1870 = n1865 & n1868;
  assign n1871 = ~n1869 & ~n1870;
  assign n1872 = n1553 & ~n1871;
  assign n1873 = pi319 & n1872;
  assign n1874 = pi319 & n1553;
  assign n1875 = n1865 & ~n1868;
  assign n1876 = ~n1865 & n1868;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = ~n1874 & ~n1877;
  assign n1879 = ~n1873 & ~n1878;
  assign n1880 = pi318 & n1582;
  assign n1881 = pi128 & n1880;
  assign n1882 = ~n1512 & ~n1881;
  assign n1883 = ~pi129 & ~n1882;
  assign n1884 = pi129 & pi318;
  assign n1885 = ~pi128 & n1884;
  assign n1886 = ~n1512 & ~n1885;
  assign n1887 = n1582 & ~n1886;
  assign n1888 = ~n1883 & ~n1887;
  assign n1889 = ~n1879 & n1888;
  assign n1890 = n1879 & ~n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = n1515 & ~n1891;
  assign n1893 = pi318 & n1892;
  assign n1894 = pi318 & n1515;
  assign n1895 = n1879 & n1888;
  assign n1896 = ~n1879 & ~n1888;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~n1894 & ~n1897;
  assign n1899 = ~n1893 & ~n1898;
  assign n1900 = pi129 & n1899;
  assign n1901 = pi317 & ~n1899;
  assign n1902 = ~pi129 & n1901;
  assign n1903 = ~n1900 & ~n1902;
  assign n1904 = n1599 & ~n1903;
  assign n1905 = pi128 & n1904;
  assign n1906 = ~pi317 & n1899;
  assign n1907 = pi128 & n1599;
  assign n1908 = ~pi129 & n1899;
  assign n1909 = pi129 & n1901;
  assign n1910 = ~n1908 & ~n1909;
  assign n1911 = ~n1907 & ~n1910;
  assign n1912 = ~n1906 & ~n1911;
  assign n1913 = ~n1905 & n1912;
  assign n1914 = pi128 & pi316;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = pi316 & n1913;
  assign n1917 = pi128 & n1916;
  assign n1918 = ~n1915 & ~n1917;
  assign n1919 = ~pi262 & ~n1791;
  assign n1920 = ~n1790 & ~n1919;
  assign n1921 = n1607 & ~n1762;
  assign n1922 = ~n1613 & ~n1730;
  assign n1923 = n1613 & n1729;
  assign n1924 = pi322 & n1923;
  assign n1925 = ~n1922 & ~n1924;
  assign n1926 = ~n1617 & ~n1925;
  assign n1927 = n1613 & ~n1730;
  assign n1928 = ~n1613 & n1729;
  assign n1929 = pi322 & n1928;
  assign n1930 = ~n1927 & ~n1929;
  assign n1931 = n1442 & ~n1930;
  assign n1932 = pi323 & n1931;
  assign n1933 = ~n1926 & ~n1932;
  assign n1934 = ~n1607 & n1762;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = ~n1921 & ~n1935;
  assign n1937 = ~n1154 & n1464;
  assign n1938 = n1156 & n1937;
  assign n1939 = n1156 & n1464;
  assign n1940 = n1154 & ~n1939;
  assign n1941 = ~n1765 & ~n1940;
  assign n1942 = ~n1938 & ~n1941;
  assign n1943 = pi325 & ~n1942;
  assign n1944 = n1936 & ~n1943;
  assign n1945 = ~n1936 & n1943;
  assign n1946 = ~n1944 & ~n1945;
  assign n1947 = n1774 & ~n1783;
  assign n1948 = ~n1765 & ~n1774;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = pi258 & ~n1949;
  assign n1951 = pi128 & n1950;
  assign n1952 = pi326 & n1951;
  assign n1953 = pi324 & n1442;
  assign n1954 = n1442 & ~n1613;
  assign n1955 = pi323 & n1954;
  assign n1956 = n1613 & ~n1617;
  assign n1957 = n1729 & ~n1956;
  assign n1958 = pi322 & n1957;
  assign n1959 = ~n1955 & ~n1958;
  assign n1960 = ~n1953 & ~n1959;
  assign n1961 = n1953 & n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = pi323 & n1729;
  assign n1964 = pi132 & pi259;
  assign n1965 = n1636 & n1640;
  assign n1966 = pi129 & pi262;
  assign n1967 = pi263 & ~n1966;
  assign n1968 = pi128 & n1967;
  assign n1969 = pi128 & pi263;
  assign n1970 = pi262 & ~n1969;
  assign n1971 = pi129 & n1970;
  assign n1972 = ~n1968 & ~n1971;
  assign n1973 = ~pi261 & ~n1972;
  assign n1974 = ~pi130 & ~n1972;
  assign n1975 = pi261 & n1972;
  assign n1976 = pi130 & n1975;
  assign n1977 = ~n1974 & ~n1976;
  assign n1978 = ~pi129 & ~n1977;
  assign n1979 = ~n1973 & ~n1978;
  assign n1980 = ~n1965 & ~n1979;
  assign n1981 = ~n1636 & n1640;
  assign n1982 = n1636 & ~n1640;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = pi129 & ~n1983;
  assign n1985 = pi261 & n1965;
  assign n1986 = ~n1984 & ~n1985;
  assign n1987 = ~n1972 & ~n1986;
  assign n1988 = pi261 & ~n1636;
  assign n1989 = ~n1640 & n1972;
  assign n1990 = n1988 & n1989;
  assign n1991 = ~n1987 & ~n1990;
  assign n1992 = pi130 & ~n1991;
  assign n1993 = ~n1640 & ~n1972;
  assign n1994 = ~n1636 & n1993;
  assign n1995 = ~n1636 & ~n1640;
  assign n1996 = pi261 & ~n1995;
  assign n1997 = pi129 & n1996;
  assign n1998 = ~n1965 & ~n1997;
  assign n1999 = n1972 & ~n1998;
  assign n2000 = ~n1994 & ~n1999;
  assign n2001 = ~pi130 & ~n2000;
  assign n2002 = n1640 & n1972;
  assign n2003 = ~pi261 & n1636;
  assign n2004 = n2002 & n2003;
  assign n2005 = ~n2001 & ~n2004;
  assign n2006 = ~n1992 & n2005;
  assign n2007 = ~n1980 & n2006;
  assign n2008 = n1647 & ~n1660;
  assign n2009 = ~n1647 & n1660;
  assign n2010 = ~n1651 & ~n2009;
  assign n2011 = ~n2008 & ~n2010;
  assign n2012 = n2007 & n2011;
  assign n2013 = ~n2007 & ~n2011;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = pi258 & ~n1620;
  assign n2016 = ~pi259 & ~n2015;
  assign n2017 = pi131 & ~n2016;
  assign n2018 = pi131 & pi260;
  assign n2019 = pi130 & ~n1625;
  assign n2020 = ~pi130 & ~n1620;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = pi259 & ~n2021;
  assign n2023 = pi258 & n2022;
  assign n2024 = pi131 & n2023;
  assign n2025 = ~n1665 & ~n2024;
  assign n2026 = ~n2018 & ~n2025;
  assign n2027 = n2017 & n2026;
  assign n2028 = n2017 & ~n2025;
  assign n2029 = n2018 & ~n2028;
  assign n2030 = ~n2027 & ~n2029;
  assign n2031 = ~n2014 & ~n2030;
  assign n2032 = n2007 & ~n2011;
  assign n2033 = ~n2007 & n2011;
  assign n2034 = ~n2032 & ~n2033;
  assign n2035 = n2018 & ~n2025;
  assign n2036 = n2017 & n2035;
  assign n2037 = ~n2018 & ~n2028;
  assign n2038 = ~n2036 & ~n2037;
  assign n2039 = ~n2034 & ~n2038;
  assign n2040 = ~n2031 & ~n2039;
  assign n2041 = ~n1964 & ~n2040;
  assign n2042 = n1964 & n2040;
  assign n2043 = ~n2041 & ~n2042;
  assign n2044 = n1679 & ~n1708;
  assign n2045 = ~n1679 & ~n1701;
  assign n2046 = n1702 & ~n1719;
  assign n2047 = ~n1668 & ~n1702;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~n2045 & ~n2048;
  assign n2050 = ~n2044 & ~n2049;
  assign n2051 = pi133 & pi258;
  assign n2052 = n2050 & ~n2051;
  assign n2053 = ~n2050 & n2051;
  assign n2054 = ~n2052 & ~n2053;
  assign n2055 = n2017 & ~n2024;
  assign n2056 = ~n1665 & n2055;
  assign n2057 = n1665 & ~n2055;
  assign n2058 = ~n2056 & ~n2057;
  assign n2059 = pi258 & ~n2058;
  assign n2060 = pi132 & n2059;
  assign n2061 = n1665 & ~n1702;
  assign n2062 = ~n1665 & n1702;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2055 & ~n2063;
  assign n2065 = n1665 & n1702;
  assign n2066 = ~n1665 & ~n1702;
  assign n2067 = ~n2065 & ~n2066;
  assign n2068 = ~n2024 & ~n2067;
  assign n2069 = n2017 & n2068;
  assign n2070 = ~n2064 & ~n2069;
  assign n2071 = n2060 & ~n2070;
  assign n2072 = ~n2060 & n2070;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2054 & ~n2073;
  assign n2075 = ~n2050 & ~n2051;
  assign n2076 = n2050 & n2051;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = ~n2060 & ~n2070;
  assign n2079 = n2060 & n2070;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n2077 & ~n2080;
  assign n2082 = ~n2074 & ~n2081;
  assign n2083 = ~n2043 & ~n2082;
  assign n2084 = ~n1964 & n2040;
  assign n2085 = n1964 & ~n2040;
  assign n2086 = ~n2084 & ~n2085;
  assign n2087 = ~n2073 & ~n2077;
  assign n2088 = ~n2054 & ~n2080;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = ~n2086 & ~n2089;
  assign n2091 = ~n2083 & ~n2090;
  assign n2092 = pi322 & n2091;
  assign n2093 = ~n1963 & ~n2092;
  assign n2094 = n1729 & n2091;
  assign n2095 = n1445 & n2094;
  assign n2096 = ~n2093 & ~n2095;
  assign n2097 = ~n1962 & ~n2096;
  assign n2098 = ~n1953 & n1959;
  assign n2099 = n1953 & ~n1959;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = ~n1963 & n2091;
  assign n2102 = pi322 & n2101;
  assign n2103 = n1729 & ~n2092;
  assign n2104 = pi323 & n2103;
  assign n2105 = ~n2102 & ~n2104;
  assign n2106 = ~n2100 & ~n2105;
  assign n2107 = ~n2097 & ~n2106;
  assign n2108 = n1952 & ~n2107;
  assign n2109 = ~n1952 & n2107;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n1256 & ~n2110;
  assign n2112 = pi325 & n2111;
  assign n2113 = pi325 & ~n1256;
  assign n2114 = ~n1952 & ~n2107;
  assign n2115 = n1952 & n2107;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = ~n2113 & ~n2116;
  assign n2118 = ~n2112 & ~n2117;
  assign n2119 = ~n1946 & ~n2118;
  assign n2120 = ~n1936 & ~n1943;
  assign n2121 = n1936 & n1943;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = ~n1256 & ~n2116;
  assign n2124 = pi325 & n2123;
  assign n2125 = ~n2110 & ~n2113;
  assign n2126 = ~n2124 & ~n2125;
  assign n2127 = ~n2122 & ~n2126;
  assign n2128 = ~n2119 & ~n2127;
  assign n2129 = pi326 & ~n1154;
  assign n2130 = ~n2128 & n2129;
  assign n2131 = n2128 & ~n2129;
  assign n2132 = ~n2130 & ~n2131;
  assign n2133 = pi327 & n1156;
  assign n2134 = n2132 & ~n2133;
  assign n2135 = pi327 & ~n2132;
  assign n2136 = n1156 & n2135;
  assign n2137 = ~n2134 & ~n2136;
  assign n2138 = ~n1920 & ~n2137;
  assign n2139 = n1920 & n2137;
  assign n2140 = ~n2138 & ~n2139;
  assign n2141 = pi263 & ~n2140;
  assign n2142 = ~n1920 & n2137;
  assign n2143 = n1920 & ~n2137;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~pi263 & ~n2144;
  assign n2146 = ~n2141 & ~n2145;
  assign n2147 = n1604 & ~n1805;
  assign n2148 = ~n1806 & ~n2147;
  assign n2149 = n2146 & ~n2148;
  assign n2150 = ~n2146 & n2148;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n1918 & ~n2151;
  assign n2153 = n2146 & n2148;
  assign n2154 = ~n2146 & ~n2148;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = n1918 & ~n2155;
  assign n2157 = ~n2152 & ~n2156;
  assign n2158 = ~n831 & ~n2157;
  assign n2159 = ~n1816 & ~n2158;
  assign n2160 = pi161 & ~n2159;
  assign n2161 = pi069 & ~pi161;
  assign n2162 = ~n2160 & ~n2161;
  assign po198 = ~pi160 & ~n2162;
  assign n2164 = pi264 & n831;
  assign n2165 = pi130 & pi133;
  assign n2166 = ~pi132 & ~n2165;
  assign n2167 = pi131 & ~n2166;
  assign n2168 = ~n1824 & ~n2167;
  assign n2169 = pi130 & pi132;
  assign n2170 = pi131 & pi133;
  assign n2171 = pi128 & n2170;
  assign n2172 = ~n2169 & ~n2171;
  assign n2173 = pi129 & ~n2172;
  assign n2174 = n2168 & ~n2173;
  assign n2175 = pi134 & n2174;
  assign n2176 = ~pi134 & ~n2174;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = pi133 & ~n2177;
  assign n2179 = pi134 & ~n2174;
  assign n2180 = ~pi134 & n2174;
  assign n2181 = ~n2179 & ~n2180;
  assign n2182 = ~pi133 & ~n2181;
  assign n2183 = ~n2178 & ~n2182;
  assign n2184 = pi321 & n2183;
  assign n2185 = n1542 & n1840;
  assign n2186 = ~n1533 & ~n2185;
  assign n2187 = n1553 & ~n2186;
  assign n2188 = n1533 & ~n1854;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = pi321 & ~n2189;
  assign n2191 = n1553 & n1841;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = pi320 & ~n2192;
  assign n2194 = n1534 & n2185;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = pi320 & n1840;
  assign n2197 = ~n2195 & ~n2196;
  assign n2198 = n1840 & n2195;
  assign n2199 = pi320 & n2198;
  assign n2200 = ~n2197 & ~n2199;
  assign n2201 = ~n2184 & ~n2200;
  assign n2202 = n2195 & ~n2196;
  assign n2203 = n1840 & ~n2195;
  assign n2204 = pi320 & n2203;
  assign n2205 = ~n2202 & ~n2204;
  assign n2206 = n2183 & ~n2205;
  assign n2207 = pi321 & n2206;
  assign n2208 = ~n2201 & ~n2207;
  assign n2209 = n1553 & ~n1870;
  assign n2210 = pi319 & n2209;
  assign n2211 = ~n1869 & ~n2210;
  assign n2212 = ~n2208 & ~n2211;
  assign n2213 = n2208 & n2211;
  assign n2214 = ~n2212 & ~n2213;
  assign n2215 = n1533 & ~n2214;
  assign n2216 = pi319 & n2215;
  assign n2217 = pi319 & n1533;
  assign n2218 = n2208 & ~n2211;
  assign n2219 = ~n2208 & n2211;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~n2217 & ~n2220;
  assign n2222 = ~n2216 & ~n2221;
  assign n2223 = n1515 & ~n1895;
  assign n2224 = pi318 & n2223;
  assign n2225 = ~n1896 & ~n2224;
  assign n2226 = n2222 & n2225;
  assign n2227 = ~n2222 & ~n2225;
  assign n2228 = ~n2226 & ~n2227;
  assign n2229 = n1553 & ~n2228;
  assign n2230 = pi318 & n2229;
  assign n2231 = pi318 & n1553;
  assign n2232 = ~n2222 & n2225;
  assign n2233 = n2222 & ~n2225;
  assign n2234 = ~n2232 & ~n2233;
  assign n2235 = ~n2231 & ~n2234;
  assign n2236 = ~n2230 & ~n2235;
  assign n2237 = n1599 & ~n1899;
  assign n2238 = ~pi129 & ~n2237;
  assign n2239 = pi128 & n2238;
  assign n2240 = n1899 & ~n1907;
  assign n2241 = pi129 & n2240;
  assign n2242 = ~n2239 & ~n2241;
  assign n2243 = pi317 & ~n2242;
  assign n2244 = ~n2236 & n2243;
  assign n2245 = n2236 & ~n2243;
  assign n2246 = ~n2244 & ~n2245;
  assign n2247 = n1515 & ~n2246;
  assign n2248 = pi317 & n2247;
  assign n2249 = pi317 & n1515;
  assign n2250 = n2236 & n2243;
  assign n2251 = ~n2236 & ~n2243;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = ~n2249 & ~n2252;
  assign n2254 = ~n2248 & ~n2253;
  assign n2255 = pi129 & n2254;
  assign n2256 = pi316 & ~n2254;
  assign n2257 = ~pi129 & n2256;
  assign n2258 = ~n2255 & ~n2257;
  assign n2259 = n1913 & ~n2258;
  assign n2260 = pi128 & n2259;
  assign n2261 = ~pi316 & n2254;
  assign n2262 = pi128 & n1913;
  assign n2263 = ~pi129 & n2254;
  assign n2264 = pi129 & n2256;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = ~n2262 & ~n2265;
  assign n2267 = ~n2261 & ~n2266;
  assign n2268 = ~n2260 & n2267;
  assign n2269 = pi315 & ~n2268;
  assign n2270 = pi128 & n2269;
  assign n2271 = pi128 & pi315;
  assign n2272 = n2268 & ~n2271;
  assign n2273 = ~n2270 & ~n2272;
  assign n2274 = ~pi263 & ~n2139;
  assign n2275 = ~n2138 & ~n2274;
  assign n2276 = ~pi326 & ~n1154;
  assign n2277 = pi258 & ~n2276;
  assign n2278 = pi128 & n2277;
  assign n2279 = ~n2128 & n2278;
  assign n2280 = ~pi326 & n2128;
  assign n2281 = n1156 & ~n2280;
  assign n2282 = ~n1154 & ~n2281;
  assign n2283 = ~n2279 & ~n2282;
  assign n2284 = pi327 & ~n2283;
  assign n2285 = n1943 & n2113;
  assign n2286 = n1936 & ~n2107;
  assign n2287 = ~n1936 & n2107;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n1943 & ~n2113;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = ~n2285 & ~n2290;
  assign n2292 = n2107 & ~n2113;
  assign n2293 = ~n2107 & n2113;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n1952 & ~n2129;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = ~n2122 & n2296;
  assign n2298 = n1952 & n2129;
  assign n2299 = n2107 & n2113;
  assign n2300 = ~n2107 & ~n2113;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2295 & ~n2301;
  assign n2303 = ~n1946 & n2302;
  assign n2304 = ~n2298 & ~n2303;
  assign n2305 = ~n2297 & n2304;
  assign n2306 = n2291 & ~n2305;
  assign n2307 = ~n2291 & n2305;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = pi324 & n1729;
  assign n2310 = n1729 & ~n1959;
  assign n2311 = pi323 & n2310;
  assign n2312 = n1959 & ~n1963;
  assign n2313 = n2091 & ~n2312;
  assign n2314 = pi322 & n2313;
  assign n2315 = ~n2311 & ~n2314;
  assign n2316 = ~n2309 & ~n2315;
  assign n2317 = n2309 & n2315;
  assign n2318 = ~n2316 & ~n2317;
  assign n2319 = pi323 & n2091;
  assign n2320 = ~n2040 & ~n2060;
  assign n2321 = n2040 & n2060;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = ~n1147 & ~n1964;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2040 & n2060;
  assign n2326 = n2040 & ~n2060;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = ~pi132 & ~n2327;
  assign n2329 = pi258 & ~n2328;
  assign n2330 = pi259 & ~n2329;
  assign n2331 = ~n2324 & ~n2330;
  assign n2332 = pi133 & ~n2331;
  assign n2333 = pi130 & pi262;
  assign n2334 = pi129 & pi263;
  assign n2335 = pi264 & ~n2334;
  assign n2336 = pi128 & n2335;
  assign n2337 = pi128 & pi264;
  assign n2338 = pi263 & ~n2337;
  assign n2339 = pi129 & n2338;
  assign n2340 = ~n2336 & ~n2339;
  assign n2341 = n1966 & n1969;
  assign n2342 = ~n1966 & ~n1969;
  assign n2343 = n1637 & n1640;
  assign n2344 = ~n1637 & ~n1640;
  assign n2345 = n1636 & ~n2344;
  assign n2346 = ~n2343 & ~n2345;
  assign n2347 = ~n2342 & ~n2346;
  assign n2348 = ~n2341 & ~n2347;
  assign n2349 = ~n2340 & ~n2348;
  assign n2350 = ~n1636 & ~n2343;
  assign n2351 = ~n2344 & ~n2350;
  assign n2352 = ~n2341 & ~n2351;
  assign n2353 = ~n2342 & ~n2352;
  assign n2354 = n2340 & ~n2353;
  assign n2355 = ~n2349 & ~n2354;
  assign n2356 = ~n2333 & n2355;
  assign n2357 = n2333 & ~n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n1972 & ~n1998;
  assign n2360 = ~pi129 & ~n1965;
  assign n2361 = ~n1995 & ~n2360;
  assign n2362 = n1972 & ~n2361;
  assign n2363 = ~n2359 & ~n2362;
  assign n2364 = ~pi130 & ~n2363;
  assign n2365 = ~n1965 & n1972;
  assign n2366 = n1640 & ~n1972;
  assign n2367 = n1636 & n2366;
  assign n2368 = ~n2365 & ~n2367;
  assign n2369 = ~pi261 & ~n2368;
  assign n2370 = ~n2364 & ~n2369;
  assign n2371 = pi131 & pi261;
  assign n2372 = pi129 & ~n1995;
  assign n2373 = ~n1965 & ~n2372;
  assign n2374 = n1972 & ~n2373;
  assign n2375 = ~n1972 & ~n2361;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = pi261 & ~n2376;
  assign n2378 = pi130 & n2377;
  assign n2379 = n2011 & ~n2378;
  assign n2380 = n2371 & ~n2379;
  assign n2381 = n2370 & n2380;
  assign n2382 = n2370 & ~n2379;
  assign n2383 = ~n2371 & ~n2382;
  assign n2384 = ~n2381 & ~n2383;
  assign n2385 = ~n2358 & ~n2384;
  assign n2386 = ~n2333 & ~n2355;
  assign n2387 = n2333 & n2355;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = ~n2371 & ~n2379;
  assign n2390 = n2370 & n2389;
  assign n2391 = n2371 & ~n2382;
  assign n2392 = ~n2390 & ~n2391;
  assign n2393 = ~n2388 & ~n2392;
  assign n2394 = ~n2385 & ~n2393;
  assign n2395 = ~n2014 & ~n2018;
  assign n2396 = n2014 & n2018;
  assign n2397 = ~n2028 & ~n2396;
  assign n2398 = ~n2395 & ~n2397;
  assign n2399 = n2394 & ~n2398;
  assign n2400 = ~n2394 & n2398;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = pi132 & pi260;
  assign n2403 = n2060 & ~n2084;
  assign n2404 = ~n2085 & ~n2403;
  assign n2405 = n2402 & ~n2404;
  assign n2406 = ~n2060 & ~n2085;
  assign n2407 = ~n2084 & ~n2406;
  assign n2408 = ~n2402 & ~n2407;
  assign n2409 = ~n2405 & ~n2408;
  assign n2410 = ~n2401 & ~n2409;
  assign n2411 = n2394 & n2398;
  assign n2412 = ~n2394 & ~n2398;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2402 & ~n2404;
  assign n2415 = n2402 & ~n2407;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = ~n2413 & ~n2416;
  assign n2418 = ~n2410 & ~n2417;
  assign n2419 = ~n2332 & ~n2418;
  assign n2420 = n2332 & n2418;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = ~n1964 & ~n2051;
  assign n2423 = n1964 & n2051;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2322 & ~n2424;
  assign n2426 = pi258 & ~n1964;
  assign n2427 = pi133 & n2426;
  assign n2428 = pi259 & ~n2051;
  assign n2429 = pi132 & n2428;
  assign n2430 = ~n2427 & ~n2429;
  assign n2431 = ~n2327 & ~n2430;
  assign n2432 = ~n2425 & ~n2431;
  assign n2433 = pi134 & pi258;
  assign n2434 = ~n2432 & ~n2433;
  assign n2435 = n2432 & n2433;
  assign n2436 = n2050 & n2435;
  assign n2437 = ~n2434 & ~n2436;
  assign n2438 = ~n2070 & ~n2437;
  assign n2439 = n2432 & ~n2433;
  assign n2440 = ~n2432 & n2433;
  assign n2441 = ~n2050 & n2440;
  assign n2442 = ~n2439 & ~n2441;
  assign n2443 = n2070 & ~n2442;
  assign n2444 = ~n2050 & n2432;
  assign n2445 = n2050 & ~n2432;
  assign n2446 = ~n2444 & ~n2445;
  assign n2447 = ~n2433 & ~n2446;
  assign n2448 = ~n2443 & ~n2447;
  assign n2449 = ~n2438 & n2448;
  assign n2450 = ~n2421 & ~n2449;
  assign n2451 = ~n2332 & n2418;
  assign n2452 = n2332 & ~n2418;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = n2050 & n2439;
  assign n2455 = ~n2440 & ~n2454;
  assign n2456 = ~n2070 & ~n2455;
  assign n2457 = ~n2050 & n2434;
  assign n2458 = ~n2435 & ~n2457;
  assign n2459 = n2070 & ~n2458;
  assign n2460 = n2433 & ~n2446;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = ~n2456 & n2461;
  assign n2463 = ~n2453 & ~n2462;
  assign n2464 = ~n2450 & ~n2463;
  assign n2465 = pi322 & n2464;
  assign n2466 = ~n2319 & ~n2465;
  assign n2467 = n2091 & n2464;
  assign n2468 = n1445 & n2467;
  assign n2469 = ~n2466 & ~n2468;
  assign n2470 = ~n2318 & ~n2469;
  assign n2471 = ~n2309 & n2315;
  assign n2472 = n2309 & ~n2315;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = ~n2319 & n2464;
  assign n2475 = pi322 & n2474;
  assign n2476 = n2091 & ~n2465;
  assign n2477 = pi323 & n2476;
  assign n2478 = ~n2475 & ~n2477;
  assign n2479 = ~n2473 & ~n2478;
  assign n2480 = ~n2470 & ~n2479;
  assign n2481 = ~n1936 & n1953;
  assign n2482 = ~n1959 & ~n2092;
  assign n2483 = n1959 & n2091;
  assign n2484 = pi322 & n2483;
  assign n2485 = ~n2482 & ~n2484;
  assign n2486 = ~n1963 & ~n2485;
  assign n2487 = n1959 & ~n2092;
  assign n2488 = ~n1959 & n2091;
  assign n2489 = pi322 & n2488;
  assign n2490 = ~n2487 & ~n2489;
  assign n2491 = n1729 & ~n2490;
  assign n2492 = pi323 & n2491;
  assign n2493 = ~n2486 & ~n2492;
  assign n2494 = n1936 & ~n1953;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = ~n2481 & ~n2495;
  assign n2497 = n2480 & ~n2496;
  assign n2498 = ~n2480 & n2496;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = pi326 & ~n1256;
  assign n2501 = pi325 & n1442;
  assign n2502 = n2500 & n2501;
  assign n2503 = ~n2500 & ~n2501;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2499 & ~n2504;
  assign n2506 = ~n2480 & ~n2496;
  assign n2507 = n2480 & n2496;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = ~n2500 & n2501;
  assign n2510 = n2500 & ~n2501;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = ~n2508 & ~n2511;
  assign n2513 = ~n2505 & ~n2512;
  assign n2514 = ~n2308 & ~n2513;
  assign n2515 = n2291 & n2305;
  assign n2516 = ~n2291 & ~n2305;
  assign n2517 = ~n2515 & ~n2516;
  assign n2518 = ~n2504 & ~n2508;
  assign n2519 = ~n2499 & ~n2511;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~n2517 & ~n2520;
  assign n2522 = ~n2514 & ~n2521;
  assign n2523 = n2284 & n2522;
  assign n2524 = ~n2284 & ~n2522;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = pi258 & ~n2525;
  assign n2527 = pi128 & n2526;
  assign n2528 = pi328 & n2527;
  assign n2529 = n2284 & ~n2522;
  assign n2530 = ~n2284 & n2522;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = pi328 & n1156;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = ~n2528 & ~n2533;
  assign n2535 = ~n2275 & ~n2534;
  assign n2536 = n2275 & n2534;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = pi264 & ~n2537;
  assign n2539 = ~n2275 & n2534;
  assign n2540 = n2275 & ~n2534;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~pi264 & ~n2541;
  assign n2543 = ~n2538 & ~n2542;
  assign n2544 = n1918 & ~n2153;
  assign n2545 = ~n2154 & ~n2544;
  assign n2546 = n2543 & ~n2545;
  assign n2547 = ~n2543 & n2545;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = ~n2273 & ~n2548;
  assign n2550 = n2543 & n2545;
  assign n2551 = ~n2543 & ~n2545;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = n2273 & ~n2552;
  assign n2554 = ~n2549 & ~n2553;
  assign n2555 = ~n831 & ~n2554;
  assign n2556 = ~n2164 & ~n2555;
  assign n2557 = pi161 & ~n2556;
  assign n2558 = pi070 & ~pi161;
  assign n2559 = ~n2557 & ~n2558;
  assign po199 = ~pi160 & ~n2559;
  assign n2561 = pi265 & n831;
  assign n2562 = ~pi135 & n2174;
  assign n2563 = pi135 & ~n2174;
  assign n2564 = ~pi134 & n2563;
  assign n2565 = ~n2562 & ~n2564;
  assign n2566 = pi133 & ~n2565;
  assign n2567 = ~pi135 & ~n2174;
  assign n2568 = pi135 & n2174;
  assign n2569 = pi134 & n2568;
  assign n2570 = ~n2567 & ~n2569;
  assign n2571 = ~pi133 & ~n2570;
  assign n2572 = ~pi135 & ~n2181;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = ~n2566 & n2573;
  assign n2575 = n2183 & ~n2195;
  assign n2576 = ~pi320 & ~n2575;
  assign n2577 = ~n1840 & ~n2183;
  assign n2578 = pi320 & n2575;
  assign n2579 = ~n2198 & ~n2578;
  assign n2580 = ~n2577 & n2579;
  assign n2581 = ~n2576 & n2580;
  assign n2582 = n2574 & ~n2581;
  assign n2583 = ~n2195 & ~n2574;
  assign n2584 = ~pi320 & n2183;
  assign n2585 = n2583 & n2584;
  assign n2586 = ~n2582 & ~n2585;
  assign n2587 = pi321 & ~n2586;
  assign n2588 = n2195 & ~n2574;
  assign n2589 = ~n1840 & n2588;
  assign n2590 = ~pi321 & ~n2203;
  assign n2591 = ~n2589 & ~n2590;
  assign n2592 = n2183 & ~n2591;
  assign n2593 = pi321 & n2574;
  assign n2594 = ~n2195 & ~n2593;
  assign n2595 = ~n2183 & n2594;
  assign n2596 = n1840 & n2595;
  assign n2597 = ~n2592 & ~n2596;
  assign n2598 = pi320 & ~n2597;
  assign n2599 = ~n2587 & ~n2598;
  assign n2600 = n1533 & ~n2213;
  assign n2601 = pi319 & n2600;
  assign n2602 = ~n2212 & ~n2601;
  assign n2603 = ~n2599 & ~n2602;
  assign n2604 = n2599 & n2602;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n1840 & ~n2605;
  assign n2607 = pi319 & n2606;
  assign n2608 = pi319 & n1840;
  assign n2609 = n2599 & ~n2602;
  assign n2610 = ~n2599 & n2602;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n2608 & ~n2611;
  assign n2613 = ~n2607 & ~n2612;
  assign n2614 = n1553 & ~n2226;
  assign n2615 = pi318 & n2614;
  assign n2616 = ~n2227 & ~n2615;
  assign n2617 = n2613 & n2616;
  assign n2618 = ~n2613 & ~n2616;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = n1533 & ~n2619;
  assign n2621 = pi318 & n2620;
  assign n2622 = pi318 & n1533;
  assign n2623 = ~n2613 & n2616;
  assign n2624 = n2613 & ~n2616;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = ~n2622 & ~n2625;
  assign n2627 = ~n2621 & ~n2626;
  assign n2628 = n1515 & ~n2245;
  assign n2629 = pi317 & n2628;
  assign n2630 = ~n2244 & ~n2629;
  assign n2631 = ~n2627 & ~n2630;
  assign n2632 = n2627 & n2630;
  assign n2633 = ~n2631 & ~n2632;
  assign n2634 = n1553 & ~n2633;
  assign n2635 = pi317 & n2634;
  assign n2636 = pi317 & n1553;
  assign n2637 = n2627 & ~n2630;
  assign n2638 = ~n2627 & n2630;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2636 & ~n2639;
  assign n2641 = ~n2635 & ~n2640;
  assign n2642 = ~n2254 & ~n2262;
  assign n2643 = pi129 & n2642;
  assign n2644 = n1913 & n2254;
  assign n2645 = ~pi129 & ~n2644;
  assign n2646 = pi128 & n2645;
  assign n2647 = ~n2643 & ~n2646;
  assign n2648 = pi316 & ~n2647;
  assign n2649 = ~n2641 & n2648;
  assign n2650 = n2641 & ~n2648;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = n1515 & ~n2651;
  assign n2653 = pi316 & n2652;
  assign n2654 = pi316 & n1515;
  assign n2655 = n2641 & n2648;
  assign n2656 = ~n2641 & ~n2648;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = ~n2654 & ~n2657;
  assign n2659 = ~n2653 & ~n2658;
  assign n2660 = pi129 & ~n2659;
  assign n2661 = pi315 & n2659;
  assign n2662 = ~pi129 & n2661;
  assign n2663 = ~n2660 & ~n2662;
  assign n2664 = ~n2268 & ~n2663;
  assign n2665 = pi128 & n2664;
  assign n2666 = ~pi315 & ~n2659;
  assign n2667 = ~pi129 & ~n2659;
  assign n2668 = pi129 & n2661;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = pi128 & ~n2268;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = ~n2666 & ~n2671;
  assign n2673 = ~n2665 & n2672;
  assign n2674 = pi128 & pi314;
  assign n2675 = ~n2673 & ~n2674;
  assign n2676 = pi314 & n2673;
  assign n2677 = pi128 & n2676;
  assign n2678 = ~n2675 & ~n2677;
  assign n2679 = ~pi264 & ~n2536;
  assign n2680 = ~n2535 & ~n2679;
  assign n2681 = pi328 & ~n1154;
  assign n2682 = ~n2291 & n2496;
  assign n2683 = n2291 & ~n2496;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = ~n2480 & n2501;
  assign n2686 = n2480 & ~n2501;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n2305 & ~n2500;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2684 & n2689;
  assign n2691 = ~n2305 & n2500;
  assign n2692 = ~n2291 & ~n2496;
  assign n2693 = n2291 & n2496;
  assign n2694 = ~n2692 & ~n2693;
  assign n2695 = n2480 & n2501;
  assign n2696 = ~n2480 & ~n2501;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = ~n2688 & ~n2697;
  assign n2699 = ~n2694 & n2698;
  assign n2700 = ~n2691 & ~n2699;
  assign n2701 = ~n2690 & n2700;
  assign n2702 = n1156 & n2132;
  assign n2703 = ~n2522 & ~n2702;
  assign n2704 = ~n1154 & ~n2703;
  assign n2705 = n2132 & n2522;
  assign n2706 = n1156 & n2705;
  assign n2707 = ~n2704 & ~n2706;
  assign n2708 = pi327 & ~n2707;
  assign n2709 = n2701 & n2708;
  assign n2710 = ~n2701 & ~n2708;
  assign n2711 = ~n2709 & ~n2710;
  assign n2712 = pi326 & n1442;
  assign n2713 = n2309 & ~n2496;
  assign n2714 = ~n2315 & ~n2465;
  assign n2715 = n2315 & n2464;
  assign n2716 = pi322 & n2715;
  assign n2717 = ~n2714 & ~n2716;
  assign n2718 = ~n2319 & ~n2717;
  assign n2719 = n2315 & ~n2465;
  assign n2720 = ~n2315 & n2464;
  assign n2721 = pi322 & n2720;
  assign n2722 = ~n2719 & ~n2721;
  assign n2723 = n2091 & ~n2722;
  assign n2724 = pi323 & n2723;
  assign n2725 = ~n2718 & ~n2724;
  assign n2726 = ~n2309 & n2496;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2713 & ~n2727;
  assign n2729 = ~n2291 & n2501;
  assign n2730 = n2291 & ~n2501;
  assign n2731 = ~n2499 & ~n2730;
  assign n2732 = ~n2729 & ~n2731;
  assign n2733 = ~n2728 & ~n2732;
  assign n2734 = n2728 & n2732;
  assign n2735 = ~n2733 & ~n2734;
  assign n2736 = pi324 & n2091;
  assign n2737 = pi323 & n2464;
  assign n2738 = n2091 & ~n2315;
  assign n2739 = pi323 & n2738;
  assign n2740 = n2315 & ~n2319;
  assign n2741 = n2464 & ~n2740;
  assign n2742 = pi322 & n2741;
  assign n2743 = ~n2739 & ~n2742;
  assign n2744 = pi130 & pi263;
  assign n2745 = pi128 & pi265;
  assign n2746 = pi264 & ~n2745;
  assign n2747 = pi129 & n2746;
  assign n2748 = pi129 & pi264;
  assign n2749 = pi265 & ~n2748;
  assign n2750 = pi128 & n2749;
  assign n2751 = ~n2747 & ~n2750;
  assign n2752 = ~n2334 & ~n2337;
  assign n2753 = pi263 & n1175;
  assign n2754 = pi264 & n2753;
  assign n2755 = ~n2353 & ~n2754;
  assign n2756 = ~n2752 & ~n2755;
  assign n2757 = ~n2751 & ~n2756;
  assign n2758 = n2751 & ~n2755;
  assign n2759 = ~n2752 & n2758;
  assign n2760 = ~n2757 & ~n2759;
  assign n2761 = ~n2744 & ~n2760;
  assign n2762 = n2751 & ~n2756;
  assign n2763 = ~n2751 & ~n2755;
  assign n2764 = ~n2752 & n2763;
  assign n2765 = ~n2762 & ~n2764;
  assign n2766 = pi263 & ~n2765;
  assign n2767 = pi130 & n2766;
  assign n2768 = ~n2761 & ~n2767;
  assign n2769 = ~n2379 & ~n2386;
  assign n2770 = n2370 & n2769;
  assign n2771 = ~n2387 & ~n2770;
  assign n2772 = n2768 & n2771;
  assign n2773 = ~n2768 & ~n2771;
  assign n2774 = ~n2772 & ~n2773;
  assign n2775 = pi131 & pi262;
  assign n2776 = n2355 & ~n2379;
  assign n2777 = n2370 & n2776;
  assign n2778 = ~n2355 & ~n2382;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = ~n2333 & ~n2779;
  assign n2781 = ~n2355 & ~n2379;
  assign n2782 = n2370 & n2781;
  assign n2783 = n2355 & ~n2382;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = pi262 & ~n2784;
  assign n2786 = pi130 & n2785;
  assign n2787 = ~n2780 & ~n2786;
  assign n2788 = n2398 & n2787;
  assign n2789 = ~n2398 & ~n2787;
  assign n2790 = n2371 & ~n2789;
  assign n2791 = ~n2788 & ~n2790;
  assign n2792 = n2775 & ~n2791;
  assign n2793 = ~n2371 & ~n2788;
  assign n2794 = ~n2789 & ~n2793;
  assign n2795 = ~n2775 & ~n2794;
  assign n2796 = ~n2792 & ~n2795;
  assign n2797 = ~n2774 & ~n2796;
  assign n2798 = n2768 & ~n2771;
  assign n2799 = ~n2768 & n2771;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = ~n2775 & ~n2791;
  assign n2802 = n2775 & ~n2794;
  assign n2803 = ~n2801 & ~n2802;
  assign n2804 = ~n2800 & ~n2803;
  assign n2805 = ~n2797 & ~n2804;
  assign n2806 = n2402 & ~n2413;
  assign n2807 = ~n2402 & n2413;
  assign n2808 = ~n2404 & ~n2807;
  assign n2809 = ~n2806 & ~n2808;
  assign n2810 = n2805 & n2809;
  assign n2811 = ~n2805 & ~n2809;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = pi133 & pi260;
  assign n2814 = pi132 & pi261;
  assign n2815 = n2813 & n2814;
  assign n2816 = ~n2813 & ~n2814;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n2812 & ~n2817;
  assign n2819 = ~n2805 & n2809;
  assign n2820 = n2805 & ~n2809;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = pi260 & ~n2814;
  assign n2823 = pi133 & n2822;
  assign n2824 = pi261 & ~n2813;
  assign n2825 = pi132 & n2824;
  assign n2826 = ~n2823 & ~n2825;
  assign n2827 = ~n2821 & ~n2826;
  assign n2828 = ~n2818 & ~n2827;
  assign n2829 = pi259 & n2418;
  assign n2830 = pi259 & ~n2322;
  assign n2831 = pi132 & n2830;
  assign n2832 = ~n1964 & ~n2327;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = ~pi259 & ~n2418;
  assign n2835 = n2833 & ~n2834;
  assign n2836 = pi258 & n2835;
  assign n2837 = ~n2829 & ~n2836;
  assign n2838 = pi133 & ~n2837;
  assign n2839 = n2828 & n2838;
  assign n2840 = ~n2828 & ~n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = pi135 & pi258;
  assign n2843 = pi134 & pi259;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = n2842 & n2843;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = pi258 & ~n2453;
  assign n2848 = pi134 & n2847;
  assign n2849 = pi258 & ~n2421;
  assign n2850 = pi134 & n2849;
  assign n2851 = ~n2433 & ~n2453;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n2848 & ~n2852;
  assign n2854 = ~n2848 & n2852;
  assign n2855 = ~n2853 & ~n2854;
  assign n2856 = ~n2846 & ~n2855;
  assign n2857 = n2842 & ~n2843;
  assign n2858 = ~n2842 & n2843;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = ~n2848 & ~n2852;
  assign n2861 = n2848 & n2852;
  assign n2862 = ~n2860 & ~n2861;
  assign n2863 = ~n2859 & ~n2862;
  assign n2864 = ~n2856 & ~n2863;
  assign n2865 = ~n2841 & ~n2864;
  assign n2866 = n2828 & ~n2838;
  assign n2867 = ~n2828 & n2838;
  assign n2868 = ~n2866 & ~n2867;
  assign n2869 = ~n2855 & ~n2859;
  assign n2870 = ~n2846 & ~n2862;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = ~n2868 & ~n2871;
  assign n2873 = ~n2865 & ~n2872;
  assign n2874 = ~n2050 & n2852;
  assign n2875 = ~n2432 & ~n2874;
  assign n2876 = n2050 & ~n2852;
  assign n2877 = n2432 & ~n2876;
  assign n2878 = ~n2070 & ~n2877;
  assign n2879 = ~n2875 & ~n2878;
  assign n2880 = n2873 & ~n2879;
  assign n2881 = ~n2873 & n2879;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = n2743 & ~n2882;
  assign n2884 = pi322 & n2883;
  assign n2885 = ~n2873 & ~n2879;
  assign n2886 = n2873 & n2879;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = pi322 & n2887;
  assign n2889 = ~n2743 & ~n2888;
  assign n2890 = ~n2884 & ~n2889;
  assign n2891 = ~n2737 & ~n2890;
  assign n2892 = ~n2743 & ~n2882;
  assign n2893 = pi322 & n2892;
  assign n2894 = n2743 & ~n2888;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = n2464 & ~n2895;
  assign n2897 = pi323 & n2896;
  assign n2898 = ~n2891 & ~n2897;
  assign n2899 = ~n2736 & n2898;
  assign n2900 = n2736 & ~n2898;
  assign n2901 = ~n2899 & ~n2900;
  assign n2902 = n1729 & ~n2901;
  assign n2903 = pi325 & n2902;
  assign n2904 = pi325 & n1729;
  assign n2905 = n2736 & n2898;
  assign n2906 = ~n2736 & ~n2898;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n2904 & ~n2907;
  assign n2909 = ~n2903 & ~n2908;
  assign n2910 = ~n2735 & ~n2909;
  assign n2911 = ~n2728 & n2732;
  assign n2912 = n2728 & ~n2732;
  assign n2913 = ~n2911 & ~n2912;
  assign n2914 = n1729 & ~n2907;
  assign n2915 = pi325 & n2914;
  assign n2916 = ~n2901 & ~n2904;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = ~n2913 & ~n2917;
  assign n2919 = ~n2910 & ~n2918;
  assign n2920 = ~n2712 & n2919;
  assign n2921 = n2712 & ~n2919;
  assign n2922 = ~n2920 & ~n2921;
  assign n2923 = pi258 & ~n2531;
  assign n2924 = pi128 & n2923;
  assign n2925 = pi328 & n2924;
  assign n2926 = pi327 & ~n1256;
  assign n2927 = n2925 & n2926;
  assign n2928 = ~n2925 & ~n2926;
  assign n2929 = ~n2927 & ~n2928;
  assign n2930 = ~n2922 & ~n2929;
  assign n2931 = n2712 & n2919;
  assign n2932 = ~n2712 & ~n2919;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = ~n2925 & n2926;
  assign n2935 = n2925 & ~n2926;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = ~n2933 & ~n2936;
  assign n2938 = ~n2930 & ~n2937;
  assign n2939 = ~n2711 & ~n2938;
  assign n2940 = n2701 & ~n2708;
  assign n2941 = ~n2701 & n2708;
  assign n2942 = ~n2940 & ~n2941;
  assign n2943 = ~n2929 & ~n2933;
  assign n2944 = ~n2922 & ~n2936;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = ~n2942 & ~n2945;
  assign n2947 = ~n2939 & ~n2946;
  assign n2948 = pi329 & n1156;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = pi329 & n2947;
  assign n2951 = n1156 & n2950;
  assign n2952 = ~n2949 & ~n2951;
  assign n2953 = ~n2681 & ~n2952;
  assign n2954 = n2947 & ~n2948;
  assign n2955 = pi329 & ~n2947;
  assign n2956 = n1156 & n2955;
  assign n2957 = ~n2954 & ~n2956;
  assign n2958 = ~n1154 & ~n2957;
  assign n2959 = pi328 & n2958;
  assign n2960 = ~n2953 & ~n2959;
  assign n2961 = ~n2680 & ~n2960;
  assign n2962 = n2680 & n2960;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = pi265 & ~n2963;
  assign n2965 = ~n2680 & n2960;
  assign n2966 = n2680 & ~n2960;
  assign n2967 = ~n2965 & ~n2966;
  assign n2968 = ~pi265 & ~n2967;
  assign n2969 = ~n2964 & ~n2968;
  assign n2970 = n2273 & ~n2550;
  assign n2971 = ~n2551 & ~n2970;
  assign n2972 = n2969 & ~n2971;
  assign n2973 = ~n2969 & n2971;
  assign n2974 = ~n2972 & ~n2973;
  assign n2975 = ~n2678 & ~n2974;
  assign n2976 = n2969 & n2971;
  assign n2977 = ~n2969 & ~n2971;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = n2678 & ~n2978;
  assign n2980 = ~n2975 & ~n2979;
  assign n2981 = ~n831 & ~n2980;
  assign n2982 = ~n2561 & ~n2981;
  assign n2983 = pi161 & ~n2982;
  assign n2984 = pi071 & ~pi161;
  assign n2985 = ~n2983 & ~n2984;
  assign po200 = ~pi160 & ~n2985;
  assign n2987 = pi266 & n831;
  assign n2988 = ~pi136 & ~n2174;
  assign n2989 = pi135 & n2988;
  assign n2990 = ~pi135 & pi136;
  assign n2991 = pi134 & n2990;
  assign n2992 = ~n2989 & ~n2991;
  assign n2993 = pi133 & ~n2992;
  assign n2994 = pi135 & pi136;
  assign n2995 = ~pi134 & n2994;
  assign n2996 = ~pi136 & n2174;
  assign n2997 = ~pi135 & n2996;
  assign n2998 = ~n2995 & ~n2997;
  assign n2999 = ~pi133 & ~n2998;
  assign n3000 = pi135 & ~pi136;
  assign n3001 = pi136 & ~n2174;
  assign n3002 = ~pi135 & n3001;
  assign n3003 = ~n3000 & ~n3002;
  assign n3004 = pi134 & ~n3003;
  assign n3005 = ~pi135 & ~pi136;
  assign n3006 = pi136 & n2174;
  assign n3007 = pi135 & n3006;
  assign n3008 = ~n3005 & ~n3007;
  assign n3009 = ~pi134 & ~n3008;
  assign n3010 = ~n3004 & ~n3009;
  assign n3011 = ~n2999 & n3010;
  assign n3012 = ~n2993 & n3011;
  assign n3013 = pi321 & n3012;
  assign n3014 = ~n2195 & n2574;
  assign n3015 = ~n2183 & ~n3014;
  assign n3016 = n1840 & ~n3015;
  assign n3017 = n2183 & ~n2588;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = pi321 & ~n3018;
  assign n3020 = n1840 & n2575;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = pi320 & ~n3021;
  assign n3023 = n2184 & n3014;
  assign n3024 = ~n3022 & ~n3023;
  assign n3025 = pi320 & n2574;
  assign n3026 = ~n3024 & ~n3025;
  assign n3027 = n2574 & n3024;
  assign n3028 = pi320 & n3027;
  assign n3029 = ~n3026 & ~n3028;
  assign n3030 = ~n3013 & ~n3029;
  assign n3031 = n3024 & ~n3025;
  assign n3032 = n2574 & ~n3024;
  assign n3033 = pi320 & n3032;
  assign n3034 = ~n3031 & ~n3033;
  assign n3035 = n3012 & ~n3034;
  assign n3036 = pi321 & n3035;
  assign n3037 = ~n3030 & ~n3036;
  assign n3038 = n1840 & ~n2604;
  assign n3039 = pi319 & n3038;
  assign n3040 = ~n2603 & ~n3039;
  assign n3041 = ~n3037 & ~n3040;
  assign n3042 = n3037 & n3040;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = n2183 & ~n3043;
  assign n3045 = pi319 & n3044;
  assign n3046 = pi319 & n2183;
  assign n3047 = n3037 & ~n3040;
  assign n3048 = ~n3037 & n3040;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = ~n3046 & ~n3049;
  assign n3051 = ~n3045 & ~n3050;
  assign n3052 = n1533 & ~n2617;
  assign n3053 = pi318 & n3052;
  assign n3054 = ~n2618 & ~n3053;
  assign n3055 = n3051 & n3054;
  assign n3056 = ~n3051 & ~n3054;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = n1840 & ~n3057;
  assign n3059 = pi318 & n3058;
  assign n3060 = pi318 & n1840;
  assign n3061 = ~n3051 & n3054;
  assign n3062 = n3051 & ~n3054;
  assign n3063 = ~n3061 & ~n3062;
  assign n3064 = ~n3060 & ~n3063;
  assign n3065 = ~n3059 & ~n3064;
  assign n3066 = n1553 & ~n2632;
  assign n3067 = pi317 & n3066;
  assign n3068 = ~n2631 & ~n3067;
  assign n3069 = ~n3065 & ~n3068;
  assign n3070 = n3065 & n3068;
  assign n3071 = ~n3069 & ~n3070;
  assign n3072 = n1533 & ~n3071;
  assign n3073 = pi317 & n3072;
  assign n3074 = pi317 & n1533;
  assign n3075 = n3065 & ~n3068;
  assign n3076 = ~n3065 & n3068;
  assign n3077 = ~n3075 & ~n3076;
  assign n3078 = ~n3074 & ~n3077;
  assign n3079 = ~n3073 & ~n3078;
  assign n3080 = n1515 & ~n2650;
  assign n3081 = pi316 & n3080;
  assign n3082 = ~n2649 & ~n3081;
  assign n3083 = ~n3079 & ~n3082;
  assign n3084 = n3079 & n3082;
  assign n3085 = ~n3083 & ~n3084;
  assign n3086 = n1553 & ~n3085;
  assign n3087 = pi316 & n3086;
  assign n3088 = pi316 & n1553;
  assign n3089 = n3079 & ~n3082;
  assign n3090 = ~n3079 & n3082;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = ~n3088 & ~n3091;
  assign n3093 = ~n3087 & ~n3092;
  assign n3094 = pi315 & n1515;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = n1515 & n3093;
  assign n3097 = pi315 & n3096;
  assign n3098 = ~n3095 & ~n3097;
  assign n3099 = ~n2268 & n2659;
  assign n3100 = ~pi129 & ~n3099;
  assign n3101 = pi128 & n3100;
  assign n3102 = ~n2659 & ~n2670;
  assign n3103 = pi129 & n3102;
  assign n3104 = ~n3101 & ~n3103;
  assign n3105 = pi315 & ~n3104;
  assign n3106 = n3098 & n3105;
  assign n3107 = ~n3098 & ~n3105;
  assign n3108 = ~n3106 & ~n3107;
  assign n3109 = pi128 & n2673;
  assign n3110 = ~pi129 & ~n3109;
  assign n3111 = pi129 & n2673;
  assign n3112 = pi128 & n3111;
  assign n3113 = pi314 & ~n3112;
  assign n3114 = ~n3110 & n3113;
  assign n3115 = ~n3108 & ~n3114;
  assign n3116 = n3098 & ~n3105;
  assign n3117 = ~n3098 & n3105;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = pi129 & ~n3109;
  assign n3120 = ~pi129 & n2673;
  assign n3121 = pi128 & n3120;
  assign n3122 = ~n3119 & ~n3121;
  assign n3123 = ~n3118 & ~n3122;
  assign n3124 = pi314 & n3123;
  assign n3125 = ~n3115 & ~n3124;
  assign n3126 = pi128 & pi313;
  assign n3127 = ~n3125 & ~n3126;
  assign n3128 = pi313 & n3125;
  assign n3129 = pi128 & n3128;
  assign n3130 = ~n3127 & ~n3129;
  assign n3131 = ~pi265 & ~n2962;
  assign n3132 = ~n2961 & ~n3131;
  assign n3133 = ~n2701 & n2712;
  assign n3134 = n2701 & ~n2712;
  assign n3135 = ~n2919 & ~n3134;
  assign n3136 = ~n3133 & ~n3135;
  assign n3137 = n2708 & n2926;
  assign n3138 = ~n2701 & ~n2919;
  assign n3139 = n2701 & n2919;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = n2712 & ~n3140;
  assign n3142 = n2701 & ~n2919;
  assign n3143 = ~n2701 & n2919;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n2712 & ~n3144;
  assign n3146 = ~n3141 & ~n3145;
  assign n3147 = ~n2708 & ~n2926;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = ~n3137 & ~n3148;
  assign n3150 = n3136 & ~n3149;
  assign n3151 = ~n3136 & n3149;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = n2464 & ~n2743;
  assign n3154 = pi323 & n3153;
  assign n3155 = ~n2737 & n2743;
  assign n3156 = n2887 & ~n3155;
  assign n3157 = pi322 & n3156;
  assign n3158 = ~n3154 & ~n3157;
  assign n3159 = ~n2728 & n2736;
  assign n3160 = n2728 & ~n2736;
  assign n3161 = ~n2898 & ~n3160;
  assign n3162 = ~n3159 & ~n3161;
  assign n3163 = ~n3158 & n3162;
  assign n3164 = n3158 & ~n3162;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = pi133 & pi261;
  assign n3167 = n2765 & ~n2771;
  assign n3168 = pi130 & pi264;
  assign n3169 = pi128 & pi266;
  assign n3170 = pi265 & ~n3169;
  assign n3171 = pi129 & n3170;
  assign n3172 = pi129 & pi265;
  assign n3173 = pi266 & ~n3172;
  assign n3174 = pi128 & n3173;
  assign n3175 = ~n3171 & ~n3174;
  assign n3176 = ~n3168 & ~n3175;
  assign n3177 = n3168 & n3175;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = ~n2745 & ~n2748;
  assign n3180 = n2745 & n2748;
  assign n3181 = ~n2756 & ~n3180;
  assign n3182 = ~n3179 & ~n3181;
  assign n3183 = ~n3178 & ~n3182;
  assign n3184 = ~n3168 & n3175;
  assign n3185 = n3168 & ~n3175;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~n2755 & ~n3179;
  assign n3188 = ~n2752 & n3187;
  assign n3189 = ~n3180 & ~n3188;
  assign n3190 = ~n3186 & ~n3189;
  assign n3191 = ~n3183 & ~n3190;
  assign n3192 = ~pi263 & ~n3191;
  assign n3193 = ~pi131 & ~n3191;
  assign n3194 = pi263 & n3191;
  assign n3195 = pi131 & n3194;
  assign n3196 = ~n3193 & ~n3195;
  assign n3197 = ~pi130 & ~n3196;
  assign n3198 = ~n3192 & ~n3197;
  assign n3199 = ~n3167 & ~n3198;
  assign n3200 = pi263 & n3167;
  assign n3201 = ~n2765 & ~n2771;
  assign n3202 = n2765 & n2771;
  assign n3203 = ~n3201 & ~n3202;
  assign n3204 = pi130 & ~n3203;
  assign n3205 = ~n3200 & ~n3204;
  assign n3206 = ~n3191 & ~n3205;
  assign n3207 = n2771 & n3191;
  assign n3208 = n2766 & n3207;
  assign n3209 = ~n3206 & ~n3208;
  assign n3210 = pi131 & ~n3209;
  assign n3211 = ~n2765 & n2771;
  assign n3212 = pi263 & ~n3211;
  assign n3213 = pi130 & n3212;
  assign n3214 = ~n3167 & ~n3213;
  assign n3215 = n3191 & ~n3214;
  assign n3216 = n2771 & ~n3191;
  assign n3217 = ~n2765 & n3216;
  assign n3218 = ~n3215 & ~n3217;
  assign n3219 = ~pi131 & ~n3218;
  assign n3220 = ~pi263 & n2765;
  assign n3221 = ~n2771 & n3191;
  assign n3222 = n3220 & n3221;
  assign n3223 = ~n3219 & ~n3222;
  assign n3224 = ~n3210 & n3223;
  assign n3225 = ~n3199 & n3224;
  assign n3226 = ~n2774 & ~n2775;
  assign n3227 = n2774 & n2775;
  assign n3228 = ~n2794 & ~n3227;
  assign n3229 = ~n3226 & ~n3228;
  assign n3230 = n3225 & ~n3229;
  assign n3231 = ~n3225 & n3229;
  assign n3232 = ~n3230 & ~n3231;
  assign n3233 = pi132 & pi262;
  assign n3234 = n2814 & ~n2819;
  assign n3235 = ~n2820 & ~n3234;
  assign n3236 = n3233 & ~n3235;
  assign n3237 = ~n2814 & ~n2820;
  assign n3238 = ~n2819 & ~n3237;
  assign n3239 = ~n3233 & ~n3238;
  assign n3240 = ~n3236 & ~n3239;
  assign n3241 = ~n3232 & ~n3240;
  assign n3242 = n3225 & n3229;
  assign n3243 = ~n3225 & ~n3229;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = ~n3233 & ~n3235;
  assign n3246 = n3233 & ~n3238;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = ~n3244 & ~n3247;
  assign n3249 = ~n3241 & ~n3248;
  assign n3250 = ~n3166 & n3249;
  assign n3251 = n3166 & ~n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = pi261 & ~n2821;
  assign n3254 = pi132 & n3253;
  assign n3255 = ~n2812 & ~n2814;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = pi260 & ~n3256;
  assign n3258 = pi133 & n3257;
  assign n3259 = pi134 & pi260;
  assign n3260 = ~n2813 & ~n3255;
  assign n3261 = ~n3254 & n3260;
  assign n3262 = n2838 & ~n3261;
  assign n3263 = ~n3259 & ~n3262;
  assign n3264 = ~n3258 & n3263;
  assign n3265 = ~n3258 & ~n3262;
  assign n3266 = n3259 & ~n3265;
  assign n3267 = ~n3264 & ~n3266;
  assign n3268 = ~n3252 & ~n3267;
  assign n3269 = ~n3166 & ~n3249;
  assign n3270 = n3166 & n3249;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = n3259 & ~n3262;
  assign n3273 = ~n3258 & n3272;
  assign n3274 = ~n3259 & ~n3265;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = ~n3271 & ~n3275;
  assign n3277 = ~n3268 & ~n3276;
  assign n3278 = n2843 & n2848;
  assign n3279 = ~n2843 & ~n2848;
  assign n3280 = ~n3258 & ~n3261;
  assign n3281 = n2838 & ~n3280;
  assign n3282 = ~n2838 & n3280;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~n3279 & ~n3283;
  assign n3285 = ~n3278 & ~n3284;
  assign n3286 = n3277 & n3285;
  assign n3287 = ~n3277 & ~n3285;
  assign n3288 = ~n3286 & ~n3287;
  assign n3289 = ~n3278 & ~n3279;
  assign n3290 = ~n2841 & ~n3289;
  assign n3291 = n2843 & ~n2848;
  assign n3292 = ~n2843 & n2848;
  assign n3293 = ~n3291 & ~n3292;
  assign n3294 = ~n2868 & ~n3293;
  assign n3295 = ~n3290 & ~n3294;
  assign n3296 = pi258 & ~n3295;
  assign n3297 = pi135 & n3296;
  assign n3298 = pi135 & pi259;
  assign n3299 = n3297 & n3298;
  assign n3300 = ~n3297 & ~n3298;
  assign n3301 = ~n3299 & ~n3300;
  assign n3302 = pi258 & ~n3301;
  assign n3303 = pi136 & n3302;
  assign n3304 = pi136 & pi258;
  assign n3305 = ~n3297 & n3298;
  assign n3306 = n3297 & ~n3298;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = ~n3304 & ~n3307;
  assign n3309 = ~n3303 & ~n3308;
  assign n3310 = ~n3288 & ~n3309;
  assign n3311 = ~n3277 & n3285;
  assign n3312 = n3277 & ~n3285;
  assign n3313 = ~n3311 & ~n3312;
  assign n3314 = pi258 & ~n3307;
  assign n3315 = pi136 & n3314;
  assign n3316 = ~n3301 & ~n3304;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = ~n3313 & ~n3317;
  assign n3319 = ~n3310 & ~n3318;
  assign n3320 = n2879 & ~n3319;
  assign n3321 = pi258 & ~n3289;
  assign n3322 = pi135 & n3321;
  assign n3323 = ~n2842 & ~n3293;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n2868 & ~n3324;
  assign n3326 = pi258 & ~n3293;
  assign n3327 = pi135 & n3326;
  assign n3328 = ~n2842 & ~n3289;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = ~n2841 & ~n3329;
  assign n3331 = ~n3325 & ~n3330;
  assign n3332 = ~n2879 & n3319;
  assign n3333 = n3331 & n3332;
  assign n3334 = ~n3320 & ~n3333;
  assign n3335 = ~n2852 & ~n3334;
  assign n3336 = ~n2879 & ~n3319;
  assign n3337 = n2879 & n3319;
  assign n3338 = ~n3331 & n3337;
  assign n3339 = ~n3336 & ~n3338;
  assign n3340 = n2852 & ~n3339;
  assign n3341 = ~n2879 & ~n3331;
  assign n3342 = n2879 & n3331;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3319 & ~n3343;
  assign n3345 = ~n3340 & ~n3344;
  assign n3346 = ~n3335 & n3345;
  assign n3347 = pi322 & ~n3346;
  assign n3348 = ~n2879 & n3331;
  assign n3349 = n2879 & ~n3331;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = n2852 & ~n3350;
  assign n3352 = ~n2852 & ~n3343;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = pi323 & ~n3353;
  assign n3355 = ~n3347 & ~n3354;
  assign n3356 = n2852 & n3348;
  assign n3357 = ~n3352 & ~n3356;
  assign n3358 = ~n3319 & ~n3357;
  assign n3359 = n2852 & ~n3331;
  assign n3360 = n3337 & n3359;
  assign n3361 = ~n3358 & ~n3360;
  assign n3362 = pi323 & ~n3361;
  assign n3363 = pi322 & n3362;
  assign n3364 = ~n3355 & ~n3363;
  assign n3365 = pi325 & n2091;
  assign n3366 = pi324 & n2464;
  assign n3367 = n3365 & n3366;
  assign n3368 = ~n3365 & ~n3366;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = ~n3364 & ~n3369;
  assign n3371 = ~n3365 & n3366;
  assign n3372 = n3365 & ~n3366;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = ~n3363 & ~n3373;
  assign n3375 = ~n3355 & n3374;
  assign n3376 = ~n3370 & ~n3375;
  assign n3377 = ~n3165 & ~n3376;
  assign n3378 = ~n3158 & ~n3162;
  assign n3379 = n3158 & n3162;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~n3364 & ~n3373;
  assign n3382 = ~n3363 & ~n3369;
  assign n3383 = ~n3355 & n3382;
  assign n3384 = ~n3381 & ~n3383;
  assign n3385 = ~n3380 & ~n3384;
  assign n3386 = ~n3377 & ~n3385;
  assign n3387 = n2728 & n2898;
  assign n3388 = ~n2728 & ~n2898;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = n2736 & ~n3389;
  assign n3391 = n2728 & ~n2898;
  assign n3392 = ~n2728 & n2898;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = ~n2736 & ~n3393;
  assign n3395 = ~n3390 & ~n3394;
  assign n3396 = n2732 & ~n2904;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = n1729 & ~n2732;
  assign n3399 = pi325 & n3398;
  assign n3400 = ~n3397 & ~n3399;
  assign n3401 = n3386 & n3400;
  assign n3402 = ~n3386 & ~n3400;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = pi327 & n1442;
  assign n3405 = pi326 & n1729;
  assign n3406 = n3404 & n3405;
  assign n3407 = ~n3404 & ~n3405;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = ~n3403 & ~n3408;
  assign n3410 = ~n3386 & n3400;
  assign n3411 = n3386 & ~n3400;
  assign n3412 = ~n3410 & ~n3411;
  assign n3413 = ~n3404 & n3405;
  assign n3414 = n3404 & ~n3405;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = ~n3412 & ~n3415;
  assign n3417 = ~n3409 & ~n3416;
  assign n3418 = ~n3152 & ~n3417;
  assign n3419 = n3136 & n3149;
  assign n3420 = ~n3136 & ~n3149;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = ~n3408 & ~n3412;
  assign n3423 = ~n3403 & ~n3415;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n3421 & ~n3424;
  assign n3426 = ~n3418 & ~n3425;
  assign n3427 = ~n1154 & n2925;
  assign n3428 = pi328 & n3427;
  assign n3429 = ~n2712 & ~n2926;
  assign n3430 = n2712 & n2926;
  assign n3431 = ~n3429 & ~n3430;
  assign n3432 = ~n3144 & ~n3431;
  assign n3433 = ~n1256 & ~n2712;
  assign n3434 = pi327 & n3433;
  assign n3435 = n1442 & ~n2926;
  assign n3436 = pi326 & n3435;
  assign n3437 = ~n3434 & ~n3436;
  assign n3438 = ~n3140 & ~n3437;
  assign n3439 = ~n3432 & ~n3438;
  assign n3440 = n2708 & n3439;
  assign n3441 = ~n2708 & ~n3439;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = ~n2681 & ~n2925;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = ~n3428 & ~n3444;
  assign n3446 = n3426 & ~n3445;
  assign n3447 = ~n3426 & n3445;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n2681 & ~n2947;
  assign n3450 = ~n1154 & n2947;
  assign n3451 = pi328 & n3450;
  assign n3452 = ~n3449 & ~n3451;
  assign n3453 = pi258 & ~n3452;
  assign n3454 = pi128 & n3453;
  assign n3455 = pi329 & n3454;
  assign n3456 = pi329 & ~n1154;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = n3455 & n3456;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = ~n1256 & ~n3459;
  assign n3461 = pi328 & n3460;
  assign n3462 = pi328 & ~n1256;
  assign n3463 = n3455 & ~n3456;
  assign n3464 = ~n3455 & n3456;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = ~n3462 & ~n3465;
  assign n3467 = ~n3461 & ~n3466;
  assign n3468 = ~n3448 & ~n3467;
  assign n3469 = n3426 & n3445;
  assign n3470 = ~n3426 & ~n3445;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = ~n1256 & ~n3465;
  assign n3473 = pi328 & n3472;
  assign n3474 = ~n3459 & ~n3462;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = ~n3471 & ~n3475;
  assign n3477 = ~n3468 & ~n3476;
  assign n3478 = pi330 & n1156;
  assign n3479 = n3477 & ~n3478;
  assign n3480 = pi330 & ~n3477;
  assign n3481 = n1156 & n3480;
  assign n3482 = ~n3479 & ~n3481;
  assign n3483 = ~n3132 & ~n3482;
  assign n3484 = n3132 & n3482;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = pi266 & ~n3485;
  assign n3487 = ~n3132 & n3482;
  assign n3488 = n3132 & ~n3482;
  assign n3489 = ~n3487 & ~n3488;
  assign n3490 = ~pi266 & ~n3489;
  assign n3491 = ~n3486 & ~n3490;
  assign n3492 = n2678 & ~n2976;
  assign n3493 = ~n2977 & ~n3492;
  assign n3494 = n3491 & ~n3493;
  assign n3495 = ~n3491 & n3493;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = ~n3130 & ~n3496;
  assign n3498 = n3491 & n3493;
  assign n3499 = ~n3491 & ~n3493;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = n3130 & ~n3500;
  assign n3502 = ~n3497 & ~n3501;
  assign n3503 = ~n831 & ~n3502;
  assign n3504 = ~n2987 & ~n3503;
  assign n3505 = pi161 & ~n3504;
  assign n3506 = pi072 & ~pi161;
  assign n3507 = ~n3505 & ~n3506;
  assign po201 = ~pi160 & ~n3507;
  assign n3509 = pi267 & n831;
  assign n3510 = ~n3093 & n3105;
  assign n3511 = n3093 & ~n3105;
  assign n3512 = n1515 & ~n3511;
  assign n3513 = pi315 & n3512;
  assign n3514 = ~n3510 & ~n3513;
  assign n3515 = ~pi129 & ~n2673;
  assign n3516 = ~n3118 & ~n3515;
  assign n3517 = ~pi128 & ~pi129;
  assign n3518 = n3113 & ~n3517;
  assign n3519 = ~n3516 & n3518;
  assign n3520 = n3514 & ~n3519;
  assign n3521 = ~n3514 & n3519;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = pi136 & ~pi137;
  assign n3524 = pi134 & n3523;
  assign n3525 = pi137 & ~n2174;
  assign n3526 = n3000 & n3525;
  assign n3527 = ~n3524 & ~n3526;
  assign n3528 = pi133 & ~n3527;
  assign n3529 = pi137 & n2174;
  assign n3530 = n2990 & n3529;
  assign n3531 = ~pi136 & ~pi137;
  assign n3532 = ~pi134 & n3531;
  assign n3533 = ~n3530 & ~n3532;
  assign n3534 = ~pi133 & ~n3533;
  assign n3535 = ~pi136 & pi137;
  assign n3536 = pi135 & n3535;
  assign n3537 = ~pi137 & ~n2174;
  assign n3538 = pi136 & n3537;
  assign n3539 = ~n3536 & ~n3538;
  assign n3540 = pi134 & ~n3539;
  assign n3541 = pi136 & pi137;
  assign n3542 = ~pi135 & n3541;
  assign n3543 = ~pi137 & n2174;
  assign n3544 = ~pi136 & n3543;
  assign n3545 = ~n3542 & ~n3544;
  assign n3546 = ~pi134 & ~n3545;
  assign n3547 = ~n2994 & ~n3005;
  assign n3548 = ~pi137 & ~n3547;
  assign n3549 = ~n3546 & ~n3548;
  assign n3550 = ~n3540 & n3549;
  assign n3551 = ~n3534 & n3550;
  assign n3552 = ~n3528 & n3551;
  assign n3553 = n3012 & ~n3024;
  assign n3554 = ~pi320 & ~n3553;
  assign n3555 = ~n2574 & ~n3012;
  assign n3556 = pi320 & n3553;
  assign n3557 = ~n3027 & ~n3556;
  assign n3558 = ~n3555 & n3557;
  assign n3559 = ~n3554 & n3558;
  assign n3560 = n3552 & ~n3559;
  assign n3561 = ~n3024 & ~n3552;
  assign n3562 = ~pi320 & n3012;
  assign n3563 = n3561 & n3562;
  assign n3564 = ~n3560 & ~n3563;
  assign n3565 = pi321 & ~n3564;
  assign n3566 = n3024 & ~n3552;
  assign n3567 = ~n2574 & n3566;
  assign n3568 = ~pi321 & ~n3032;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = n3012 & ~n3569;
  assign n3571 = pi321 & n3552;
  assign n3572 = ~n3024 & ~n3571;
  assign n3573 = ~n3012 & n3572;
  assign n3574 = n2574 & n3573;
  assign n3575 = ~n3570 & ~n3574;
  assign n3576 = pi320 & ~n3575;
  assign n3577 = ~n3565 & ~n3576;
  assign n3578 = n2183 & ~n3042;
  assign n3579 = pi319 & n3578;
  assign n3580 = ~n3041 & ~n3579;
  assign n3581 = ~n3577 & ~n3580;
  assign n3582 = n3577 & n3580;
  assign n3583 = ~n3581 & ~n3582;
  assign n3584 = n2574 & ~n3583;
  assign n3585 = pi319 & n3584;
  assign n3586 = pi319 & n2574;
  assign n3587 = n3577 & ~n3580;
  assign n3588 = ~n3577 & n3580;
  assign n3589 = ~n3587 & ~n3588;
  assign n3590 = ~n3586 & ~n3589;
  assign n3591 = ~n3585 & ~n3590;
  assign n3592 = n1840 & ~n3055;
  assign n3593 = pi318 & n3592;
  assign n3594 = ~n3056 & ~n3593;
  assign n3595 = n3591 & n3594;
  assign n3596 = ~n3591 & ~n3594;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = n2183 & ~n3597;
  assign n3599 = pi318 & n3598;
  assign n3600 = pi318 & n2183;
  assign n3601 = ~n3591 & n3594;
  assign n3602 = n3591 & ~n3594;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = ~n3600 & ~n3603;
  assign n3605 = ~n3599 & ~n3604;
  assign n3606 = n1533 & ~n3070;
  assign n3607 = pi317 & n3606;
  assign n3608 = ~n3069 & ~n3607;
  assign n3609 = ~n3605 & ~n3608;
  assign n3610 = n3605 & n3608;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = n1840 & ~n3611;
  assign n3613 = pi317 & n3612;
  assign n3614 = pi317 & n1840;
  assign n3615 = n3605 & ~n3608;
  assign n3616 = ~n3605 & n3608;
  assign n3617 = ~n3615 & ~n3616;
  assign n3618 = ~n3614 & ~n3617;
  assign n3619 = ~n3613 & ~n3618;
  assign n3620 = pi316 & n1533;
  assign n3621 = ~n3619 & ~n3620;
  assign n3622 = n1533 & n3619;
  assign n3623 = pi316 & n3622;
  assign n3624 = ~n3621 & ~n3623;
  assign n3625 = n1553 & ~n3084;
  assign n3626 = pi316 & n3625;
  assign n3627 = ~n3083 & ~n3626;
  assign n3628 = ~n3624 & ~n3627;
  assign n3629 = n3624 & n3627;
  assign n3630 = ~n3628 & ~n3629;
  assign n3631 = n1553 & ~n3630;
  assign n3632 = pi315 & n3631;
  assign n3633 = pi315 & n1553;
  assign n3634 = n3624 & ~n3627;
  assign n3635 = ~n3624 & n3627;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = ~n3633 & ~n3636;
  assign n3638 = ~n3632 & ~n3637;
  assign n3639 = pi314 & n1515;
  assign n3640 = n3638 & ~n3639;
  assign n3641 = n1515 & ~n3638;
  assign n3642 = pi314 & n3641;
  assign n3643 = ~n3640 & ~n3642;
  assign n3644 = ~n3522 & ~n3643;
  assign n3645 = ~n3514 & ~n3519;
  assign n3646 = n3514 & n3519;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n3638 & ~n3639;
  assign n3649 = n1515 & n3638;
  assign n3650 = pi314 & n3649;
  assign n3651 = ~n3648 & ~n3650;
  assign n3652 = ~n3647 & ~n3651;
  assign n3653 = ~n3644 & ~n3652;
  assign n3654 = pi129 & n3653;
  assign n3655 = pi313 & ~n3653;
  assign n3656 = ~pi129 & n3655;
  assign n3657 = ~n3654 & ~n3656;
  assign n3658 = n3125 & ~n3657;
  assign n3659 = pi128 & n3658;
  assign n3660 = ~pi313 & n3653;
  assign n3661 = pi128 & n3125;
  assign n3662 = ~pi129 & n3653;
  assign n3663 = pi129 & n3655;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = ~n3661 & ~n3664;
  assign n3666 = ~n3660 & ~n3665;
  assign n3667 = ~n3659 & n3666;
  assign n3668 = pi128 & pi312;
  assign n3669 = ~n3667 & ~n3668;
  assign n3670 = pi312 & n3667;
  assign n3671 = pi128 & n3670;
  assign n3672 = ~n3669 & ~n3671;
  assign n3673 = ~pi266 & ~n3484;
  assign n3674 = ~n3483 & ~n3673;
  assign n3675 = n1156 & n3477;
  assign n3676 = ~n1154 & ~n3675;
  assign n3677 = n1154 & n3477;
  assign n3678 = n1156 & n3677;
  assign n3679 = ~n3676 & ~n3678;
  assign n3680 = pi330 & ~n3679;
  assign n3681 = ~n1256 & ~n3469;
  assign n3682 = pi328 & n3681;
  assign n3683 = ~n3470 & ~n3682;
  assign n3684 = ~n1256 & ~n3448;
  assign n3685 = pi328 & n3684;
  assign n3686 = ~n3462 & ~n3471;
  assign n3687 = ~n3685 & ~n3686;
  assign n3688 = ~n3458 & ~n3687;
  assign n3689 = ~n3457 & ~n3688;
  assign n3690 = n3683 & n3689;
  assign n3691 = ~n3683 & ~n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = pi329 & ~n1256;
  assign n3694 = ~n3136 & n3405;
  assign n3695 = n3136 & ~n3405;
  assign n3696 = ~n3412 & ~n3695;
  assign n3697 = ~n3694 & ~n3696;
  assign n3698 = ~n3136 & ~n3400;
  assign n3699 = n3136 & n3400;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3149 & n3404;
  assign n3702 = ~n3386 & n3405;
  assign n3703 = n3386 & ~n3405;
  assign n3704 = ~n3702 & ~n3703;
  assign n3705 = ~n3701 & ~n3704;
  assign n3706 = ~n3700 & n3705;
  assign n3707 = ~n3136 & n3400;
  assign n3708 = n3136 & ~n3400;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n3386 & n3405;
  assign n3711 = ~n3386 & ~n3405;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~n3701 & ~n3712;
  assign n3714 = ~n3709 & n3713;
  assign n3715 = n3149 & ~n3404;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = ~n3706 & n3716;
  assign n3718 = n3697 & n3717;
  assign n3719 = ~n3697 & ~n3717;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = ~n3158 & ~n3355;
  assign n3722 = ~n3363 & ~n3721;
  assign n3723 = ~n3162 & n3366;
  assign n3724 = ~n3158 & ~n3364;
  assign n3725 = n3158 & ~n3363;
  assign n3726 = ~n3355 & n3725;
  assign n3727 = ~n3724 & ~n3726;
  assign n3728 = n3162 & ~n3366;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~n3723 & ~n3729;
  assign n3731 = ~n3722 & n3730;
  assign n3732 = n3722 & ~n3730;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n2852 & ~n3342;
  assign n3735 = ~n3341 & ~n3734;
  assign n3736 = n3169 & n3172;
  assign n3737 = ~n3169 & ~n3172;
  assign n3738 = ~n3189 & ~n3737;
  assign n3739 = ~n3736 & ~n3738;
  assign n3740 = pi128 & pi267;
  assign n3741 = pi266 & ~n3740;
  assign n3742 = pi129 & n3741;
  assign n3743 = pi129 & pi266;
  assign n3744 = pi267 & ~n3743;
  assign n3745 = pi128 & n3744;
  assign n3746 = ~n3742 & ~n3745;
  assign n3747 = ~n3739 & ~n3746;
  assign n3748 = n3739 & n3746;
  assign n3749 = ~n3747 & ~n3748;
  assign n3750 = pi265 & ~n3749;
  assign n3751 = pi130 & n3750;
  assign n3752 = pi130 & pi265;
  assign n3753 = n3739 & ~n3746;
  assign n3754 = ~n3739 & n3746;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n3752 & ~n3755;
  assign n3757 = ~n3751 & ~n3756;
  assign n3758 = ~n3175 & n3189;
  assign n3759 = n3175 & ~n3189;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = n3168 & ~n3760;
  assign n3762 = ~n3168 & n3760;
  assign n3763 = n2744 & ~n3211;
  assign n3764 = ~n3167 & ~n3763;
  assign n3765 = ~n3762 & ~n3764;
  assign n3766 = ~n3761 & ~n3765;
  assign n3767 = n3757 & n3766;
  assign n3768 = ~n3757 & ~n3766;
  assign n3769 = ~n3767 & ~n3768;
  assign n3770 = pi130 & ~n3211;
  assign n3771 = ~n3167 & ~n3770;
  assign n3772 = n3191 & ~n3771;
  assign n3773 = ~pi130 & ~n3167;
  assign n3774 = ~n3211 & ~n3773;
  assign n3775 = ~n3191 & ~n3774;
  assign n3776 = ~n3772 & ~n3775;
  assign n3777 = pi263 & ~n3776;
  assign n3778 = pi131 & n3777;
  assign n3779 = pi131 & pi264;
  assign n3780 = ~n3191 & ~n3214;
  assign n3781 = n3191 & ~n3774;
  assign n3782 = ~n3780 & ~n3781;
  assign n3783 = ~pi131 & ~n3782;
  assign n3784 = ~n2771 & ~n3191;
  assign n3785 = n2765 & n3784;
  assign n3786 = ~n3167 & n3191;
  assign n3787 = ~n3785 & ~n3786;
  assign n3788 = ~pi263 & ~n3787;
  assign n3789 = ~n3783 & ~n3788;
  assign n3790 = n3229 & n3789;
  assign n3791 = ~n3779 & ~n3790;
  assign n3792 = ~n3778 & n3791;
  assign n3793 = ~n3778 & ~n3790;
  assign n3794 = n3779 & ~n3793;
  assign n3795 = ~n3792 & ~n3794;
  assign n3796 = ~n3769 & ~n3795;
  assign n3797 = n3757 & ~n3766;
  assign n3798 = ~n3757 & n3766;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = n3779 & ~n3790;
  assign n3801 = ~n3778 & n3800;
  assign n3802 = ~n3779 & ~n3793;
  assign n3803 = ~n3801 & ~n3802;
  assign n3804 = ~n3799 & ~n3803;
  assign n3805 = ~n3796 & ~n3804;
  assign n3806 = n3233 & ~n3244;
  assign n3807 = ~n3233 & n3244;
  assign n3808 = ~n3235 & ~n3807;
  assign n3809 = ~n3806 & ~n3808;
  assign n3810 = n3805 & n3809;
  assign n3811 = ~n3805 & ~n3809;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = pi133 & pi262;
  assign n3814 = pi132 & pi263;
  assign n3815 = n3813 & n3814;
  assign n3816 = ~n3813 & ~n3814;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3812 & ~n3817;
  assign n3819 = ~n3805 & n3809;
  assign n3820 = n3805 & ~n3809;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = pi262 & ~n3814;
  assign n3823 = pi133 & n3822;
  assign n3824 = pi263 & ~n3813;
  assign n3825 = pi132 & n3824;
  assign n3826 = ~n3823 & ~n3825;
  assign n3827 = ~n3821 & ~n3826;
  assign n3828 = ~n3818 & ~n3827;
  assign n3829 = ~n3265 & ~n3269;
  assign n3830 = ~n3270 & ~n3829;
  assign n3831 = n3828 & n3830;
  assign n3832 = ~n3828 & ~n3830;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = pi134 & pi261;
  assign n3835 = n3249 & ~n3262;
  assign n3836 = ~n3258 & n3835;
  assign n3837 = ~n3249 & ~n3265;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n3166 & ~n3838;
  assign n3840 = ~n3249 & ~n3262;
  assign n3841 = ~n3258 & n3840;
  assign n3842 = n3249 & ~n3265;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = pi261 & ~n3843;
  assign n3845 = pi133 & n3844;
  assign n3846 = ~n3839 & ~n3845;
  assign n3847 = ~n3285 & ~n3846;
  assign n3848 = n3285 & n3846;
  assign n3849 = n3259 & ~n3848;
  assign n3850 = ~n3847 & ~n3849;
  assign n3851 = n3834 & ~n3850;
  assign n3852 = ~n3259 & ~n3847;
  assign n3853 = ~n3848 & ~n3852;
  assign n3854 = ~n3834 & ~n3853;
  assign n3855 = ~n3851 & ~n3854;
  assign n3856 = ~n3833 & ~n3855;
  assign n3857 = n3828 & ~n3830;
  assign n3858 = ~n3828 & n3830;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = ~n3834 & ~n3850;
  assign n3861 = n3834 & ~n3853;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = ~n3859 & ~n3862;
  assign n3864 = ~n3856 & ~n3863;
  assign n3865 = ~n3300 & ~n3313;
  assign n3866 = ~n3299 & ~n3865;
  assign n3867 = n3864 & n3866;
  assign n3868 = ~n3864 & ~n3866;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = pi136 & pi259;
  assign n3871 = ~n3288 & ~n3301;
  assign n3872 = ~n3307 & ~n3313;
  assign n3873 = n3304 & ~n3872;
  assign n3874 = ~n3871 & n3873;
  assign n3875 = ~n3870 & ~n3874;
  assign n3876 = pi135 & n3297;
  assign n3877 = ~pi135 & ~n3297;
  assign n3878 = ~n3876 & ~n3877;
  assign n3879 = ~n3313 & ~n3878;
  assign n3880 = pi135 & ~n3297;
  assign n3881 = ~pi135 & n3297;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = ~n3288 & ~n3882;
  assign n3884 = ~n3879 & ~n3883;
  assign n3885 = n3304 & ~n3884;
  assign n3886 = pi259 & n3885;
  assign n3887 = ~n3875 & ~n3886;
  assign n3888 = pi137 & pi258;
  assign n3889 = pi135 & pi260;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = n3888 & n3889;
  assign n3892 = ~n3890 & ~n3891;
  assign n3893 = ~n3887 & ~n3892;
  assign n3894 = ~n3888 & n3889;
  assign n3895 = n3888 & ~n3889;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3886 & ~n3896;
  assign n3898 = ~n3875 & n3897;
  assign n3899 = ~n3893 & ~n3898;
  assign n3900 = ~n3869 & ~n3899;
  assign n3901 = n3864 & ~n3866;
  assign n3902 = ~n3864 & n3866;
  assign n3903 = ~n3901 & ~n3902;
  assign n3904 = ~n3887 & ~n3896;
  assign n3905 = ~n3886 & ~n3892;
  assign n3906 = ~n3875 & n3905;
  assign n3907 = ~n3904 & ~n3906;
  assign n3908 = ~n3903 & ~n3907;
  assign n3909 = ~n3900 & ~n3908;
  assign n3910 = n3735 & ~n3909;
  assign n3911 = ~n3735 & n3909;
  assign n3912 = n3319 & n3911;
  assign n3913 = ~n3910 & ~n3912;
  assign n3914 = ~n3331 & ~n3913;
  assign n3915 = ~n3735 & ~n3909;
  assign n3916 = n3735 & n3909;
  assign n3917 = ~n3319 & n3916;
  assign n3918 = ~n3915 & ~n3917;
  assign n3919 = n3331 & ~n3918;
  assign n3920 = ~n3319 & ~n3735;
  assign n3921 = n3319 & n3735;
  assign n3922 = ~n3920 & ~n3921;
  assign n3923 = ~n3909 & ~n3922;
  assign n3924 = ~n3919 & ~n3923;
  assign n3925 = ~n3914 & n3924;
  assign n3926 = pi322 & ~n3925;
  assign n3927 = n3319 & ~n3735;
  assign n3928 = ~n3319 & n3735;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = n3331 & ~n3929;
  assign n3931 = ~n3331 & ~n3922;
  assign n3932 = ~n3930 & ~n3931;
  assign n3933 = pi323 & ~n3932;
  assign n3934 = ~n3926 & ~n3933;
  assign n3935 = n3331 & n3927;
  assign n3936 = ~n3931 & ~n3935;
  assign n3937 = ~n3909 & ~n3936;
  assign n3938 = ~n3319 & n3331;
  assign n3939 = n3916 & n3938;
  assign n3940 = ~n3937 & ~n3939;
  assign n3941 = pi323 & ~n3940;
  assign n3942 = pi322 & n3941;
  assign n3943 = ~n3934 & ~n3942;
  assign n3944 = pi325 & n2464;
  assign n3945 = pi324 & n2887;
  assign n3946 = n3944 & n3945;
  assign n3947 = ~n3944 & ~n3945;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = ~n3943 & ~n3948;
  assign n3950 = ~n3944 & n3945;
  assign n3951 = n3944 & ~n3945;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = ~n3942 & ~n3952;
  assign n3954 = ~n3934 & n3953;
  assign n3955 = ~n3949 & ~n3954;
  assign n3956 = ~n3733 & ~n3955;
  assign n3957 = ~n3722 & ~n3730;
  assign n3958 = n3722 & n3730;
  assign n3959 = ~n3957 & ~n3958;
  assign n3960 = ~n3943 & ~n3952;
  assign n3961 = ~n3942 & ~n3948;
  assign n3962 = ~n3934 & n3961;
  assign n3963 = ~n3960 & ~n3962;
  assign n3964 = ~n3959 & ~n3963;
  assign n3965 = ~n3956 & ~n3964;
  assign n3966 = n3365 & ~n3400;
  assign n3967 = ~n3162 & ~n3727;
  assign n3968 = n3162 & n3727;
  assign n3969 = ~n3967 & ~n3968;
  assign n3970 = n3366 & ~n3969;
  assign n3971 = n3162 & ~n3727;
  assign n3972 = ~n3162 & n3727;
  assign n3973 = ~n3971 & ~n3972;
  assign n3974 = ~n3366 & ~n3973;
  assign n3975 = ~n3970 & ~n3974;
  assign n3976 = ~n3365 & n3400;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3966 & ~n3977;
  assign n3979 = n3965 & n3978;
  assign n3980 = ~n3965 & ~n3978;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = pi327 & n1729;
  assign n3983 = pi326 & n2091;
  assign n3984 = n3982 & n3983;
  assign n3985 = ~n3982 & ~n3983;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = ~n3981 & ~n3986;
  assign n3988 = ~n3965 & n3978;
  assign n3989 = n3965 & ~n3978;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = ~n3982 & n3983;
  assign n3992 = n3982 & ~n3983;
  assign n3993 = ~n3991 & ~n3992;
  assign n3994 = ~n3990 & ~n3993;
  assign n3995 = ~n3987 & ~n3994;
  assign n3996 = ~n3720 & ~n3995;
  assign n3997 = n3697 & ~n3717;
  assign n3998 = ~n3697 & n3717;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = ~n3986 & ~n3990;
  assign n4001 = ~n3981 & ~n3993;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = ~n3999 & ~n4002;
  assign n4004 = ~n3996 & ~n4003;
  assign n4005 = ~n3693 & n4004;
  assign n4006 = n3693 & ~n4004;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = n1442 & ~n4007;
  assign n4009 = pi328 & n4008;
  assign n4010 = pi328 & n1442;
  assign n4011 = n3693 & n4004;
  assign n4012 = ~n3693 & ~n4004;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = ~n4010 & ~n4013;
  assign n4015 = ~n4009 & ~n4014;
  assign n4016 = ~n3692 & ~n4015;
  assign n4017 = n3683 & ~n3689;
  assign n4018 = ~n3683 & n3689;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = n1442 & ~n4013;
  assign n4021 = pi328 & n4020;
  assign n4022 = ~n4007 & ~n4010;
  assign n4023 = ~n4021 & ~n4022;
  assign n4024 = ~n4019 & ~n4023;
  assign n4025 = ~n4016 & ~n4024;
  assign n4026 = n3680 & n4025;
  assign n4027 = ~n3680 & ~n4025;
  assign n4028 = ~n4026 & ~n4027;
  assign n4029 = pi258 & ~n4028;
  assign n4030 = pi128 & n4029;
  assign n4031 = pi331 & n4030;
  assign n4032 = n3680 & ~n4025;
  assign n4033 = ~n3680 & n4025;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = pi331 & n1156;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n4031 & ~n4036;
  assign n4038 = ~n3674 & ~n4037;
  assign n4039 = n3674 & n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = pi267 & ~n4040;
  assign n4042 = ~n3674 & n4037;
  assign n4043 = n3674 & ~n4037;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = ~pi267 & ~n4044;
  assign n4046 = ~n4041 & ~n4045;
  assign n4047 = n3130 & ~n3498;
  assign n4048 = ~n3499 & ~n4047;
  assign n4049 = n4046 & ~n4048;
  assign n4050 = ~n4046 & n4048;
  assign n4051 = ~n4049 & ~n4050;
  assign n4052 = ~n3672 & ~n4051;
  assign n4053 = n4046 & n4048;
  assign n4054 = ~n4046 & ~n4048;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = n3672 & ~n4055;
  assign n4057 = ~n4052 & ~n4056;
  assign n4058 = ~n831 & ~n4057;
  assign n4059 = ~n3509 & ~n4058;
  assign n4060 = pi161 & ~n4059;
  assign n4061 = pi073 & ~pi161;
  assign n4062 = ~n4060 & ~n4061;
  assign po202 = ~pi160 & ~n4062;
  assign n4064 = pi268 & n831;
  assign n4065 = pi312 & ~n1568;
  assign n4066 = ~n3619 & ~n3627;
  assign n4067 = pi134 & pi136;
  assign n4068 = pi135 & n3525;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = pi133 & ~n4069;
  assign n4071 = pi135 & pi137;
  assign n4072 = ~n3001 & ~n4071;
  assign n4073 = pi134 & ~n4072;
  assign n4074 = ~pi135 & ~pi137;
  assign n4075 = pi136 & ~n4074;
  assign n4076 = ~n4073 & ~n4075;
  assign n4077 = ~n4070 & n4076;
  assign n4078 = pi138 & n4077;
  assign n4079 = ~pi138 & ~n4077;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = pi137 & ~n4080;
  assign n4082 = pi138 & ~n4077;
  assign n4083 = ~pi138 & n4077;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~pi137 & ~n4084;
  assign n4086 = ~n4081 & ~n4085;
  assign n4087 = pi321 & n4086;
  assign n4088 = ~n3024 & n3552;
  assign n4089 = ~n3012 & ~n4088;
  assign n4090 = n2574 & ~n4089;
  assign n4091 = n3012 & ~n3566;
  assign n4092 = ~n4090 & ~n4091;
  assign n4093 = pi321 & ~n4092;
  assign n4094 = n2574 & n3553;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = pi320 & ~n4095;
  assign n4097 = n3013 & n4088;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = pi320 & n3552;
  assign n4100 = ~n4098 & ~n4099;
  assign n4101 = n3552 & n4098;
  assign n4102 = pi320 & n4101;
  assign n4103 = ~n4100 & ~n4102;
  assign n4104 = ~n4087 & ~n4103;
  assign n4105 = n4098 & ~n4099;
  assign n4106 = n3552 & ~n4098;
  assign n4107 = pi320 & n4106;
  assign n4108 = ~n4105 & ~n4107;
  assign n4109 = n4086 & ~n4108;
  assign n4110 = pi321 & n4109;
  assign n4111 = ~n4104 & ~n4110;
  assign n4112 = n2574 & ~n3582;
  assign n4113 = pi319 & n4112;
  assign n4114 = ~n3581 & ~n4113;
  assign n4115 = ~n4111 & ~n4114;
  assign n4116 = n4111 & n4114;
  assign n4117 = ~n4115 & ~n4116;
  assign n4118 = n3012 & ~n4117;
  assign n4119 = pi319 & n4118;
  assign n4120 = pi319 & n3012;
  assign n4121 = n4111 & ~n4114;
  assign n4122 = ~n4111 & n4114;
  assign n4123 = ~n4121 & ~n4122;
  assign n4124 = ~n4120 & ~n4123;
  assign n4125 = ~n4119 & ~n4124;
  assign n4126 = n2183 & ~n3595;
  assign n4127 = pi318 & n4126;
  assign n4128 = ~n3596 & ~n4127;
  assign n4129 = n4125 & n4128;
  assign n4130 = ~n4125 & ~n4128;
  assign n4131 = ~n4129 & ~n4130;
  assign n4132 = n2574 & ~n4131;
  assign n4133 = pi318 & n4132;
  assign n4134 = pi318 & n2574;
  assign n4135 = ~n4125 & n4128;
  assign n4136 = n4125 & ~n4128;
  assign n4137 = ~n4135 & ~n4136;
  assign n4138 = ~n4134 & ~n4137;
  assign n4139 = ~n4133 & ~n4138;
  assign n4140 = ~pi317 & ~n4139;
  assign n4141 = ~n2183 & ~n4139;
  assign n4142 = n2183 & n4139;
  assign n4143 = pi317 & n4142;
  assign n4144 = ~n4141 & ~n4143;
  assign n4145 = ~n1840 & ~n4144;
  assign n4146 = ~n4140 & ~n4145;
  assign n4147 = ~n3609 & ~n4146;
  assign n4148 = n3608 & n4139;
  assign n4149 = n3605 & n4148;
  assign n4150 = ~n3608 & ~n4139;
  assign n4151 = ~n3605 & n4150;
  assign n4152 = ~n4149 & ~n4151;
  assign n4153 = pi317 & ~n4152;
  assign n4154 = ~n3617 & ~n4139;
  assign n4155 = n1840 & n4154;
  assign n4156 = ~n4153 & ~n4155;
  assign n4157 = n2183 & ~n4156;
  assign n4158 = n3608 & ~n4139;
  assign n4159 = n3605 & n4158;
  assign n4160 = n1840 & ~n3610;
  assign n4161 = pi317 & n4160;
  assign n4162 = ~n3609 & ~n4161;
  assign n4163 = n4139 & ~n4162;
  assign n4164 = ~n4159 & ~n4163;
  assign n4165 = ~n2183 & ~n4164;
  assign n4166 = ~pi317 & ~n3605;
  assign n4167 = ~n3608 & n4139;
  assign n4168 = n4166 & n4167;
  assign n4169 = ~n4165 & ~n4168;
  assign n4170 = ~n4157 & n4169;
  assign n4171 = ~n4147 & n4170;
  assign n4172 = ~pi316 & ~n4171;
  assign n4173 = ~n1840 & ~n4171;
  assign n4174 = n1840 & n4171;
  assign n4175 = pi316 & n4174;
  assign n4176 = ~n4173 & ~n4175;
  assign n4177 = ~n1533 & ~n4176;
  assign n4178 = ~n4172 & ~n4177;
  assign n4179 = ~n4066 & ~n4178;
  assign n4180 = n3627 & n4171;
  assign n4181 = n3619 & n4180;
  assign n4182 = ~n3627 & ~n4171;
  assign n4183 = ~n3619 & n4182;
  assign n4184 = ~n4181 & ~n4183;
  assign n4185 = pi316 & ~n4184;
  assign n4186 = ~n3619 & n3627;
  assign n4187 = n3619 & ~n3627;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~n4171 & ~n4188;
  assign n4190 = n1533 & n4189;
  assign n4191 = ~n4185 & ~n4190;
  assign n4192 = n1840 & ~n4191;
  assign n4193 = n3627 & ~n4171;
  assign n4194 = n3619 & n4193;
  assign n4195 = n3619 & n3627;
  assign n4196 = n1533 & ~n4195;
  assign n4197 = pi316 & n4196;
  assign n4198 = ~n4066 & ~n4197;
  assign n4199 = n4171 & ~n4198;
  assign n4200 = ~n4194 & ~n4199;
  assign n4201 = ~n1840 & ~n4200;
  assign n4202 = ~pi316 & ~n3619;
  assign n4203 = ~n3627 & n4171;
  assign n4204 = n4202 & n4203;
  assign n4205 = ~n4201 & ~n4204;
  assign n4206 = ~n4192 & n4205;
  assign n4207 = ~n4179 & n4206;
  assign n4208 = n3514 & ~n3633;
  assign n4209 = ~n3636 & ~n4208;
  assign n4210 = n1553 & ~n3514;
  assign n4211 = pi315 & n4210;
  assign n4212 = ~n4209 & ~n4211;
  assign n4213 = ~n4207 & n4212;
  assign n4214 = n4207 & ~n4212;
  assign n4215 = ~n4213 & ~n4214;
  assign n4216 = n1533 & ~n4215;
  assign n4217 = pi315 & n4216;
  assign n4218 = pi315 & n1533;
  assign n4219 = n4207 & n4212;
  assign n4220 = ~n4207 & ~n4212;
  assign n4221 = ~n4219 & ~n4220;
  assign n4222 = ~n4218 & ~n4221;
  assign n4223 = ~n4217 & ~n4222;
  assign n4224 = n3514 & ~n3638;
  assign n4225 = ~n3514 & n3638;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = ~n3519 & ~n3639;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = n1515 & n3519;
  assign n4230 = pi314 & n4229;
  assign n4231 = ~n4228 & ~n4230;
  assign n4232 = ~n4223 & ~n4231;
  assign n4233 = n4223 & n4231;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = n1553 & ~n4234;
  assign n4236 = pi314 & n4235;
  assign n4237 = pi314 & n1553;
  assign n4238 = n4223 & ~n4231;
  assign n4239 = ~n4223 & n4231;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = ~n4237 & ~n4240;
  assign n4242 = ~n4236 & ~n4241;
  assign n4243 = n4065 & ~n4242;
  assign n4244 = ~n4065 & n4242;
  assign n4245 = ~n4243 & ~n4244;
  assign n4246 = ~n3667 & n3668;
  assign n4247 = n3125 & ~n3653;
  assign n4248 = ~pi129 & ~n4247;
  assign n4249 = pi128 & n4248;
  assign n4250 = n3653 & ~n3661;
  assign n4251 = pi129 & n4250;
  assign n4252 = ~n4249 & ~n4251;
  assign n4253 = pi313 & ~n4252;
  assign n4254 = pi313 & n1515;
  assign n4255 = n4253 & n4254;
  assign n4256 = ~n4253 & ~n4254;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = n4246 & ~n4257;
  assign n4259 = ~n4246 & n4257;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = ~n4245 & ~n4260;
  assign n4262 = n4065 & n4242;
  assign n4263 = ~n4065 & ~n4242;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = n4246 & n4257;
  assign n4266 = ~n4246 & ~n4257;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~n4264 & ~n4267;
  assign n4269 = ~n4261 & ~n4268;
  assign n4270 = pi311 & ~n4269;
  assign n4271 = pi128 & n4270;
  assign n4272 = pi128 & pi311;
  assign n4273 = n4269 & ~n4272;
  assign n4274 = ~n4271 & ~n4273;
  assign n4275 = ~pi267 & ~n4039;
  assign n4276 = ~n4038 & ~n4275;
  assign n4277 = ~n1154 & n4025;
  assign n4278 = n1154 & ~n4025;
  assign n4279 = n3477 & ~n4278;
  assign n4280 = n1156 & n4279;
  assign n4281 = ~n4277 & ~n4280;
  assign n4282 = n1256 & ~n4281;
  assign n4283 = ~n3675 & ~n4277;
  assign n4284 = ~n4278 & ~n4283;
  assign n4285 = ~n1256 & ~n4284;
  assign n4286 = ~n4282 & ~n4285;
  assign n4287 = pi330 & ~n4286;
  assign n4288 = ~n3683 & ~n4004;
  assign n4289 = n3683 & n4004;
  assign n4290 = n1442 & ~n4289;
  assign n4291 = pi328 & n4290;
  assign n4292 = ~n4288 & ~n4291;
  assign n4293 = ~n3689 & ~n3693;
  assign n4294 = n3689 & n3693;
  assign n4295 = ~n3683 & n4004;
  assign n4296 = n3683 & ~n4004;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = n1442 & ~n4297;
  assign n4299 = pi328 & n4298;
  assign n4300 = ~n4288 & ~n4289;
  assign n4301 = ~n4010 & ~n4300;
  assign n4302 = ~n4299 & ~n4301;
  assign n4303 = ~n4294 & ~n4302;
  assign n4304 = ~n4293 & ~n4303;
  assign n4305 = n4292 & n4304;
  assign n4306 = ~n4292 & ~n4304;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = pi329 & n1442;
  assign n4309 = ~n3697 & n3983;
  assign n4310 = n3697 & ~n3983;
  assign n4311 = ~n3990 & ~n4310;
  assign n4312 = ~n4309 & ~n4311;
  assign n4313 = ~n3697 & ~n3978;
  assign n4314 = n3697 & n3978;
  assign n4315 = ~n4313 & ~n4314;
  assign n4316 = n3717 & n3982;
  assign n4317 = ~n3965 & n3983;
  assign n4318 = n3965 & ~n3983;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = ~n4316 & ~n4319;
  assign n4321 = ~n4315 & n4320;
  assign n4322 = ~n3697 & n3978;
  assign n4323 = n3697 & ~n3978;
  assign n4324 = ~n4322 & ~n4323;
  assign n4325 = n3965 & n3983;
  assign n4326 = ~n3965 & ~n3983;
  assign n4327 = ~n4325 & ~n4326;
  assign n4328 = ~n4316 & ~n4327;
  assign n4329 = ~n4324 & n4328;
  assign n4330 = ~n3717 & ~n3982;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~n4321 & n4331;
  assign n4333 = n4312 & n4332;
  assign n4334 = ~n4312 & ~n4332;
  assign n4335 = ~n4333 & ~n4334;
  assign n4336 = ~n3722 & ~n3934;
  assign n4337 = ~n3942 & ~n4336;
  assign n4338 = ~n3730 & n3945;
  assign n4339 = ~n3722 & ~n3943;
  assign n4340 = n3722 & ~n3942;
  assign n4341 = ~n3934 & n4340;
  assign n4342 = ~n4339 & ~n4341;
  assign n4343 = n3730 & ~n3945;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = ~n4338 & ~n4344;
  assign n4346 = ~n4337 & n4345;
  assign n4347 = n4337 & ~n4345;
  assign n4348 = ~n4346 & ~n4347;
  assign n4349 = ~n3331 & ~n3921;
  assign n4350 = ~n3920 & ~n4349;
  assign n4351 = pi136 & pi260;
  assign n4352 = n3889 & n4351;
  assign n4353 = ~n3886 & n4352;
  assign n4354 = ~n3889 & ~n4351;
  assign n4355 = ~n3875 & n4354;
  assign n4356 = ~n4353 & ~n4355;
  assign n4357 = ~n3869 & ~n4356;
  assign n4358 = ~n3889 & n4351;
  assign n4359 = ~n3886 & n4358;
  assign n4360 = n3889 & ~n4351;
  assign n4361 = ~n3875 & n4360;
  assign n4362 = ~n4359 & ~n4361;
  assign n4363 = ~n3903 & ~n4362;
  assign n4364 = n3875 & n4351;
  assign n4365 = n3886 & ~n4351;
  assign n4366 = ~n3875 & n4365;
  assign n4367 = ~n4364 & ~n4366;
  assign n4368 = ~n4363 & n4367;
  assign n4369 = ~n4357 & n4368;
  assign n4370 = pi133 & pi263;
  assign n4371 = n3749 & ~n3766;
  assign n4372 = ~n3739 & n3740;
  assign n4373 = pi128 & pi268;
  assign n4374 = pi267 & ~n4373;
  assign n4375 = pi129 & n4374;
  assign n4376 = pi129 & pi267;
  assign n4377 = pi268 & ~n4376;
  assign n4378 = pi128 & n4377;
  assign n4379 = ~n4375 & ~n4378;
  assign n4380 = ~pi129 & n4379;
  assign n4381 = pi130 & pi266;
  assign n4382 = n4380 & n4381;
  assign n4383 = pi266 & ~n1328;
  assign n4384 = ~n4379 & ~n4383;
  assign n4385 = ~n4382 & ~n4384;
  assign n4386 = ~n4372 & ~n4385;
  assign n4387 = ~pi130 & ~n4379;
  assign n4388 = n4379 & n4381;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390 = ~n3740 & ~n4389;
  assign n4391 = n3739 & n4390;
  assign n4392 = ~pi129 & ~n3740;
  assign n4393 = pi130 & ~n4392;
  assign n4394 = ~n4379 & n4393;
  assign n4395 = n1319 & n4379;
  assign n4396 = ~n4394 & ~n4395;
  assign n4397 = pi266 & ~n4396;
  assign n4398 = n4379 & ~n4381;
  assign n4399 = n3740 & n4398;
  assign n4400 = ~n4397 & ~n4399;
  assign n4401 = ~n3739 & ~n4400;
  assign n4402 = pi130 & ~n4379;
  assign n4403 = ~pi130 & n4379;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = pi266 & ~n4404;
  assign n4406 = pi129 & n4405;
  assign n4407 = n3740 & n4406;
  assign n4408 = ~n4401 & ~n4407;
  assign n4409 = ~n4391 & n4408;
  assign n4410 = ~n4386 & n4409;
  assign n4411 = ~pi265 & ~n4410;
  assign n4412 = ~pi131 & ~n4410;
  assign n4413 = pi265 & n4410;
  assign n4414 = pi131 & n4413;
  assign n4415 = ~n4412 & ~n4414;
  assign n4416 = ~pi130 & ~n4415;
  assign n4417 = ~n4411 & ~n4416;
  assign n4418 = ~n4371 & ~n4417;
  assign n4419 = pi265 & n4371;
  assign n4420 = ~n3749 & ~n3766;
  assign n4421 = n3749 & n3766;
  assign n4422 = ~n4420 & ~n4421;
  assign n4423 = pi130 & ~n4422;
  assign n4424 = ~n4419 & ~n4423;
  assign n4425 = ~n4410 & ~n4424;
  assign n4426 = n3766 & n4410;
  assign n4427 = n3750 & n4426;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = pi131 & ~n4428;
  assign n4430 = ~n3749 & n3766;
  assign n4431 = pi265 & ~n4430;
  assign n4432 = pi130 & n4431;
  assign n4433 = ~n4371 & ~n4432;
  assign n4434 = n4410 & ~n4433;
  assign n4435 = n3766 & ~n4410;
  assign n4436 = ~n3749 & n4435;
  assign n4437 = ~n4434 & ~n4436;
  assign n4438 = ~pi131 & ~n4437;
  assign n4439 = ~pi265 & n3749;
  assign n4440 = ~n3766 & n4410;
  assign n4441 = n4439 & n4440;
  assign n4442 = ~n4438 & ~n4441;
  assign n4443 = ~n4429 & n4442;
  assign n4444 = ~n4418 & n4443;
  assign n4445 = ~n3769 & ~n3779;
  assign n4446 = n3769 & n3779;
  assign n4447 = ~n3790 & ~n4446;
  assign n4448 = ~n3778 & n4447;
  assign n4449 = ~n4445 & ~n4448;
  assign n4450 = n4444 & ~n4449;
  assign n4451 = ~n4444 & n4449;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = pi132 & pi264;
  assign n4454 = n3814 & ~n3819;
  assign n4455 = ~n3820 & ~n4454;
  assign n4456 = n4453 & ~n4455;
  assign n4457 = ~n3814 & ~n3820;
  assign n4458 = ~n3819 & ~n4457;
  assign n4459 = ~n4453 & ~n4458;
  assign n4460 = ~n4456 & ~n4459;
  assign n4461 = ~n4452 & ~n4460;
  assign n4462 = n4444 & n4449;
  assign n4463 = ~n4444 & ~n4449;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = ~n4453 & ~n4455;
  assign n4466 = n4453 & ~n4458;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = ~n4464 & ~n4467;
  assign n4469 = ~n4461 & ~n4468;
  assign n4470 = ~n4370 & n4469;
  assign n4471 = n4370 & ~n4469;
  assign n4472 = ~n4470 & ~n4471;
  assign n4473 = pi263 & ~n3821;
  assign n4474 = pi132 & n4473;
  assign n4475 = ~n3812 & ~n3814;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = pi262 & ~n4476;
  assign n4478 = pi133 & n4477;
  assign n4479 = pi134 & pi262;
  assign n4480 = ~n3813 & ~n4475;
  assign n4481 = ~n4474 & n4480;
  assign n4482 = ~n3830 & ~n4481;
  assign n4483 = ~n4479 & ~n4482;
  assign n4484 = ~n4478 & n4483;
  assign n4485 = ~n4478 & ~n4482;
  assign n4486 = n4479 & ~n4485;
  assign n4487 = ~n4484 & ~n4486;
  assign n4488 = ~n4472 & ~n4487;
  assign n4489 = ~n4370 & ~n4469;
  assign n4490 = n4370 & n4469;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = n4479 & ~n4482;
  assign n4493 = ~n4478 & n4492;
  assign n4494 = ~n4479 & ~n4485;
  assign n4495 = ~n4493 & ~n4494;
  assign n4496 = ~n4491 & ~n4495;
  assign n4497 = ~n4488 & ~n4496;
  assign n4498 = n3834 & ~n3859;
  assign n4499 = ~n3834 & n3859;
  assign n4500 = ~n3850 & ~n4499;
  assign n4501 = ~n4498 & ~n4500;
  assign n4502 = n4497 & n4501;
  assign n4503 = ~n4497 & ~n4501;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = pi135 & pi261;
  assign n4506 = n3889 & ~n3902;
  assign n4507 = ~n3901 & ~n4506;
  assign n4508 = n4505 & ~n4507;
  assign n4509 = ~n3889 & ~n3901;
  assign n4510 = ~n3902 & ~n4509;
  assign n4511 = ~n4505 & ~n4510;
  assign n4512 = ~n4508 & ~n4511;
  assign n4513 = ~n4504 & ~n4512;
  assign n4514 = n4497 & ~n4501;
  assign n4515 = ~n4497 & n4501;
  assign n4516 = ~n4514 & ~n4515;
  assign n4517 = ~n4505 & ~n4507;
  assign n4518 = n4505 & ~n4510;
  assign n4519 = ~n4517 & ~n4518;
  assign n4520 = ~n4516 & ~n4519;
  assign n4521 = ~n4513 & ~n4520;
  assign n4522 = ~n4369 & n4521;
  assign n4523 = n4369 & ~n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = ~n3886 & ~n3889;
  assign n4526 = ~n3875 & n4525;
  assign n4527 = ~n3887 & n3889;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = ~n3903 & ~n4528;
  assign n4530 = ~n3886 & n3889;
  assign n4531 = ~n3875 & n4530;
  assign n4532 = ~n3887 & ~n3889;
  assign n4533 = ~n4531 & ~n4532;
  assign n4534 = ~n3869 & ~n4533;
  assign n4535 = ~n4529 & ~n4534;
  assign n4536 = n3888 & ~n4535;
  assign n4537 = pi137 & pi259;
  assign n4538 = n4536 & n4537;
  assign n4539 = ~n4536 & ~n4537;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = pi258 & ~n4540;
  assign n4542 = pi138 & n4541;
  assign n4543 = pi138 & pi258;
  assign n4544 = ~n4536 & n4537;
  assign n4545 = n4536 & ~n4537;
  assign n4546 = ~n4544 & ~n4545;
  assign n4547 = ~n4543 & ~n4546;
  assign n4548 = ~n4542 & ~n4547;
  assign n4549 = ~n4524 & ~n4548;
  assign n4550 = n4369 & n4521;
  assign n4551 = ~n4369 & ~n4521;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = pi258 & ~n4546;
  assign n4554 = pi138 & n4553;
  assign n4555 = ~n4540 & ~n4543;
  assign n4556 = ~n4554 & ~n4555;
  assign n4557 = ~n4552 & ~n4556;
  assign n4558 = ~n4549 & ~n4557;
  assign n4559 = n4350 & ~n4558;
  assign n4560 = ~n4350 & n4558;
  assign n4561 = n3909 & n4560;
  assign n4562 = ~n4559 & ~n4561;
  assign n4563 = ~n3319 & ~n4562;
  assign n4564 = ~n4350 & ~n4558;
  assign n4565 = n4350 & n4558;
  assign n4566 = ~n3909 & n4565;
  assign n4567 = ~n4564 & ~n4566;
  assign n4568 = n3319 & ~n4567;
  assign n4569 = ~n3909 & ~n4350;
  assign n4570 = n3909 & n4350;
  assign n4571 = ~n4569 & ~n4570;
  assign n4572 = ~n4558 & ~n4571;
  assign n4573 = ~n4568 & ~n4572;
  assign n4574 = ~n4563 & n4573;
  assign n4575 = pi322 & ~n4574;
  assign n4576 = n3909 & ~n4350;
  assign n4577 = ~n3909 & n4350;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = n3319 & ~n4578;
  assign n4580 = ~n3319 & ~n4571;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = pi323 & ~n4581;
  assign n4583 = ~n4575 & ~n4582;
  assign n4584 = n3319 & n4576;
  assign n4585 = ~n4580 & ~n4584;
  assign n4586 = ~n4558 & ~n4585;
  assign n4587 = n3319 & ~n3909;
  assign n4588 = n4565 & n4587;
  assign n4589 = ~n4586 & ~n4588;
  assign n4590 = pi323 & ~n4589;
  assign n4591 = pi322 & n4590;
  assign n4592 = ~n4583 & ~n4591;
  assign n4593 = pi325 & n2887;
  assign n4594 = ~n3331 & ~n3929;
  assign n4595 = n3331 & ~n3922;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = pi324 & n4596;
  assign n4598 = n4593 & n4597;
  assign n4599 = ~n4593 & ~n4597;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = ~n4592 & ~n4600;
  assign n4602 = ~n4593 & n4597;
  assign n4603 = n4593 & ~n4597;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = ~n4591 & ~n4604;
  assign n4606 = ~n4583 & n4605;
  assign n4607 = ~n4601 & ~n4606;
  assign n4608 = ~n4348 & ~n4607;
  assign n4609 = ~n4337 & ~n4345;
  assign n4610 = n4337 & n4345;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n4592 & ~n4604;
  assign n4613 = ~n4591 & ~n4600;
  assign n4614 = ~n4583 & n4613;
  assign n4615 = ~n4612 & ~n4614;
  assign n4616 = ~n4611 & ~n4615;
  assign n4617 = ~n4608 & ~n4616;
  assign n4618 = n3944 & ~n3978;
  assign n4619 = ~n3942 & ~n3945;
  assign n4620 = ~n3934 & n4619;
  assign n4621 = n2887 & ~n3943;
  assign n4622 = pi324 & n4621;
  assign n4623 = ~n4620 & ~n4622;
  assign n4624 = ~n3959 & ~n4623;
  assign n4625 = ~n3943 & ~n3945;
  assign n4626 = n3943 & n3945;
  assign n4627 = ~n4625 & ~n4626;
  assign n4628 = ~n3733 & ~n4627;
  assign n4629 = ~n4624 & ~n4628;
  assign n4630 = ~n3944 & n3978;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n4618 & ~n4631;
  assign n4633 = n4617 & n4632;
  assign n4634 = ~n4617 & ~n4632;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = pi327 & n2091;
  assign n4637 = pi326 & n2464;
  assign n4638 = n4636 & n4637;
  assign n4639 = ~n4636 & ~n4637;
  assign n4640 = ~n4638 & ~n4639;
  assign n4641 = ~n4635 & ~n4640;
  assign n4642 = ~n4617 & n4632;
  assign n4643 = n4617 & ~n4632;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = ~n4636 & n4637;
  assign n4646 = n4636 & ~n4637;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = ~n4644 & ~n4647;
  assign n4649 = ~n4641 & ~n4648;
  assign n4650 = ~n4335 & ~n4649;
  assign n4651 = n4312 & ~n4332;
  assign n4652 = ~n4312 & n4332;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = ~n4640 & ~n4644;
  assign n4655 = ~n4635 & ~n4647;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = ~n4653 & ~n4656;
  assign n4658 = ~n4650 & ~n4657;
  assign n4659 = ~n4308 & n4658;
  assign n4660 = n4308 & ~n4658;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = n1729 & ~n4661;
  assign n4663 = pi328 & n4662;
  assign n4664 = pi328 & n1729;
  assign n4665 = n4308 & n4658;
  assign n4666 = ~n4308 & ~n4658;
  assign n4667 = ~n4665 & ~n4666;
  assign n4668 = ~n4664 & ~n4667;
  assign n4669 = ~n4663 & ~n4668;
  assign n4670 = ~n4307 & ~n4669;
  assign n4671 = n4292 & ~n4304;
  assign n4672 = ~n4292 & n4304;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = n1729 & ~n4667;
  assign n4675 = pi328 & n4674;
  assign n4676 = ~n4661 & ~n4664;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = ~n4673 & ~n4677;
  assign n4679 = ~n4670 & ~n4678;
  assign n4680 = ~n4287 & ~n4679;
  assign n4681 = n4287 & n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = pi258 & ~n4034;
  assign n4684 = pi128 & n4683;
  assign n4685 = pi331 & n4684;
  assign n4686 = pi331 & ~n1154;
  assign n4687 = ~n4685 & ~n4686;
  assign n4688 = ~n1154 & n4685;
  assign n4689 = pi331 & n4688;
  assign n4690 = ~n4687 & ~n4689;
  assign n4691 = ~n4682 & ~n4690;
  assign n4692 = n4287 & ~n4679;
  assign n4693 = ~n4287 & n4679;
  assign n4694 = ~n4692 & ~n4693;
  assign n4695 = n4685 & ~n4686;
  assign n4696 = ~n1154 & ~n4685;
  assign n4697 = pi331 & n4696;
  assign n4698 = ~n4695 & ~n4697;
  assign n4699 = ~n4694 & ~n4698;
  assign n4700 = ~n4691 & ~n4699;
  assign n4701 = pi332 & n1156;
  assign n4702 = n4700 & ~n4701;
  assign n4703 = pi332 & ~n4700;
  assign n4704 = n1156 & n4703;
  assign n4705 = ~n4702 & ~n4704;
  assign n4706 = ~n4276 & ~n4705;
  assign n4707 = n4276 & n4705;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = pi268 & ~n4708;
  assign n4710 = ~n4276 & n4705;
  assign n4711 = n4276 & ~n4705;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = ~pi268 & ~n4712;
  assign n4714 = ~n4709 & ~n4713;
  assign n4715 = n3672 & ~n4053;
  assign n4716 = ~n4054 & ~n4715;
  assign n4717 = n4714 & ~n4716;
  assign n4718 = ~n4714 & n4716;
  assign n4719 = ~n4717 & ~n4718;
  assign n4720 = ~n4274 & ~n4719;
  assign n4721 = n4714 & n4716;
  assign n4722 = ~n4714 & ~n4716;
  assign n4723 = ~n4721 & ~n4722;
  assign n4724 = n4274 & ~n4723;
  assign n4725 = ~n4720 & ~n4724;
  assign n4726 = ~n831 & ~n4725;
  assign n4727 = ~n4064 & ~n4726;
  assign n4728 = pi161 & ~n4727;
  assign n4729 = pi074 & ~pi161;
  assign n4730 = ~n4728 & ~n4729;
  assign po203 = ~pi160 & ~n4730;
  assign n4732 = pi269 & n831;
  assign n4733 = ~n4242 & ~n4253;
  assign n4734 = n4242 & n4253;
  assign n4735 = ~n1515 & ~n4734;
  assign n4736 = ~n4733 & ~n4735;
  assign n4737 = n1553 & ~n4736;
  assign n4738 = ~n1553 & ~n4733;
  assign n4739 = n1515 & n4738;
  assign n4740 = ~n4737 & ~n4739;
  assign n4741 = pi313 & ~n4740;
  assign n4742 = pi313 & n1553;
  assign n4743 = n4242 & ~n4742;
  assign n4744 = n4253 & n4743;
  assign n4745 = ~n4741 & ~n4744;
  assign n4746 = ~n1840 & n4171;
  assign n4747 = ~n4195 & ~n4746;
  assign n4748 = n1533 & n4747;
  assign n4749 = ~n4066 & n4171;
  assign n4750 = n1840 & ~n4749;
  assign n4751 = ~n4748 & ~n4750;
  assign n4752 = pi316 & ~n4751;
  assign n4753 = ~n4183 & ~n4752;
  assign n4754 = n1533 & ~n4219;
  assign n4755 = pi315 & n4754;
  assign n4756 = ~n4220 & ~n4755;
  assign n4757 = ~n4753 & ~n4756;
  assign n4758 = n4753 & n4756;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = ~pi139 & n4077;
  assign n4761 = pi139 & ~n4077;
  assign n4762 = ~pi138 & n4761;
  assign n4763 = ~n4760 & ~n4762;
  assign n4764 = pi137 & ~n4763;
  assign n4765 = ~pi139 & ~n4077;
  assign n4766 = pi139 & n4077;
  assign n4767 = pi138 & n4766;
  assign n4768 = ~n4765 & ~n4767;
  assign n4769 = ~pi137 & ~n4768;
  assign n4770 = ~pi139 & ~n4084;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4764 & n4771;
  assign n4773 = n4086 & ~n4098;
  assign n4774 = ~pi320 & ~n4773;
  assign n4775 = ~n3552 & ~n4086;
  assign n4776 = pi320 & n4773;
  assign n4777 = ~n4101 & ~n4776;
  assign n4778 = ~n4775 & n4777;
  assign n4779 = ~n4774 & n4778;
  assign n4780 = n4772 & ~n4779;
  assign n4781 = ~n4098 & ~n4772;
  assign n4782 = ~pi320 & n4086;
  assign n4783 = n4781 & n4782;
  assign n4784 = ~n4780 & ~n4783;
  assign n4785 = pi321 & ~n4784;
  assign n4786 = n4098 & ~n4772;
  assign n4787 = ~n3552 & n4786;
  assign n4788 = ~pi321 & ~n4106;
  assign n4789 = ~n4787 & ~n4788;
  assign n4790 = n4086 & ~n4789;
  assign n4791 = pi321 & n4772;
  assign n4792 = ~n4098 & ~n4791;
  assign n4793 = ~n4086 & n4792;
  assign n4794 = n3552 & n4793;
  assign n4795 = ~n4790 & ~n4794;
  assign n4796 = pi320 & ~n4795;
  assign n4797 = ~n4785 & ~n4796;
  assign n4798 = n3012 & ~n4116;
  assign n4799 = pi319 & n4798;
  assign n4800 = ~n4115 & ~n4799;
  assign n4801 = ~n4797 & ~n4800;
  assign n4802 = n4797 & n4800;
  assign n4803 = ~n4801 & ~n4802;
  assign n4804 = n3552 & ~n4803;
  assign n4805 = pi319 & n4804;
  assign n4806 = pi319 & n3552;
  assign n4807 = n4797 & ~n4800;
  assign n4808 = ~n4797 & n4800;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = ~n4806 & ~n4809;
  assign n4811 = ~n4805 & ~n4810;
  assign n4812 = n2574 & ~n4129;
  assign n4813 = pi318 & n4812;
  assign n4814 = ~n4130 & ~n4813;
  assign n4815 = n4811 & n4814;
  assign n4816 = ~n4811 & ~n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = n3012 & ~n4817;
  assign n4819 = pi318 & n4818;
  assign n4820 = pi318 & n3012;
  assign n4821 = ~n4811 & n4814;
  assign n4822 = n4811 & ~n4814;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = ~n4820 & ~n4823;
  assign n4825 = ~n4819 & ~n4824;
  assign n4826 = ~n2183 & n4139;
  assign n4827 = ~n3610 & ~n4826;
  assign n4828 = n1840 & n4827;
  assign n4829 = ~n3609 & n4139;
  assign n4830 = n2183 & ~n4829;
  assign n4831 = ~n4828 & ~n4830;
  assign n4832 = pi317 & ~n4831;
  assign n4833 = ~n4151 & ~n4832;
  assign n4834 = ~n4825 & ~n4833;
  assign n4835 = n4825 & n4833;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = n2574 & ~n4836;
  assign n4838 = pi317 & n4837;
  assign n4839 = pi317 & n2574;
  assign n4840 = n4825 & ~n4833;
  assign n4841 = ~n4825 & n4833;
  assign n4842 = ~n4840 & ~n4841;
  assign n4843 = ~n4839 & ~n4842;
  assign n4844 = ~n4838 & ~n4843;
  assign n4845 = pi316 & n2183;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = n2183 & n4844;
  assign n4848 = pi316 & n4847;
  assign n4849 = ~n4846 & ~n4848;
  assign n4850 = pi315 & n1840;
  assign n4851 = n4849 & ~n4850;
  assign n4852 = n1840 & ~n4849;
  assign n4853 = pi315 & n4852;
  assign n4854 = ~n4851 & ~n4853;
  assign n4855 = ~n4759 & ~n4854;
  assign n4856 = n4753 & ~n4756;
  assign n4857 = ~n4753 & n4756;
  assign n4858 = ~n4856 & ~n4857;
  assign n4859 = ~n4849 & ~n4850;
  assign n4860 = n1840 & n4849;
  assign n4861 = pi315 & n4860;
  assign n4862 = ~n4859 & ~n4861;
  assign n4863 = ~n4858 & ~n4862;
  assign n4864 = ~n4855 & ~n4863;
  assign n4865 = n1553 & ~n4239;
  assign n4866 = pi314 & n4865;
  assign n4867 = ~n4238 & ~n4866;
  assign n4868 = ~n4864 & ~n4867;
  assign n4869 = n4864 & n4867;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = n1533 & ~n4870;
  assign n4872 = pi314 & n4871;
  assign n4873 = pi314 & n1533;
  assign n4874 = n4864 & ~n4867;
  assign n4875 = ~n4864 & n4867;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = ~n4873 & ~n4876;
  assign n4878 = ~n4872 & ~n4877;
  assign n4879 = ~n4745 & ~n4878;
  assign n4880 = n4745 & n4878;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = pi312 & n1515;
  assign n4883 = n4881 & n4882;
  assign n4884 = ~n4881 & ~n4882;
  assign n4885 = ~n4883 & ~n4884;
  assign n4886 = n4065 & n4246;
  assign n4887 = ~n4065 & ~n4246;
  assign n4888 = ~n4242 & ~n4256;
  assign n4889 = ~n4255 & n4888;
  assign n4890 = n4242 & ~n4257;
  assign n4891 = ~n4889 & ~n4890;
  assign n4892 = ~n4887 & ~n4891;
  assign n4893 = ~n4886 & ~n4892;
  assign n4894 = ~n4885 & ~n4893;
  assign n4895 = n4885 & n4893;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = n4269 & n4272;
  assign n4898 = pi129 & n4897;
  assign n4899 = pi311 & ~n1568;
  assign n4900 = ~n4897 & n4899;
  assign n4901 = ~n4898 & ~n4900;
  assign n4902 = ~n4896 & ~n4901;
  assign n4903 = n4885 & ~n4893;
  assign n4904 = ~n4885 & n4893;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = ~pi129 & n4897;
  assign n4907 = ~n4897 & ~n4899;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = ~n4905 & ~n4908;
  assign n4910 = ~n4902 & ~n4909;
  assign n4911 = pi128 & pi310;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = pi310 & n4910;
  assign n4914 = pi128 & n4913;
  assign n4915 = ~n4912 & ~n4914;
  assign n4916 = ~pi268 & ~n4707;
  assign n4917 = ~n4706 & ~n4916;
  assign n4918 = n1156 & n4700;
  assign n4919 = ~n1154 & ~n4918;
  assign n4920 = n1154 & n4700;
  assign n4921 = n1156 & n4920;
  assign n4922 = ~n4919 & ~n4921;
  assign n4923 = pi332 & ~n4922;
  assign n4924 = ~n4292 & ~n4658;
  assign n4925 = n4292 & n4658;
  assign n4926 = n1729 & ~n4925;
  assign n4927 = pi328 & n4926;
  assign n4928 = ~n4924 & ~n4927;
  assign n4929 = ~n4304 & ~n4308;
  assign n4930 = n4304 & n4308;
  assign n4931 = ~n4292 & n4658;
  assign n4932 = n4292 & ~n4658;
  assign n4933 = ~n4931 & ~n4932;
  assign n4934 = n1729 & ~n4933;
  assign n4935 = pi328 & n4934;
  assign n4936 = ~n4924 & ~n4925;
  assign n4937 = ~n4664 & ~n4936;
  assign n4938 = ~n4935 & ~n4937;
  assign n4939 = ~n4930 & ~n4938;
  assign n4940 = ~n4929 & ~n4939;
  assign n4941 = n4928 & n4940;
  assign n4942 = ~n4928 & ~n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = pi328 & n2091;
  assign n4945 = ~n4312 & n4637;
  assign n4946 = n4312 & ~n4637;
  assign n4947 = ~n4644 & ~n4946;
  assign n4948 = ~n4945 & ~n4947;
  assign n4949 = ~n4312 & ~n4632;
  assign n4950 = n4312 & n4632;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = n4332 & n4636;
  assign n4953 = ~n4617 & n4637;
  assign n4954 = n4617 & ~n4637;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = ~n4952 & ~n4955;
  assign n4957 = ~n4951 & n4956;
  assign n4958 = ~n4312 & n4632;
  assign n4959 = n4312 & ~n4632;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = n4617 & n4637;
  assign n4962 = ~n4617 & ~n4637;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = ~n4952 & ~n4963;
  assign n4965 = ~n4960 & n4964;
  assign n4966 = ~n4332 & ~n4636;
  assign n4967 = ~n4965 & ~n4966;
  assign n4968 = ~n4957 & n4967;
  assign n4969 = n4948 & n4968;
  assign n4970 = ~n4948 & ~n4968;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = ~n4337 & ~n4583;
  assign n4973 = ~n4591 & ~n4972;
  assign n4974 = ~n4345 & n4597;
  assign n4975 = ~n4337 & ~n4592;
  assign n4976 = n4337 & ~n4591;
  assign n4977 = ~n4583 & n4976;
  assign n4978 = ~n4975 & ~n4977;
  assign n4979 = n4345 & ~n4597;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~n4974 & ~n4980;
  assign n4982 = ~n4973 & n4981;
  assign n4983 = n4973 & ~n4981;
  assign n4984 = ~n4982 & ~n4983;
  assign n4985 = ~n3319 & ~n4570;
  assign n4986 = ~n4569 & ~n4985;
  assign n4987 = n4558 & n4986;
  assign n4988 = ~n4558 & ~n4986;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = ~n3909 & ~n4989;
  assign n4991 = ~n4558 & n4986;
  assign n4992 = n4558 & ~n4986;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = n3909 & ~n4993;
  assign n4995 = ~n4990 & ~n4994;
  assign n4996 = pi323 & ~n4995;
  assign n4997 = pi139 & pi258;
  assign n4998 = ~n4558 & n4997;
  assign n4999 = n4558 & ~n4997;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = n4351 & n4521;
  assign n5002 = pi260 & ~n3869;
  assign n5003 = pi135 & n5002;
  assign n5004 = ~n3889 & ~n3903;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = ~n3886 & ~n5005;
  assign n5007 = ~n4351 & ~n4521;
  assign n5008 = ~n5006 & ~n5007;
  assign n5009 = ~n3875 & n5008;
  assign n5010 = ~n5001 & ~n5009;
  assign n5011 = ~n4539 & ~n4552;
  assign n5012 = ~n4538 & ~n5011;
  assign n5013 = ~n5010 & n5012;
  assign n5014 = n5010 & ~n5012;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = pi137 & pi260;
  assign n5017 = ~n3740 & ~n3743;
  assign n5018 = ~n3739 & ~n5017;
  assign n5019 = n3740 & n3743;
  assign n5020 = ~n5018 & ~n5019;
  assign n5021 = n4373 & ~n5020;
  assign n5022 = pi129 & pi268;
  assign n5023 = pi128 & pi269;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = pi268 & n1175;
  assign n5026 = pi269 & n5025;
  assign n5027 = ~n5024 & ~n5026;
  assign n5028 = ~pi267 & n5027;
  assign n5029 = ~pi130 & n5027;
  assign n5030 = pi267 & ~n5027;
  assign n5031 = pi130 & n5030;
  assign n5032 = ~n5029 & ~n5031;
  assign n5033 = ~pi129 & ~n5032;
  assign n5034 = ~n5028 & ~n5033;
  assign n5035 = ~n5021 & ~n5034;
  assign n5036 = n4373 & n5020;
  assign n5037 = ~n4373 & ~n5020;
  assign n5038 = ~n5036 & ~n5037;
  assign n5039 = pi129 & ~n5038;
  assign n5040 = pi267 & n5021;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n5027 & ~n5041;
  assign n5043 = pi267 & n5020;
  assign n5044 = ~n4373 & ~n5027;
  assign n5045 = n5043 & n5044;
  assign n5046 = ~n5042 & ~n5045;
  assign n5047 = pi130 & ~n5046;
  assign n5048 = ~n4373 & n5027;
  assign n5049 = n5020 & n5048;
  assign n5050 = ~n4373 & n5020;
  assign n5051 = pi267 & ~n5050;
  assign n5052 = pi129 & n5051;
  assign n5053 = ~n5021 & ~n5052;
  assign n5054 = ~n5027 & ~n5053;
  assign n5055 = ~n5049 & ~n5054;
  assign n5056 = ~pi130 & ~n5055;
  assign n5057 = n4373 & ~n5027;
  assign n5058 = ~pi267 & ~n5020;
  assign n5059 = n5057 & n5058;
  assign n5060 = ~n5056 & ~n5059;
  assign n5061 = ~n5047 & n5060;
  assign n5062 = ~n5035 & n5061;
  assign n5063 = ~n4379 & n5020;
  assign n5064 = n4379 & ~n5020;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = n4381 & ~n5065;
  assign n5067 = ~n4381 & n5065;
  assign n5068 = n3752 & ~n4430;
  assign n5069 = ~n4371 & ~n5068;
  assign n5070 = ~n5067 & ~n5069;
  assign n5071 = ~n5066 & ~n5070;
  assign n5072 = n5062 & n5071;
  assign n5073 = ~n5062 & ~n5071;
  assign n5074 = ~n5072 & ~n5073;
  assign n5075 = pi130 & ~n4430;
  assign n5076 = ~n4371 & ~n5075;
  assign n5077 = n4410 & ~n5076;
  assign n5078 = ~pi130 & ~n4371;
  assign n5079 = ~n4430 & ~n5078;
  assign n5080 = ~n4410 & ~n5079;
  assign n5081 = ~n5077 & ~n5080;
  assign n5082 = pi265 & ~n5081;
  assign n5083 = pi131 & n5082;
  assign n5084 = pi131 & pi266;
  assign n5085 = ~n4410 & ~n4433;
  assign n5086 = n4410 & ~n5079;
  assign n5087 = ~n5085 & ~n5086;
  assign n5088 = ~pi131 & ~n5087;
  assign n5089 = ~n3766 & ~n4410;
  assign n5090 = n3749 & n5089;
  assign n5091 = ~n4371 & n4410;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~pi265 & ~n5092;
  assign n5094 = ~n5088 & ~n5093;
  assign n5095 = n4449 & n5094;
  assign n5096 = ~n5084 & ~n5095;
  assign n5097 = ~n5083 & n5096;
  assign n5098 = ~n5083 & ~n5095;
  assign n5099 = n5084 & ~n5098;
  assign n5100 = ~n5097 & ~n5099;
  assign n5101 = ~n5074 & ~n5100;
  assign n5102 = n5062 & ~n5071;
  assign n5103 = ~n5062 & n5071;
  assign n5104 = ~n5102 & ~n5103;
  assign n5105 = n5084 & ~n5095;
  assign n5106 = ~n5083 & n5105;
  assign n5107 = ~n5084 & ~n5098;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = ~n5104 & ~n5108;
  assign n5110 = ~n5101 & ~n5109;
  assign n5111 = n4453 & ~n4464;
  assign n5112 = ~n4453 & n4464;
  assign n5113 = ~n4455 & ~n5112;
  assign n5114 = ~n5111 & ~n5113;
  assign n5115 = n5110 & n5114;
  assign n5116 = ~n5110 & ~n5114;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = pi133 & pi264;
  assign n5119 = pi132 & pi265;
  assign n5120 = n5118 & n5119;
  assign n5121 = ~n5118 & ~n5119;
  assign n5122 = ~n5120 & ~n5121;
  assign n5123 = ~n5117 & ~n5122;
  assign n5124 = ~n5110 & n5114;
  assign n5125 = n5110 & ~n5114;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = pi264 & ~n5119;
  assign n5128 = pi133 & n5127;
  assign n5129 = pi265 & ~n5118;
  assign n5130 = pi132 & n5129;
  assign n5131 = ~n5128 & ~n5130;
  assign n5132 = ~n5126 & ~n5131;
  assign n5133 = ~n5123 & ~n5132;
  assign n5134 = ~n4485 & ~n4489;
  assign n5135 = ~n4490 & ~n5134;
  assign n5136 = n5133 & n5135;
  assign n5137 = ~n5133 & ~n5135;
  assign n5138 = ~n5136 & ~n5137;
  assign n5139 = pi134 & pi263;
  assign n5140 = n4469 & ~n4482;
  assign n5141 = ~n4478 & n5140;
  assign n5142 = ~n4469 & ~n4485;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = ~n4370 & ~n5143;
  assign n5145 = ~n4469 & ~n4482;
  assign n5146 = ~n4478 & n5145;
  assign n5147 = n4469 & ~n4485;
  assign n5148 = ~n5146 & ~n5147;
  assign n5149 = pi263 & ~n5148;
  assign n5150 = pi133 & n5149;
  assign n5151 = ~n5144 & ~n5150;
  assign n5152 = ~n4501 & ~n5151;
  assign n5153 = n4501 & n5151;
  assign n5154 = n4479 & ~n5153;
  assign n5155 = ~n5152 & ~n5154;
  assign n5156 = n5139 & ~n5155;
  assign n5157 = ~n4479 & ~n5152;
  assign n5158 = ~n5153 & ~n5157;
  assign n5159 = ~n5139 & ~n5158;
  assign n5160 = ~n5156 & ~n5159;
  assign n5161 = ~n5138 & ~n5160;
  assign n5162 = n5133 & ~n5135;
  assign n5163 = ~n5133 & n5135;
  assign n5164 = ~n5162 & ~n5163;
  assign n5165 = ~n5139 & ~n5155;
  assign n5166 = n5139 & ~n5158;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = ~n5164 & ~n5167;
  assign n5169 = ~n5161 & ~n5168;
  assign n5170 = ~n4504 & ~n4505;
  assign n5171 = n4504 & n4505;
  assign n5172 = ~n4510 & ~n5171;
  assign n5173 = ~n5170 & ~n5172;
  assign n5174 = ~n5169 & n5173;
  assign n5175 = n5169 & ~n5173;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = pi136 & pi261;
  assign n5178 = pi135 & pi262;
  assign n5179 = n5177 & n5178;
  assign n5180 = ~n5177 & ~n5178;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = ~n5176 & ~n5181;
  assign n5183 = n5169 & n5173;
  assign n5184 = ~n5169 & ~n5173;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = pi261 & ~n5178;
  assign n5187 = pi136 & n5186;
  assign n5188 = pi262 & ~n5177;
  assign n5189 = pi135 & n5188;
  assign n5190 = ~n5187 & ~n5189;
  assign n5191 = ~n5185 & ~n5190;
  assign n5192 = ~n5182 & ~n5191;
  assign n5193 = ~n5016 & n5192;
  assign n5194 = n5016 & ~n5192;
  assign n5195 = ~n5193 & ~n5194;
  assign n5196 = pi138 & pi259;
  assign n5197 = ~n4524 & ~n4540;
  assign n5198 = ~n4546 & ~n4552;
  assign n5199 = n4543 & ~n5198;
  assign n5200 = ~n5197 & n5199;
  assign n5201 = ~n5196 & ~n5200;
  assign n5202 = pi137 & n4536;
  assign n5203 = ~pi137 & ~n4536;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n4552 & ~n5204;
  assign n5206 = pi137 & ~n4536;
  assign n5207 = ~pi137 & n4536;
  assign n5208 = ~n5206 & ~n5207;
  assign n5209 = ~n4524 & ~n5208;
  assign n5210 = ~n5205 & ~n5209;
  assign n5211 = n4543 & ~n5210;
  assign n5212 = pi259 & n5211;
  assign n5213 = ~n5201 & ~n5212;
  assign n5214 = ~n5195 & ~n5213;
  assign n5215 = n5016 & n5192;
  assign n5216 = ~n5016 & ~n5192;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5212 & ~n5217;
  assign n5219 = ~n5201 & n5218;
  assign n5220 = ~n5214 & ~n5219;
  assign n5221 = ~n5015 & ~n5220;
  assign n5222 = ~n5010 & ~n5012;
  assign n5223 = n5010 & n5012;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5213 & ~n5217;
  assign n5226 = ~n5195 & ~n5212;
  assign n5227 = ~n5201 & n5226;
  assign n5228 = ~n5225 & ~n5227;
  assign n5229 = ~n5224 & ~n5228;
  assign n5230 = ~n5221 & ~n5229;
  assign n5231 = ~n3909 & ~n4987;
  assign n5232 = ~n4988 & ~n5231;
  assign n5233 = n5230 & n5232;
  assign n5234 = ~n5230 & ~n5232;
  assign n5235 = ~n5233 & ~n5234;
  assign n5236 = ~n5000 & ~n5235;
  assign n5237 = n5230 & ~n5232;
  assign n5238 = ~n5230 & n5232;
  assign n5239 = ~n5237 & ~n5238;
  assign n5240 = n4558 & n4997;
  assign n5241 = ~n4558 & ~n4997;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~n5239 & ~n5242;
  assign n5244 = pi322 & ~n5243;
  assign n5245 = ~n5236 & n5244;
  assign n5246 = ~n4996 & ~n5245;
  assign n5247 = pi322 & ~n4995;
  assign n5248 = ~n5000 & ~n5239;
  assign n5249 = ~n5235 & ~n5242;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = n5247 & ~n5250;
  assign n5252 = pi323 & n5251;
  assign n5253 = ~n5246 & ~n5252;
  assign n5254 = pi325 & n4596;
  assign n5255 = ~n3319 & ~n4578;
  assign n5256 = n3319 & ~n4571;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = pi324 & n5257;
  assign n5259 = n5254 & n5258;
  assign n5260 = ~n5254 & ~n5258;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~n5253 & ~n5261;
  assign n5263 = ~n5254 & n5258;
  assign n5264 = n5254 & ~n5258;
  assign n5265 = ~n5263 & ~n5264;
  assign n5266 = ~n5252 & ~n5265;
  assign n5267 = ~n5246 & n5266;
  assign n5268 = ~n5262 & ~n5267;
  assign n5269 = ~n4984 & ~n5268;
  assign n5270 = ~n4973 & ~n4981;
  assign n5271 = n4973 & n4981;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = ~n5253 & ~n5265;
  assign n5274 = ~n5252 & ~n5261;
  assign n5275 = ~n5246 & n5274;
  assign n5276 = ~n5273 & ~n5275;
  assign n5277 = ~n5272 & ~n5276;
  assign n5278 = ~n5269 & ~n5277;
  assign n5279 = n4593 & ~n4632;
  assign n5280 = ~n4597 & ~n4978;
  assign n5281 = n4337 & ~n4592;
  assign n5282 = ~n4337 & ~n4591;
  assign n5283 = ~n4583 & n5282;
  assign n5284 = ~n5281 & ~n5283;
  assign n5285 = n4596 & ~n5284;
  assign n5286 = pi324 & n5285;
  assign n5287 = ~n5280 & ~n5286;
  assign n5288 = n4345 & ~n5287;
  assign n5289 = ~n4345 & n5287;
  assign n5290 = ~n5288 & ~n5289;
  assign n5291 = ~n4593 & n4632;
  assign n5292 = ~n5290 & ~n5291;
  assign n5293 = ~n5279 & ~n5292;
  assign n5294 = n5278 & n5293;
  assign n5295 = ~n5278 & ~n5293;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = pi327 & n2464;
  assign n5298 = pi326 & n2887;
  assign n5299 = n5297 & n5298;
  assign n5300 = ~n5297 & ~n5298;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~n5296 & ~n5301;
  assign n5303 = ~n5278 & n5293;
  assign n5304 = n5278 & ~n5293;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5297 & n5298;
  assign n5307 = n5297 & ~n5298;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = ~n5305 & ~n5308;
  assign n5310 = ~n5302 & ~n5309;
  assign n5311 = ~n4971 & ~n5310;
  assign n5312 = n4948 & ~n4968;
  assign n5313 = ~n4948 & n4968;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = ~n5301 & ~n5305;
  assign n5316 = ~n5296 & ~n5308;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = ~n5314 & ~n5317;
  assign n5319 = ~n5311 & ~n5318;
  assign n5320 = ~n4944 & n5319;
  assign n5321 = n4944 & ~n5319;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = n1729 & ~n5322;
  assign n5324 = pi329 & n5323;
  assign n5325 = pi329 & n1729;
  assign n5326 = n4944 & n5319;
  assign n5327 = ~n4944 & ~n5319;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = ~n5325 & ~n5328;
  assign n5330 = ~n5324 & ~n5329;
  assign n5331 = ~n4943 & ~n5330;
  assign n5332 = n4928 & ~n4940;
  assign n5333 = ~n4928 & n4940;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = n1729 & ~n5328;
  assign n5336 = pi329 & n5335;
  assign n5337 = ~n5322 & ~n5325;
  assign n5338 = ~n5336 & ~n5337;
  assign n5339 = ~n5334 & ~n5338;
  assign n5340 = ~n5331 & ~n5339;
  assign n5341 = ~n4687 & ~n4694;
  assign n5342 = ~n4689 & ~n5341;
  assign n5343 = n5340 & n5342;
  assign n5344 = ~n5340 & ~n5342;
  assign n5345 = ~n5343 & ~n5344;
  assign n5346 = ~n3675 & ~n4025;
  assign n5347 = ~n1154 & ~n5346;
  assign n5348 = n3477 & n4025;
  assign n5349 = n1156 & n5348;
  assign n5350 = ~n5347 & ~n5349;
  assign n5351 = pi330 & ~n5350;
  assign n5352 = n4679 & n5351;
  assign n5353 = ~n4679 & ~n5351;
  assign n5354 = ~n1256 & ~n5353;
  assign n5355 = ~n5352 & ~n5354;
  assign n5356 = n1442 & ~n5355;
  assign n5357 = pi330 & n5356;
  assign n5358 = ~n1442 & ~n5354;
  assign n5359 = pi330 & ~n5358;
  assign n5360 = ~n5352 & ~n5359;
  assign n5361 = ~n5357 & ~n5360;
  assign n5362 = ~n1256 & ~n5361;
  assign n5363 = pi331 & n5362;
  assign n5364 = pi331 & ~n1256;
  assign n5365 = ~n5360 & ~n5364;
  assign n5366 = ~n5357 & n5365;
  assign n5367 = ~n5363 & ~n5366;
  assign n5368 = ~n5345 & ~n5367;
  assign n5369 = n5340 & ~n5342;
  assign n5370 = ~n5340 & n5342;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = ~n5361 & ~n5364;
  assign n5373 = n5361 & n5364;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n5371 & ~n5374;
  assign n5376 = ~n5368 & ~n5375;
  assign n5377 = n4923 & n5376;
  assign n5378 = ~n4923 & ~n5376;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = pi258 & ~n5379;
  assign n5381 = pi128 & n5380;
  assign n5382 = pi333 & n5381;
  assign n5383 = n4923 & ~n5376;
  assign n5384 = ~n4923 & n5376;
  assign n5385 = ~n5383 & ~n5384;
  assign n5386 = pi333 & n1156;
  assign n5387 = ~n5385 & ~n5386;
  assign n5388 = ~n5382 & ~n5387;
  assign n5389 = ~n4917 & ~n5388;
  assign n5390 = n4917 & n5388;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = pi269 & ~n5391;
  assign n5393 = ~n4917 & n5388;
  assign n5394 = n4917 & ~n5388;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~pi269 & ~n5395;
  assign n5397 = ~n5392 & ~n5396;
  assign n5398 = n4274 & ~n4721;
  assign n5399 = ~n4722 & ~n5398;
  assign n5400 = n5397 & ~n5399;
  assign n5401 = ~n5397 & n5399;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~n4915 & ~n5402;
  assign n5404 = n5397 & n5399;
  assign n5405 = ~n5397 & ~n5399;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = n4915 & ~n5406;
  assign n5408 = ~n5403 & ~n5407;
  assign n5409 = ~n831 & ~n5408;
  assign n5410 = ~n4732 & ~n5409;
  assign n5411 = pi161 & ~n5410;
  assign n5412 = pi075 & ~pi161;
  assign n5413 = ~n5411 & ~n5412;
  assign po204 = ~pi160 & ~n5413;
  assign n5415 = pi270 & n831;
  assign n5416 = ~n4905 & ~n4907;
  assign n5417 = ~n4906 & ~n5416;
  assign n5418 = pi311 & n1515;
  assign n5419 = n5417 & n5418;
  assign n5420 = ~n5417 & ~n5418;
  assign n5421 = ~n5419 & ~n5420;
  assign n5422 = n4242 & n4878;
  assign n5423 = n4253 & n5422;
  assign n5424 = ~n1553 & ~n4878;
  assign n5425 = ~n4733 & ~n5424;
  assign n5426 = n1515 & n5425;
  assign n5427 = ~n4734 & ~n4878;
  assign n5428 = n1553 & ~n5427;
  assign n5429 = ~n5426 & ~n5428;
  assign n5430 = pi313 & ~n5429;
  assign n5431 = ~n5423 & ~n5430;
  assign n5432 = pi313 & n1533;
  assign n5433 = n5431 & n5432;
  assign n5434 = ~n5431 & ~n5432;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = n1533 & ~n4875;
  assign n5437 = pi314 & n5436;
  assign n5438 = ~n4874 & ~n5437;
  assign n5439 = ~pi140 & ~n4077;
  assign n5440 = pi139 & n5439;
  assign n5441 = ~pi139 & pi140;
  assign n5442 = pi138 & n5441;
  assign n5443 = ~n5440 & ~n5442;
  assign n5444 = pi137 & ~n5443;
  assign n5445 = pi139 & pi140;
  assign n5446 = ~pi138 & n5445;
  assign n5447 = ~pi140 & n4077;
  assign n5448 = ~pi139 & n5447;
  assign n5449 = ~n5446 & ~n5448;
  assign n5450 = ~pi137 & ~n5449;
  assign n5451 = pi139 & ~pi140;
  assign n5452 = pi140 & ~n4077;
  assign n5453 = ~pi139 & n5452;
  assign n5454 = ~n5451 & ~n5453;
  assign n5455 = pi138 & ~n5454;
  assign n5456 = ~pi139 & ~pi140;
  assign n5457 = pi140 & n4077;
  assign n5458 = pi139 & n5457;
  assign n5459 = ~n5456 & ~n5458;
  assign n5460 = ~pi138 & ~n5459;
  assign n5461 = ~n5455 & ~n5460;
  assign n5462 = ~n5450 & n5461;
  assign n5463 = ~n5444 & n5462;
  assign n5464 = pi321 & n5463;
  assign n5465 = ~n4098 & n4772;
  assign n5466 = ~n4086 & ~n5465;
  assign n5467 = n3552 & ~n5466;
  assign n5468 = n4086 & ~n4786;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = pi321 & ~n5469;
  assign n5471 = n3552 & n4773;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = pi320 & ~n5472;
  assign n5474 = n4087 & n5465;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = pi320 & n4772;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = n4772 & n5475;
  assign n5479 = pi320 & n5478;
  assign n5480 = ~n5477 & ~n5479;
  assign n5481 = ~n5464 & ~n5480;
  assign n5482 = n5475 & ~n5476;
  assign n5483 = n4772 & ~n5475;
  assign n5484 = pi320 & n5483;
  assign n5485 = ~n5482 & ~n5484;
  assign n5486 = n5463 & ~n5485;
  assign n5487 = pi321 & n5486;
  assign n5488 = ~n5481 & ~n5487;
  assign n5489 = n3552 & ~n4802;
  assign n5490 = pi319 & n5489;
  assign n5491 = ~n4801 & ~n5490;
  assign n5492 = ~n5488 & ~n5491;
  assign n5493 = n5488 & n5491;
  assign n5494 = ~n5492 & ~n5493;
  assign n5495 = n4086 & ~n5494;
  assign n5496 = pi319 & n5495;
  assign n5497 = pi319 & n4086;
  assign n5498 = n5488 & ~n5491;
  assign n5499 = ~n5488 & n5491;
  assign n5500 = ~n5498 & ~n5499;
  assign n5501 = ~n5497 & ~n5500;
  assign n5502 = ~n5496 & ~n5501;
  assign n5503 = n3012 & ~n4815;
  assign n5504 = pi318 & n5503;
  assign n5505 = ~n4816 & ~n5504;
  assign n5506 = n5502 & n5505;
  assign n5507 = ~n5502 & ~n5505;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = n3552 & ~n5508;
  assign n5510 = pi318 & n5509;
  assign n5511 = pi318 & n3552;
  assign n5512 = ~n5502 & n5505;
  assign n5513 = n5502 & ~n5505;
  assign n5514 = ~n5512 & ~n5513;
  assign n5515 = ~n5511 & ~n5514;
  assign n5516 = ~n5510 & ~n5515;
  assign n5517 = n2574 & ~n4835;
  assign n5518 = pi317 & n5517;
  assign n5519 = ~n4834 & ~n5518;
  assign n5520 = ~n5516 & ~n5519;
  assign n5521 = n5516 & n5519;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = n3012 & ~n5522;
  assign n5524 = pi317 & n5523;
  assign n5525 = pi317 & n3012;
  assign n5526 = n5516 & ~n5519;
  assign n5527 = ~n5516 & n5519;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = ~n5525 & ~n5528;
  assign n5530 = ~n5524 & ~n5529;
  assign n5531 = ~n4753 & ~n4844;
  assign n5532 = n4753 & n4844;
  assign n5533 = n2183 & ~n5532;
  assign n5534 = pi316 & n5533;
  assign n5535 = ~n5531 & ~n5534;
  assign n5536 = ~n5530 & ~n5535;
  assign n5537 = n5530 & n5535;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = n2574 & ~n5538;
  assign n5540 = pi316 & n5539;
  assign n5541 = pi316 & n2574;
  assign n5542 = n5530 & ~n5535;
  assign n5543 = ~n5530 & n5535;
  assign n5544 = ~n5542 & ~n5543;
  assign n5545 = ~n5541 & ~n5544;
  assign n5546 = ~n5540 & ~n5545;
  assign n5547 = pi315 & n2183;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = n2183 & n5546;
  assign n5550 = pi315 & n5549;
  assign n5551 = ~n5548 & ~n5550;
  assign n5552 = ~n4753 & n4849;
  assign n5553 = n4753 & ~n4849;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = n4756 & ~n4850;
  assign n5556 = ~n5554 & ~n5555;
  assign n5557 = n1840 & ~n4756;
  assign n5558 = pi315 & n5557;
  assign n5559 = ~n5556 & ~n5558;
  assign n5560 = ~n5551 & n5559;
  assign n5561 = n5551 & ~n5559;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = n1840 & ~n5562;
  assign n5564 = pi314 & n5563;
  assign n5565 = pi314 & n1840;
  assign n5566 = ~n5561 & ~n5565;
  assign n5567 = ~n5560 & n5566;
  assign n5568 = ~n5564 & ~n5567;
  assign n5569 = n5438 & ~n5568;
  assign n5570 = ~n5438 & ~n5567;
  assign n5571 = ~n5564 & n5570;
  assign n5572 = ~n5569 & ~n5571;
  assign n5573 = n5435 & ~n5572;
  assign n5574 = ~n5435 & n5572;
  assign n5575 = ~n5573 & ~n5574;
  assign n5576 = pi312 & n1553;
  assign n5577 = ~n4881 & ~n4893;
  assign n5578 = n4881 & n4893;
  assign n5579 = n4882 & ~n5578;
  assign n5580 = ~n5577 & ~n5579;
  assign n5581 = n5576 & ~n5580;
  assign n5582 = ~n4882 & ~n5577;
  assign n5583 = ~n5578 & ~n5582;
  assign n5584 = ~n5576 & ~n5583;
  assign n5585 = ~n5581 & ~n5584;
  assign n5586 = ~n5575 & ~n5585;
  assign n5587 = n5435 & n5572;
  assign n5588 = ~n5435 & ~n5572;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = ~n5576 & ~n5580;
  assign n5591 = n5576 & ~n5583;
  assign n5592 = ~n5590 & ~n5591;
  assign n5593 = ~n5589 & ~n5592;
  assign n5594 = ~n5586 & ~n5593;
  assign n5595 = n5421 & ~n5594;
  assign n5596 = ~n5421 & n5594;
  assign n5597 = ~n5595 & ~n5596;
  assign n5598 = pi128 & n4910;
  assign n5599 = ~pi129 & ~n5598;
  assign n5600 = pi129 & n4910;
  assign n5601 = pi128 & n5600;
  assign n5602 = pi310 & ~n5601;
  assign n5603 = ~n5599 & n5602;
  assign n5604 = ~n5597 & ~n5603;
  assign n5605 = n5421 & n5594;
  assign n5606 = ~n5421 & ~n5594;
  assign n5607 = ~n5605 & ~n5606;
  assign n5608 = pi129 & ~n5598;
  assign n5609 = ~pi129 & n4910;
  assign n5610 = pi128 & n5609;
  assign n5611 = ~n5608 & ~n5610;
  assign n5612 = ~n5607 & ~n5611;
  assign n5613 = pi310 & n5612;
  assign n5614 = ~n5604 & ~n5613;
  assign n5615 = pi309 & ~n5614;
  assign n5616 = pi128 & n5615;
  assign n5617 = pi128 & pi309;
  assign n5618 = n5614 & ~n5617;
  assign n5619 = ~n5616 & ~n5618;
  assign n5620 = ~pi269 & ~n5390;
  assign n5621 = ~n5389 & ~n5620;
  assign n5622 = pi258 & ~n5385;
  assign n5623 = pi128 & n5622;
  assign n5624 = pi333 & n5623;
  assign n5625 = ~n4928 & n5319;
  assign n5626 = n4928 & ~n5319;
  assign n5627 = ~n5625 & ~n5626;
  assign n5628 = ~n4944 & ~n5627;
  assign n5629 = ~n4928 & ~n5319;
  assign n5630 = n4928 & n5319;
  assign n5631 = ~n5629 & ~n5630;
  assign n5632 = n4944 & ~n5631;
  assign n5633 = ~n5628 & ~n5632;
  assign n5634 = ~n4940 & ~n5325;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = n1729 & n4940;
  assign n5637 = pi329 & n5636;
  assign n5638 = ~n5635 & ~n5637;
  assign n5639 = ~n1256 & ~n5342;
  assign n5640 = pi331 & n5639;
  assign n5641 = n5342 & ~n5364;
  assign n5642 = ~n5340 & ~n5360;
  assign n5643 = ~n5357 & n5642;
  assign n5644 = n5340 & ~n5361;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = ~n5641 & ~n5645;
  assign n5647 = ~n5640 & ~n5646;
  assign n5648 = ~n5638 & n5647;
  assign n5649 = n5638 & ~n5647;
  assign n5650 = ~n5648 & ~n5649;
  assign n5651 = n5340 & ~n5360;
  assign n5652 = ~n5357 & ~n5651;
  assign n5653 = n1729 & n5652;
  assign n5654 = pi330 & n5653;
  assign n5655 = pi330 & n1729;
  assign n5656 = ~n5652 & ~n5655;
  assign n5657 = ~n5654 & ~n5656;
  assign n5658 = ~n4948 & ~n5293;
  assign n5659 = n4948 & n5293;
  assign n5660 = ~n5658 & ~n5659;
  assign n5661 = n4968 & n5297;
  assign n5662 = ~n5278 & n5298;
  assign n5663 = n5278 & ~n5298;
  assign n5664 = ~n5662 & ~n5663;
  assign n5665 = ~n5661 & ~n5664;
  assign n5666 = ~n5660 & n5665;
  assign n5667 = ~n4948 & n5293;
  assign n5668 = n4948 & ~n5293;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = n5278 & n5298;
  assign n5671 = ~n5278 & ~n5298;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = ~n5661 & ~n5672;
  assign n5674 = ~n5669 & n5673;
  assign n5675 = ~n4968 & ~n5297;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~n5666 & n5676;
  assign n5678 = ~n4928 & n4944;
  assign n5679 = n4928 & ~n4944;
  assign n5680 = ~n5319 & ~n5679;
  assign n5681 = ~n5678 & ~n5680;
  assign n5682 = n5677 & ~n5681;
  assign n5683 = ~n5677 & n5681;
  assign n5684 = ~n5682 & ~n5683;
  assign n5685 = pi327 & n2887;
  assign n5686 = n5254 & ~n5293;
  assign n5687 = ~n4973 & ~n5253;
  assign n5688 = n4973 & ~n5252;
  assign n5689 = ~n5246 & n5688;
  assign n5690 = ~n5687 & ~n5689;
  assign n5691 = ~n5258 & ~n5690;
  assign n5692 = n4973 & ~n5253;
  assign n5693 = ~n4973 & ~n5252;
  assign n5694 = ~n5246 & n5693;
  assign n5695 = ~n5692 & ~n5694;
  assign n5696 = n5257 & ~n5695;
  assign n5697 = pi324 & n5696;
  assign n5698 = ~n5691 & ~n5697;
  assign n5699 = n4981 & ~n5698;
  assign n5700 = ~n4981 & n5698;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = ~n5254 & n5293;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = ~n5686 & ~n5703;
  assign n5705 = ~n4948 & n5298;
  assign n5706 = n4948 & ~n5298;
  assign n5707 = ~n5305 & ~n5706;
  assign n5708 = ~n5705 & ~n5707;
  assign n5709 = n5704 & ~n5708;
  assign n5710 = ~n5704 & n5708;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = ~n3909 & ~n4993;
  assign n5713 = n3909 & ~n4989;
  assign n5714 = ~n5712 & ~n5713;
  assign n5715 = pi324 & n5714;
  assign n5716 = ~n4973 & ~n5246;
  assign n5717 = ~n5252 & ~n5716;
  assign n5718 = ~n5715 & ~n5717;
  assign n5719 = n5715 & n5717;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = n4997 & n5230;
  assign n5722 = ~n4997 & ~n5230;
  assign n5723 = ~n5721 & ~n5722;
  assign n5724 = n5232 & ~n5723;
  assign n5725 = ~n5232 & n5723;
  assign n5726 = ~n5724 & ~n5725;
  assign n5727 = ~n4558 & ~n5726;
  assign n5728 = ~n5232 & ~n5723;
  assign n5729 = n5232 & n5723;
  assign n5730 = ~n5728 & ~n5729;
  assign n5731 = n4558 & ~n5730;
  assign n5732 = ~n5727 & ~n5731;
  assign n5733 = pi323 & n5732;
  assign n5734 = ~n5012 & n5016;
  assign n5735 = n5012 & ~n5016;
  assign n5736 = pi262 & ~n5185;
  assign n5737 = pi135 & n5736;
  assign n5738 = ~n5176 & ~n5178;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = pi261 & ~n5739;
  assign n5741 = pi136 & n5740;
  assign n5742 = ~n5177 & ~n5738;
  assign n5743 = ~n5737 & n5742;
  assign n5744 = ~n5741 & ~n5743;
  assign n5745 = ~n5010 & ~n5744;
  assign n5746 = n5010 & n5744;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~n5735 & ~n5747;
  assign n5749 = ~n5734 & ~n5748;
  assign n5750 = ~n5015 & ~n5195;
  assign n5751 = ~n5217 & ~n5224;
  assign n5752 = ~n5212 & ~n5751;
  assign n5753 = ~n5750 & n5752;
  assign n5754 = ~n5201 & ~n5753;
  assign n5755 = n5749 & ~n5754;
  assign n5756 = ~n5749 & n5754;
  assign n5757 = ~n5755 & ~n5756;
  assign n5758 = pi137 & pi261;
  assign n5759 = pi133 & pi265;
  assign n5760 = n4373 & n4376;
  assign n5761 = ~n4373 & ~n4376;
  assign n5762 = ~n5020 & ~n5761;
  assign n5763 = ~n5760 & ~n5762;
  assign n5764 = n5027 & ~n5763;
  assign n5765 = ~n4376 & ~n5021;
  assign n5766 = ~n5050 & ~n5765;
  assign n5767 = ~n5027 & ~n5766;
  assign n5768 = ~n5764 & ~n5767;
  assign n5769 = ~n5071 & n5768;
  assign n5770 = n3739 & ~n5019;
  assign n5771 = ~n5017 & ~n5770;
  assign n5772 = ~n5760 & ~n5771;
  assign n5773 = ~n5761 & ~n5772;
  assign n5774 = ~n5026 & ~n5773;
  assign n5775 = ~n5024 & ~n5774;
  assign n5776 = pi128 & pi270;
  assign n5777 = pi269 & ~n5776;
  assign n5778 = pi129 & n5777;
  assign n5779 = pi129 & pi269;
  assign n5780 = pi270 & ~n5779;
  assign n5781 = pi128 & n5780;
  assign n5782 = ~n5778 & ~n5781;
  assign n5783 = pi130 & pi268;
  assign n5784 = ~n5782 & ~n5783;
  assign n5785 = pi268 & n5782;
  assign n5786 = pi130 & n5785;
  assign n5787 = ~n5784 & ~n5786;
  assign n5788 = ~n5775 & ~n5787;
  assign n5789 = n5782 & ~n5783;
  assign n5790 = pi268 & ~n5782;
  assign n5791 = pi130 & n5790;
  assign n5792 = ~n5789 & ~n5791;
  assign n5793 = ~n5774 & ~n5792;
  assign n5794 = ~n5024 & n5793;
  assign n5795 = ~n5788 & ~n5794;
  assign n5796 = ~pi267 & ~n5795;
  assign n5797 = ~pi131 & ~n5795;
  assign n5798 = pi267 & n5795;
  assign n5799 = pi131 & n5798;
  assign n5800 = ~n5797 & ~n5799;
  assign n5801 = ~pi130 & ~n5800;
  assign n5802 = ~n5796 & ~n5801;
  assign n5803 = ~n5769 & ~n5802;
  assign n5804 = pi267 & n5769;
  assign n5805 = ~n5071 & ~n5768;
  assign n5806 = n5071 & n5768;
  assign n5807 = ~n5805 & ~n5806;
  assign n5808 = pi130 & ~n5807;
  assign n5809 = ~n5804 & ~n5808;
  assign n5810 = ~n5795 & ~n5809;
  assign n5811 = n5071 & n5795;
  assign n5812 = pi267 & ~n5768;
  assign n5813 = n5811 & n5812;
  assign n5814 = ~n5810 & ~n5813;
  assign n5815 = pi131 & ~n5814;
  assign n5816 = n5071 & ~n5768;
  assign n5817 = pi267 & ~n5816;
  assign n5818 = pi130 & n5817;
  assign n5819 = ~n5769 & ~n5818;
  assign n5820 = n5795 & ~n5819;
  assign n5821 = n5071 & ~n5795;
  assign n5822 = ~n5768 & n5821;
  assign n5823 = ~n5820 & ~n5822;
  assign n5824 = ~pi131 & ~n5823;
  assign n5825 = ~pi267 & n5768;
  assign n5826 = ~n5071 & n5795;
  assign n5827 = n5825 & n5826;
  assign n5828 = ~n5824 & ~n5827;
  assign n5829 = ~n5815 & n5828;
  assign n5830 = ~n5803 & n5829;
  assign n5831 = ~n5074 & ~n5084;
  assign n5832 = n5074 & n5084;
  assign n5833 = ~n5095 & ~n5832;
  assign n5834 = ~n5083 & n5833;
  assign n5835 = ~n5831 & ~n5834;
  assign n5836 = n5830 & ~n5835;
  assign n5837 = ~n5830 & n5835;
  assign n5838 = ~n5836 & ~n5837;
  assign n5839 = pi132 & pi266;
  assign n5840 = n5119 & ~n5124;
  assign n5841 = ~n5125 & ~n5840;
  assign n5842 = n5839 & ~n5841;
  assign n5843 = ~n5119 & ~n5125;
  assign n5844 = ~n5124 & ~n5843;
  assign n5845 = ~n5839 & ~n5844;
  assign n5846 = ~n5842 & ~n5845;
  assign n5847 = ~n5838 & ~n5846;
  assign n5848 = n5830 & n5835;
  assign n5849 = ~n5830 & ~n5835;
  assign n5850 = ~n5848 & ~n5849;
  assign n5851 = ~n5839 & ~n5841;
  assign n5852 = n5839 & ~n5844;
  assign n5853 = ~n5851 & ~n5852;
  assign n5854 = ~n5850 & ~n5853;
  assign n5855 = ~n5847 & ~n5854;
  assign n5856 = ~n5759 & n5855;
  assign n5857 = n5759 & ~n5855;
  assign n5858 = ~n5856 & ~n5857;
  assign n5859 = pi265 & ~n5126;
  assign n5860 = pi132 & n5859;
  assign n5861 = ~n5117 & ~n5119;
  assign n5862 = ~n5860 & ~n5861;
  assign n5863 = pi264 & ~n5862;
  assign n5864 = pi133 & n5863;
  assign n5865 = pi134 & pi264;
  assign n5866 = ~n5118 & ~n5861;
  assign n5867 = ~n5860 & n5866;
  assign n5868 = ~n5135 & ~n5867;
  assign n5869 = ~n5865 & ~n5868;
  assign n5870 = ~n5864 & n5869;
  assign n5871 = ~n5864 & ~n5868;
  assign n5872 = n5865 & ~n5871;
  assign n5873 = ~n5870 & ~n5872;
  assign n5874 = ~n5858 & ~n5873;
  assign n5875 = ~n5759 & ~n5855;
  assign n5876 = n5759 & n5855;
  assign n5877 = ~n5875 & ~n5876;
  assign n5878 = n5865 & ~n5868;
  assign n5879 = ~n5864 & n5878;
  assign n5880 = ~n5865 & ~n5871;
  assign n5881 = ~n5879 & ~n5880;
  assign n5882 = ~n5877 & ~n5881;
  assign n5883 = ~n5874 & ~n5882;
  assign n5884 = n5139 & ~n5164;
  assign n5885 = ~n5139 & n5164;
  assign n5886 = ~n5155 & ~n5885;
  assign n5887 = ~n5884 & ~n5886;
  assign n5888 = ~n5883 & ~n5887;
  assign n5889 = n5883 & n5887;
  assign n5890 = ~n5888 & ~n5889;
  assign n5891 = pi263 & ~n5890;
  assign n5892 = pi135 & n5891;
  assign n5893 = pi135 & pi263;
  assign n5894 = n5883 & ~n5887;
  assign n5895 = ~n5883 & n5887;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = ~n5893 & ~n5896;
  assign n5898 = ~n5892 & ~n5897;
  assign n5899 = n5173 & n5178;
  assign n5900 = ~n5173 & ~n5178;
  assign n5901 = n5169 & ~n5900;
  assign n5902 = ~n5899 & ~n5901;
  assign n5903 = n5898 & ~n5902;
  assign n5904 = ~n5898 & n5902;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = pi136 & pi262;
  assign n5907 = ~n5010 & ~n5743;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = ~n5741 & n5908;
  assign n5910 = ~n5741 & ~n5907;
  assign n5911 = n5906 & ~n5910;
  assign n5912 = ~n5909 & ~n5911;
  assign n5913 = ~n5905 & ~n5912;
  assign n5914 = n5898 & n5902;
  assign n5915 = ~n5898 & ~n5902;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = n5906 & ~n5907;
  assign n5918 = ~n5741 & n5917;
  assign n5919 = ~n5906 & ~n5910;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n5916 & ~n5920;
  assign n5922 = ~n5913 & ~n5921;
  assign n5923 = ~n5758 & n5922;
  assign n5924 = n5758 & ~n5922;
  assign n5925 = ~n5923 & ~n5924;
  assign n5926 = pi260 & ~n5925;
  assign n5927 = pi138 & n5926;
  assign n5928 = pi138 & pi260;
  assign n5929 = n5758 & n5922;
  assign n5930 = ~n5758 & ~n5922;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = ~n5928 & ~n5931;
  assign n5933 = ~n5927 & ~n5932;
  assign n5934 = ~n5757 & ~n5933;
  assign n5935 = n5749 & n5754;
  assign n5936 = ~n5749 & ~n5754;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = pi260 & ~n5931;
  assign n5939 = pi138 & n5938;
  assign n5940 = ~n5925 & ~n5928;
  assign n5941 = ~n5939 & ~n5940;
  assign n5942 = ~n5937 & ~n5941;
  assign n5943 = ~n5934 & ~n5942;
  assign n5944 = ~n4558 & ~n5232;
  assign n5945 = n4558 & n5232;
  assign n5946 = ~n5723 & ~n5945;
  assign n5947 = ~n5944 & ~n5946;
  assign n5948 = n5943 & ~n5947;
  assign n5949 = ~n5943 & n5947;
  assign n5950 = ~n5948 & ~n5949;
  assign n5951 = pi140 & pi258;
  assign n5952 = pi139 & pi259;
  assign n5953 = ~n5951 & ~n5952;
  assign n5954 = n5951 & n5952;
  assign n5955 = ~n5953 & ~n5954;
  assign n5956 = ~n4997 & n5230;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = n5951 & ~n5952;
  assign n5959 = ~n5951 & n5952;
  assign n5960 = ~n5958 & ~n5959;
  assign n5961 = n5230 & ~n5960;
  assign n5962 = ~n4997 & n5961;
  assign n5963 = ~n5957 & ~n5962;
  assign n5964 = ~n5950 & ~n5963;
  assign n5965 = n5943 & n5947;
  assign n5966 = ~n5943 & ~n5947;
  assign n5967 = ~n5965 & ~n5966;
  assign n5968 = ~n5956 & ~n5960;
  assign n5969 = n5230 & ~n5955;
  assign n5970 = ~n4997 & n5969;
  assign n5971 = ~n5968 & ~n5970;
  assign n5972 = ~n5967 & ~n5971;
  assign n5973 = ~n5964 & ~n5972;
  assign n5974 = pi322 & n5973;
  assign n5975 = ~n5733 & ~n5974;
  assign n5976 = n5732 & n5973;
  assign n5977 = n1445 & n5976;
  assign n5978 = ~n5975 & ~n5977;
  assign n5979 = ~n5720 & ~n5978;
  assign n5980 = ~n5715 & n5717;
  assign n5981 = n5715 & ~n5717;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~n5733 & n5973;
  assign n5984 = pi322 & n5983;
  assign n5985 = n5732 & ~n5974;
  assign n5986 = pi323 & n5985;
  assign n5987 = ~n5984 & ~n5986;
  assign n5988 = ~n5982 & ~n5987;
  assign n5989 = ~n5979 & ~n5988;
  assign n5990 = ~n4981 & n5258;
  assign n5991 = n4981 & ~n5258;
  assign n5992 = ~n5690 & ~n5991;
  assign n5993 = ~n5990 & ~n5992;
  assign n5994 = n5989 & ~n5993;
  assign n5995 = ~n5989 & n5993;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = pi326 & n4596;
  assign n5998 = pi325 & n5257;
  assign n5999 = n5997 & n5998;
  assign n6000 = ~n5997 & ~n5998;
  assign n6001 = ~n5999 & ~n6000;
  assign n6002 = ~n5996 & ~n6001;
  assign n6003 = ~n5989 & ~n5993;
  assign n6004 = n5989 & n5993;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = ~n5997 & n5998;
  assign n6007 = n5997 & ~n5998;
  assign n6008 = ~n6006 & ~n6007;
  assign n6009 = ~n6005 & ~n6008;
  assign n6010 = ~n6002 & ~n6009;
  assign n6011 = ~n5711 & ~n6010;
  assign n6012 = n5704 & n5708;
  assign n6013 = ~n5704 & ~n5708;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = ~n6001 & ~n6005;
  assign n6016 = ~n5996 & ~n6008;
  assign n6017 = ~n6015 & ~n6016;
  assign n6018 = ~n6014 & ~n6017;
  assign n6019 = ~n6011 & ~n6018;
  assign n6020 = ~n5685 & n6019;
  assign n6021 = n5685 & ~n6019;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = pi329 & n2091;
  assign n6024 = pi328 & n2464;
  assign n6025 = n6023 & n6024;
  assign n6026 = ~n6023 & ~n6024;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = ~n6022 & ~n6027;
  assign n6029 = n5685 & n6019;
  assign n6030 = ~n5685 & ~n6019;
  assign n6031 = ~n6029 & ~n6030;
  assign n6032 = ~n6023 & n6024;
  assign n6033 = n6023 & ~n6024;
  assign n6034 = ~n6032 & ~n6033;
  assign n6035 = ~n6031 & ~n6034;
  assign n6036 = ~n6028 & ~n6035;
  assign n6037 = ~n5684 & ~n6036;
  assign n6038 = n5677 & n5681;
  assign n6039 = ~n5677 & ~n5681;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n6027 & ~n6031;
  assign n6042 = ~n6022 & ~n6034;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = ~n6040 & ~n6043;
  assign n6045 = ~n6037 & ~n6044;
  assign n6046 = n5657 & n6045;
  assign n6047 = ~n5657 & ~n6045;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = n1442 & ~n6048;
  assign n6050 = pi331 & n6049;
  assign n6051 = pi331 & n1442;
  assign n6052 = ~n5657 & n6045;
  assign n6053 = n5657 & ~n6045;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = ~n6051 & ~n6054;
  assign n6056 = ~n6050 & ~n6055;
  assign n6057 = ~n5650 & ~n6056;
  assign n6058 = ~n5638 & ~n5647;
  assign n6059 = n5638 & n5647;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = n1442 & ~n6054;
  assign n6062 = pi331 & n6061;
  assign n6063 = ~n6048 & ~n6051;
  assign n6064 = ~n6062 & ~n6063;
  assign n6065 = ~n6060 & ~n6064;
  assign n6066 = ~n6057 & ~n6065;
  assign n6067 = n5624 & n6066;
  assign n6068 = ~n5624 & ~n6066;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n1154 & n5376;
  assign n6071 = n1154 & ~n5376;
  assign n6072 = n4700 & ~n6071;
  assign n6073 = n1156 & n6072;
  assign n6074 = ~n6070 & ~n6073;
  assign n6075 = ~n1256 & ~n6074;
  assign n6076 = pi332 & n6075;
  assign n6077 = n1256 & ~n6070;
  assign n6078 = ~n6073 & n6077;
  assign n6079 = pi332 & ~n6078;
  assign n6080 = ~n6076 & n6079;
  assign n6081 = ~n1154 & ~n6080;
  assign n6082 = pi333 & n6081;
  assign n6083 = pi333 & ~n1154;
  assign n6084 = n6079 & ~n6083;
  assign n6085 = ~n6076 & n6084;
  assign n6086 = ~n6082 & ~n6085;
  assign n6087 = ~n6069 & ~n6086;
  assign n6088 = n5624 & ~n6066;
  assign n6089 = ~n5624 & n6066;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = ~n6080 & ~n6083;
  assign n6092 = n6080 & n6083;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = ~n6090 & ~n6093;
  assign n6095 = ~n6087 & ~n6094;
  assign n6096 = ~n5621 & n6095;
  assign n6097 = n5621 & ~n6095;
  assign n6098 = ~n6096 & ~n6097;
  assign n6099 = pi270 & pi334;
  assign n6100 = n1156 & n6099;
  assign n6101 = pi334 & n1156;
  assign n6102 = ~pi270 & ~n6101;
  assign n6103 = ~n6100 & ~n6102;
  assign n6104 = ~n6098 & ~n6103;
  assign n6105 = n5621 & n6095;
  assign n6106 = ~n5621 & ~n6095;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = pi270 & ~n6101;
  assign n6109 = ~pi270 & pi334;
  assign n6110 = n1156 & n6109;
  assign n6111 = ~n6108 & ~n6110;
  assign n6112 = ~n6107 & ~n6111;
  assign n6113 = ~n6104 & ~n6112;
  assign n6114 = n4915 & ~n5404;
  assign n6115 = ~n5405 & ~n6114;
  assign n6116 = n6113 & ~n6115;
  assign n6117 = ~n6113 & n6115;
  assign n6118 = ~n6116 & ~n6117;
  assign n6119 = ~n5619 & ~n6118;
  assign n6120 = n6113 & n6115;
  assign n6121 = ~n6113 & ~n6115;
  assign n6122 = ~n6120 & ~n6121;
  assign n6123 = n5619 & ~n6122;
  assign n6124 = ~n6119 & ~n6123;
  assign n6125 = ~n831 & ~n6124;
  assign n6126 = ~n5415 & ~n6125;
  assign n6127 = pi161 & ~n6126;
  assign n6128 = pi076 & ~pi161;
  assign n6129 = ~n6127 & ~n6128;
  assign po205 = ~pi160 & ~n6129;
  assign n6131 = pi077 & ~pi161;
  assign n6132 = ~pi270 & ~n5621;
  assign n6133 = pi270 & n5621;
  assign n6134 = ~n6095 & ~n6101;
  assign n6135 = pi334 & n6095;
  assign n6136 = n1156 & n6135;
  assign n6137 = ~n6134 & ~n6136;
  assign n6138 = ~n6133 & ~n6137;
  assign n6139 = ~n6132 & ~n6138;
  assign n6140 = n1154 & ~n6095;
  assign n6141 = n1156 & n6140;
  assign n6142 = n1156 & ~n6095;
  assign n6143 = ~n1154 & ~n6142;
  assign n6144 = ~n6141 & ~n6143;
  assign n6145 = pi334 & ~n6144;
  assign n6146 = ~n5638 & n6023;
  assign n6147 = n2464 & ~n6022;
  assign n6148 = pi328 & n6147;
  assign n6149 = ~n6024 & ~n6031;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n5684 & ~n6150;
  assign n6152 = n2464 & ~n6031;
  assign n6153 = pi328 & n6152;
  assign n6154 = ~n6022 & ~n6024;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6040 & ~n6155;
  assign n6157 = ~n6151 & ~n6156;
  assign n6158 = n5638 & ~n6023;
  assign n6159 = n6157 & ~n6158;
  assign n6160 = ~n6146 & ~n6159;
  assign n6161 = n5638 & n6045;
  assign n6162 = ~n5638 & ~n6045;
  assign n6163 = ~n6161 & ~n6162;
  assign n6164 = ~n5657 & ~n6163;
  assign n6165 = ~n5638 & n6045;
  assign n6166 = n5638 & ~n6045;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = n5657 & ~n6167;
  assign n6169 = ~n6164 & ~n6168;
  assign n6170 = n5647 & ~n6051;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = n1442 & ~n5647;
  assign n6173 = pi331 & n6172;
  assign n6174 = ~n6171 & ~n6173;
  assign n6175 = ~n6160 & n6174;
  assign n6176 = n6160 & ~n6174;
  assign n6177 = ~n6175 & ~n6176;
  assign n6178 = pi329 & n2464;
  assign n6179 = n5677 & n5685;
  assign n6180 = ~n5677 & ~n5685;
  assign n6181 = n6019 & ~n6180;
  assign n6182 = ~n6179 & ~n6181;
  assign n6183 = ~n5681 & n6024;
  assign n6184 = ~n5677 & ~n6019;
  assign n6185 = n5677 & n6019;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = n5685 & ~n6186;
  assign n6188 = n5677 & ~n6019;
  assign n6189 = ~n5677 & n6019;
  assign n6190 = ~n6188 & ~n6189;
  assign n6191 = ~n5685 & ~n6190;
  assign n6192 = ~n6187 & ~n6191;
  assign n6193 = n5681 & ~n6024;
  assign n6194 = ~n6192 & ~n6193;
  assign n6195 = ~n6183 & ~n6194;
  assign n6196 = ~n6182 & ~n6195;
  assign n6197 = n6182 & n6195;
  assign n6198 = ~n6196 & ~n6197;
  assign n6199 = n5715 & ~n5993;
  assign n6200 = ~n5717 & ~n5974;
  assign n6201 = n5717 & n5973;
  assign n6202 = pi322 & n6201;
  assign n6203 = ~n6200 & ~n6202;
  assign n6204 = ~n5733 & ~n6203;
  assign n6205 = n5717 & ~n5974;
  assign n6206 = ~n5717 & n5973;
  assign n6207 = pi322 & n6206;
  assign n6208 = ~n6205 & ~n6207;
  assign n6209 = n5732 & ~n6208;
  assign n6210 = pi323 & n6209;
  assign n6211 = ~n6204 & ~n6210;
  assign n6212 = ~n5715 & n5993;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = ~n6199 & ~n6213;
  assign n6215 = ~n5704 & n5998;
  assign n6216 = n5704 & ~n5998;
  assign n6217 = ~n5996 & ~n6216;
  assign n6218 = ~n6215 & ~n6217;
  assign n6219 = ~n6214 & n6218;
  assign n6220 = n6214 & ~n6218;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = pi324 & n5732;
  assign n6223 = pi323 & n5973;
  assign n6224 = ~n5717 & n5732;
  assign n6225 = pi323 & n6224;
  assign n6226 = n5717 & ~n5733;
  assign n6227 = n5973 & ~n6226;
  assign n6228 = pi322 & n6227;
  assign n6229 = ~n6225 & ~n6228;
  assign n6230 = pi130 & pi269;
  assign n6231 = pi128 & pi271;
  assign n6232 = pi270 & ~n6231;
  assign n6233 = pi129 & n6232;
  assign n6234 = pi129 & pi270;
  assign n6235 = pi271 & ~n6234;
  assign n6236 = pi128 & n6235;
  assign n6237 = ~n6233 & ~n6236;
  assign n6238 = ~n5776 & ~n5779;
  assign n6239 = n5776 & n5779;
  assign n6240 = ~n5775 & ~n6239;
  assign n6241 = ~n6238 & ~n6240;
  assign n6242 = ~n6237 & ~n6241;
  assign n6243 = ~n5774 & ~n6238;
  assign n6244 = ~n5024 & n6243;
  assign n6245 = ~n6239 & ~n6244;
  assign n6246 = n6237 & ~n6245;
  assign n6247 = ~n6242 & ~n6246;
  assign n6248 = n6230 & ~n6247;
  assign n6249 = n6237 & ~n6241;
  assign n6250 = ~n6237 & ~n6245;
  assign n6251 = ~n6249 & ~n6250;
  assign n6252 = ~n6230 & ~n6251;
  assign n6253 = ~n6248 & ~n6252;
  assign n6254 = ~n5775 & ~n5782;
  assign n6255 = ~n5774 & n5782;
  assign n6256 = ~n5024 & n6255;
  assign n6257 = ~n5783 & ~n6256;
  assign n6258 = ~n6254 & n6257;
  assign n6259 = ~n6254 & ~n6256;
  assign n6260 = pi268 & ~n6259;
  assign n6261 = pi130 & n6260;
  assign n6262 = n5027 & ~n5053;
  assign n6263 = ~pi129 & ~n5021;
  assign n6264 = ~n5050 & ~n6263;
  assign n6265 = ~n5027 & ~n6264;
  assign n6266 = ~n6262 & ~n6265;
  assign n6267 = ~pi130 & ~n6266;
  assign n6268 = ~n5021 & ~n5027;
  assign n6269 = n4373 & n5027;
  assign n6270 = ~n5020 & n6269;
  assign n6271 = ~n6268 & ~n6270;
  assign n6272 = ~pi267 & ~n6271;
  assign n6273 = ~n6267 & ~n6272;
  assign n6274 = pi129 & ~n5050;
  assign n6275 = ~n5021 & ~n6274;
  assign n6276 = ~n5027 & ~n6275;
  assign n6277 = n5027 & ~n6264;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = pi267 & ~n6278;
  assign n6280 = pi130 & n6279;
  assign n6281 = n5071 & ~n6280;
  assign n6282 = n6273 & ~n6281;
  assign n6283 = ~n6261 & ~n6282;
  assign n6284 = ~n6258 & ~n6283;
  assign n6285 = ~n6253 & ~n6284;
  assign n6286 = n6253 & n6284;
  assign n6287 = ~n6285 & ~n6286;
  assign n6288 = pi130 & ~n5816;
  assign n6289 = ~n5769 & ~n6288;
  assign n6290 = n5795 & ~n6289;
  assign n6291 = ~pi130 & ~n5769;
  assign n6292 = ~n5816 & ~n6291;
  assign n6293 = ~n5795 & ~n6292;
  assign n6294 = ~n6290 & ~n6293;
  assign n6295 = pi267 & ~n6294;
  assign n6296 = pi131 & n6295;
  assign n6297 = pi131 & pi268;
  assign n6298 = ~n5795 & ~n5819;
  assign n6299 = n5795 & ~n6292;
  assign n6300 = ~n6298 & ~n6299;
  assign n6301 = ~pi131 & ~n6300;
  assign n6302 = ~n5071 & ~n5795;
  assign n6303 = n5768 & n6302;
  assign n6304 = ~n5769 & n5795;
  assign n6305 = ~n6303 & ~n6304;
  assign n6306 = ~pi267 & ~n6305;
  assign n6307 = ~n6301 & ~n6306;
  assign n6308 = n5835 & n6307;
  assign n6309 = ~n6297 & ~n6308;
  assign n6310 = ~n6296 & n6309;
  assign n6311 = ~n6296 & ~n6308;
  assign n6312 = n6297 & ~n6311;
  assign n6313 = ~n6310 & ~n6312;
  assign n6314 = ~n6287 & ~n6313;
  assign n6315 = ~n6253 & n6284;
  assign n6316 = n6253 & ~n6284;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = n6297 & ~n6308;
  assign n6319 = ~n6296 & n6318;
  assign n6320 = ~n6297 & ~n6311;
  assign n6321 = ~n6319 & ~n6320;
  assign n6322 = ~n6317 & ~n6321;
  assign n6323 = ~n6314 & ~n6322;
  assign n6324 = n5839 & ~n5850;
  assign n6325 = ~n5839 & n5850;
  assign n6326 = ~n5841 & ~n6325;
  assign n6327 = ~n6324 & ~n6326;
  assign n6328 = n6323 & n6327;
  assign n6329 = ~n6323 & ~n6327;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = pi133 & pi266;
  assign n6332 = pi132 & pi267;
  assign n6333 = n6331 & n6332;
  assign n6334 = ~n6331 & ~n6332;
  assign n6335 = ~n6333 & ~n6334;
  assign n6336 = ~n6330 & ~n6335;
  assign n6337 = ~n6323 & n6327;
  assign n6338 = n6323 & ~n6327;
  assign n6339 = ~n6337 & ~n6338;
  assign n6340 = pi266 & ~n6332;
  assign n6341 = pi133 & n6340;
  assign n6342 = pi267 & ~n6331;
  assign n6343 = pi132 & n6342;
  assign n6344 = ~n6341 & ~n6343;
  assign n6345 = ~n6339 & ~n6344;
  assign n6346 = ~n6336 & ~n6345;
  assign n6347 = ~n5871 & ~n5875;
  assign n6348 = ~n5876 & ~n6347;
  assign n6349 = n6346 & n6348;
  assign n6350 = ~n6346 & ~n6348;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = pi134 & pi265;
  assign n6353 = n5855 & ~n5868;
  assign n6354 = ~n5864 & n6353;
  assign n6355 = ~n5855 & ~n5871;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n5759 & ~n6356;
  assign n6358 = ~n5855 & ~n5868;
  assign n6359 = ~n5864 & n6358;
  assign n6360 = n5855 & ~n5871;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = pi265 & ~n6361;
  assign n6363 = pi133 & n6362;
  assign n6364 = ~n6357 & ~n6363;
  assign n6365 = ~n5887 & ~n6364;
  assign n6366 = n5887 & n6364;
  assign n6367 = n5865 & ~n6366;
  assign n6368 = ~n6365 & ~n6367;
  assign n6369 = n6352 & ~n6368;
  assign n6370 = ~n5865 & ~n6365;
  assign n6371 = ~n6366 & ~n6370;
  assign n6372 = ~n6352 & ~n6371;
  assign n6373 = ~n6369 & ~n6372;
  assign n6374 = ~n6351 & ~n6373;
  assign n6375 = n6346 & ~n6348;
  assign n6376 = ~n6346 & n6348;
  assign n6377 = ~n6375 & ~n6376;
  assign n6378 = ~n6352 & ~n6368;
  assign n6379 = n6352 & ~n6371;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6377 & ~n6380;
  assign n6382 = ~n6374 & ~n6381;
  assign n6383 = ~n5890 & ~n5893;
  assign n6384 = ~n5178 & ~n5183;
  assign n6385 = ~n5184 & ~n6384;
  assign n6386 = n5890 & n5893;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = ~n6383 & ~n6387;
  assign n6389 = ~n6382 & n6388;
  assign n6390 = n6382 & ~n6388;
  assign n6391 = ~n6389 & ~n6390;
  assign n6392 = pi136 & pi263;
  assign n6393 = pi135 & pi264;
  assign n6394 = n6392 & n6393;
  assign n6395 = ~n6392 & ~n6393;
  assign n6396 = ~n6394 & ~n6395;
  assign n6397 = ~n6391 & ~n6396;
  assign n6398 = n6382 & n6388;
  assign n6399 = ~n6382 & ~n6388;
  assign n6400 = ~n6398 & ~n6399;
  assign n6401 = pi263 & ~n6393;
  assign n6402 = pi136 & n6401;
  assign n6403 = pi264 & ~n6392;
  assign n6404 = pi135 & n6403;
  assign n6405 = ~n6402 & ~n6404;
  assign n6406 = ~n6400 & ~n6405;
  assign n6407 = ~n6397 & ~n6406;
  assign n6408 = ~n5906 & ~n5916;
  assign n6409 = n5906 & n5916;
  assign n6410 = ~n5907 & ~n6409;
  assign n6411 = ~n5741 & n6410;
  assign n6412 = ~n6408 & ~n6411;
  assign n6413 = n6407 & ~n6412;
  assign n6414 = ~n6407 & n6412;
  assign n6415 = ~n6413 & ~n6414;
  assign n6416 = pi137 & pi262;
  assign n6417 = ~n5749 & ~n5922;
  assign n6418 = n5749 & n5922;
  assign n6419 = n5758 & ~n6418;
  assign n6420 = ~n6417 & ~n6419;
  assign n6421 = n6416 & ~n6420;
  assign n6422 = ~n5758 & ~n6417;
  assign n6423 = ~n6418 & ~n6422;
  assign n6424 = ~n6416 & ~n6423;
  assign n6425 = ~n6421 & ~n6424;
  assign n6426 = ~n6415 & ~n6425;
  assign n6427 = n6407 & n6412;
  assign n6428 = ~n6407 & ~n6412;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n6416 & ~n6420;
  assign n6431 = n6416 & ~n6423;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n6429 & ~n6432;
  assign n6434 = ~n6426 & ~n6433;
  assign n6435 = ~n5749 & n5922;
  assign n6436 = n5749 & ~n5922;
  assign n6437 = ~n6435 & ~n6436;
  assign n6438 = ~n5758 & ~n6437;
  assign n6439 = ~n6417 & ~n6418;
  assign n6440 = n5758 & ~n6439;
  assign n6441 = ~n6438 & ~n6440;
  assign n6442 = ~n5754 & ~n5928;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = pi260 & n5754;
  assign n6445 = pi138 & n6444;
  assign n6446 = ~n6443 & ~n6445;
  assign n6447 = ~n6434 & ~n6446;
  assign n6448 = n6434 & n6446;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = pi139 & pi260;
  assign n6451 = pi138 & pi261;
  assign n6452 = n6450 & n6451;
  assign n6453 = ~n6450 & ~n6451;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n6449 & ~n6454;
  assign n6456 = n6434 & ~n6446;
  assign n6457 = ~n6434 & n6446;
  assign n6458 = ~n6456 & ~n6457;
  assign n6459 = pi260 & ~n6451;
  assign n6460 = pi139 & n6459;
  assign n6461 = pi261 & ~n6450;
  assign n6462 = pi138 & n6461;
  assign n6463 = ~n6460 & ~n6462;
  assign n6464 = ~n6458 & ~n6463;
  assign n6465 = ~n6455 & ~n6464;
  assign n6466 = pi259 & ~n5943;
  assign n6467 = ~pi259 & n5943;
  assign n6468 = pi258 & ~n6467;
  assign n6469 = ~n5230 & n6468;
  assign n6470 = ~n6466 & ~n6469;
  assign n6471 = pi139 & ~n6470;
  assign n6472 = n6465 & n6471;
  assign n6473 = ~n6465 & ~n6471;
  assign n6474 = ~n6472 & ~n6473;
  assign n6475 = pi140 & pi259;
  assign n6476 = pi141 & pi258;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = n6475 & n6476;
  assign n6479 = ~n6477 & ~n6478;
  assign n6480 = pi139 & ~pi259;
  assign n6481 = n5943 & n6480;
  assign n6482 = ~n6466 & ~n6481;
  assign n6483 = ~n5230 & ~n6482;
  assign n6484 = ~pi139 & ~n5943;
  assign n6485 = ~pi259 & ~n5943;
  assign n6486 = n5943 & n5952;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = n5230 & ~n6487;
  assign n6489 = ~n6484 & ~n6488;
  assign n6490 = ~n6483 & n6489;
  assign n6491 = pi140 & ~n6490;
  assign n6492 = pi258 & n6491;
  assign n6493 = pi140 & ~pi259;
  assign n6494 = pi139 & n6493;
  assign n6495 = ~pi140 & pi259;
  assign n6496 = pi258 & n6495;
  assign n6497 = ~n6494 & ~n6496;
  assign n6498 = ~n5230 & ~n6497;
  assign n6499 = ~pi140 & ~pi259;
  assign n6500 = n4997 & n6475;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = n5230 & ~n6501;
  assign n6503 = ~pi258 & ~pi259;
  assign n6504 = ~pi139 & ~n5951;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = ~n6502 & n6505;
  assign n6507 = ~n6498 & n6506;
  assign n6508 = ~n5943 & ~n6507;
  assign n6509 = pi139 & n6499;
  assign n6510 = ~n6475 & ~n6509;
  assign n6511 = ~n5230 & ~n6510;
  assign n6512 = ~pi259 & n5230;
  assign n6513 = pi139 & ~n6512;
  assign n6514 = pi140 & ~n6513;
  assign n6515 = ~n6511 & ~n6514;
  assign n6516 = pi258 & ~n6515;
  assign n6517 = ~pi140 & n5230;
  assign n6518 = pi258 & ~n6517;
  assign n6519 = pi259 & ~n6518;
  assign n6520 = pi139 & n6519;
  assign n6521 = ~n6516 & ~n6520;
  assign n6522 = n5943 & ~n6521;
  assign n6523 = ~n6508 & ~n6522;
  assign n6524 = n6492 & ~n6523;
  assign n6525 = ~n6492 & n6523;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = ~n6479 & ~n6526;
  assign n6528 = ~n6475 & n6476;
  assign n6529 = n6475 & ~n6476;
  assign n6530 = ~n6528 & ~n6529;
  assign n6531 = ~n6492 & ~n6523;
  assign n6532 = n6492 & n6523;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = ~n6530 & ~n6533;
  assign n6535 = ~n6527 & ~n6534;
  assign n6536 = ~n6474 & ~n6535;
  assign n6537 = n6465 & ~n6471;
  assign n6538 = ~n6465 & n6471;
  assign n6539 = ~n6537 & ~n6538;
  assign n6540 = ~n6526 & ~n6530;
  assign n6541 = ~n6479 & ~n6533;
  assign n6542 = ~n6540 & ~n6541;
  assign n6543 = ~n6539 & ~n6542;
  assign n6544 = ~n6536 & ~n6543;
  assign n6545 = ~n5947 & ~n6523;
  assign n6546 = n5947 & n6523;
  assign n6547 = ~n5723 & ~n6546;
  assign n6548 = ~n6545 & ~n6547;
  assign n6549 = n6544 & ~n6548;
  assign n6550 = ~n6544 & n6548;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = n6229 & ~n6551;
  assign n6553 = pi322 & n6552;
  assign n6554 = ~n6544 & ~n6548;
  assign n6555 = n6544 & n6548;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = pi322 & n6556;
  assign n6558 = ~n6229 & ~n6557;
  assign n6559 = ~n6553 & ~n6558;
  assign n6560 = ~n6223 & ~n6559;
  assign n6561 = ~n6229 & ~n6551;
  assign n6562 = pi322 & n6561;
  assign n6563 = n6229 & ~n6557;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = n5973 & ~n6564;
  assign n6566 = pi323 & n6565;
  assign n6567 = ~n6560 & ~n6566;
  assign n6568 = ~n6222 & n6567;
  assign n6569 = n6222 & ~n6567;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = pi326 & n5257;
  assign n6572 = pi325 & n5714;
  assign n6573 = n6571 & n6572;
  assign n6574 = ~n6571 & ~n6572;
  assign n6575 = ~n6573 & ~n6574;
  assign n6576 = ~n6570 & ~n6575;
  assign n6577 = n6222 & n6567;
  assign n6578 = ~n6222 & ~n6567;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = ~n6571 & n6572;
  assign n6581 = n6571 & ~n6572;
  assign n6582 = ~n6580 & ~n6581;
  assign n6583 = ~n6579 & ~n6582;
  assign n6584 = ~n6576 & ~n6583;
  assign n6585 = ~n6221 & ~n6584;
  assign n6586 = ~n6214 & ~n6218;
  assign n6587 = n6214 & n6218;
  assign n6588 = ~n6586 & ~n6587;
  assign n6589 = ~n6575 & ~n6579;
  assign n6590 = ~n6570 & ~n6582;
  assign n6591 = ~n6589 & ~n6590;
  assign n6592 = ~n6588 & ~n6591;
  assign n6593 = ~n6585 & ~n6592;
  assign n6594 = ~n5704 & n5993;
  assign n6595 = n5704 & ~n5993;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = ~n5989 & n5998;
  assign n6598 = n5989 & ~n5998;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = n5708 & ~n5997;
  assign n6601 = ~n6599 & ~n6600;
  assign n6602 = ~n6596 & n6601;
  assign n6603 = ~n5708 & n5997;
  assign n6604 = ~n5704 & ~n5993;
  assign n6605 = n5704 & n5993;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = n5989 & n5998;
  assign n6608 = ~n5989 & ~n5998;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = ~n6600 & ~n6609;
  assign n6611 = ~n6606 & n6610;
  assign n6612 = ~n6603 & ~n6611;
  assign n6613 = ~n6602 & n6612;
  assign n6614 = n6593 & n6613;
  assign n6615 = ~n6593 & ~n6613;
  assign n6616 = ~n6614 & ~n6615;
  assign n6617 = pi328 & n2887;
  assign n6618 = pi327 & n4596;
  assign n6619 = n6617 & n6618;
  assign n6620 = ~n6617 & ~n6618;
  assign n6621 = ~n6619 & ~n6620;
  assign n6622 = ~n6616 & ~n6621;
  assign n6623 = ~n6593 & n6613;
  assign n6624 = n6593 & ~n6613;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = ~n6617 & n6618;
  assign n6627 = n6617 & ~n6618;
  assign n6628 = ~n6626 & ~n6627;
  assign n6629 = ~n6625 & ~n6628;
  assign n6630 = ~n6622 & ~n6629;
  assign n6631 = ~n6198 & ~n6630;
  assign n6632 = ~n6182 & n6195;
  assign n6633 = n6182 & ~n6195;
  assign n6634 = ~n6632 & ~n6633;
  assign n6635 = ~n6621 & ~n6625;
  assign n6636 = ~n6616 & ~n6628;
  assign n6637 = ~n6635 & ~n6636;
  assign n6638 = ~n6634 & ~n6637;
  assign n6639 = ~n6631 & ~n6638;
  assign n6640 = ~n6178 & n6639;
  assign n6641 = n6178 & ~n6639;
  assign n6642 = ~n6640 & ~n6641;
  assign n6643 = pi331 & n1729;
  assign n6644 = ~pi330 & ~n5652;
  assign n6645 = n5652 & ~n5655;
  assign n6646 = ~n2091 & ~n6645;
  assign n6647 = ~n6644 & ~n6646;
  assign n6648 = ~n6167 & ~n6647;
  assign n6649 = ~n2091 & ~n5652;
  assign n6650 = n1729 & n6649;
  assign n6651 = ~n1729 & n5652;
  assign n6652 = n1729 & ~n5652;
  assign n6653 = ~n6163 & ~n6652;
  assign n6654 = ~n6651 & ~n6653;
  assign n6655 = n2091 & ~n6654;
  assign n6656 = ~n6650 & ~n6655;
  assign n6657 = pi330 & ~n6656;
  assign n6658 = ~n6648 & ~n6657;
  assign n6659 = n6643 & ~n6658;
  assign n6660 = ~n6643 & n6658;
  assign n6661 = ~n6659 & ~n6660;
  assign n6662 = ~n6642 & ~n6661;
  assign n6663 = n6178 & n6639;
  assign n6664 = ~n6178 & ~n6639;
  assign n6665 = ~n6663 & ~n6664;
  assign n6666 = ~n6643 & ~n6658;
  assign n6667 = n6643 & n6658;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = ~n6665 & ~n6668;
  assign n6670 = ~n6662 & ~n6669;
  assign n6671 = ~n6177 & ~n6670;
  assign n6672 = ~n6160 & ~n6174;
  assign n6673 = n6160 & n6174;
  assign n6674 = ~n6672 & ~n6673;
  assign n6675 = ~n6661 & ~n6665;
  assign n6676 = ~n6642 & ~n6668;
  assign n6677 = ~n6675 & ~n6676;
  assign n6678 = ~n6674 & ~n6677;
  assign n6679 = ~n6671 & ~n6678;
  assign n6680 = ~n1154 & n5624;
  assign n6681 = pi333 & n6680;
  assign n6682 = ~n5624 & ~n6083;
  assign n6683 = ~n6066 & n6079;
  assign n6684 = ~n6076 & n6683;
  assign n6685 = n6066 & ~n6080;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = ~n6682 & ~n6686;
  assign n6688 = ~n6681 & ~n6687;
  assign n6689 = n6679 & ~n6688;
  assign n6690 = ~n6679 & n6688;
  assign n6691 = ~n6689 & ~n6690;
  assign n6692 = n6066 & n6079;
  assign n6693 = ~n6076 & ~n6692;
  assign n6694 = n1442 & ~n6693;
  assign n6695 = pi332 & n6694;
  assign n6696 = pi332 & n1442;
  assign n6697 = ~n6692 & ~n6696;
  assign n6698 = ~n6076 & n6697;
  assign n6699 = ~n6695 & ~n6698;
  assign n6700 = ~n1256 & ~n6699;
  assign n6701 = pi333 & n6700;
  assign n6702 = pi333 & ~n1256;
  assign n6703 = ~n6698 & ~n6702;
  assign n6704 = ~n6695 & n6703;
  assign n6705 = ~n6701 & ~n6704;
  assign n6706 = ~n6691 & ~n6705;
  assign n6707 = n6679 & n6688;
  assign n6708 = ~n6679 & ~n6688;
  assign n6709 = ~n6707 & ~n6708;
  assign n6710 = ~n6699 & ~n6702;
  assign n6711 = n6699 & n6702;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n6709 & ~n6712;
  assign n6714 = ~n6706 & ~n6713;
  assign n6715 = n6145 & ~n6714;
  assign n6716 = ~n6145 & n6714;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = pi258 & ~n6717;
  assign n6719 = pi128 & n6718;
  assign n6720 = pi335 & n6719;
  assign n6721 = n6145 & n6714;
  assign n6722 = ~n6145 & ~n6714;
  assign n6723 = ~n6721 & ~n6722;
  assign n6724 = pi335 & n1156;
  assign n6725 = ~n6723 & ~n6724;
  assign n6726 = ~n6720 & ~n6725;
  assign n6727 = ~n6139 & ~n6726;
  assign n6728 = n6139 & n6726;
  assign n6729 = ~n6727 & ~n6728;
  assign n6730 = pi271 & ~n6729;
  assign n6731 = ~n6139 & n6726;
  assign n6732 = n6139 & ~n6726;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~pi271 & ~n6733;
  assign n6735 = ~n6730 & ~n6734;
  assign n6736 = n5619 & ~n6120;
  assign n6737 = ~n6121 & ~n6736;
  assign n6738 = n6735 & ~n6737;
  assign n6739 = ~n6735 & n6737;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = pi128 & ~n5614;
  assign n6742 = pi129 & ~n6741;
  assign n6743 = ~pi129 & ~n5614;
  assign n6744 = pi128 & n6743;
  assign n6745 = ~n6742 & ~n6744;
  assign n6746 = pi309 & ~n6745;
  assign n6747 = ~n5431 & n5572;
  assign n6748 = pi140 & ~pi141;
  assign n6749 = pi138 & n6748;
  assign n6750 = pi141 & ~n4077;
  assign n6751 = n5451 & n6750;
  assign n6752 = ~n6749 & ~n6751;
  assign n6753 = pi137 & ~n6752;
  assign n6754 = pi141 & n4077;
  assign n6755 = n5441 & n6754;
  assign n6756 = ~pi140 & ~pi141;
  assign n6757 = ~pi138 & n6756;
  assign n6758 = ~n6755 & ~n6757;
  assign n6759 = ~pi137 & ~n6758;
  assign n6760 = ~pi140 & pi141;
  assign n6761 = pi139 & n6760;
  assign n6762 = ~pi141 & ~n4077;
  assign n6763 = pi140 & n6762;
  assign n6764 = ~n6761 & ~n6763;
  assign n6765 = pi138 & ~n6764;
  assign n6766 = pi140 & pi141;
  assign n6767 = ~pi139 & n6766;
  assign n6768 = ~pi141 & n4077;
  assign n6769 = ~pi140 & n6768;
  assign n6770 = ~n6767 & ~n6769;
  assign n6771 = ~pi138 & ~n6770;
  assign n6772 = ~n5445 & ~n5456;
  assign n6773 = ~pi141 & ~n6772;
  assign n6774 = ~n6771 & ~n6773;
  assign n6775 = ~n6765 & n6774;
  assign n6776 = ~n6759 & n6775;
  assign n6777 = ~n6753 & n6776;
  assign n6778 = pi321 & n6777;
  assign n6779 = ~n5464 & n5475;
  assign n6780 = n4772 & ~n6779;
  assign n6781 = pi320 & n6780;
  assign n6782 = n5463 & ~n5475;
  assign n6783 = pi321 & n6782;
  assign n6784 = ~n6781 & ~n6783;
  assign n6785 = pi320 & n5463;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = n5463 & n6784;
  assign n6788 = pi320 & n6787;
  assign n6789 = ~n6786 & ~n6788;
  assign n6790 = ~n6778 & ~n6789;
  assign n6791 = n6784 & ~n6785;
  assign n6792 = n5463 & ~n6784;
  assign n6793 = pi320 & n6792;
  assign n6794 = ~n6791 & ~n6793;
  assign n6795 = n6777 & ~n6794;
  assign n6796 = pi321 & n6795;
  assign n6797 = ~n6790 & ~n6796;
  assign n6798 = n4086 & ~n5493;
  assign n6799 = pi319 & n6798;
  assign n6800 = ~n5492 & ~n6799;
  assign n6801 = ~n6797 & ~n6800;
  assign n6802 = n6797 & n6800;
  assign n6803 = ~n6801 & ~n6802;
  assign n6804 = n4772 & ~n6803;
  assign n6805 = pi319 & n6804;
  assign n6806 = pi319 & n4772;
  assign n6807 = n6797 & ~n6800;
  assign n6808 = ~n6797 & n6800;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = ~n6806 & ~n6809;
  assign n6811 = ~n6805 & ~n6810;
  assign n6812 = n3552 & ~n5506;
  assign n6813 = pi318 & n6812;
  assign n6814 = ~n5507 & ~n6813;
  assign n6815 = n6811 & n6814;
  assign n6816 = ~n6811 & ~n6814;
  assign n6817 = ~n6815 & ~n6816;
  assign n6818 = n4086 & ~n6817;
  assign n6819 = pi318 & n6818;
  assign n6820 = pi318 & n4086;
  assign n6821 = ~n6811 & n6814;
  assign n6822 = n6811 & ~n6814;
  assign n6823 = ~n6821 & ~n6822;
  assign n6824 = ~n6820 & ~n6823;
  assign n6825 = ~n6819 & ~n6824;
  assign n6826 = n3012 & ~n5521;
  assign n6827 = pi317 & n6826;
  assign n6828 = ~n5520 & ~n6827;
  assign n6829 = ~n6825 & ~n6828;
  assign n6830 = n6825 & n6828;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = n3552 & ~n6831;
  assign n6833 = pi317 & n6832;
  assign n6834 = pi317 & n3552;
  assign n6835 = n6825 & ~n6828;
  assign n6836 = ~n6825 & n6828;
  assign n6837 = ~n6835 & ~n6836;
  assign n6838 = ~n6834 & ~n6837;
  assign n6839 = ~n6833 & ~n6838;
  assign n6840 = pi316 & n3012;
  assign n6841 = ~n6839 & ~n6840;
  assign n6842 = n3012 & n6839;
  assign n6843 = pi316 & n6842;
  assign n6844 = ~n6841 & ~n6843;
  assign n6845 = n2574 & ~n5537;
  assign n6846 = pi316 & n6845;
  assign n6847 = ~n5536 & ~n6846;
  assign n6848 = ~n6844 & ~n6847;
  assign n6849 = n6844 & n6847;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = n2574 & ~n6850;
  assign n6852 = pi315 & n6851;
  assign n6853 = pi315 & n2574;
  assign n6854 = n6844 & ~n6847;
  assign n6855 = ~n6844 & n6847;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = ~n6853 & ~n6856;
  assign n6858 = ~n6852 & ~n6857;
  assign n6859 = ~n5546 & ~n5559;
  assign n6860 = n5546 & n5559;
  assign n6861 = n2183 & ~n6860;
  assign n6862 = pi315 & n6861;
  assign n6863 = ~n6859 & ~n6862;
  assign n6864 = n6858 & n6863;
  assign n6865 = ~n6858 & ~n6863;
  assign n6866 = ~n6864 & ~n6865;
  assign n6867 = pi314 & n2183;
  assign n6868 = ~n5570 & ~n6867;
  assign n6869 = ~n5564 & n6868;
  assign n6870 = ~n5564 & ~n5570;
  assign n6871 = n6867 & ~n6870;
  assign n6872 = ~n6869 & ~n6871;
  assign n6873 = ~n6866 & ~n6872;
  assign n6874 = n6858 & ~n6863;
  assign n6875 = ~n6858 & n6863;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = ~n5570 & n6867;
  assign n6878 = ~n5564 & n6877;
  assign n6879 = ~n6867 & ~n6870;
  assign n6880 = ~n6878 & ~n6879;
  assign n6881 = ~n6876 & ~n6880;
  assign n6882 = ~n6873 & ~n6881;
  assign n6883 = ~n1533 & ~n1840;
  assign n6884 = pi313 & ~n6883;
  assign n6885 = n6882 & ~n6884;
  assign n6886 = ~n1533 & n1840;
  assign n6887 = pi313 & ~n6882;
  assign n6888 = n6886 & n6887;
  assign n6889 = ~n6885 & ~n6888;
  assign n6890 = ~n6747 & ~n6889;
  assign n6891 = ~n1840 & n6882;
  assign n6892 = pi313 & n1840;
  assign n6893 = ~n6882 & n6892;
  assign n6894 = ~n6891 & ~n6893;
  assign n6895 = ~n5572 & ~n6894;
  assign n6896 = n5431 & n6895;
  assign n6897 = n1533 & ~n1840;
  assign n6898 = ~n6882 & n6897;
  assign n6899 = ~n1533 & ~n5572;
  assign n6900 = n1840 & ~n6899;
  assign n6901 = n6882 & n6900;
  assign n6902 = ~n6898 & ~n6901;
  assign n6903 = pi313 & ~n6902;
  assign n6904 = ~n6882 & ~n6892;
  assign n6905 = n5572 & n6904;
  assign n6906 = ~n6903 & ~n6905;
  assign n6907 = ~n5431 & ~n6906;
  assign n6908 = ~n1840 & ~n6882;
  assign n6909 = n1840 & n6882;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = n1533 & ~n6910;
  assign n6912 = pi313 & n6911;
  assign n6913 = n5572 & n6912;
  assign n6914 = ~n6907 & ~n6913;
  assign n6915 = ~n6896 & n6914;
  assign n6916 = ~n6890 & n6915;
  assign n6917 = pi312 & n1533;
  assign n6918 = n6916 & n6917;
  assign n6919 = ~n6916 & ~n6917;
  assign n6920 = ~n6918 & ~n6919;
  assign n6921 = n5576 & ~n5589;
  assign n6922 = ~n5576 & n5589;
  assign n6923 = ~n5580 & ~n6922;
  assign n6924 = ~n6921 & ~n6923;
  assign n6925 = ~n6920 & ~n6924;
  assign n6926 = n6920 & n6924;
  assign n6927 = ~n6925 & ~n6926;
  assign n6928 = ~pi129 & ~n4910;
  assign n6929 = pi128 & n6928;
  assign n6930 = ~n1567 & ~n5608;
  assign n6931 = ~n5607 & ~n6930;
  assign n6932 = ~n6929 & ~n6931;
  assign n6933 = pi310 & ~n6932;
  assign n6934 = n6927 & n6933;
  assign n6935 = ~n6927 & ~n6933;
  assign n6936 = ~n6934 & ~n6935;
  assign n6937 = ~n1515 & ~n5594;
  assign n6938 = n1515 & n5594;
  assign n6939 = n5417 & ~n6938;
  assign n6940 = ~n6937 & ~n6939;
  assign n6941 = n1553 & ~n6940;
  assign n6942 = n5417 & ~n5594;
  assign n6943 = ~n1553 & ~n6942;
  assign n6944 = n1515 & n6943;
  assign n6945 = ~n6941 & ~n6944;
  assign n6946 = pi311 & ~n6945;
  assign n6947 = pi311 & n1553;
  assign n6948 = n5594 & ~n6947;
  assign n6949 = ~n5417 & n6948;
  assign n6950 = ~n6946 & ~n6949;
  assign n6951 = pi310 & n1515;
  assign n6952 = n6950 & ~n6951;
  assign n6953 = n1515 & ~n6950;
  assign n6954 = pi310 & n6953;
  assign n6955 = ~n6952 & ~n6954;
  assign n6956 = ~n6936 & ~n6955;
  assign n6957 = ~n6927 & n6933;
  assign n6958 = n6927 & ~n6933;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6950 & ~n6951;
  assign n6961 = n1515 & n6950;
  assign n6962 = pi310 & n6961;
  assign n6963 = ~n6960 & ~n6962;
  assign n6964 = ~n6959 & ~n6963;
  assign n6965 = ~n6956 & ~n6964;
  assign n6966 = n6746 & ~n6965;
  assign n6967 = ~n6746 & n6965;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = pi128 & pi308;
  assign n6970 = n6968 & ~n6969;
  assign n6971 = pi308 & ~n6968;
  assign n6972 = pi128 & n6971;
  assign n6973 = ~n6970 & ~n6972;
  assign n6974 = ~n6740 & ~n6973;
  assign n6975 = n6735 & n6737;
  assign n6976 = ~n6735 & ~n6737;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = ~n6968 & ~n6969;
  assign n6979 = pi308 & n6968;
  assign n6980 = pi128 & n6979;
  assign n6981 = ~n6978 & ~n6980;
  assign n6982 = ~n6977 & ~n6981;
  assign n6983 = ~n6974 & ~n6982;
  assign n6984 = ~n831 & ~n6983;
  assign n6985 = ~pi271 & n831;
  assign n6986 = ~n6984 & ~n6985;
  assign n6987 = pi161 & n6986;
  assign n6988 = ~n6131 & ~n6987;
  assign po206 = ~pi160 & ~n6988;
  assign n6990 = pi272 & n831;
  assign n6991 = pi308 & ~n1568;
  assign n6992 = n6927 & n6950;
  assign n6993 = ~n6927 & ~n6950;
  assign n6994 = ~n6992 & ~n6993;
  assign n6995 = ~n6933 & ~n6951;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = n1515 & n6933;
  assign n6998 = pi310 & n6997;
  assign n6999 = ~n6996 & ~n6998;
  assign n7000 = ~n6927 & ~n6947;
  assign n7001 = ~n5417 & n5594;
  assign n7002 = ~n5418 & ~n7001;
  assign n7003 = ~n6942 & ~n7002;
  assign n7004 = n6927 & n6947;
  assign n7005 = ~n7003 & ~n7004;
  assign n7006 = ~n7000 & ~n7005;
  assign n7007 = n5572 & ~n6904;
  assign n7008 = n1533 & ~n6908;
  assign n7009 = pi313 & n7008;
  assign n7010 = ~n7007 & ~n7009;
  assign n7011 = ~n5431 & ~n7010;
  assign n7012 = n5572 & n7008;
  assign n7013 = ~n6909 & ~n7012;
  assign n7014 = pi313 & ~n7013;
  assign n7015 = ~n7011 & ~n7014;
  assign n7016 = pi313 & n2183;
  assign n7017 = n7015 & n7016;
  assign n7018 = ~n7015 & ~n7016;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = ~n6866 & ~n6867;
  assign n7021 = n6866 & n6867;
  assign n7022 = ~n5570 & ~n7021;
  assign n7023 = ~n5564 & n7022;
  assign n7024 = ~n7020 & ~n7023;
  assign n7025 = pi138 & pi140;
  assign n7026 = pi139 & n6750;
  assign n7027 = ~n7025 & ~n7026;
  assign n7028 = pi137 & ~n7027;
  assign n7029 = pi139 & pi141;
  assign n7030 = ~n5452 & ~n7029;
  assign n7031 = pi138 & ~n7030;
  assign n7032 = ~pi139 & ~pi141;
  assign n7033 = pi140 & ~n7032;
  assign n7034 = ~n7031 & ~n7033;
  assign n7035 = ~n7028 & n7034;
  assign n7036 = pi142 & n7035;
  assign n7037 = ~pi142 & ~n7035;
  assign n7038 = ~n7036 & ~n7037;
  assign n7039 = pi141 & ~n7038;
  assign n7040 = pi142 & ~n7035;
  assign n7041 = ~pi142 & n7035;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = ~pi141 & ~n7042;
  assign n7044 = ~n7039 & ~n7043;
  assign n7045 = pi321 & n7044;
  assign n7046 = ~n6778 & n6784;
  assign n7047 = n5463 & ~n7046;
  assign n7048 = pi320 & n7047;
  assign n7049 = n6777 & ~n6784;
  assign n7050 = pi321 & n7049;
  assign n7051 = ~n7048 & ~n7050;
  assign n7052 = pi320 & n6777;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = n6777 & n7051;
  assign n7055 = pi320 & n7054;
  assign n7056 = ~n7053 & ~n7055;
  assign n7057 = ~n7045 & ~n7056;
  assign n7058 = n7051 & ~n7052;
  assign n7059 = n6777 & ~n7051;
  assign n7060 = pi320 & n7059;
  assign n7061 = ~n7058 & ~n7060;
  assign n7062 = n7044 & ~n7061;
  assign n7063 = pi321 & n7062;
  assign n7064 = ~n7057 & ~n7063;
  assign n7065 = n4772 & ~n6802;
  assign n7066 = pi319 & n7065;
  assign n7067 = ~n6801 & ~n7066;
  assign n7068 = ~n7064 & ~n7067;
  assign n7069 = n7064 & n7067;
  assign n7070 = ~n7068 & ~n7069;
  assign n7071 = n5463 & ~n7070;
  assign n7072 = pi319 & n7071;
  assign n7073 = pi319 & n5463;
  assign n7074 = n7064 & ~n7067;
  assign n7075 = ~n7064 & n7067;
  assign n7076 = ~n7074 & ~n7075;
  assign n7077 = ~n7073 & ~n7076;
  assign n7078 = ~n7072 & ~n7077;
  assign n7079 = n4086 & ~n6815;
  assign n7080 = pi318 & n7079;
  assign n7081 = ~n6816 & ~n7080;
  assign n7082 = n7078 & n7081;
  assign n7083 = ~n7078 & ~n7081;
  assign n7084 = ~n7082 & ~n7083;
  assign n7085 = n4772 & ~n7084;
  assign n7086 = pi318 & n7085;
  assign n7087 = pi318 & n4772;
  assign n7088 = ~n7078 & n7081;
  assign n7089 = n7078 & ~n7081;
  assign n7090 = ~n7088 & ~n7089;
  assign n7091 = ~n7087 & ~n7090;
  assign n7092 = ~n7086 & ~n7091;
  assign n7093 = ~pi317 & ~n7092;
  assign n7094 = ~n4086 & ~n7092;
  assign n7095 = n4086 & n7092;
  assign n7096 = pi317 & n7095;
  assign n7097 = ~n7094 & ~n7096;
  assign n7098 = ~n3552 & ~n7097;
  assign n7099 = ~n7093 & ~n7098;
  assign n7100 = ~n6829 & ~n7099;
  assign n7101 = n6828 & n7092;
  assign n7102 = n6825 & n7101;
  assign n7103 = ~n6828 & ~n7092;
  assign n7104 = ~n6825 & n7103;
  assign n7105 = ~n7102 & ~n7104;
  assign n7106 = pi317 & ~n7105;
  assign n7107 = ~n6837 & ~n7092;
  assign n7108 = n3552 & n7107;
  assign n7109 = ~n7106 & ~n7108;
  assign n7110 = n4086 & ~n7109;
  assign n7111 = n6828 & ~n7092;
  assign n7112 = n6825 & n7111;
  assign n7113 = n3552 & ~n6830;
  assign n7114 = pi317 & n7113;
  assign n7115 = ~n6829 & ~n7114;
  assign n7116 = n7092 & ~n7115;
  assign n7117 = ~n7112 & ~n7116;
  assign n7118 = ~n4086 & ~n7117;
  assign n7119 = ~pi317 & ~n6825;
  assign n7120 = ~n6828 & n7092;
  assign n7121 = n7119 & n7120;
  assign n7122 = ~n7118 & ~n7121;
  assign n7123 = ~n7110 & n7122;
  assign n7124 = ~n7100 & n7123;
  assign n7125 = ~n6839 & ~n6847;
  assign n7126 = n6839 & n6847;
  assign n7127 = n3012 & ~n7126;
  assign n7128 = pi316 & n7127;
  assign n7129 = ~n7125 & ~n7128;
  assign n7130 = ~n7124 & ~n7129;
  assign n7131 = n7124 & n7129;
  assign n7132 = ~n7130 & ~n7131;
  assign n7133 = n3552 & ~n7132;
  assign n7134 = pi316 & n7133;
  assign n7135 = pi316 & n3552;
  assign n7136 = n7124 & ~n7129;
  assign n7137 = ~n7124 & n7129;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = ~n7135 & ~n7138;
  assign n7140 = ~n7134 & ~n7139;
  assign n7141 = ~n6853 & n6863;
  assign n7142 = ~n6856 & ~n7141;
  assign n7143 = n2574 & ~n6863;
  assign n7144 = pi315 & n7143;
  assign n7145 = ~n7142 & ~n7144;
  assign n7146 = n7140 & n7145;
  assign n7147 = ~n7140 & ~n7145;
  assign n7148 = ~n7146 & ~n7147;
  assign n7149 = n3012 & ~n7148;
  assign n7150 = pi315 & n7149;
  assign n7151 = pi315 & n3012;
  assign n7152 = ~n7140 & n7145;
  assign n7153 = n7140 & ~n7145;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = ~n7151 & ~n7154;
  assign n7156 = ~n7150 & ~n7155;
  assign n7157 = n2574 & ~n7156;
  assign n7158 = pi314 & n7157;
  assign n7159 = pi314 & n2574;
  assign n7160 = ~n7155 & ~n7159;
  assign n7161 = ~n7150 & n7160;
  assign n7162 = ~n7158 & ~n7161;
  assign n7163 = ~n7024 & ~n7162;
  assign n7164 = n7024 & ~n7161;
  assign n7165 = ~n7158 & n7164;
  assign n7166 = ~n7163 & ~n7165;
  assign n7167 = n7019 & ~n7166;
  assign n7168 = ~n7019 & n7166;
  assign n7169 = ~n7167 & ~n7168;
  assign n7170 = pi312 & n1840;
  assign n7171 = ~n6916 & ~n6924;
  assign n7172 = n6916 & n6924;
  assign n7173 = n6917 & ~n7172;
  assign n7174 = ~n7171 & ~n7173;
  assign n7175 = n7170 & ~n7174;
  assign n7176 = ~n6917 & ~n7171;
  assign n7177 = ~n7172 & ~n7176;
  assign n7178 = ~n7170 & ~n7177;
  assign n7179 = ~n7175 & ~n7178;
  assign n7180 = ~n7169 & ~n7179;
  assign n7181 = n7019 & n7166;
  assign n7182 = ~n7019 & ~n7166;
  assign n7183 = ~n7181 & ~n7182;
  assign n7184 = ~n7170 & ~n7174;
  assign n7185 = n7170 & ~n7177;
  assign n7186 = ~n7184 & ~n7185;
  assign n7187 = ~n7183 & ~n7186;
  assign n7188 = ~n7180 & ~n7187;
  assign n7189 = n7006 & n7188;
  assign n7190 = ~n7006 & ~n7188;
  assign n7191 = ~n7189 & ~n7190;
  assign n7192 = n1533 & ~n7191;
  assign n7193 = pi311 & n7192;
  assign n7194 = pi311 & n1533;
  assign n7195 = ~n7006 & n7188;
  assign n7196 = n7006 & ~n7188;
  assign n7197 = ~n7195 & ~n7196;
  assign n7198 = ~n7194 & ~n7197;
  assign n7199 = ~n7193 & ~n7198;
  assign n7200 = n1553 & ~n7199;
  assign n7201 = pi310 & n7200;
  assign n7202 = pi310 & n1553;
  assign n7203 = ~n7198 & ~n7202;
  assign n7204 = ~n7193 & n7203;
  assign n7205 = ~n7201 & ~n7204;
  assign n7206 = ~n6999 & ~n7205;
  assign n7207 = n6999 & ~n7204;
  assign n7208 = ~n7201 & n7207;
  assign n7209 = ~n7206 & ~n7208;
  assign n7210 = n6991 & ~n7209;
  assign n7211 = ~n6991 & n7209;
  assign n7212 = ~n7210 & ~n7211;
  assign n7213 = n5614 & n6965;
  assign n7214 = ~n5614 & ~n6965;
  assign n7215 = ~pi129 & ~n7214;
  assign n7216 = ~n7213 & ~n7215;
  assign n7217 = pi130 & ~n7216;
  assign n7218 = pi128 & n7217;
  assign n7219 = ~pi130 & n6965;
  assign n7220 = n1335 & n7219;
  assign n7221 = ~n7218 & ~n7220;
  assign n7222 = pi309 & ~n7221;
  assign n7223 = pi129 & ~n7213;
  assign n7224 = pi128 & n7223;
  assign n7225 = pi128 & ~n7214;
  assign n7226 = ~pi129 & ~n7225;
  assign n7227 = ~n7224 & ~n7226;
  assign n7228 = ~pi130 & ~n7227;
  assign n7229 = pi130 & ~n6965;
  assign n7230 = n1335 & n7229;
  assign n7231 = pi309 & ~n7230;
  assign n7232 = ~n7228 & n7231;
  assign n7233 = ~n7222 & n7232;
  assign n7234 = n6972 & ~n7233;
  assign n7235 = ~n6972 & n7233;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = ~n7212 & ~n7236;
  assign n7238 = n6991 & n7209;
  assign n7239 = ~n6991 & ~n7209;
  assign n7240 = ~n7238 & ~n7239;
  assign n7241 = n6972 & n7233;
  assign n7242 = ~n6972 & ~n7233;
  assign n7243 = ~n7241 & ~n7242;
  assign n7244 = ~n7240 & ~n7243;
  assign n7245 = ~n7237 & ~n7244;
  assign n7246 = ~pi271 & ~n6728;
  assign n7247 = ~n6727 & ~n7246;
  assign n7248 = pi258 & ~n6723;
  assign n7249 = pi128 & n7248;
  assign n7250 = pi335 & n7249;
  assign n7251 = n6160 & n6639;
  assign n7252 = ~n6160 & ~n6639;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = n6178 & ~n6658;
  assign n7255 = ~n6178 & n6658;
  assign n7256 = ~n7254 & ~n7255;
  assign n7257 = n6174 & ~n6643;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = ~n7253 & n7258;
  assign n7260 = ~n6174 & n6643;
  assign n7261 = n6160 & ~n6639;
  assign n7262 = ~n6160 & n6639;
  assign n7263 = ~n7261 & ~n7262;
  assign n7264 = ~n6178 & ~n6658;
  assign n7265 = n6178 & n6658;
  assign n7266 = ~n7264 & ~n7265;
  assign n7267 = ~n7257 & ~n7266;
  assign n7268 = ~n7263 & n7267;
  assign n7269 = ~n7260 & ~n7268;
  assign n7270 = ~n7259 & n7269;
  assign n7271 = ~n1256 & ~n6688;
  assign n7272 = pi333 & n7271;
  assign n7273 = ~n6679 & ~n6698;
  assign n7274 = ~n6695 & n7273;
  assign n7275 = n6679 & ~n6699;
  assign n7276 = ~n7274 & ~n7275;
  assign n7277 = n6688 & ~n6702;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = ~n7272 & ~n7278;
  assign n7280 = n7270 & ~n7279;
  assign n7281 = ~n7270 & n7279;
  assign n7282 = ~n7280 & ~n7281;
  assign n7283 = pi331 & n2091;
  assign n7284 = n6182 & ~n6613;
  assign n7285 = ~n6182 & n6613;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = ~n6593 & n6618;
  assign n7288 = n6593 & ~n6618;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = n6195 & ~n6617;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = ~n7286 & n7291;
  assign n7293 = ~n6195 & n6617;
  assign n7294 = n6182 & n6613;
  assign n7295 = ~n6182 & ~n6613;
  assign n7296 = ~n7294 & ~n7295;
  assign n7297 = n6593 & n6618;
  assign n7298 = ~n6593 & ~n6618;
  assign n7299 = ~n7297 & ~n7298;
  assign n7300 = ~n7290 & ~n7299;
  assign n7301 = ~n7296 & n7300;
  assign n7302 = ~n7293 & ~n7301;
  assign n7303 = ~n7292 & n7302;
  assign n7304 = ~n6160 & n6178;
  assign n7305 = n6160 & ~n6178;
  assign n7306 = n6639 & ~n7305;
  assign n7307 = ~n7304 & ~n7306;
  assign n7308 = n7303 & ~n7307;
  assign n7309 = ~n7303 & n7307;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = pi328 & n4596;
  assign n7312 = n6571 & ~n6613;
  assign n7313 = n5714 & ~n6570;
  assign n7314 = pi325 & n7313;
  assign n7315 = ~n6572 & ~n6579;
  assign n7316 = ~n7314 & ~n7315;
  assign n7317 = ~n6588 & ~n7316;
  assign n7318 = n5714 & ~n6579;
  assign n7319 = pi325 & n7318;
  assign n7320 = ~n6570 & ~n6572;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = ~n6221 & ~n7321;
  assign n7323 = ~n7317 & ~n7322;
  assign n7324 = ~n6571 & n6613;
  assign n7325 = ~n7323 & ~n7324;
  assign n7326 = ~n7312 & ~n7325;
  assign n7327 = n6182 & ~n6618;
  assign n7328 = ~n6625 & ~n7327;
  assign n7329 = ~n6182 & n6618;
  assign n7330 = ~n7328 & ~n7329;
  assign n7331 = n7326 & ~n7330;
  assign n7332 = ~n7326 & n7330;
  assign n7333 = ~n7331 & ~n7332;
  assign n7334 = n5973 & ~n6229;
  assign n7335 = pi323 & n7334;
  assign n7336 = ~n6223 & n6229;
  assign n7337 = n6556 & ~n7336;
  assign n7338 = pi322 & n7337;
  assign n7339 = ~n7335 & ~n7338;
  assign n7340 = ~n6214 & n6222;
  assign n7341 = n6214 & ~n6222;
  assign n7342 = ~n6567 & ~n7341;
  assign n7343 = ~n7340 & ~n7342;
  assign n7344 = ~n7339 & n7343;
  assign n7345 = n7339 & ~n7343;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = pi323 & n6556;
  assign n7348 = n6475 & n6492;
  assign n7349 = ~n6475 & ~n6492;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = pi258 & ~n7350;
  assign n7352 = pi141 & n7351;
  assign n7353 = n6475 & ~n6492;
  assign n7354 = ~n6475 & n6492;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = ~n6476 & ~n7355;
  assign n7357 = ~n7352 & ~n7356;
  assign n7358 = ~n6539 & ~n7357;
  assign n7359 = pi258 & ~n7355;
  assign n7360 = pi141 & n7359;
  assign n7361 = ~n6476 & ~n7350;
  assign n7362 = ~n7360 & ~n7361;
  assign n7363 = ~n6474 & ~n7362;
  assign n7364 = ~n7358 & ~n7363;
  assign n7365 = pi139 & pi261;
  assign n7366 = pi136 & pi264;
  assign n7367 = pi133 & pi267;
  assign n7368 = n6231 & n6234;
  assign n7369 = ~n6231 & ~n6234;
  assign n7370 = ~n6245 & ~n7369;
  assign n7371 = ~n7368 & ~n7370;
  assign n7372 = pi128 & pi272;
  assign n7373 = pi271 & ~n7372;
  assign n7374 = pi129 & n7373;
  assign n7375 = pi129 & pi271;
  assign n7376 = pi272 & ~n7375;
  assign n7377 = pi128 & n7376;
  assign n7378 = ~n7374 & ~n7377;
  assign n7379 = ~n7371 & n7378;
  assign n7380 = n7371 & ~n7378;
  assign n7381 = ~n7379 & ~n7380;
  assign n7382 = pi270 & ~n7381;
  assign n7383 = pi130 & n7382;
  assign n7384 = pi130 & pi270;
  assign n7385 = ~n7380 & ~n7384;
  assign n7386 = ~n7379 & n7385;
  assign n7387 = ~n7383 & ~n7386;
  assign n7388 = ~n6248 & ~n6284;
  assign n7389 = ~n6252 & ~n7388;
  assign n7390 = pi269 & ~n7389;
  assign n7391 = pi131 & n7390;
  assign n7392 = pi131 & pi269;
  assign n7393 = ~n7388 & ~n7392;
  assign n7394 = ~n6252 & n7393;
  assign n7395 = ~n7391 & ~n7394;
  assign n7396 = ~n7387 & ~n7395;
  assign n7397 = ~n7389 & ~n7392;
  assign n7398 = n7389 & n7392;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = ~n7386 & ~n7399;
  assign n7401 = ~n7383 & n7400;
  assign n7402 = ~n7396 & ~n7401;
  assign n7403 = ~n6287 & ~n6297;
  assign n7404 = n6287 & n6297;
  assign n7405 = ~n6308 & ~n7404;
  assign n7406 = ~n6296 & n7405;
  assign n7407 = ~n7403 & ~n7406;
  assign n7408 = n7402 & ~n7407;
  assign n7409 = ~n7402 & n7407;
  assign n7410 = ~n7408 & ~n7409;
  assign n7411 = pi132 & pi268;
  assign n7412 = n6332 & ~n6337;
  assign n7413 = ~n6338 & ~n7412;
  assign n7414 = n7411 & ~n7413;
  assign n7415 = ~n6332 & ~n6338;
  assign n7416 = ~n6337 & ~n7415;
  assign n7417 = ~n7411 & ~n7416;
  assign n7418 = ~n7414 & ~n7417;
  assign n7419 = ~n7410 & ~n7418;
  assign n7420 = n7402 & n7407;
  assign n7421 = ~n7402 & ~n7407;
  assign n7422 = ~n7420 & ~n7421;
  assign n7423 = ~n7411 & ~n7413;
  assign n7424 = n7411 & ~n7416;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = ~n7422 & ~n7425;
  assign n7427 = ~n7419 & ~n7426;
  assign n7428 = ~n7367 & n7427;
  assign n7429 = n7367 & ~n7427;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = pi267 & ~n6339;
  assign n7432 = pi132 & n7431;
  assign n7433 = ~n6330 & ~n6332;
  assign n7434 = ~n7432 & ~n7433;
  assign n7435 = pi266 & ~n7434;
  assign n7436 = pi133 & n7435;
  assign n7437 = pi134 & pi266;
  assign n7438 = ~n6331 & ~n7433;
  assign n7439 = ~n7432 & n7438;
  assign n7440 = ~n6348 & ~n7439;
  assign n7441 = ~n7437 & ~n7440;
  assign n7442 = ~n7436 & n7441;
  assign n7443 = ~n7436 & ~n7440;
  assign n7444 = n7437 & ~n7443;
  assign n7445 = ~n7442 & ~n7444;
  assign n7446 = ~n7430 & ~n7445;
  assign n7447 = ~n7367 & ~n7427;
  assign n7448 = n7367 & n7427;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = n7437 & ~n7440;
  assign n7451 = ~n7436 & n7450;
  assign n7452 = ~n7437 & ~n7443;
  assign n7453 = ~n7451 & ~n7452;
  assign n7454 = ~n7449 & ~n7453;
  assign n7455 = ~n7446 & ~n7454;
  assign n7456 = n6352 & ~n6377;
  assign n7457 = ~n6352 & n6377;
  assign n7458 = ~n6368 & ~n7457;
  assign n7459 = ~n7456 & ~n7458;
  assign n7460 = n7455 & n7459;
  assign n7461 = ~n7455 & ~n7459;
  assign n7462 = ~n7460 & ~n7461;
  assign n7463 = pi135 & pi265;
  assign n7464 = n6393 & ~n6399;
  assign n7465 = ~n6398 & ~n7464;
  assign n7466 = n7463 & ~n7465;
  assign n7467 = ~n6393 & ~n6398;
  assign n7468 = ~n6399 & ~n7467;
  assign n7469 = ~n7463 & ~n7468;
  assign n7470 = ~n7466 & ~n7469;
  assign n7471 = ~n7462 & ~n7470;
  assign n7472 = n7455 & ~n7459;
  assign n7473 = ~n7455 & n7459;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = ~n7463 & ~n7465;
  assign n7476 = n7463 & ~n7468;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n7474 & ~n7477;
  assign n7479 = ~n7471 & ~n7478;
  assign n7480 = ~n7366 & n7479;
  assign n7481 = n7366 & ~n7479;
  assign n7482 = ~n7480 & ~n7481;
  assign n7483 = pi264 & ~n6400;
  assign n7484 = pi135 & n7483;
  assign n7485 = ~n6391 & ~n6393;
  assign n7486 = ~n7484 & ~n7485;
  assign n7487 = pi263 & ~n7486;
  assign n7488 = pi136 & n7487;
  assign n7489 = pi137 & pi263;
  assign n7490 = ~n6392 & ~n7485;
  assign n7491 = ~n7484 & n7490;
  assign n7492 = n6412 & ~n7491;
  assign n7493 = ~n7489 & ~n7492;
  assign n7494 = ~n7488 & n7493;
  assign n7495 = ~n7488 & ~n7492;
  assign n7496 = n7489 & ~n7495;
  assign n7497 = ~n7494 & ~n7496;
  assign n7498 = ~n7482 & ~n7497;
  assign n7499 = ~n7366 & ~n7479;
  assign n7500 = n7366 & n7479;
  assign n7501 = ~n7499 & ~n7500;
  assign n7502 = n7489 & ~n7492;
  assign n7503 = ~n7488 & n7502;
  assign n7504 = ~n7489 & ~n7495;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n7501 & ~n7505;
  assign n7507 = ~n7498 & ~n7506;
  assign n7508 = n6416 & ~n6429;
  assign n7509 = ~n6416 & n6429;
  assign n7510 = ~n6420 & ~n7509;
  assign n7511 = ~n7508 & ~n7510;
  assign n7512 = n7507 & ~n7511;
  assign n7513 = ~n7507 & n7511;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 = pi138 & pi262;
  assign n7516 = n6451 & ~n6457;
  assign n7517 = ~n6456 & ~n7516;
  assign n7518 = n7515 & ~n7517;
  assign n7519 = ~n6451 & ~n6456;
  assign n7520 = ~n6457 & ~n7519;
  assign n7521 = ~n7515 & ~n7520;
  assign n7522 = ~n7518 & ~n7521;
  assign n7523 = ~n7514 & ~n7522;
  assign n7524 = n7507 & n7511;
  assign n7525 = ~n7507 & ~n7511;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = ~n7515 & ~n7517;
  assign n7528 = n7515 & ~n7520;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = ~n7526 & ~n7529;
  assign n7531 = ~n7523 & ~n7530;
  assign n7532 = ~n7365 & ~n7531;
  assign n7533 = n7365 & n7531;
  assign n7534 = ~n7532 & ~n7533;
  assign n7535 = pi261 & ~n6458;
  assign n7536 = pi138 & n7535;
  assign n7537 = ~n6449 & ~n6451;
  assign n7538 = ~n6450 & ~n7537;
  assign n7539 = ~n7536 & n7538;
  assign n7540 = pi140 & pi260;
  assign n7541 = ~n7536 & ~n7537;
  assign n7542 = pi260 & ~n7541;
  assign n7543 = pi139 & n7542;
  assign n7544 = ~n6471 & ~n7543;
  assign n7545 = n7540 & ~n7544;
  assign n7546 = ~n7539 & n7545;
  assign n7547 = ~n7539 & ~n7544;
  assign n7548 = ~n7540 & ~n7547;
  assign n7549 = ~n7546 & ~n7548;
  assign n7550 = ~n7534 & ~n7549;
  assign n7551 = ~n7365 & n7531;
  assign n7552 = n7365 & ~n7531;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7540 & ~n7544;
  assign n7555 = ~n7539 & n7554;
  assign n7556 = n7540 & ~n7547;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = ~n7553 & ~n7557;
  assign n7559 = ~n7550 & ~n7558;
  assign n7560 = ~n7539 & ~n7543;
  assign n7561 = n6471 & ~n7560;
  assign n7562 = ~n6471 & n7560;
  assign n7563 = ~n7561 & ~n7562;
  assign n7564 = ~n7349 & ~n7563;
  assign n7565 = ~n7348 & ~n7564;
  assign n7566 = n7559 & n7565;
  assign n7567 = ~n7559 & ~n7565;
  assign n7568 = ~n7566 & ~n7567;
  assign n7569 = pi141 & pi259;
  assign n7570 = ~n6539 & ~n7350;
  assign n7571 = ~n6474 & ~n7355;
  assign n7572 = n6476 & ~n7571;
  assign n7573 = ~n7570 & n7572;
  assign n7574 = ~n7569 & ~n7573;
  assign n7575 = pi140 & n6492;
  assign n7576 = ~pi140 & ~n6492;
  assign n7577 = ~n7575 & ~n7576;
  assign n7578 = ~n6474 & ~n7577;
  assign n7579 = pi140 & ~n6492;
  assign n7580 = ~pi140 & n6492;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~n6539 & ~n7581;
  assign n7583 = ~n7578 & ~n7582;
  assign n7584 = n6476 & ~n7583;
  assign n7585 = pi259 & n7584;
  assign n7586 = ~n7574 & ~n7585;
  assign n7587 = pi258 & ~n7586;
  assign n7588 = pi142 & n7587;
  assign n7589 = pi142 & pi258;
  assign n7590 = ~n7585 & ~n7589;
  assign n7591 = ~n7574 & n7590;
  assign n7592 = ~n7588 & ~n7591;
  assign n7593 = ~n7568 & ~n7592;
  assign n7594 = n7559 & ~n7565;
  assign n7595 = ~n7559 & n7565;
  assign n7596 = ~n7594 & ~n7595;
  assign n7597 = ~n7586 & ~n7589;
  assign n7598 = n7586 & n7589;
  assign n7599 = ~n7597 & ~n7598;
  assign n7600 = ~n7596 & ~n7599;
  assign n7601 = ~n7593 & ~n7600;
  assign n7602 = ~n6548 & ~n7364;
  assign n7603 = n6548 & n7364;
  assign n7604 = ~n6523 & ~n7603;
  assign n7605 = ~n7602 & ~n7604;
  assign n7606 = n7601 & n7605;
  assign n7607 = ~n7601 & ~n7605;
  assign n7608 = ~n7606 & ~n7607;
  assign n7609 = ~n7364 & ~n7608;
  assign n7610 = n7601 & ~n7605;
  assign n7611 = ~n7601 & n7605;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = n7364 & ~n7612;
  assign n7614 = ~n7609 & ~n7613;
  assign n7615 = pi322 & ~n7614;
  assign n7616 = ~n7347 & ~n7615;
  assign n7617 = n6556 & ~n7614;
  assign n7618 = pi323 & n7617;
  assign n7619 = pi322 & n7618;
  assign n7620 = ~n7616 & ~n7619;
  assign n7621 = pi325 & n5732;
  assign n7622 = pi324 & n5973;
  assign n7623 = n7621 & n7622;
  assign n7624 = ~n7621 & ~n7622;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n7620 & ~n7625;
  assign n7627 = ~n7621 & n7622;
  assign n7628 = n7621 & ~n7622;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~n7619 & ~n7629;
  assign n7631 = ~n7616 & n7630;
  assign n7632 = ~n7626 & ~n7631;
  assign n7633 = ~n7346 & ~n7632;
  assign n7634 = ~n7339 & ~n7343;
  assign n7635 = n7339 & n7343;
  assign n7636 = ~n7634 & ~n7635;
  assign n7637 = ~n7620 & ~n7629;
  assign n7638 = ~n7619 & ~n7625;
  assign n7639 = ~n7616 & n7638;
  assign n7640 = ~n7637 & ~n7639;
  assign n7641 = ~n7636 & ~n7640;
  assign n7642 = ~n7633 & ~n7641;
  assign n7643 = ~n6218 & n6572;
  assign n7644 = ~n6214 & ~n6567;
  assign n7645 = n6214 & n6567;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = n6222 & ~n7646;
  assign n7648 = n6214 & ~n6567;
  assign n7649 = ~n6214 & n6567;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = ~n6222 & ~n7650;
  assign n7652 = ~n7647 & ~n7651;
  assign n7653 = n6218 & ~n6572;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~n7643 & ~n7654;
  assign n7656 = n7642 & n7655;
  assign n7657 = ~n7642 & ~n7655;
  assign n7658 = ~n7656 & ~n7657;
  assign n7659 = pi327 & n5257;
  assign n7660 = pi326 & n5714;
  assign n7661 = n7659 & n7660;
  assign n7662 = ~n7659 & ~n7660;
  assign n7663 = ~n7661 & ~n7662;
  assign n7664 = ~n7658 & ~n7663;
  assign n7665 = ~n7642 & n7655;
  assign n7666 = n7642 & ~n7655;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = ~n7659 & n7660;
  assign n7669 = n7659 & ~n7660;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7667 & ~n7670;
  assign n7672 = ~n7664 & ~n7671;
  assign n7673 = ~n7333 & ~n7672;
  assign n7674 = n7326 & n7330;
  assign n7675 = ~n7326 & ~n7330;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = ~n7663 & ~n7667;
  assign n7678 = ~n7658 & ~n7670;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7676 & ~n7679;
  assign n7681 = ~n7673 & ~n7680;
  assign n7682 = ~n7311 & n7681;
  assign n7683 = n7311 & ~n7681;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = ~n6167 & ~n6645;
  assign n7686 = ~n2091 & ~n6652;
  assign n7687 = pi330 & ~n7686;
  assign n7688 = ~n7685 & ~n7687;
  assign n7689 = pi330 & n2464;
  assign n7690 = n6178 & ~n7689;
  assign n7691 = ~n7688 & n7690;
  assign n7692 = ~n6167 & ~n6651;
  assign n7693 = ~n6652 & ~n7692;
  assign n7694 = n2091 & ~n7693;
  assign n7695 = pi330 & n7694;
  assign n7696 = ~n6178 & n7689;
  assign n7697 = ~n7695 & n7696;
  assign n7698 = ~n7691 & ~n7697;
  assign n7699 = ~n7263 & ~n7698;
  assign n7700 = n6178 & n7689;
  assign n7701 = ~n7695 & n7700;
  assign n7702 = ~n6178 & ~n7689;
  assign n7703 = ~n7688 & n7702;
  assign n7704 = ~n7701 & ~n7703;
  assign n7705 = ~n7253 & ~n7704;
  assign n7706 = ~n7689 & n7695;
  assign n7707 = n7688 & n7689;
  assign n7708 = ~n7695 & n7707;
  assign n7709 = ~n7706 & ~n7708;
  assign n7710 = ~n7705 & n7709;
  assign n7711 = ~n7699 & n7710;
  assign n7712 = pi329 & n2887;
  assign n7713 = ~n7711 & n7712;
  assign n7714 = n7711 & ~n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = ~n7684 & ~n7715;
  assign n7717 = n7311 & n7681;
  assign n7718 = ~n7311 & ~n7681;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = n7711 & n7712;
  assign n7721 = ~n7711 & ~n7712;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = ~n7719 & ~n7722;
  assign n7724 = ~n7716 & ~n7723;
  assign n7725 = ~n7310 & ~n7724;
  assign n7726 = n7303 & n7307;
  assign n7727 = ~n7303 & ~n7307;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = ~n7715 & ~n7719;
  assign n7730 = ~n7684 & ~n7722;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = ~n7728 & ~n7731;
  assign n7733 = ~n7725 & ~n7732;
  assign n7734 = ~n7283 & n7733;
  assign n7735 = n7283 & ~n7733;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = pi333 & n1442;
  assign n7738 = n6679 & ~n6698;
  assign n7739 = ~n6695 & ~n7738;
  assign n7740 = n1729 & n7739;
  assign n7741 = pi332 & n7740;
  assign n7742 = pi332 & n1729;
  assign n7743 = ~n7739 & ~n7742;
  assign n7744 = ~n7741 & ~n7743;
  assign n7745 = n7737 & ~n7744;
  assign n7746 = ~n7737 & n7744;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = ~n7736 & ~n7747;
  assign n7749 = n7283 & n7733;
  assign n7750 = ~n7283 & ~n7733;
  assign n7751 = ~n7749 & ~n7750;
  assign n7752 = ~n7737 & ~n7744;
  assign n7753 = n7737 & n7744;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = ~n7751 & ~n7754;
  assign n7756 = ~n7748 & ~n7755;
  assign n7757 = ~n7282 & ~n7756;
  assign n7758 = n7270 & n7279;
  assign n7759 = ~n7270 & ~n7279;
  assign n7760 = ~n7758 & ~n7759;
  assign n7761 = ~n7747 & ~n7751;
  assign n7762 = ~n7736 & ~n7754;
  assign n7763 = ~n7761 & ~n7762;
  assign n7764 = ~n7760 & ~n7763;
  assign n7765 = ~n7757 & ~n7764;
  assign n7766 = ~n7250 & ~n7765;
  assign n7767 = n7250 & n7765;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = ~n1154 & ~n6714;
  assign n7770 = n1154 & n6714;
  assign n7771 = ~n6095 & ~n7770;
  assign n7772 = n1156 & n7771;
  assign n7773 = ~n7769 & ~n7772;
  assign n7774 = ~n1256 & ~n7773;
  assign n7775 = pi334 & n7774;
  assign n7776 = n1256 & ~n7769;
  assign n7777 = ~n7772 & n7776;
  assign n7778 = pi334 & ~n7777;
  assign n7779 = ~n7775 & n7778;
  assign n7780 = ~n1154 & ~n7779;
  assign n7781 = pi335 & n7780;
  assign n7782 = pi335 & ~n1154;
  assign n7783 = n7778 & ~n7782;
  assign n7784 = ~n7775 & n7783;
  assign n7785 = ~n7781 & ~n7784;
  assign n7786 = ~n7768 & ~n7785;
  assign n7787 = n7250 & ~n7765;
  assign n7788 = ~n7250 & n7765;
  assign n7789 = ~n7787 & ~n7788;
  assign n7790 = n7779 & n7782;
  assign n7791 = ~n7779 & ~n7782;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = ~n7789 & ~n7792;
  assign n7794 = ~n7786 & ~n7793;
  assign n7795 = n7247 & n7794;
  assign n7796 = ~n7247 & ~n7794;
  assign n7797 = ~n7795 & ~n7796;
  assign n7798 = pi272 & pi336;
  assign n7799 = n1156 & n7798;
  assign n7800 = pi336 & n1156;
  assign n7801 = ~pi272 & ~n7800;
  assign n7802 = ~n7799 & ~n7801;
  assign n7803 = ~n7797 & ~n7802;
  assign n7804 = ~n7247 & n7794;
  assign n7805 = n7247 & ~n7794;
  assign n7806 = ~n7804 & ~n7805;
  assign n7807 = pi272 & ~n7800;
  assign n7808 = ~pi272 & pi336;
  assign n7809 = n1156 & n7808;
  assign n7810 = ~n7807 & ~n7809;
  assign n7811 = ~n7806 & ~n7810;
  assign n7812 = ~n7803 & ~n7811;
  assign n7813 = ~n7245 & n7812;
  assign n7814 = n7245 & ~n7812;
  assign n7815 = ~n7813 & ~n7814;
  assign n7816 = pi307 & ~n7815;
  assign n7817 = pi128 & n7816;
  assign n7818 = pi128 & pi307;
  assign n7819 = n7245 & n7812;
  assign n7820 = ~n7245 & ~n7812;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~n7818 & ~n7821;
  assign n7823 = ~n7817 & ~n7822;
  assign n7824 = ~n6968 & n6969;
  assign n7825 = ~n6970 & ~n7824;
  assign n7826 = ~n6975 & ~n7825;
  assign n7827 = ~n6976 & ~n7826;
  assign n7828 = n7823 & ~n7827;
  assign n7829 = ~n7823 & n7827;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = ~n831 & ~n7830;
  assign n7832 = ~n6990 & ~n7831;
  assign n7833 = pi161 & ~n7832;
  assign n7834 = pi078 & ~pi161;
  assign n7835 = ~n7833 & ~n7834;
  assign po207 = ~pi160 & ~n7835;
  assign n7837 = pi273 & n831;
  assign n7838 = pi309 & n1553;
  assign n7839 = ~n1533 & ~n7188;
  assign n7840 = n1533 & n7188;
  assign n7841 = ~n7006 & ~n7840;
  assign n7842 = ~n7839 & ~n7841;
  assign n7843 = n1840 & ~n7842;
  assign n7844 = ~n1840 & ~n7190;
  assign n7845 = n1533 & n7844;
  assign n7846 = ~n7843 & ~n7845;
  assign n7847 = pi311 & ~n7846;
  assign n7848 = pi311 & n1840;
  assign n7849 = n7188 & ~n7848;
  assign n7850 = n7006 & n7849;
  assign n7851 = ~n7847 & ~n7850;
  assign n7852 = pi313 & n2574;
  assign n7853 = pi316 & n4086;
  assign n7854 = ~n4086 & n7092;
  assign n7855 = ~n6830 & ~n7854;
  assign n7856 = n3552 & n7855;
  assign n7857 = ~n6829 & n7092;
  assign n7858 = n4086 & ~n7857;
  assign n7859 = ~n7856 & ~n7858;
  assign n7860 = pi317 & ~n7859;
  assign n7861 = ~n7104 & ~n7860;
  assign n7862 = ~pi143 & n7035;
  assign n7863 = pi143 & ~n7035;
  assign n7864 = ~pi142 & n7863;
  assign n7865 = ~n7862 & ~n7864;
  assign n7866 = pi141 & ~n7865;
  assign n7867 = ~pi143 & ~n7035;
  assign n7868 = pi143 & n7035;
  assign n7869 = pi142 & n7868;
  assign n7870 = ~n7867 & ~n7869;
  assign n7871 = ~pi141 & ~n7870;
  assign n7872 = ~pi143 & ~n7042;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = ~n7866 & n7873;
  assign n7875 = pi321 & n7874;
  assign n7876 = ~n7045 & n7051;
  assign n7877 = n6777 & ~n7876;
  assign n7878 = pi320 & n7877;
  assign n7879 = n7044 & ~n7051;
  assign n7880 = pi321 & n7879;
  assign n7881 = ~n7878 & ~n7880;
  assign n7882 = pi320 & n7044;
  assign n7883 = ~n7881 & ~n7882;
  assign n7884 = n7044 & n7881;
  assign n7885 = pi320 & n7884;
  assign n7886 = ~n7883 & ~n7885;
  assign n7887 = ~n7875 & ~n7886;
  assign n7888 = n7881 & ~n7882;
  assign n7889 = n7044 & ~n7881;
  assign n7890 = pi320 & n7889;
  assign n7891 = ~n7888 & ~n7890;
  assign n7892 = n7874 & ~n7891;
  assign n7893 = pi321 & n7892;
  assign n7894 = ~n7887 & ~n7893;
  assign n7895 = n5463 & ~n7069;
  assign n7896 = pi319 & n7895;
  assign n7897 = ~n7068 & ~n7896;
  assign n7898 = ~n7894 & ~n7897;
  assign n7899 = n7894 & n7897;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = n6777 & ~n7900;
  assign n7902 = pi319 & n7901;
  assign n7903 = pi319 & n6777;
  assign n7904 = n7894 & ~n7897;
  assign n7905 = ~n7894 & n7897;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = ~n7903 & ~n7906;
  assign n7908 = ~n7902 & ~n7907;
  assign n7909 = pi318 & n5463;
  assign n7910 = ~n7908 & ~n7909;
  assign n7911 = n5463 & n7908;
  assign n7912 = pi318 & n7911;
  assign n7913 = ~n7910 & ~n7912;
  assign n7914 = n4772 & ~n7082;
  assign n7915 = pi318 & n7914;
  assign n7916 = ~n7083 & ~n7915;
  assign n7917 = ~n7913 & n7916;
  assign n7918 = n7913 & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = n4772 & ~n7919;
  assign n7921 = pi317 & n7920;
  assign n7922 = pi317 & n4772;
  assign n7923 = ~n7918 & ~n7922;
  assign n7924 = ~n7917 & n7923;
  assign n7925 = ~n7921 & ~n7924;
  assign n7926 = ~n7861 & ~n7925;
  assign n7927 = n7861 & ~n7924;
  assign n7928 = ~n7921 & n7927;
  assign n7929 = ~n7926 & ~n7928;
  assign n7930 = ~n7853 & ~n7929;
  assign n7931 = n7861 & ~n7925;
  assign n7932 = ~n7861 & ~n7924;
  assign n7933 = ~n7921 & n7932;
  assign n7934 = ~n7931 & ~n7933;
  assign n7935 = n4086 & ~n7934;
  assign n7936 = pi316 & n7935;
  assign n7937 = ~n7930 & ~n7936;
  assign n7938 = n3552 & ~n7131;
  assign n7939 = pi316 & n7938;
  assign n7940 = ~n7130 & ~n7939;
  assign n7941 = n7937 & n7940;
  assign n7942 = ~n7937 & ~n7940;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = n3552 & ~n7943;
  assign n7945 = pi315 & n7944;
  assign n7946 = pi315 & n3552;
  assign n7947 = ~n7937 & n7940;
  assign n7948 = n7937 & ~n7940;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = ~n7946 & ~n7949;
  assign n7951 = ~n7945 & ~n7950;
  assign n7952 = ~n7145 & n7151;
  assign n7953 = n7145 & ~n7151;
  assign n7954 = ~n7140 & ~n7953;
  assign n7955 = ~n7952 & ~n7954;
  assign n7956 = n7951 & n7955;
  assign n7957 = ~n7951 & ~n7955;
  assign n7958 = ~n7956 & ~n7957;
  assign n7959 = pi314 & n3012;
  assign n7960 = ~n7164 & ~n7959;
  assign n7961 = ~n7158 & n7960;
  assign n7962 = ~n7158 & ~n7164;
  assign n7963 = n7959 & ~n7962;
  assign n7964 = ~n7961 & ~n7963;
  assign n7965 = ~n7958 & ~n7964;
  assign n7966 = n7951 & ~n7955;
  assign n7967 = ~n7951 & n7955;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = ~n7164 & n7959;
  assign n7970 = ~n7158 & n7969;
  assign n7971 = ~n7959 & ~n7962;
  assign n7972 = ~n7970 & ~n7971;
  assign n7973 = ~n7968 & ~n7972;
  assign n7974 = ~n7965 & ~n7973;
  assign n7975 = ~n7852 & n7974;
  assign n7976 = n7852 & ~n7974;
  assign n7977 = ~n7975 & ~n7976;
  assign n7978 = pi312 & n2183;
  assign n7979 = ~n7015 & n7166;
  assign n7980 = n7015 & ~n7166;
  assign n7981 = n7016 & ~n7980;
  assign n7982 = ~n7979 & ~n7981;
  assign n7983 = n7978 & ~n7982;
  assign n7984 = ~n7016 & ~n7979;
  assign n7985 = ~n7980 & ~n7984;
  assign n7986 = ~n7978 & ~n7985;
  assign n7987 = ~n7983 & ~n7986;
  assign n7988 = ~n7977 & ~n7987;
  assign n7989 = ~n7852 & ~n7974;
  assign n7990 = n7852 & n7974;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = ~n7978 & ~n7982;
  assign n7993 = n7978 & ~n7985;
  assign n7994 = ~n7992 & ~n7993;
  assign n7995 = ~n7991 & ~n7994;
  assign n7996 = ~n7988 & ~n7995;
  assign n7997 = n7170 & ~n7183;
  assign n7998 = ~n7170 & n7183;
  assign n7999 = ~n7174 & ~n7998;
  assign n8000 = ~n7997 & ~n7999;
  assign n8001 = ~n7996 & ~n8000;
  assign n8002 = n7996 & n8000;
  assign n8003 = ~n8001 & ~n8002;
  assign n8004 = n7851 & n8003;
  assign n8005 = ~n7851 & ~n8003;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = pi310 & n1533;
  assign n8008 = ~n6999 & ~n7204;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~n7201 & n8009;
  assign n8011 = ~n7201 & ~n8008;
  assign n8012 = n8007 & ~n8011;
  assign n8013 = ~n8010 & ~n8012;
  assign n8014 = ~n8006 & ~n8013;
  assign n8015 = n7851 & ~n8003;
  assign n8016 = ~n7851 & n8003;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = n8007 & ~n8008;
  assign n8019 = ~n7201 & n8018;
  assign n8020 = ~n8007 & ~n8011;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = ~n8017 & ~n8021;
  assign n8023 = ~n8014 & ~n8022;
  assign n8024 = ~n7838 & ~n8023;
  assign n8025 = n7838 & n8023;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = pi308 & n1515;
  assign n8028 = ~n7209 & n7232;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = ~n7222 & n8029;
  assign n8031 = ~n7222 & ~n8028;
  assign n8032 = n8027 & ~n8031;
  assign n8033 = ~n8030 & ~n8032;
  assign n8034 = ~n8026 & ~n8033;
  assign n8035 = ~n7838 & n8023;
  assign n8036 = n7838 & ~n8023;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = n8027 & ~n8028;
  assign n8039 = ~n7222 & n8038;
  assign n8040 = ~n8027 & ~n8031;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = ~n8037 & ~n8041;
  assign n8043 = ~n8034 & ~n8042;
  assign n8044 = n6972 & n6991;
  assign n8045 = ~n6972 & ~n6991;
  assign n8046 = ~n7209 & ~n7233;
  assign n8047 = n7209 & n7233;
  assign n8048 = ~n8046 & ~n8047;
  assign n8049 = ~n8045 & ~n8048;
  assign n8050 = ~n8044 & ~n8049;
  assign n8051 = n8043 & ~n8050;
  assign n8052 = ~n8043 & n8050;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = pi129 & ~n6965;
  assign n8055 = ~pi128 & ~n8054;
  assign n8056 = ~n5614 & n6965;
  assign n8057 = pi128 & ~n6965;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = pi129 & ~n8058;
  assign n8060 = ~pi129 & n7214;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = ~n8055 & n8061;
  assign n8063 = pi130 & ~n8062;
  assign n8064 = ~pi128 & n8054;
  assign n8065 = pi128 & ~n7216;
  assign n8066 = ~n8064 & ~n8065;
  assign n8067 = ~pi130 & ~n8066;
  assign n8068 = ~n8063 & ~n8067;
  assign n8069 = pi309 & ~n8068;
  assign n8070 = ~n7209 & ~n8069;
  assign n8071 = n7209 & n8069;
  assign n8072 = ~n8070 & ~n8071;
  assign n8073 = ~n8044 & ~n8045;
  assign n8074 = ~n8072 & ~n8073;
  assign n8075 = n7209 & ~n8069;
  assign n8076 = ~n7209 & n8069;
  assign n8077 = ~n8075 & ~n8076;
  assign n8078 = n6972 & ~n6991;
  assign n8079 = ~n6972 & n6991;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = ~n8077 & ~n8080;
  assign n8082 = ~n8074 & ~n8081;
  assign n8083 = pi307 & ~n8082;
  assign n8084 = pi128 & n8083;
  assign n8085 = pi128 & pi306;
  assign n8086 = pi307 & ~n1568;
  assign n8087 = ~n8085 & ~n8086;
  assign n8088 = n8085 & n8086;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~n8084 & ~n8089;
  assign n8091 = pi129 & n8085;
  assign n8092 = ~pi129 & ~n8085;
  assign n8093 = ~n8091 & ~n8092;
  assign n8094 = n8084 & ~n8093;
  assign n8095 = ~n8090 & ~n8094;
  assign n8096 = ~n8053 & ~n8095;
  assign n8097 = n8043 & n8050;
  assign n8098 = ~n8043 & ~n8050;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = n8085 & ~n8086;
  assign n8101 = ~n8085 & n8086;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n8084 & ~n8102;
  assign n8104 = pi129 & ~n8085;
  assign n8105 = ~pi129 & n8085;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = n8084 & ~n8106;
  assign n8108 = ~n8103 & ~n8107;
  assign n8109 = ~n8099 & ~n8108;
  assign n8110 = ~n8096 & ~n8109;
  assign n8111 = n1256 & ~n7773;
  assign n8112 = ~n6142 & ~n7769;
  assign n8113 = ~n7770 & ~n8112;
  assign n8114 = ~n1256 & ~n8113;
  assign n8115 = ~n8111 & ~n8114;
  assign n8116 = pi334 & ~n8115;
  assign n8117 = ~n7765 & ~n8116;
  assign n8118 = n7765 & n8116;
  assign n8119 = ~n8117 & ~n8118;
  assign n8120 = ~n7250 & ~n7782;
  assign n8121 = n7250 & n7782;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n8119 & ~n8122;
  assign n8124 = n7765 & ~n8116;
  assign n8125 = ~n7765 & n8116;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = n7250 & ~n7782;
  assign n8128 = ~n7250 & n7782;
  assign n8129 = ~n8127 & ~n8128;
  assign n8130 = ~n8126 & ~n8129;
  assign n8131 = ~n8123 & ~n8130;
  assign n8132 = n1156 & ~n8131;
  assign n8133 = pi336 & n8132;
  assign n8134 = n1154 & n8133;
  assign n8135 = ~n1154 & ~n8133;
  assign n8136 = pi336 & n8135;
  assign n8137 = ~n8134 & ~n8136;
  assign n8138 = n7270 & n7733;
  assign n8139 = ~n7270 & ~n7733;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = ~n7279 & n7737;
  assign n8142 = n7283 & ~n7744;
  assign n8143 = ~n7283 & n7744;
  assign n8144 = ~n8142 & ~n8143;
  assign n8145 = ~n8141 & ~n8144;
  assign n8146 = ~n8140 & n8145;
  assign n8147 = ~n7270 & n7733;
  assign n8148 = n7270 & ~n7733;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = ~n7283 & ~n7744;
  assign n8151 = n7283 & n7744;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = ~n8141 & ~n8152;
  assign n8154 = ~n8149 & n8153;
  assign n8155 = n7279 & ~n7737;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n8146 & n8156;
  assign n8158 = ~n7765 & ~n7779;
  assign n8159 = n7765 & n7779;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = ~n8120 & ~n8160;
  assign n8162 = ~n8121 & ~n8161;
  assign n8163 = n8157 & n8162;
  assign n8164 = ~n8157 & ~n8162;
  assign n8165 = ~n8163 & ~n8164;
  assign n8166 = pi333 & n1729;
  assign n8167 = ~n7303 & n7311;
  assign n8168 = n7303 & ~n7311;
  assign n8169 = ~n7681 & ~n8168;
  assign n8170 = ~n8167 & ~n8169;
  assign n8171 = ~n7307 & n7712;
  assign n8172 = ~n7303 & ~n7681;
  assign n8173 = n7303 & n7681;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = n7311 & ~n8174;
  assign n8176 = n7303 & ~n7681;
  assign n8177 = ~n7303 & n7681;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = ~n7311 & ~n8178;
  assign n8180 = ~n8175 & ~n8179;
  assign n8181 = n7307 & ~n7712;
  assign n8182 = ~n8180 & ~n8181;
  assign n8183 = ~n8171 & ~n8182;
  assign n8184 = n8170 & ~n8183;
  assign n8185 = ~n8170 & n8183;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = pi329 & n4596;
  assign n8188 = ~n7326 & n7660;
  assign n8189 = n7326 & ~n7660;
  assign n8190 = ~n7667 & ~n8189;
  assign n8191 = ~n8188 & ~n8190;
  assign n8192 = ~n7326 & ~n7655;
  assign n8193 = n7326 & n7655;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = ~n7330 & n7659;
  assign n8196 = ~n7642 & n7660;
  assign n8197 = n7642 & ~n7660;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = ~n8195 & ~n8198;
  assign n8200 = ~n8194 & n8199;
  assign n8201 = ~n7326 & n7655;
  assign n8202 = n7326 & ~n7655;
  assign n8203 = ~n8201 & ~n8202;
  assign n8204 = n7642 & n7660;
  assign n8205 = ~n7642 & ~n7660;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = ~n8195 & ~n8206;
  assign n8208 = ~n8203 & n8207;
  assign n8209 = n7330 & ~n7659;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8200 & n8210;
  assign n8212 = n8191 & n8211;
  assign n8213 = ~n8191 & ~n8211;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~n7339 & ~n7616;
  assign n8216 = ~n7619 & ~n8215;
  assign n8217 = ~n7343 & n7622;
  assign n8218 = ~n7339 & ~n7620;
  assign n8219 = n7339 & ~n7619;
  assign n8220 = ~n7616 & n8219;
  assign n8221 = ~n8218 & ~n8220;
  assign n8222 = n7343 & ~n7622;
  assign n8223 = ~n8221 & ~n8222;
  assign n8224 = ~n8217 & ~n8223;
  assign n8225 = ~n8216 & n8224;
  assign n8226 = n8216 & ~n8224;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = pi141 & pi260;
  assign n8229 = ~n7585 & n7596;
  assign n8230 = ~n8228 & ~n8229;
  assign n8231 = ~n7574 & n8230;
  assign n8232 = ~n7568 & ~n7585;
  assign n8233 = ~n7574 & ~n8232;
  assign n8234 = pi260 & ~n8233;
  assign n8235 = pi141 & n8234;
  assign n8236 = ~n8231 & ~n8235;
  assign n8237 = pi131 & pi270;
  assign n8238 = ~n7387 & ~n7388;
  assign n8239 = ~n6252 & n8238;
  assign n8240 = ~n7386 & ~n7389;
  assign n8241 = ~n7383 & n8240;
  assign n8242 = ~n8239 & ~n8241;
  assign n8243 = pi269 & ~n8242;
  assign n8244 = pi131 & n8243;
  assign n8245 = ~n7371 & n7372;
  assign n8246 = pi128 & pi273;
  assign n8247 = pi272 & ~n8246;
  assign n8248 = pi129 & n8247;
  assign n8249 = pi129 & pi272;
  assign n8250 = pi273 & ~n8249;
  assign n8251 = pi128 & n8250;
  assign n8252 = ~n8248 & ~n8251;
  assign n8253 = ~pi129 & n8252;
  assign n8254 = pi130 & pi271;
  assign n8255 = n8253 & n8254;
  assign n8256 = pi271 & ~n1328;
  assign n8257 = ~n8252 & ~n8256;
  assign n8258 = ~n8255 & ~n8257;
  assign n8259 = ~n8245 & ~n8258;
  assign n8260 = ~pi130 & ~n8252;
  assign n8261 = n8252 & n8254;
  assign n8262 = ~n8260 & ~n8261;
  assign n8263 = ~n7372 & ~n8262;
  assign n8264 = n7371 & n8263;
  assign n8265 = ~pi129 & ~n7372;
  assign n8266 = pi130 & ~n8265;
  assign n8267 = ~n8252 & n8266;
  assign n8268 = n1319 & n8252;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = pi271 & ~n8269;
  assign n8271 = n8252 & ~n8254;
  assign n8272 = n7372 & n8271;
  assign n8273 = ~n8270 & ~n8272;
  assign n8274 = ~n7371 & ~n8273;
  assign n8275 = pi130 & ~n8252;
  assign n8276 = ~pi130 & n8252;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = pi271 & ~n8277;
  assign n8279 = pi129 & n8278;
  assign n8280 = n7372 & n8279;
  assign n8281 = ~n8274 & ~n8280;
  assign n8282 = ~n8264 & n8281;
  assign n8283 = ~n8259 & n8282;
  assign n8284 = ~n7383 & ~n7389;
  assign n8285 = ~n8283 & ~n8284;
  assign n8286 = ~n7386 & n8285;
  assign n8287 = ~n7386 & ~n8284;
  assign n8288 = n8283 & ~n8287;
  assign n8289 = ~n8286 & ~n8288;
  assign n8290 = ~n7392 & ~n8241;
  assign n8291 = ~n8239 & n8290;
  assign n8292 = n7407 & ~n8291;
  assign n8293 = ~n8289 & ~n8292;
  assign n8294 = ~n8244 & n8293;
  assign n8295 = ~n8244 & ~n8292;
  assign n8296 = n8289 & ~n8295;
  assign n8297 = ~n8294 & ~n8296;
  assign n8298 = ~n8237 & ~n8297;
  assign n8299 = n8289 & ~n8292;
  assign n8300 = ~n8244 & n8299;
  assign n8301 = ~n8289 & ~n8295;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = pi270 & ~n8302;
  assign n8304 = pi131 & n8303;
  assign n8305 = ~n8298 & ~n8304;
  assign n8306 = n7411 & ~n7422;
  assign n8307 = ~n7411 & n7422;
  assign n8308 = ~n7413 & ~n8307;
  assign n8309 = ~n8306 & ~n8308;
  assign n8310 = n8305 & n8309;
  assign n8311 = ~n8305 & ~n8309;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = pi133 & pi268;
  assign n8314 = pi132 & pi269;
  assign n8315 = n8313 & n8314;
  assign n8316 = ~n8313 & ~n8314;
  assign n8317 = ~n8315 & ~n8316;
  assign n8318 = ~n8312 & ~n8317;
  assign n8319 = ~n8305 & n8309;
  assign n8320 = n8305 & ~n8309;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = pi268 & ~n8314;
  assign n8323 = pi133 & n8322;
  assign n8324 = pi269 & ~n8313;
  assign n8325 = pi132 & n8324;
  assign n8326 = ~n8323 & ~n8325;
  assign n8327 = ~n8321 & ~n8326;
  assign n8328 = ~n8318 & ~n8327;
  assign n8329 = ~n7443 & ~n7447;
  assign n8330 = ~n7448 & ~n8329;
  assign n8331 = n8328 & n8330;
  assign n8332 = ~n8328 & ~n8330;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = pi134 & pi267;
  assign n8335 = n7427 & ~n7440;
  assign n8336 = ~n7436 & n8335;
  assign n8337 = ~n7427 & ~n7443;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = ~n7367 & ~n8338;
  assign n8340 = ~n7427 & ~n7440;
  assign n8341 = ~n7436 & n8340;
  assign n8342 = n7427 & ~n7443;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = pi267 & ~n8343;
  assign n8345 = pi133 & n8344;
  assign n8346 = ~n8339 & ~n8345;
  assign n8347 = ~n7459 & ~n8346;
  assign n8348 = n7459 & n8346;
  assign n8349 = n7437 & ~n8348;
  assign n8350 = ~n8347 & ~n8349;
  assign n8351 = n8334 & ~n8350;
  assign n8352 = ~n7437 & ~n8347;
  assign n8353 = ~n8348 & ~n8352;
  assign n8354 = ~n8334 & ~n8353;
  assign n8355 = ~n8351 & ~n8354;
  assign n8356 = ~n8333 & ~n8355;
  assign n8357 = n8328 & ~n8330;
  assign n8358 = ~n8328 & n8330;
  assign n8359 = ~n8357 & ~n8358;
  assign n8360 = ~n8334 & ~n8350;
  assign n8361 = n8334 & ~n8353;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = ~n8359 & ~n8362;
  assign n8364 = ~n8356 & ~n8363;
  assign n8365 = ~n7462 & ~n7463;
  assign n8366 = n7462 & n7463;
  assign n8367 = ~n7468 & ~n8366;
  assign n8368 = ~n8365 & ~n8367;
  assign n8369 = ~n8364 & n8368;
  assign n8370 = n8364 & ~n8368;
  assign n8371 = ~n8369 & ~n8370;
  assign n8372 = pi136 & pi265;
  assign n8373 = pi135 & pi266;
  assign n8374 = n8372 & n8373;
  assign n8375 = ~n8372 & ~n8373;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = ~n8371 & ~n8376;
  assign n8378 = n8364 & n8368;
  assign n8379 = ~n8364 & ~n8368;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = pi265 & ~n8373;
  assign n8382 = pi136 & n8381;
  assign n8383 = pi266 & ~n8372;
  assign n8384 = pi135 & n8383;
  assign n8385 = ~n8382 & ~n8384;
  assign n8386 = ~n8380 & ~n8385;
  assign n8387 = ~n8377 & ~n8386;
  assign n8388 = ~n7495 & ~n7499;
  assign n8389 = ~n7500 & ~n8388;
  assign n8390 = n8387 & n8389;
  assign n8391 = ~n8387 & ~n8389;
  assign n8392 = ~n8390 & ~n8391;
  assign n8393 = pi137 & pi264;
  assign n8394 = n7479 & ~n7492;
  assign n8395 = ~n7488 & n8394;
  assign n8396 = ~n7479 & ~n7495;
  assign n8397 = ~n8395 & ~n8396;
  assign n8398 = ~n7366 & ~n8397;
  assign n8399 = ~n7479 & ~n7492;
  assign n8400 = ~n7488 & n8399;
  assign n8401 = n7479 & ~n7495;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = pi264 & ~n8402;
  assign n8404 = pi136 & n8403;
  assign n8405 = ~n8398 & ~n8404;
  assign n8406 = ~n7511 & ~n8405;
  assign n8407 = n7511 & n8405;
  assign n8408 = n7489 & ~n8407;
  assign n8409 = ~n8406 & ~n8408;
  assign n8410 = n8393 & ~n8409;
  assign n8411 = ~n7489 & ~n8406;
  assign n8412 = ~n8407 & ~n8411;
  assign n8413 = ~n8393 & ~n8412;
  assign n8414 = ~n8410 & ~n8413;
  assign n8415 = ~n8392 & ~n8414;
  assign n8416 = n8387 & ~n8389;
  assign n8417 = ~n8387 & n8389;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = ~n8393 & ~n8409;
  assign n8420 = n8393 & ~n8412;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = ~n8418 & ~n8421;
  assign n8423 = ~n8415 & ~n8422;
  assign n8424 = ~n7515 & ~n7526;
  assign n8425 = n7515 & n7526;
  assign n8426 = ~n7520 & ~n8425;
  assign n8427 = ~n8424 & ~n8426;
  assign n8428 = ~n8423 & n8427;
  assign n8429 = n8423 & ~n8427;
  assign n8430 = ~n8428 & ~n8429;
  assign n8431 = pi139 & pi262;
  assign n8432 = pi138 & pi263;
  assign n8433 = n8431 & n8432;
  assign n8434 = ~n8431 & ~n8432;
  assign n8435 = ~n8433 & ~n8434;
  assign n8436 = ~n8430 & ~n8435;
  assign n8437 = n8423 & n8427;
  assign n8438 = ~n8423 & ~n8427;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = pi262 & ~n8432;
  assign n8441 = pi139 & n8440;
  assign n8442 = pi263 & ~n8431;
  assign n8443 = pi138 & n8442;
  assign n8444 = ~n8441 & ~n8443;
  assign n8445 = ~n8439 & ~n8444;
  assign n8446 = ~n8436 & ~n8445;
  assign n8447 = ~n7544 & ~n7551;
  assign n8448 = ~n7539 & n8447;
  assign n8449 = ~n7552 & ~n8448;
  assign n8450 = n8446 & n8449;
  assign n8451 = ~n8446 & ~n8449;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = pi140 & pi261;
  assign n8454 = ~n7531 & ~n7544;
  assign n8455 = ~n7539 & n8454;
  assign n8456 = n7531 & ~n7547;
  assign n8457 = ~n8455 & ~n8456;
  assign n8458 = ~n7365 & ~n8457;
  assign n8459 = n7531 & ~n7544;
  assign n8460 = ~n7539 & n8459;
  assign n8461 = ~n7531 & ~n7547;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = pi261 & ~n8462;
  assign n8464 = pi139 & n8463;
  assign n8465 = ~n8458 & ~n8464;
  assign n8466 = ~n7565 & n8465;
  assign n8467 = n7565 & ~n8465;
  assign n8468 = n7540 & ~n8467;
  assign n8469 = ~n8466 & ~n8468;
  assign n8470 = n8453 & ~n8469;
  assign n8471 = ~n7540 & ~n8466;
  assign n8472 = ~n8467 & ~n8471;
  assign n8473 = ~n8453 & ~n8472;
  assign n8474 = ~n8470 & ~n8473;
  assign n8475 = ~n8452 & ~n8474;
  assign n8476 = n8446 & ~n8449;
  assign n8477 = ~n8446 & n8449;
  assign n8478 = ~n8476 & ~n8477;
  assign n8479 = ~n8453 & ~n8469;
  assign n8480 = n8453 & ~n8472;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n8478 & ~n8481;
  assign n8483 = ~n8475 & ~n8482;
  assign n8484 = ~n8236 & n8483;
  assign n8485 = n8236 & ~n8483;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = ~n7586 & ~n7596;
  assign n8488 = ~n7574 & n8232;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = pi258 & ~n8489;
  assign n8491 = pi142 & n8490;
  assign n8492 = pi142 & pi259;
  assign n8493 = n8491 & n8492;
  assign n8494 = ~n8491 & ~n8492;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = pi258 & ~n8495;
  assign n8497 = pi143 & n8496;
  assign n8498 = pi143 & pi258;
  assign n8499 = ~n8491 & n8492;
  assign n8500 = n8491 & ~n8492;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = ~n8498 & ~n8501;
  assign n8503 = ~n8497 & ~n8502;
  assign n8504 = ~n8486 & ~n8503;
  assign n8505 = n8236 & n8483;
  assign n8506 = ~n8236 & ~n8483;
  assign n8507 = ~n8505 & ~n8506;
  assign n8508 = pi258 & ~n8501;
  assign n8509 = pi143 & n8508;
  assign n8510 = ~n8495 & ~n8498;
  assign n8511 = ~n8509 & ~n8510;
  assign n8512 = ~n8507 & ~n8511;
  assign n8513 = ~n8504 & ~n8512;
  assign n8514 = n7605 & ~n8513;
  assign n8515 = ~n7605 & n8513;
  assign n8516 = n7601 & n8515;
  assign n8517 = ~n8514 & ~n8516;
  assign n8518 = ~n7364 & ~n8517;
  assign n8519 = ~n7605 & ~n8513;
  assign n8520 = n7605 & n8513;
  assign n8521 = ~n7601 & n8520;
  assign n8522 = ~n8519 & ~n8521;
  assign n8523 = n7364 & ~n8522;
  assign n8524 = ~n7608 & ~n8513;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = ~n8518 & n8525;
  assign n8527 = pi322 & ~n8526;
  assign n8528 = pi323 & ~n7614;
  assign n8529 = ~n8527 & ~n8528;
  assign n8530 = n7364 & n7610;
  assign n8531 = ~n7609 & ~n8530;
  assign n8532 = ~n8513 & ~n8531;
  assign n8533 = n7364 & ~n7601;
  assign n8534 = n8520 & n8533;
  assign n8535 = ~n8532 & ~n8534;
  assign n8536 = pi323 & ~n8535;
  assign n8537 = pi322 & n8536;
  assign n8538 = ~n8529 & ~n8537;
  assign n8539 = pi325 & n5973;
  assign n8540 = pi324 & n6556;
  assign n8541 = n8539 & n8540;
  assign n8542 = ~n8539 & ~n8540;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = ~n8538 & ~n8543;
  assign n8545 = ~n8539 & n8540;
  assign n8546 = n8539 & ~n8540;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = ~n8537 & ~n8547;
  assign n8549 = ~n8529 & n8548;
  assign n8550 = ~n8544 & ~n8549;
  assign n8551 = ~n8227 & ~n8550;
  assign n8552 = ~n8216 & ~n8224;
  assign n8553 = n8216 & n8224;
  assign n8554 = ~n8552 & ~n8553;
  assign n8555 = ~n8538 & ~n8547;
  assign n8556 = ~n8537 & ~n8543;
  assign n8557 = ~n8529 & n8556;
  assign n8558 = ~n8555 & ~n8557;
  assign n8559 = ~n8554 & ~n8558;
  assign n8560 = ~n8551 & ~n8559;
  assign n8561 = n7621 & ~n7655;
  assign n8562 = ~n7622 & ~n8221;
  assign n8563 = n7339 & ~n7620;
  assign n8564 = ~n7339 & ~n7619;
  assign n8565 = ~n7616 & n8564;
  assign n8566 = ~n8563 & ~n8565;
  assign n8567 = n5973 & ~n8566;
  assign n8568 = pi324 & n8567;
  assign n8569 = ~n8562 & ~n8568;
  assign n8570 = n7343 & ~n8569;
  assign n8571 = ~n7343 & n8569;
  assign n8572 = ~n8570 & ~n8571;
  assign n8573 = ~n7621 & n7655;
  assign n8574 = ~n8572 & ~n8573;
  assign n8575 = ~n8561 & ~n8574;
  assign n8576 = n8560 & n8575;
  assign n8577 = ~n8560 & ~n8575;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = pi327 & n5714;
  assign n8580 = pi326 & n5732;
  assign n8581 = n8579 & n8580;
  assign n8582 = ~n8579 & ~n8580;
  assign n8583 = ~n8581 & ~n8582;
  assign n8584 = ~n8578 & ~n8583;
  assign n8585 = ~n8560 & n8575;
  assign n8586 = n8560 & ~n8575;
  assign n8587 = ~n8585 & ~n8586;
  assign n8588 = ~n8579 & n8580;
  assign n8589 = n8579 & ~n8580;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n8587 & ~n8590;
  assign n8592 = ~n8584 & ~n8591;
  assign n8593 = ~n8214 & ~n8592;
  assign n8594 = n8191 & ~n8211;
  assign n8595 = ~n8191 & n8211;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~n8583 & ~n8587;
  assign n8598 = ~n8578 & ~n8590;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8596 & ~n8599;
  assign n8601 = ~n8593 & ~n8600;
  assign n8602 = ~n8187 & n8601;
  assign n8603 = n8187 & ~n8601;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = n5257 & ~n8604;
  assign n8606 = pi328 & n8605;
  assign n8607 = pi328 & n5257;
  assign n8608 = n8187 & n8601;
  assign n8609 = ~n8187 & ~n8601;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = ~n8607 & ~n8610;
  assign n8612 = ~n8606 & ~n8611;
  assign n8613 = ~n8186 & ~n8612;
  assign n8614 = n8170 & n8183;
  assign n8615 = ~n8170 & ~n8183;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = n5257 & ~n8610;
  assign n8618 = pi328 & n8617;
  assign n8619 = ~n8604 & ~n8607;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = ~n8616 & ~n8620;
  assign n8622 = ~n8613 & ~n8621;
  assign n8623 = ~n7270 & n7283;
  assign n8624 = n7270 & ~n7283;
  assign n8625 = ~n7733 & ~n8624;
  assign n8626 = ~n8623 & ~n8625;
  assign n8627 = n8622 & n8626;
  assign n8628 = ~n8622 & ~n8626;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = pi331 & n2464;
  assign n8631 = n2464 & ~n7253;
  assign n8632 = pi329 & n8631;
  assign n8633 = ~n6178 & ~n7263;
  assign n8634 = ~n7688 & ~n8633;
  assign n8635 = ~n8632 & n8634;
  assign n8636 = ~n7695 & ~n8635;
  assign n8637 = n2887 & ~n7684;
  assign n8638 = pi329 & n8637;
  assign n8639 = ~n7712 & ~n7719;
  assign n8640 = ~n8638 & ~n8639;
  assign n8641 = ~n7310 & ~n8640;
  assign n8642 = n2887 & ~n7719;
  assign n8643 = pi329 & n8642;
  assign n8644 = ~n7684 & ~n7712;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = ~n7728 & ~n8645;
  assign n8647 = ~n8641 & ~n8646;
  assign n8648 = pi330 & n2887;
  assign n8649 = n8647 & ~n8648;
  assign n8650 = ~n8636 & n8649;
  assign n8651 = n8636 & ~n8647;
  assign n8652 = n2464 & ~n8651;
  assign n8653 = ~n2887 & n8652;
  assign n8654 = ~n2464 & ~n8647;
  assign n8655 = n2464 & n8647;
  assign n8656 = n8636 & ~n8655;
  assign n8657 = ~n8654 & ~n8656;
  assign n8658 = n2887 & ~n8657;
  assign n8659 = ~n8653 & ~n8658;
  assign n8660 = pi330 & ~n8659;
  assign n8661 = ~n8650 & ~n8660;
  assign n8662 = ~n8630 & n8661;
  assign n8663 = n8630 & ~n8661;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = pi332 & n2091;
  assign n8666 = n1729 & ~n7739;
  assign n8667 = pi332 & n8666;
  assign n8668 = n7283 & ~n8140;
  assign n8669 = ~n7283 & ~n8149;
  assign n8670 = ~n8668 & ~n8669;
  assign n8671 = n7739 & ~n7742;
  assign n8672 = ~n8670 & ~n8671;
  assign n8673 = ~n8667 & ~n8672;
  assign n8674 = n8665 & n8673;
  assign n8675 = ~n8665 & ~n8673;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = ~n8664 & ~n8676;
  assign n8678 = n8630 & n8661;
  assign n8679 = ~n8630 & ~n8661;
  assign n8680 = ~n8678 & ~n8679;
  assign n8681 = ~n8665 & n8673;
  assign n8682 = n8665 & ~n8673;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = ~n8680 & ~n8683;
  assign n8685 = ~n8677 & ~n8684;
  assign n8686 = ~n8629 & ~n8685;
  assign n8687 = n8622 & ~n8626;
  assign n8688 = ~n8622 & n8626;
  assign n8689 = ~n8687 & ~n8688;
  assign n8690 = ~n8676 & ~n8680;
  assign n8691 = ~n8664 & ~n8683;
  assign n8692 = ~n8690 & ~n8691;
  assign n8693 = ~n8689 & ~n8692;
  assign n8694 = ~n8686 & ~n8693;
  assign n8695 = ~n8166 & n8694;
  assign n8696 = n8166 & ~n8694;
  assign n8697 = ~n8695 & ~n8696;
  assign n8698 = pi335 & ~n1256;
  assign n8699 = ~n7765 & n7778;
  assign n8700 = ~n7775 & ~n8699;
  assign n8701 = n1442 & n8700;
  assign n8702 = pi334 & n8701;
  assign n8703 = pi334 & n1442;
  assign n8704 = ~n8700 & ~n8703;
  assign n8705 = ~n8702 & ~n8704;
  assign n8706 = n8698 & ~n8705;
  assign n8707 = ~n8698 & n8705;
  assign n8708 = ~n8706 & ~n8707;
  assign n8709 = ~n8697 & ~n8708;
  assign n8710 = n8166 & n8694;
  assign n8711 = ~n8166 & ~n8694;
  assign n8712 = ~n8710 & ~n8711;
  assign n8713 = ~n8698 & ~n8705;
  assign n8714 = n8698 & n8705;
  assign n8715 = ~n8713 & ~n8714;
  assign n8716 = ~n8712 & ~n8715;
  assign n8717 = ~n8709 & ~n8716;
  assign n8718 = ~n8165 & ~n8717;
  assign n8719 = n8157 & ~n8162;
  assign n8720 = ~n8157 & n8162;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = ~n8708 & ~n8712;
  assign n8723 = ~n8697 & ~n8715;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = ~n8721 & ~n8724;
  assign n8726 = ~n8718 & ~n8725;
  assign n8727 = ~n8137 & ~n8726;
  assign n8728 = n8137 & n8726;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = pi258 & ~n8729;
  assign n8731 = pi128 & n8730;
  assign n8732 = pi337 & n8731;
  assign n8733 = pi337 & n1156;
  assign n8734 = ~n8727 & ~n8733;
  assign n8735 = ~n8728 & n8734;
  assign n8736 = ~n8732 & ~n8735;
  assign n8737 = ~pi272 & ~n7247;
  assign n8738 = pi272 & n7247;
  assign n8739 = n7794 & ~n7800;
  assign n8740 = pi336 & ~n7794;
  assign n8741 = n1156 & n8740;
  assign n8742 = ~n8739 & ~n8741;
  assign n8743 = ~n8738 & ~n8742;
  assign n8744 = ~n8737 & ~n8743;
  assign n8745 = ~pi273 & ~n8744;
  assign n8746 = pi273 & n8744;
  assign n8747 = ~n8745 & ~n8746;
  assign n8748 = ~n8736 & ~n8747;
  assign n8749 = pi273 & ~n8744;
  assign n8750 = ~pi273 & n8744;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8735 & ~n8751;
  assign n8753 = ~n8732 & n8752;
  assign n8754 = ~n8748 & ~n8753;
  assign n8755 = ~n7812 & ~n7827;
  assign n8756 = n7812 & n7827;
  assign n8757 = pi307 & ~n7245;
  assign n8758 = pi128 & n8757;
  assign n8759 = n7245 & ~n7818;
  assign n8760 = ~n8758 & ~n8759;
  assign n8761 = ~n8756 & ~n8760;
  assign n8762 = ~n8755 & ~n8761;
  assign n8763 = n8754 & ~n8762;
  assign n8764 = ~n8754 & n8762;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = ~n8110 & ~n8765;
  assign n8767 = n8754 & n8762;
  assign n8768 = ~n8754 & ~n8762;
  assign n8769 = ~n8767 & ~n8768;
  assign n8770 = n8110 & ~n8769;
  assign n8771 = ~n8766 & ~n8770;
  assign n8772 = ~n831 & ~n8771;
  assign n8773 = ~n7837 & ~n8772;
  assign n8774 = pi161 & ~n8773;
  assign n8775 = pi079 & ~pi161;
  assign n8776 = ~n8774 & ~n8775;
  assign po208 = ~pi160 & ~n8776;
  assign n8778 = pi274 & n831;
  assign n8779 = n8736 & ~n8744;
  assign n8780 = ~n8736 & n8744;
  assign n8781 = ~pi273 & ~n8780;
  assign n8782 = ~n8779 & ~n8781;
  assign n8783 = n8157 & n8166;
  assign n8784 = ~n8157 & ~n8166;
  assign n8785 = n8694 & ~n8784;
  assign n8786 = ~n8783 & ~n8785;
  assign n8787 = ~n8157 & ~n8694;
  assign n8788 = n8157 & n8694;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~n8162 & n8698;
  assign n8791 = n8166 & ~n8705;
  assign n8792 = ~n8166 & n8705;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = ~n8790 & ~n8793;
  assign n8795 = ~n8789 & n8794;
  assign n8796 = ~n8157 & n8694;
  assign n8797 = n8157 & ~n8694;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = ~n8166 & ~n8705;
  assign n8800 = n8166 & n8705;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8790 & ~n8801;
  assign n8803 = ~n8798 & n8802;
  assign n8804 = n8162 & ~n8698;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = ~n8795 & n8805;
  assign n8807 = ~n8786 & ~n8806;
  assign n8808 = n8786 & n8806;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = pi333 & n2091;
  assign n8811 = ~n8170 & ~n8601;
  assign n8812 = n8170 & n8601;
  assign n8813 = n5257 & ~n8812;
  assign n8814 = pi328 & n8813;
  assign n8815 = ~n8811 & ~n8814;
  assign n8816 = n8183 & ~n8187;
  assign n8817 = ~n8183 & n8187;
  assign n8818 = ~n8170 & n8601;
  assign n8819 = n8170 & ~n8601;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = n5257 & ~n8820;
  assign n8822 = pi328 & n8821;
  assign n8823 = ~n8811 & ~n8812;
  assign n8824 = ~n8607 & ~n8823;
  assign n8825 = ~n8822 & ~n8824;
  assign n8826 = ~n8817 & ~n8825;
  assign n8827 = ~n8816 & ~n8826;
  assign n8828 = n8815 & n8827;
  assign n8829 = ~n8815 & ~n8827;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = pi329 & n5257;
  assign n8832 = ~n8191 & n8580;
  assign n8833 = n8191 & ~n8580;
  assign n8834 = ~n8587 & ~n8833;
  assign n8835 = ~n8832 & ~n8834;
  assign n8836 = ~n8191 & ~n8575;
  assign n8837 = n8191 & n8575;
  assign n8838 = ~n8836 & ~n8837;
  assign n8839 = n8211 & n8579;
  assign n8840 = ~n8560 & n8580;
  assign n8841 = n8560 & ~n8580;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = ~n8839 & ~n8842;
  assign n8844 = ~n8838 & n8843;
  assign n8845 = ~n8191 & n8575;
  assign n8846 = n8191 & ~n8575;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = n8560 & n8580;
  assign n8849 = ~n8560 & ~n8580;
  assign n8850 = ~n8848 & ~n8849;
  assign n8851 = ~n8839 & ~n8850;
  assign n8852 = ~n8847 & n8851;
  assign n8853 = ~n8211 & ~n8579;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = ~n8844 & n8854;
  assign n8856 = n8835 & n8855;
  assign n8857 = ~n8835 & ~n8855;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8216 & ~n8529;
  assign n8860 = ~n8537 & ~n8859;
  assign n8861 = ~n8224 & n8540;
  assign n8862 = ~n8216 & ~n8538;
  assign n8863 = n8216 & ~n8537;
  assign n8864 = ~n8529 & n8863;
  assign n8865 = ~n8862 & ~n8864;
  assign n8866 = n8224 & ~n8540;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = ~n8861 & ~n8867;
  assign n8869 = ~n8860 & n8868;
  assign n8870 = n8860 & ~n8868;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = ~n7364 & ~n7606;
  assign n8873 = ~n7607 & ~n8872;
  assign n8874 = pi139 & pi263;
  assign n8875 = pi136 & pi266;
  assign n8876 = pi133 & pi269;
  assign n8877 = pi271 & pi272;
  assign n8878 = ~n7371 & n8877;
  assign n8879 = ~pi271 & ~pi273;
  assign n8880 = pi272 & ~n8879;
  assign n8881 = pi271 & pi273;
  assign n8882 = ~pi272 & ~n8881;
  assign n8883 = ~n7371 & ~n8882;
  assign n8884 = ~n8880 & ~n8883;
  assign n8885 = pi128 & ~n8884;
  assign n8886 = ~n8878 & ~n8885;
  assign n8887 = pi129 & ~n8886;
  assign n8888 = pi272 & ~n7371;
  assign n8889 = n8246 & n8888;
  assign n8890 = ~n8887 & ~n8889;
  assign n8891 = pi129 & pi273;
  assign n8892 = pi128 & pi274;
  assign n8893 = ~n8891 & ~n8892;
  assign n8894 = pi273 & n1175;
  assign n8895 = pi274 & n8894;
  assign n8896 = ~n8893 & ~n8895;
  assign n8897 = ~n8890 & ~n8896;
  assign n8898 = n8890 & n8896;
  assign n8899 = ~n8897 & ~n8898;
  assign n8900 = pi272 & ~n8899;
  assign n8901 = pi130 & n8900;
  assign n8902 = pi130 & pi272;
  assign n8903 = ~n8898 & ~n8902;
  assign n8904 = ~n8897 & n8903;
  assign n8905 = ~n8901 & ~n8904;
  assign n8906 = n7372 & n7375;
  assign n8907 = ~n7372 & ~n7375;
  assign n8908 = ~n7371 & ~n8907;
  assign n8909 = ~n8906 & ~n8908;
  assign n8910 = ~n8252 & ~n8909;
  assign n8911 = ~n7375 & ~n8245;
  assign n8912 = n7371 & ~n7372;
  assign n8913 = ~n8911 & ~n8912;
  assign n8914 = n8252 & ~n8913;
  assign n8915 = ~n8910 & ~n8914;
  assign n8916 = n8254 & n8915;
  assign n8917 = ~n8254 & ~n8915;
  assign n8918 = ~n8284 & ~n8917;
  assign n8919 = ~n7386 & n8918;
  assign n8920 = ~n8916 & ~n8919;
  assign n8921 = pi131 & pi271;
  assign n8922 = ~n8920 & ~n8921;
  assign n8923 = pi271 & n8920;
  assign n8924 = pi131 & n8923;
  assign n8925 = ~n8922 & ~n8924;
  assign n8926 = ~n8905 & ~n8925;
  assign n8927 = pi271 & ~n8920;
  assign n8928 = pi131 & n8927;
  assign n8929 = n8920 & ~n8921;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = ~n8904 & ~n8930;
  assign n8932 = ~n8901 & n8931;
  assign n8933 = ~n8926 & ~n8932;
  assign n8934 = ~n8237 & ~n8289;
  assign n8935 = ~n8295 & ~n8934;
  assign n8936 = pi270 & n8289;
  assign n8937 = pi131 & n8936;
  assign n8938 = ~n8935 & ~n8937;
  assign n8939 = n8933 & n8938;
  assign n8940 = ~n8933 & ~n8938;
  assign n8941 = ~n8939 & ~n8940;
  assign n8942 = pi132 & pi270;
  assign n8943 = n8314 & ~n8319;
  assign n8944 = ~n8320 & ~n8943;
  assign n8945 = n8942 & ~n8944;
  assign n8946 = ~n8314 & ~n8320;
  assign n8947 = ~n8319 & ~n8946;
  assign n8948 = ~n8942 & ~n8947;
  assign n8949 = ~n8945 & ~n8948;
  assign n8950 = ~n8941 & ~n8949;
  assign n8951 = n8933 & ~n8938;
  assign n8952 = ~n8933 & n8938;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = ~n8942 & ~n8944;
  assign n8955 = n8942 & ~n8947;
  assign n8956 = ~n8954 & ~n8955;
  assign n8957 = ~n8953 & ~n8956;
  assign n8958 = ~n8950 & ~n8957;
  assign n8959 = ~n8876 & n8958;
  assign n8960 = n8876 & ~n8958;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = pi269 & ~n8321;
  assign n8963 = pi132 & n8962;
  assign n8964 = ~n8312 & ~n8314;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = pi268 & ~n8965;
  assign n8967 = pi133 & n8966;
  assign n8968 = pi134 & pi268;
  assign n8969 = ~n8313 & ~n8964;
  assign n8970 = ~n8963 & n8969;
  assign n8971 = ~n8330 & ~n8970;
  assign n8972 = ~n8968 & ~n8971;
  assign n8973 = ~n8967 & n8972;
  assign n8974 = ~n8967 & ~n8971;
  assign n8975 = n8968 & ~n8974;
  assign n8976 = ~n8973 & ~n8975;
  assign n8977 = ~n8961 & ~n8976;
  assign n8978 = ~n8876 & ~n8958;
  assign n8979 = n8876 & n8958;
  assign n8980 = ~n8978 & ~n8979;
  assign n8981 = n8968 & ~n8971;
  assign n8982 = ~n8967 & n8981;
  assign n8983 = ~n8968 & ~n8974;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = ~n8980 & ~n8984;
  assign n8986 = ~n8977 & ~n8985;
  assign n8987 = n8334 & ~n8359;
  assign n8988 = ~n8334 & n8359;
  assign n8989 = ~n8350 & ~n8988;
  assign n8990 = ~n8987 & ~n8989;
  assign n8991 = n8986 & n8990;
  assign n8992 = ~n8986 & ~n8990;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = pi135 & pi267;
  assign n8995 = n8373 & ~n8379;
  assign n8996 = ~n8378 & ~n8995;
  assign n8997 = n8994 & ~n8996;
  assign n8998 = ~n8373 & ~n8378;
  assign n8999 = ~n8379 & ~n8998;
  assign n9000 = ~n8994 & ~n8999;
  assign n9001 = ~n8997 & ~n9000;
  assign n9002 = ~n8993 & ~n9001;
  assign n9003 = n8986 & ~n8990;
  assign n9004 = ~n8986 & n8990;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n8994 & ~n8996;
  assign n9007 = n8994 & ~n8999;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = ~n9005 & ~n9008;
  assign n9010 = ~n9002 & ~n9009;
  assign n9011 = ~n8875 & n9010;
  assign n9012 = n8875 & ~n9010;
  assign n9013 = ~n9011 & ~n9012;
  assign n9014 = pi266 & ~n8380;
  assign n9015 = pi135 & n9014;
  assign n9016 = ~n8371 & ~n8373;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = pi265 & ~n9017;
  assign n9019 = pi136 & n9018;
  assign n9020 = pi137 & pi265;
  assign n9021 = ~n8372 & ~n9016;
  assign n9022 = ~n9015 & n9021;
  assign n9023 = ~n8389 & ~n9022;
  assign n9024 = ~n9020 & ~n9023;
  assign n9025 = ~n9019 & n9024;
  assign n9026 = ~n9019 & ~n9023;
  assign n9027 = n9020 & ~n9026;
  assign n9028 = ~n9025 & ~n9027;
  assign n9029 = ~n9013 & ~n9028;
  assign n9030 = ~n8875 & ~n9010;
  assign n9031 = n8875 & n9010;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = n9020 & ~n9023;
  assign n9034 = ~n9019 & n9033;
  assign n9035 = ~n9020 & ~n9026;
  assign n9036 = ~n9034 & ~n9035;
  assign n9037 = ~n9032 & ~n9036;
  assign n9038 = ~n9029 & ~n9037;
  assign n9039 = n8393 & ~n8418;
  assign n9040 = ~n8393 & n8418;
  assign n9041 = ~n8409 & ~n9040;
  assign n9042 = ~n9039 & ~n9041;
  assign n9043 = n9038 & ~n9042;
  assign n9044 = ~n9038 & n9042;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = pi138 & pi264;
  assign n9047 = n8432 & ~n8438;
  assign n9048 = ~n8437 & ~n9047;
  assign n9049 = n9046 & ~n9048;
  assign n9050 = ~n8432 & ~n8437;
  assign n9051 = ~n8438 & ~n9050;
  assign n9052 = ~n9046 & ~n9051;
  assign n9053 = ~n9049 & ~n9052;
  assign n9054 = ~n9045 & ~n9053;
  assign n9055 = n9038 & n9042;
  assign n9056 = ~n9038 & ~n9042;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n9046 & ~n9048;
  assign n9059 = n9046 & ~n9051;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = ~n9057 & ~n9060;
  assign n9062 = ~n9054 & ~n9061;
  assign n9063 = ~n8874 & ~n9062;
  assign n9064 = n8874 & n9062;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = pi263 & ~n8439;
  assign n9067 = pi138 & n9066;
  assign n9068 = ~n8430 & ~n8432;
  assign n9069 = ~n8431 & ~n9068;
  assign n9070 = ~n9067 & n9069;
  assign n9071 = pi140 & pi262;
  assign n9072 = ~n9067 & ~n9068;
  assign n9073 = pi262 & ~n9072;
  assign n9074 = pi139 & n9073;
  assign n9075 = n8449 & ~n9074;
  assign n9076 = n9071 & ~n9075;
  assign n9077 = ~n9070 & n9076;
  assign n9078 = ~n9070 & ~n9075;
  assign n9079 = ~n9071 & ~n9078;
  assign n9080 = ~n9077 & ~n9079;
  assign n9081 = ~n9065 & ~n9080;
  assign n9082 = ~n8874 & n9062;
  assign n9083 = n8874 & ~n9062;
  assign n9084 = ~n9082 & ~n9083;
  assign n9085 = ~n9071 & ~n9075;
  assign n9086 = ~n9070 & n9085;
  assign n9087 = n9071 & ~n9078;
  assign n9088 = ~n9086 & ~n9087;
  assign n9089 = ~n9084 & ~n9088;
  assign n9090 = ~n9081 & ~n9089;
  assign n9091 = ~n8452 & ~n8453;
  assign n9092 = n8452 & n8453;
  assign n9093 = ~n8472 & ~n9092;
  assign n9094 = ~n9091 & ~n9093;
  assign n9095 = n9090 & n9094;
  assign n9096 = ~n9090 & ~n9094;
  assign n9097 = ~n9095 & ~n9096;
  assign n9098 = ~n7574 & ~n8229;
  assign n9099 = pi260 & n9098;
  assign n9100 = pi141 & n9099;
  assign n9101 = pi141 & pi261;
  assign n9102 = ~n8228 & ~n9098;
  assign n9103 = n8483 & ~n9102;
  assign n9104 = ~n9101 & ~n9103;
  assign n9105 = ~n9100 & n9104;
  assign n9106 = ~n9100 & ~n9103;
  assign n9107 = n9101 & ~n9106;
  assign n9108 = ~n9105 & ~n9107;
  assign n9109 = ~n9097 & ~n9108;
  assign n9110 = n9090 & ~n9094;
  assign n9111 = ~n9090 & n9094;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = n9101 & ~n9103;
  assign n9114 = ~n9100 & n9113;
  assign n9115 = ~n9101 & ~n9106;
  assign n9116 = ~n9114 & ~n9115;
  assign n9117 = ~n9112 & ~n9116;
  assign n9118 = ~n9109 & ~n9117;
  assign n9119 = ~n9100 & ~n9102;
  assign n9120 = n8483 & ~n9119;
  assign n9121 = ~n8483 & n9119;
  assign n9122 = ~n9120 & ~n9121;
  assign n9123 = ~n8494 & ~n9122;
  assign n9124 = ~n8493 & ~n9123;
  assign n9125 = n9118 & ~n9124;
  assign n9126 = ~n9118 & n9124;
  assign n9127 = ~n9125 & ~n9126;
  assign n9128 = pi143 & pi259;
  assign n9129 = ~n8486 & ~n8495;
  assign n9130 = ~n8501 & ~n8507;
  assign n9131 = n8498 & ~n9130;
  assign n9132 = ~n9129 & n9131;
  assign n9133 = ~n9128 & ~n9132;
  assign n9134 = pi142 & n8491;
  assign n9135 = ~pi142 & ~n8491;
  assign n9136 = ~n9134 & ~n9135;
  assign n9137 = ~n8507 & ~n9136;
  assign n9138 = pi142 & ~n8491;
  assign n9139 = ~pi142 & n8491;
  assign n9140 = ~n9138 & ~n9139;
  assign n9141 = ~n8486 & ~n9140;
  assign n9142 = ~n9137 & ~n9141;
  assign n9143 = n8498 & ~n9142;
  assign n9144 = pi259 & n9143;
  assign n9145 = ~n9133 & ~n9144;
  assign n9146 = pi144 & pi258;
  assign n9147 = pi142 & pi260;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = n9146 & n9147;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = ~n9145 & ~n9150;
  assign n9152 = ~n9146 & n9147;
  assign n9153 = n9146 & ~n9147;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = ~n9144 & ~n9154;
  assign n9156 = ~n9133 & n9155;
  assign n9157 = ~n9151 & ~n9156;
  assign n9158 = ~n9127 & ~n9157;
  assign n9159 = n9118 & n9124;
  assign n9160 = ~n9118 & ~n9124;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = ~n9145 & ~n9154;
  assign n9163 = ~n9144 & ~n9150;
  assign n9164 = ~n9133 & n9163;
  assign n9165 = ~n9162 & ~n9164;
  assign n9166 = ~n9161 & ~n9165;
  assign n9167 = ~n9158 & ~n9166;
  assign n9168 = n8873 & ~n9167;
  assign n9169 = ~n8873 & n9167;
  assign n9170 = n8513 & n9169;
  assign n9171 = ~n9168 & ~n9170;
  assign n9172 = ~n7601 & ~n9171;
  assign n9173 = ~n8873 & ~n9167;
  assign n9174 = n8873 & n9167;
  assign n9175 = ~n8513 & n9174;
  assign n9176 = ~n9173 & ~n9175;
  assign n9177 = n7601 & ~n9176;
  assign n9178 = ~n8513 & ~n8873;
  assign n9179 = n8513 & n8873;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = ~n9167 & ~n9180;
  assign n9182 = ~n9177 & ~n9181;
  assign n9183 = ~n9172 & n9182;
  assign n9184 = pi322 & ~n9183;
  assign n9185 = n8513 & ~n8873;
  assign n9186 = ~n8513 & n8873;
  assign n9187 = ~n9185 & ~n9186;
  assign n9188 = n7601 & ~n9187;
  assign n9189 = ~n7601 & ~n9180;
  assign n9190 = ~n9188 & ~n9189;
  assign n9191 = pi323 & ~n9190;
  assign n9192 = ~n9184 & ~n9191;
  assign n9193 = n7601 & n9185;
  assign n9194 = ~n9189 & ~n9193;
  assign n9195 = ~n9167 & ~n9194;
  assign n9196 = n7601 & ~n8513;
  assign n9197 = n9174 & n9196;
  assign n9198 = ~n9195 & ~n9197;
  assign n9199 = pi323 & ~n9198;
  assign n9200 = pi322 & n9199;
  assign n9201 = ~n9192 & ~n9200;
  assign n9202 = pi325 & n6556;
  assign n9203 = ~n7364 & ~n7612;
  assign n9204 = n7364 & ~n7608;
  assign n9205 = ~n9203 & ~n9204;
  assign n9206 = pi324 & n9205;
  assign n9207 = n9202 & n9206;
  assign n9208 = ~n9202 & ~n9206;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = ~n9201 & ~n9209;
  assign n9211 = ~n9202 & n9206;
  assign n9212 = n9202 & ~n9206;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = ~n9200 & ~n9213;
  assign n9215 = ~n9192 & n9214;
  assign n9216 = ~n9210 & ~n9215;
  assign n9217 = ~n8871 & ~n9216;
  assign n9218 = ~n8860 & ~n8868;
  assign n9219 = n8860 & n8868;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = ~n9201 & ~n9213;
  assign n9222 = ~n9200 & ~n9209;
  assign n9223 = ~n9192 & n9222;
  assign n9224 = ~n9221 & ~n9223;
  assign n9225 = ~n9220 & ~n9224;
  assign n9226 = ~n9217 & ~n9225;
  assign n9227 = n8539 & ~n8575;
  assign n9228 = ~n8540 & ~n8865;
  assign n9229 = n8216 & ~n8538;
  assign n9230 = ~n8216 & ~n8537;
  assign n9231 = ~n8529 & n9230;
  assign n9232 = ~n9229 & ~n9231;
  assign n9233 = n6556 & ~n9232;
  assign n9234 = pi324 & n9233;
  assign n9235 = ~n9228 & ~n9234;
  assign n9236 = n8224 & ~n9235;
  assign n9237 = ~n8224 & n9235;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = ~n8539 & n8575;
  assign n9240 = ~n9238 & ~n9239;
  assign n9241 = ~n9227 & ~n9240;
  assign n9242 = n9226 & n9241;
  assign n9243 = ~n9226 & ~n9241;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = pi327 & n5732;
  assign n9246 = pi326 & n5973;
  assign n9247 = n9245 & n9246;
  assign n9248 = ~n9245 & ~n9246;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = ~n9244 & ~n9249;
  assign n9251 = ~n9226 & n9241;
  assign n9252 = n9226 & ~n9241;
  assign n9253 = ~n9251 & ~n9252;
  assign n9254 = ~n9245 & n9246;
  assign n9255 = n9245 & ~n9246;
  assign n9256 = ~n9254 & ~n9255;
  assign n9257 = ~n9253 & ~n9256;
  assign n9258 = ~n9250 & ~n9257;
  assign n9259 = ~n8858 & ~n9258;
  assign n9260 = n8835 & ~n8855;
  assign n9261 = ~n8835 & n8855;
  assign n9262 = ~n9260 & ~n9261;
  assign n9263 = ~n9249 & ~n9253;
  assign n9264 = ~n9244 & ~n9256;
  assign n9265 = ~n9263 & ~n9264;
  assign n9266 = ~n9262 & ~n9265;
  assign n9267 = ~n9259 & ~n9266;
  assign n9268 = ~n8831 & n9267;
  assign n9269 = n8831 & ~n9267;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = n5714 & ~n9270;
  assign n9272 = pi328 & n9271;
  assign n9273 = pi328 & n5714;
  assign n9274 = n8831 & n9267;
  assign n9275 = ~n8831 & ~n9267;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = ~n9273 & ~n9276;
  assign n9278 = ~n9272 & ~n9277;
  assign n9279 = ~n8830 & ~n9278;
  assign n9280 = n8815 & ~n8827;
  assign n9281 = ~n8815 & n8827;
  assign n9282 = ~n9280 & ~n9281;
  assign n9283 = n5714 & ~n9276;
  assign n9284 = pi328 & n9283;
  assign n9285 = ~n9270 & ~n9273;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n9282 & ~n9286;
  assign n9288 = ~n9279 & ~n9287;
  assign n9289 = ~n8626 & n8630;
  assign n9290 = n8626 & ~n8630;
  assign n9291 = ~n8636 & ~n8654;
  assign n9292 = ~n8655 & ~n9291;
  assign n9293 = n2887 & ~n9292;
  assign n9294 = pi330 & n9293;
  assign n9295 = ~n7689 & ~n8647;
  assign n9296 = ~n8636 & ~n9295;
  assign n9297 = ~n2887 & ~n8655;
  assign n9298 = pi330 & ~n9297;
  assign n9299 = ~n9296 & ~n9298;
  assign n9300 = ~n9294 & ~n9299;
  assign n9301 = n8622 & ~n9300;
  assign n9302 = ~n8622 & n9300;
  assign n9303 = ~n9301 & ~n9302;
  assign n9304 = ~n9290 & ~n9303;
  assign n9305 = ~n9289 & ~n9304;
  assign n9306 = n9288 & n9305;
  assign n9307 = ~n9288 & ~n9305;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = pi331 & n2887;
  assign n9310 = n8622 & ~n9299;
  assign n9311 = ~n9294 & ~n9310;
  assign n9312 = n4596 & n9311;
  assign n9313 = pi330 & n9312;
  assign n9314 = pi330 & n4596;
  assign n9315 = ~n9311 & ~n9314;
  assign n9316 = ~n9313 & ~n9315;
  assign n9317 = ~n9309 & n9316;
  assign n9318 = n9309 & ~n9316;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = pi332 & n2464;
  assign n9321 = ~n8664 & ~n8682;
  assign n9322 = ~n8689 & n9321;
  assign n9323 = ~n8680 & ~n8682;
  assign n9324 = ~n8629 & n9323;
  assign n9325 = ~n8681 & ~n9324;
  assign n9326 = ~n9322 & n9325;
  assign n9327 = n9320 & ~n9326;
  assign n9328 = ~n9320 & n9326;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n9319 & ~n9329;
  assign n9331 = n9309 & n9316;
  assign n9332 = ~n9309 & ~n9316;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = ~n9320 & ~n9326;
  assign n9335 = n9320 & n9326;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = ~n9333 & ~n9336;
  assign n9338 = ~n9330 & ~n9337;
  assign n9339 = ~n9308 & ~n9338;
  assign n9340 = n9288 & ~n9305;
  assign n9341 = ~n9288 & n9305;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = ~n9329 & ~n9333;
  assign n9344 = ~n9319 & ~n9336;
  assign n9345 = ~n9343 & ~n9344;
  assign n9346 = ~n9342 & ~n9345;
  assign n9347 = ~n9339 & ~n9346;
  assign n9348 = ~n8810 & n9347;
  assign n9349 = n8810 & ~n9347;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = pi335 & n1442;
  assign n9352 = ~n8699 & ~n8703;
  assign n9353 = ~n7775 & n9352;
  assign n9354 = pi334 & n1729;
  assign n9355 = n8166 & ~n9354;
  assign n9356 = ~n9353 & n9355;
  assign n9357 = n1442 & ~n8700;
  assign n9358 = pi334 & n9357;
  assign n9359 = ~n8166 & n9354;
  assign n9360 = ~n9358 & n9359;
  assign n9361 = ~n9356 & ~n9360;
  assign n9362 = ~n8789 & ~n9361;
  assign n9363 = n8166 & n9354;
  assign n9364 = ~n9358 & n9363;
  assign n9365 = ~n8166 & ~n9354;
  assign n9366 = ~n9353 & n9365;
  assign n9367 = ~n9364 & ~n9366;
  assign n9368 = ~n8798 & ~n9367;
  assign n9369 = ~n9354 & n9358;
  assign n9370 = n9353 & n9354;
  assign n9371 = ~n9358 & n9370;
  assign n9372 = ~n9369 & ~n9371;
  assign n9373 = ~n9368 & n9372;
  assign n9374 = ~n9362 & n9373;
  assign n9375 = n9351 & ~n9374;
  assign n9376 = ~n9351 & n9374;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = ~n9350 & ~n9377;
  assign n9379 = n8810 & n9347;
  assign n9380 = ~n8810 & ~n9347;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = ~n9351 & ~n9374;
  assign n9383 = n9351 & n9374;
  assign n9384 = ~n9382 & ~n9383;
  assign n9385 = ~n9381 & ~n9384;
  assign n9386 = ~n9378 & ~n9385;
  assign n9387 = ~n8809 & ~n9386;
  assign n9388 = ~n8786 & n8806;
  assign n9389 = n8786 & ~n8806;
  assign n9390 = ~n9388 & ~n9389;
  assign n9391 = ~n9377 & ~n9381;
  assign n9392 = ~n9350 & ~n9384;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = ~n9390 & ~n9393;
  assign n9395 = ~n9387 & ~n9394;
  assign n9396 = n8732 & ~n9395;
  assign n9397 = ~n8732 & n9395;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = n8133 & n8726;
  assign n9400 = ~n8133 & ~n8726;
  assign n9401 = ~n1154 & ~n9400;
  assign n9402 = ~n9399 & ~n9401;
  assign n9403 = ~n1256 & ~n9402;
  assign n9404 = pi336 & n9403;
  assign n9405 = ~n1154 & n8726;
  assign n9406 = n1256 & ~n9405;
  assign n9407 = pi336 & ~n9406;
  assign n9408 = n1154 & ~n8726;
  assign n9409 = n8133 & ~n9408;
  assign n9410 = ~n9407 & ~n9409;
  assign n9411 = ~n9404 & ~n9410;
  assign n9412 = ~n1154 & ~n9411;
  assign n9413 = pi337 & n9412;
  assign n9414 = pi337 & ~n1154;
  assign n9415 = ~n9410 & ~n9414;
  assign n9416 = ~n9404 & n9415;
  assign n9417 = ~n9413 & ~n9416;
  assign n9418 = ~n9398 & ~n9417;
  assign n9419 = n8732 & n9395;
  assign n9420 = ~n8732 & ~n9395;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n9411 & ~n9414;
  assign n9423 = n9411 & n9414;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = ~n9421 & ~n9424;
  assign n9426 = ~n9418 & ~n9425;
  assign n9427 = pi274 & ~n9426;
  assign n9428 = ~pi274 & n9426;
  assign n9429 = ~n9427 & ~n9428;
  assign n9430 = pi258 & ~n9429;
  assign n9431 = pi128 & n9430;
  assign n9432 = pi338 & n9431;
  assign n9433 = pi274 & n9426;
  assign n9434 = ~pi274 & ~n9426;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = pi338 & n1156;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = ~n9432 & ~n9437;
  assign n9439 = ~n8782 & ~n9438;
  assign n9440 = n8782 & n9438;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = ~n8084 & n8086;
  assign n9443 = pi129 & n8084;
  assign n9444 = ~n9442 & ~n9443;
  assign n9445 = ~n8099 & ~n9444;
  assign n9446 = ~n8084 & ~n8086;
  assign n9447 = ~pi129 & n8084;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n8053 & ~n9448;
  assign n9450 = ~n9445 & ~n9449;
  assign n9451 = n8085 & ~n9450;
  assign n9452 = pi306 & ~n1568;
  assign n9453 = n9451 & n9452;
  assign n9454 = ~n9451 & ~n9452;
  assign n9455 = ~n9453 & ~n9454;
  assign n9456 = pi307 & n1515;
  assign n9457 = ~n8099 & ~n9447;
  assign n9458 = ~n9446 & ~n9457;
  assign n9459 = n9456 & ~n9458;
  assign n9460 = ~n8053 & ~n9446;
  assign n9461 = ~n9447 & ~n9460;
  assign n9462 = ~n9456 & ~n9461;
  assign n9463 = ~n9459 & ~n9462;
  assign n9464 = pi309 & n1533;
  assign n9465 = ~n8031 & ~n8035;
  assign n9466 = ~n8036 & ~n9465;
  assign n9467 = ~n9464 & ~n9466;
  assign n9468 = ~n8028 & ~n8036;
  assign n9469 = ~n7222 & n9468;
  assign n9470 = ~n8035 & ~n9469;
  assign n9471 = n9464 & ~n9470;
  assign n9472 = ~n9467 & ~n9471;
  assign n9473 = ~n7848 & ~n8003;
  assign n9474 = ~n7189 & ~n7194;
  assign n9475 = ~n7190 & ~n9474;
  assign n9476 = n7848 & n8003;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = ~n9473 & ~n9477;
  assign n9479 = pi313 & n3012;
  assign n9480 = ~n7982 & ~n7989;
  assign n9481 = ~n7990 & ~n9480;
  assign n9482 = ~n9479 & ~n9481;
  assign n9483 = ~n7985 & ~n7990;
  assign n9484 = ~n7989 & ~n9483;
  assign n9485 = n9479 & ~n9484;
  assign n9486 = ~n9482 & ~n9485;
  assign n9487 = ~n7958 & ~n7959;
  assign n9488 = n7958 & n7959;
  assign n9489 = ~n7164 & ~n9488;
  assign n9490 = ~n7158 & n9489;
  assign n9491 = ~n9487 & ~n9490;
  assign n9492 = pi316 & n4772;
  assign n9493 = ~pi144 & ~n7035;
  assign n9494 = pi143 & n9493;
  assign n9495 = ~pi143 & pi144;
  assign n9496 = pi142 & n9495;
  assign n9497 = ~n9494 & ~n9496;
  assign n9498 = pi141 & ~n9497;
  assign n9499 = pi143 & pi144;
  assign n9500 = ~pi142 & n9499;
  assign n9501 = ~pi144 & n7035;
  assign n9502 = ~pi143 & n9501;
  assign n9503 = ~n9500 & ~n9502;
  assign n9504 = ~pi141 & ~n9503;
  assign n9505 = pi143 & ~pi144;
  assign n9506 = pi144 & ~n7035;
  assign n9507 = ~pi143 & n9506;
  assign n9508 = ~n9505 & ~n9507;
  assign n9509 = pi142 & ~n9508;
  assign n9510 = ~pi143 & ~pi144;
  assign n9511 = pi144 & n7035;
  assign n9512 = pi143 & n9511;
  assign n9513 = ~n9510 & ~n9512;
  assign n9514 = ~pi142 & ~n9513;
  assign n9515 = ~n9509 & ~n9514;
  assign n9516 = ~n9504 & n9515;
  assign n9517 = ~n9498 & n9516;
  assign n9518 = pi321 & n9517;
  assign n9519 = ~n7875 & n7881;
  assign n9520 = n7044 & ~n9519;
  assign n9521 = pi320 & n9520;
  assign n9522 = n7874 & ~n7881;
  assign n9523 = pi321 & n9522;
  assign n9524 = ~n9521 & ~n9523;
  assign n9525 = pi320 & n7874;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = n7874 & n9524;
  assign n9528 = pi320 & n9527;
  assign n9529 = ~n9526 & ~n9528;
  assign n9530 = ~n9518 & ~n9529;
  assign n9531 = n9524 & ~n9525;
  assign n9532 = n7874 & ~n9524;
  assign n9533 = pi320 & n9532;
  assign n9534 = ~n9531 & ~n9533;
  assign n9535 = n9517 & ~n9534;
  assign n9536 = pi321 & n9535;
  assign n9537 = ~n9530 & ~n9536;
  assign n9538 = n6777 & ~n7899;
  assign n9539 = pi319 & n9538;
  assign n9540 = ~n7898 & ~n9539;
  assign n9541 = ~n9537 & ~n9540;
  assign n9542 = n9537 & n9540;
  assign n9543 = ~n9541 & ~n9542;
  assign n9544 = n7044 & ~n9543;
  assign n9545 = pi319 & n9544;
  assign n9546 = pi319 & n7044;
  assign n9547 = n9537 & ~n9540;
  assign n9548 = ~n9537 & n9540;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~n9546 & ~n9549;
  assign n9551 = ~n9545 & ~n9550;
  assign n9552 = pi318 & n6777;
  assign n9553 = ~n9551 & ~n9552;
  assign n9554 = n6777 & n9551;
  assign n9555 = pi318 & n9554;
  assign n9556 = ~n9553 & ~n9555;
  assign n9557 = ~n7908 & ~n7916;
  assign n9558 = n7908 & n7916;
  assign n9559 = n5463 & ~n9558;
  assign n9560 = pi318 & n9559;
  assign n9561 = ~n9557 & ~n9560;
  assign n9562 = n9556 & ~n9561;
  assign n9563 = ~n9556 & n9561;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = pi317 & n5463;
  assign n9566 = ~n7932 & ~n9565;
  assign n9567 = ~n7921 & n9566;
  assign n9568 = ~n7921 & ~n7932;
  assign n9569 = n9565 & ~n9568;
  assign n9570 = ~n9567 & ~n9569;
  assign n9571 = ~n9564 & ~n9570;
  assign n9572 = n9556 & n9561;
  assign n9573 = ~n9556 & ~n9561;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = ~n7932 & n9565;
  assign n9576 = ~n7921 & n9575;
  assign n9577 = ~n9565 & ~n9568;
  assign n9578 = ~n9576 & ~n9577;
  assign n9579 = ~n9574 & ~n9578;
  assign n9580 = ~n9571 & ~n9579;
  assign n9581 = ~n9492 & ~n9580;
  assign n9582 = n9492 & n9580;
  assign n9583 = ~n9581 & ~n9582;
  assign n9584 = pi315 & n4086;
  assign n9585 = ~n7929 & ~n7940;
  assign n9586 = n7929 & n7940;
  assign n9587 = n7853 & ~n9586;
  assign n9588 = ~n9585 & ~n9587;
  assign n9589 = n9584 & ~n9588;
  assign n9590 = ~n7853 & ~n9585;
  assign n9591 = ~n9586 & ~n9590;
  assign n9592 = ~n9584 & ~n9591;
  assign n9593 = ~n9589 & ~n9592;
  assign n9594 = ~n9583 & ~n9593;
  assign n9595 = ~n9492 & n9580;
  assign n9596 = n9492 & ~n9580;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = ~n9584 & ~n9588;
  assign n9599 = n9584 & ~n9591;
  assign n9600 = ~n9598 & ~n9599;
  assign n9601 = ~n9597 & ~n9600;
  assign n9602 = ~n9594 & ~n9601;
  assign n9603 = n7946 & ~n7955;
  assign n9604 = ~n7946 & n7955;
  assign n9605 = ~n7949 & ~n9604;
  assign n9606 = ~n9603 & ~n9605;
  assign n9607 = ~n9602 & n9606;
  assign n9608 = n9602 & ~n9606;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = n3552 & ~n9609;
  assign n9611 = pi314 & n9610;
  assign n9612 = pi314 & n3552;
  assign n9613 = ~n9608 & ~n9612;
  assign n9614 = ~n9607 & n9613;
  assign n9615 = ~n9611 & ~n9614;
  assign n9616 = ~n9491 & ~n9615;
  assign n9617 = n9491 & ~n9614;
  assign n9618 = ~n9611 & n9617;
  assign n9619 = ~n9616 & ~n9618;
  assign n9620 = n9486 & ~n9619;
  assign n9621 = ~n9486 & n9619;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = pi312 & n2574;
  assign n9624 = ~n2183 & ~n2574;
  assign n9625 = pi313 & ~n9624;
  assign n9626 = n7974 & ~n9625;
  assign n9627 = ~n2183 & n2574;
  assign n9628 = pi313 & ~n7974;
  assign n9629 = n9627 & n9628;
  assign n9630 = ~n9626 & ~n9629;
  assign n9631 = ~n7979 & ~n9630;
  assign n9632 = ~n2574 & n7974;
  assign n9633 = ~n7976 & ~n9632;
  assign n9634 = ~n7166 & ~n9633;
  assign n9635 = n7015 & n9634;
  assign n9636 = n2183 & ~n2574;
  assign n9637 = ~n7974 & n9636;
  assign n9638 = ~n2183 & ~n7166;
  assign n9639 = n2574 & ~n9638;
  assign n9640 = n7974 & n9639;
  assign n9641 = ~n9637 & ~n9640;
  assign n9642 = pi313 & ~n9641;
  assign n9643 = n7166 & n7989;
  assign n9644 = ~n9642 & ~n9643;
  assign n9645 = ~n7015 & ~n9644;
  assign n9646 = ~n2574 & ~n7974;
  assign n9647 = n2574 & n7974;
  assign n9648 = ~n9646 & ~n9647;
  assign n9649 = n2183 & ~n9648;
  assign n9650 = pi313 & n9649;
  assign n9651 = n7166 & n9650;
  assign n9652 = ~n9645 & ~n9651;
  assign n9653 = ~n9635 & n9652;
  assign n9654 = ~n9631 & n9653;
  assign n9655 = ~n8000 & ~n9654;
  assign n9656 = n8000 & n9654;
  assign n9657 = n7978 & ~n9656;
  assign n9658 = ~n9655 & ~n9657;
  assign n9659 = n9623 & ~n9658;
  assign n9660 = ~n7978 & ~n9655;
  assign n9661 = ~n9656 & ~n9660;
  assign n9662 = ~n9623 & ~n9661;
  assign n9663 = ~n9659 & ~n9662;
  assign n9664 = ~n9622 & ~n9663;
  assign n9665 = n9486 & n9619;
  assign n9666 = ~n9486 & ~n9619;
  assign n9667 = ~n9665 & ~n9666;
  assign n9668 = ~n9623 & ~n9658;
  assign n9669 = n9623 & ~n9661;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = ~n9667 & ~n9670;
  assign n9672 = ~n9664 & ~n9671;
  assign n9673 = n9478 & ~n9672;
  assign n9674 = ~n9478 & n9672;
  assign n9675 = ~n9673 & ~n9674;
  assign n9676 = n2183 & ~n9675;
  assign n9677 = pi311 & n9676;
  assign n9678 = pi311 & n2183;
  assign n9679 = ~n9478 & ~n9672;
  assign n9680 = n9478 & n9672;
  assign n9681 = ~n9679 & ~n9680;
  assign n9682 = ~n9678 & ~n9681;
  assign n9683 = ~n9677 & ~n9682;
  assign n9684 = ~n8007 & ~n8017;
  assign n9685 = n8007 & n8017;
  assign n9686 = ~n8008 & ~n9685;
  assign n9687 = ~n7201 & n9686;
  assign n9688 = ~n9684 & ~n9687;
  assign n9689 = n9683 & n9688;
  assign n9690 = ~n9683 & ~n9688;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n1840 & ~n9691;
  assign n9693 = pi310 & n9692;
  assign n9694 = pi310 & n1840;
  assign n9695 = ~n9683 & n9688;
  assign n9696 = n9683 & ~n9688;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n9694 & ~n9697;
  assign n9699 = ~n9693 & ~n9698;
  assign n9700 = n9472 & n9699;
  assign n9701 = ~n9472 & ~n9699;
  assign n9702 = ~n9700 & ~n9701;
  assign n9703 = pi308 & n1553;
  assign n9704 = n8023 & ~n8028;
  assign n9705 = ~n7222 & n9704;
  assign n9706 = ~n8023 & ~n8031;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = ~n7838 & ~n9707;
  assign n9709 = ~n8023 & ~n8028;
  assign n9710 = ~n7222 & n9709;
  assign n9711 = n8023 & ~n8031;
  assign n9712 = ~n9710 & ~n9711;
  assign n9713 = n1553 & ~n9712;
  assign n9714 = pi309 & n9713;
  assign n9715 = ~n9708 & ~n9714;
  assign n9716 = ~n8050 & n9715;
  assign n9717 = n8050 & ~n9715;
  assign n9718 = n8027 & ~n9717;
  assign n9719 = ~n9716 & ~n9718;
  assign n9720 = n9703 & ~n9719;
  assign n9721 = ~n8027 & ~n9716;
  assign n9722 = ~n9717 & ~n9721;
  assign n9723 = ~n9703 & ~n9722;
  assign n9724 = ~n9720 & ~n9723;
  assign n9725 = ~n9702 & ~n9724;
  assign n9726 = n9472 & ~n9699;
  assign n9727 = ~n9472 & n9699;
  assign n9728 = ~n9726 & ~n9727;
  assign n9729 = ~n9703 & ~n9719;
  assign n9730 = n9703 & ~n9722;
  assign n9731 = ~n9729 & ~n9730;
  assign n9732 = ~n9728 & ~n9731;
  assign n9733 = ~n9725 & ~n9732;
  assign n9734 = ~n9463 & n9733;
  assign n9735 = n9463 & ~n9733;
  assign n9736 = ~n9734 & ~n9735;
  assign n9737 = ~n9455 & ~n9736;
  assign n9738 = n9463 & n9733;
  assign n9739 = ~n9463 & ~n9733;
  assign n9740 = ~n9738 & ~n9739;
  assign n9741 = ~n9451 & n9452;
  assign n9742 = n9451 & ~n9452;
  assign n9743 = ~n9741 & ~n9742;
  assign n9744 = ~n9740 & ~n9743;
  assign n9745 = ~n9737 & ~n9744;
  assign n9746 = pi305 & ~n9745;
  assign n9747 = pi128 & n9746;
  assign n9748 = pi128 & pi305;
  assign n9749 = n9745 & ~n9748;
  assign n9750 = ~n9747 & ~n9749;
  assign n9751 = ~n9441 & ~n9750;
  assign n9752 = n8782 & ~n9438;
  assign n9753 = ~n8782 & n9438;
  assign n9754 = ~n9752 & ~n9753;
  assign n9755 = ~n9745 & ~n9748;
  assign n9756 = pi305 & n9745;
  assign n9757 = pi128 & n9756;
  assign n9758 = ~n9755 & ~n9757;
  assign n9759 = ~n9754 & ~n9758;
  assign n9760 = ~n9751 & ~n9759;
  assign n9761 = n8110 & ~n8767;
  assign n9762 = ~n8768 & ~n9761;
  assign n9763 = n9760 & ~n9762;
  assign n9764 = ~n9760 & n9762;
  assign n9765 = ~n9763 & ~n9764;
  assign n9766 = ~n831 & ~n9765;
  assign n9767 = ~n8778 & ~n9766;
  assign n9768 = pi161 & ~n9767;
  assign n9769 = pi080 & ~pi161;
  assign n9770 = ~n9768 & ~n9769;
  assign po209 = ~pi160 & ~n9770;
  assign n9772 = pi275 & n831;
  assign n9773 = ~n9455 & ~n9740;
  assign n9774 = ~n9736 & ~n9743;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = pi305 & ~n9775;
  assign n9777 = pi128 & n9776;
  assign n9778 = ~pi128 & pi305;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = pi129 & ~n9779;
  assign n9781 = pi305 & ~n9777;
  assign n9782 = n1567 & n9781;
  assign n9783 = ~n9780 & ~n9782;
  assign n9784 = pi309 & n1840;
  assign n9785 = pi313 & n3552;
  assign n9786 = pi144 & ~pi145;
  assign n9787 = pi142 & n9786;
  assign n9788 = pi145 & ~n7035;
  assign n9789 = n9505 & n9788;
  assign n9790 = ~n9787 & ~n9789;
  assign n9791 = pi141 & ~n9790;
  assign n9792 = pi145 & n7035;
  assign n9793 = n9495 & n9792;
  assign n9794 = ~pi144 & ~pi145;
  assign n9795 = ~pi142 & n9794;
  assign n9796 = ~n9793 & ~n9795;
  assign n9797 = ~pi141 & ~n9796;
  assign n9798 = ~pi144 & pi145;
  assign n9799 = pi143 & n9798;
  assign n9800 = ~pi145 & ~n7035;
  assign n9801 = pi144 & n9800;
  assign n9802 = ~n9799 & ~n9801;
  assign n9803 = pi142 & ~n9802;
  assign n9804 = pi144 & pi145;
  assign n9805 = ~pi143 & n9804;
  assign n9806 = ~pi145 & n7035;
  assign n9807 = ~pi144 & n9806;
  assign n9808 = ~n9805 & ~n9807;
  assign n9809 = ~pi142 & ~n9808;
  assign n9810 = ~n9499 & ~n9510;
  assign n9811 = ~pi145 & ~n9810;
  assign n9812 = ~n9809 & ~n9811;
  assign n9813 = ~n9803 & n9812;
  assign n9814 = ~n9797 & n9813;
  assign n9815 = ~n9791 & n9814;
  assign n9816 = pi321 & n9815;
  assign n9817 = ~n9518 & n9524;
  assign n9818 = n7874 & ~n9817;
  assign n9819 = pi320 & n9818;
  assign n9820 = n9517 & ~n9524;
  assign n9821 = pi321 & n9820;
  assign n9822 = ~n9819 & ~n9821;
  assign n9823 = pi320 & n9517;
  assign n9824 = ~n9822 & ~n9823;
  assign n9825 = n9517 & n9822;
  assign n9826 = pi320 & n9825;
  assign n9827 = ~n9824 & ~n9826;
  assign n9828 = ~n9816 & ~n9827;
  assign n9829 = n9822 & ~n9823;
  assign n9830 = n9517 & ~n9822;
  assign n9831 = pi320 & n9830;
  assign n9832 = ~n9829 & ~n9831;
  assign n9833 = n9815 & ~n9832;
  assign n9834 = pi321 & n9833;
  assign n9835 = ~n9828 & ~n9834;
  assign n9836 = pi319 & n7874;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = n7874 & n9835;
  assign n9839 = pi319 & n9838;
  assign n9840 = ~n9837 & ~n9839;
  assign n9841 = n7044 & ~n9542;
  assign n9842 = pi319 & n9841;
  assign n9843 = ~n9541 & ~n9842;
  assign n9844 = n9840 & n9843;
  assign n9845 = ~n9840 & ~n9843;
  assign n9846 = ~n9844 & ~n9845;
  assign n9847 = n7044 & ~n9846;
  assign n9848 = pi318 & n9847;
  assign n9849 = pi318 & n7044;
  assign n9850 = ~n9840 & n9843;
  assign n9851 = n9840 & ~n9843;
  assign n9852 = ~n9850 & ~n9851;
  assign n9853 = ~n9849 & ~n9852;
  assign n9854 = ~n9848 & ~n9853;
  assign n9855 = ~n9551 & ~n9561;
  assign n9856 = n9551 & n9561;
  assign n9857 = n6777 & ~n9856;
  assign n9858 = pi318 & n9857;
  assign n9859 = ~n9855 & ~n9858;
  assign n9860 = n9854 & ~n9859;
  assign n9861 = ~n9854 & n9859;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = n6777 & ~n9862;
  assign n9864 = pi317 & n9863;
  assign n9865 = pi317 & n6777;
  assign n9866 = n9862 & ~n9865;
  assign n9867 = ~n9864 & ~n9866;
  assign n9868 = ~n9565 & ~n9574;
  assign n9869 = n9565 & n9574;
  assign n9870 = ~n7932 & ~n9869;
  assign n9871 = ~n7921 & n9870;
  assign n9872 = ~n9868 & ~n9871;
  assign n9873 = pi316 & n5463;
  assign n9874 = n9872 & ~n9873;
  assign n9875 = n5463 & ~n9872;
  assign n9876 = pi316 & n9875;
  assign n9877 = ~n9874 & ~n9876;
  assign n9878 = ~n9867 & ~n9877;
  assign n9879 = ~n9872 & ~n9873;
  assign n9880 = n5463 & n9872;
  assign n9881 = pi316 & n9880;
  assign n9882 = ~n9879 & ~n9881;
  assign n9883 = ~n9866 & ~n9882;
  assign n9884 = ~n9864 & n9883;
  assign n9885 = ~n9878 & ~n9884;
  assign n9886 = ~n7940 & ~n9595;
  assign n9887 = ~n4772 & n9580;
  assign n9888 = n4086 & ~n9887;
  assign n9889 = pi316 & n9888;
  assign n9890 = ~n9886 & ~n9889;
  assign n9891 = ~n7929 & ~n9890;
  assign n9892 = n4772 & ~n9580;
  assign n9893 = ~n7940 & n9888;
  assign n9894 = ~n9892 & ~n9893;
  assign n9895 = pi316 & ~n9894;
  assign n9896 = ~n9891 & ~n9895;
  assign n9897 = n9885 & n9896;
  assign n9898 = ~n9885 & ~n9896;
  assign n9899 = ~n9897 & ~n9898;
  assign n9900 = n4772 & ~n9899;
  assign n9901 = pi315 & n9900;
  assign n9902 = pi315 & n4772;
  assign n9903 = ~n9885 & n9896;
  assign n9904 = n9885 & ~n9896;
  assign n9905 = ~n9903 & ~n9904;
  assign n9906 = ~n9902 & ~n9905;
  assign n9907 = ~n9901 & ~n9906;
  assign n9908 = n9584 & ~n9606;
  assign n9909 = ~n4086 & n4772;
  assign n9910 = pi316 & n9580;
  assign n9911 = n9909 & n9910;
  assign n9912 = ~n4086 & ~n4772;
  assign n9913 = pi316 & ~n9912;
  assign n9914 = ~n9580 & ~n9913;
  assign n9915 = ~n9911 & ~n9914;
  assign n9916 = ~n9585 & ~n9915;
  assign n9917 = ~n4772 & ~n9580;
  assign n9918 = ~n9582 & ~n9917;
  assign n9919 = n7940 & ~n9918;
  assign n9920 = n7929 & n9919;
  assign n9921 = ~n4086 & n7940;
  assign n9922 = n4772 & ~n9921;
  assign n9923 = ~n9580 & n9922;
  assign n9924 = n4086 & ~n4772;
  assign n9925 = n9580 & n9924;
  assign n9926 = ~n9923 & ~n9925;
  assign n9927 = pi316 & ~n9926;
  assign n9928 = ~n7940 & n9595;
  assign n9929 = ~n9927 & ~n9928;
  assign n9930 = ~n7929 & ~n9929;
  assign n9931 = ~n9887 & ~n9892;
  assign n9932 = n4086 & ~n9931;
  assign n9933 = pi316 & n9932;
  assign n9934 = ~n7940 & n9933;
  assign n9935 = ~n9930 & ~n9934;
  assign n9936 = ~n9920 & n9935;
  assign n9937 = ~n9916 & n9936;
  assign n9938 = ~n9584 & n9606;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = ~n9908 & ~n9939;
  assign n9941 = n9907 & n9940;
  assign n9942 = ~n9907 & ~n9940;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = pi314 & n4086;
  assign n9945 = ~n9617 & ~n9944;
  assign n9946 = ~n9611 & n9945;
  assign n9947 = ~n9611 & ~n9617;
  assign n9948 = n9944 & ~n9947;
  assign n9949 = ~n9946 & ~n9948;
  assign n9950 = ~n9943 & ~n9949;
  assign n9951 = n9907 & ~n9940;
  assign n9952 = ~n9907 & n9940;
  assign n9953 = ~n9951 & ~n9952;
  assign n9954 = ~n9617 & n9944;
  assign n9955 = ~n9611 & n9954;
  assign n9956 = ~n9944 & ~n9947;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~n9953 & ~n9957;
  assign n9959 = ~n9950 & ~n9958;
  assign n9960 = ~n9785 & n9959;
  assign n9961 = n9785 & ~n9959;
  assign n9962 = ~n9960 & ~n9961;
  assign n9963 = pi312 & n3012;
  assign n9964 = n7166 & ~n7989;
  assign n9965 = n2183 & ~n9646;
  assign n9966 = pi313 & n9965;
  assign n9967 = ~n9964 & ~n9966;
  assign n9968 = ~n7015 & ~n9967;
  assign n9969 = n7166 & n9965;
  assign n9970 = ~n9647 & ~n9969;
  assign n9971 = pi313 & ~n9970;
  assign n9972 = ~n9968 & ~n9971;
  assign n9973 = n9619 & ~n9972;
  assign n9974 = ~n9619 & n9972;
  assign n9975 = n9479 & ~n9974;
  assign n9976 = ~n9973 & ~n9975;
  assign n9977 = n9963 & ~n9976;
  assign n9978 = ~n9479 & ~n9973;
  assign n9979 = ~n9974 & ~n9978;
  assign n9980 = ~n9963 & ~n9979;
  assign n9981 = ~n9977 & ~n9980;
  assign n9982 = ~n9962 & ~n9981;
  assign n9983 = ~n9785 & ~n9959;
  assign n9984 = n9785 & n9959;
  assign n9985 = ~n9983 & ~n9984;
  assign n9986 = ~n9963 & ~n9976;
  assign n9987 = n9963 & ~n9979;
  assign n9988 = ~n9986 & ~n9987;
  assign n9989 = ~n9985 & ~n9988;
  assign n9990 = ~n9982 & ~n9989;
  assign n9991 = n9623 & ~n9667;
  assign n9992 = ~n9623 & n9667;
  assign n9993 = ~n9658 & ~n9992;
  assign n9994 = ~n9991 & ~n9993;
  assign n9995 = n9990 & n9994;
  assign n9996 = ~n9990 & ~n9994;
  assign n9997 = ~n9995 & ~n9996;
  assign n9998 = pi311 & n2574;
  assign n9999 = n9678 & ~n9679;
  assign n10000 = ~n9680 & ~n9999;
  assign n10001 = n9998 & ~n10000;
  assign n10002 = ~n9678 & ~n9680;
  assign n10003 = ~n9679 & ~n10002;
  assign n10004 = ~n9998 & ~n10003;
  assign n10005 = ~n10001 & ~n10004;
  assign n10006 = ~n9997 & ~n10005;
  assign n10007 = n9990 & ~n9994;
  assign n10008 = ~n9990 & n9994;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = ~n9998 & ~n10000;
  assign n10011 = n9998 & ~n10003;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = ~n10009 & ~n10012;
  assign n10014 = ~n10006 & ~n10013;
  assign n10015 = ~pi310 & n10014;
  assign n10016 = ~n2183 & n10014;
  assign n10017 = n2183 & ~n10014;
  assign n10018 = pi310 & n10017;
  assign n10019 = ~n10016 & ~n10018;
  assign n10020 = ~n1840 & ~n10019;
  assign n10021 = ~n10015 & ~n10020;
  assign n10022 = ~n9689 & ~n10021;
  assign n10023 = ~n9688 & ~n10019;
  assign n10024 = n1840 & n9688;
  assign n10025 = n2183 & n10014;
  assign n10026 = n10024 & n10025;
  assign n10027 = ~n10023 & ~n10026;
  assign n10028 = ~n9683 & ~n10027;
  assign n10029 = n9688 & n10025;
  assign n10030 = ~n2183 & ~n10014;
  assign n10031 = n1840 & n10030;
  assign n10032 = ~n10029 & ~n10031;
  assign n10033 = pi310 & ~n10032;
  assign n10034 = pi310 & n2183;
  assign n10035 = ~n10014 & ~n10034;
  assign n10036 = n9688 & n10035;
  assign n10037 = n1840 & ~n9688;
  assign n10038 = n10025 & n10037;
  assign n10039 = ~n10036 & ~n10038;
  assign n10040 = ~n10033 & n10039;
  assign n10041 = n9683 & ~n10040;
  assign n10042 = n9688 & n10030;
  assign n10043 = n9694 & n10042;
  assign n10044 = ~n10041 & ~n10043;
  assign n10045 = ~n10028 & n10044;
  assign n10046 = ~n10022 & n10045;
  assign n10047 = ~n9784 & ~n10046;
  assign n10048 = n9784 & n10046;
  assign n10049 = ~n10047 & ~n10048;
  assign n10050 = pi308 & n1533;
  assign n10051 = ~n9466 & ~n9699;
  assign n10052 = n9466 & n9699;
  assign n10053 = n9464 & ~n10052;
  assign n10054 = ~n10051 & ~n10053;
  assign n10055 = n10050 & ~n10054;
  assign n10056 = ~n9464 & ~n10051;
  assign n10057 = ~n10052 & ~n10056;
  assign n10058 = ~n10050 & ~n10057;
  assign n10059 = ~n10055 & ~n10058;
  assign n10060 = ~n10049 & ~n10059;
  assign n10061 = ~n9784 & n10046;
  assign n10062 = n9784 & ~n10046;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10050 & ~n10054;
  assign n10065 = n10050 & ~n10057;
  assign n10066 = ~n10064 & ~n10065;
  assign n10067 = ~n10063 & ~n10066;
  assign n10068 = ~n10060 & ~n10067;
  assign n10069 = ~n9702 & ~n9703;
  assign n10070 = n9702 & n9703;
  assign n10071 = ~n9722 & ~n10070;
  assign n10072 = ~n10069 & ~n10071;
  assign n10073 = n10068 & ~n10072;
  assign n10074 = ~n10068 & n10072;
  assign n10075 = ~n10073 & ~n10074;
  assign n10076 = ~n9454 & ~n9740;
  assign n10077 = ~n9453 & ~n10076;
  assign n10078 = n10075 & ~n10077;
  assign n10079 = ~n10075 & n10077;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = ~n1515 & ~n9733;
  assign n10082 = n1515 & n9733;
  assign n10083 = n9461 & ~n10082;
  assign n10084 = ~n10081 & ~n10083;
  assign n10085 = n1553 & ~n10084;
  assign n10086 = n9461 & ~n9733;
  assign n10087 = ~n1553 & ~n10086;
  assign n10088 = n1515 & n10087;
  assign n10089 = ~n10085 & ~n10088;
  assign n10090 = pi307 & ~n10089;
  assign n10091 = pi307 & n1553;
  assign n10092 = n9733 & ~n10091;
  assign n10093 = ~n9461 & n10092;
  assign n10094 = ~n10090 & ~n10093;
  assign n10095 = pi306 & n1515;
  assign n10096 = n10094 & ~n10095;
  assign n10097 = n1515 & ~n10094;
  assign n10098 = pi306 & n10097;
  assign n10099 = ~n10096 & ~n10098;
  assign n10100 = ~n10080 & ~n10099;
  assign n10101 = ~n10075 & ~n10077;
  assign n10102 = n10075 & n10077;
  assign n10103 = ~n10101 & ~n10102;
  assign n10104 = ~n10094 & ~n10095;
  assign n10105 = n1515 & n10094;
  assign n10106 = pi306 & n10105;
  assign n10107 = ~n10104 & ~n10106;
  assign n10108 = ~n10103 & ~n10107;
  assign n10109 = ~n10100 & ~n10108;
  assign n10110 = ~n9783 & n10109;
  assign n10111 = n9783 & ~n10109;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = pi304 & ~n10112;
  assign n10114 = pi128 & n10113;
  assign n10115 = pi128 & pi304;
  assign n10116 = n9783 & n10109;
  assign n10117 = ~n9783 & ~n10109;
  assign n10118 = ~n10116 & ~n10117;
  assign n10119 = ~n10115 & ~n10118;
  assign n10120 = ~n10114 & ~n10119;
  assign n10121 = n1156 & n9426;
  assign n10122 = ~n1154 & ~n10121;
  assign n10123 = n1154 & n9426;
  assign n10124 = n1156 & n10123;
  assign n10125 = ~n10122 & ~n10124;
  assign n10126 = pi338 & ~n10125;
  assign n10127 = ~n8786 & n8810;
  assign n10128 = n8786 & ~n8810;
  assign n10129 = n9347 & ~n10128;
  assign n10130 = ~n10127 & ~n10129;
  assign n10131 = n8786 & ~n9347;
  assign n10132 = ~n8786 & n9347;
  assign n10133 = ~n10131 & ~n10132;
  assign n10134 = n8806 & n9351;
  assign n10135 = n8810 & ~n9374;
  assign n10136 = ~n8810 & n9374;
  assign n10137 = ~n10135 & ~n10136;
  assign n10138 = ~n10134 & ~n10137;
  assign n10139 = ~n10133 & n10138;
  assign n10140 = n8786 & n9347;
  assign n10141 = ~n8786 & ~n9347;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = ~n8810 & ~n9374;
  assign n10144 = n8810 & n9374;
  assign n10145 = ~n10143 & ~n10144;
  assign n10146 = ~n10134 & ~n10145;
  assign n10147 = ~n10142 & n10146;
  assign n10148 = ~n8806 & ~n9351;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = ~n10139 & n10149;
  assign n10151 = ~n10130 & ~n10150;
  assign n10152 = n10130 & n10150;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = pi333 & n2464;
  assign n10155 = ~n8815 & ~n9267;
  assign n10156 = n8815 & n9267;
  assign n10157 = n5714 & ~n10156;
  assign n10158 = pi328 & n10157;
  assign n10159 = ~n10155 & ~n10158;
  assign n10160 = ~n8827 & ~n8831;
  assign n10161 = n8827 & n8831;
  assign n10162 = ~n8815 & n9267;
  assign n10163 = n8815 & ~n9267;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = n5714 & ~n10164;
  assign n10166 = pi328 & n10165;
  assign n10167 = ~n10155 & ~n10156;
  assign n10168 = ~n9273 & ~n10167;
  assign n10169 = ~n10166 & ~n10168;
  assign n10170 = ~n10161 & ~n10169;
  assign n10171 = ~n10160 & ~n10170;
  assign n10172 = n10159 & n10171;
  assign n10173 = ~n10159 & ~n10171;
  assign n10174 = ~n10172 & ~n10173;
  assign n10175 = pi329 & n5714;
  assign n10176 = ~n8835 & n9246;
  assign n10177 = n8835 & ~n9246;
  assign n10178 = ~n9253 & ~n10177;
  assign n10179 = ~n10176 & ~n10178;
  assign n10180 = ~n8835 & ~n9241;
  assign n10181 = n8835 & n9241;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = n8855 & n9245;
  assign n10184 = ~n9226 & n9246;
  assign n10185 = n9226 & ~n9246;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = ~n10183 & ~n10186;
  assign n10188 = ~n10182 & n10187;
  assign n10189 = ~n8835 & n9241;
  assign n10190 = n8835 & ~n9241;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = n9226 & n9246;
  assign n10193 = ~n9226 & ~n9246;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = ~n10183 & ~n10194;
  assign n10196 = ~n10191 & n10195;
  assign n10197 = ~n8855 & ~n9245;
  assign n10198 = ~n10196 & ~n10197;
  assign n10199 = ~n10188 & n10198;
  assign n10200 = n10179 & n10199;
  assign n10201 = ~n10179 & ~n10199;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = ~n8860 & ~n9192;
  assign n10204 = ~n9200 & ~n10203;
  assign n10205 = ~n8868 & n9206;
  assign n10206 = ~n8860 & ~n9201;
  assign n10207 = n8860 & ~n9200;
  assign n10208 = ~n9192 & n10207;
  assign n10209 = ~n10206 & ~n10208;
  assign n10210 = n8868 & ~n9206;
  assign n10211 = ~n10209 & ~n10210;
  assign n10212 = ~n10205 & ~n10211;
  assign n10213 = ~n10204 & n10212;
  assign n10214 = n10204 & ~n10212;
  assign n10215 = ~n10213 & ~n10214;
  assign n10216 = ~n7601 & ~n9179;
  assign n10217 = ~n9178 & ~n10216;
  assign n10218 = n9167 & n10217;
  assign n10219 = ~n9167 & ~n10217;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = ~n8513 & ~n10220;
  assign n10222 = ~n9167 & n10217;
  assign n10223 = n9167 & ~n10217;
  assign n10224 = ~n10222 & ~n10223;
  assign n10225 = n8513 & ~n10224;
  assign n10226 = ~n10221 & ~n10225;
  assign n10227 = pi323 & ~n10226;
  assign n10228 = pi145 & pi258;
  assign n10229 = ~n9167 & n10228;
  assign n10230 = n9167 & ~n10228;
  assign n10231 = ~n10229 & ~n10230;
  assign n10232 = ~n9124 & n9147;
  assign n10233 = n9124 & ~n9147;
  assign n10234 = ~n9118 & ~n10233;
  assign n10235 = ~n10232 & ~n10234;
  assign n10236 = pi260 & ~n9161;
  assign n10237 = pi142 & n10236;
  assign n10238 = ~n9127 & ~n9147;
  assign n10239 = ~n9144 & ~n10238;
  assign n10240 = ~n10237 & n10239;
  assign n10241 = ~n9133 & ~n10240;
  assign n10242 = n10235 & ~n10241;
  assign n10243 = ~n10235 & n10241;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = pi143 & pi260;
  assign n10246 = pi131 & pi272;
  assign n10247 = ~n8905 & ~n8920;
  assign n10248 = n8905 & n8920;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = pi271 & ~n10249;
  assign n10251 = pi131 & n10250;
  assign n10252 = pi130 & pi273;
  assign n10253 = pi128 & pi275;
  assign n10254 = pi274 & ~n10253;
  assign n10255 = pi129 & n10254;
  assign n10256 = pi129 & pi274;
  assign n10257 = pi275 & ~n10256;
  assign n10258 = pi128 & n10257;
  assign n10259 = ~n10255 & ~n10258;
  assign n10260 = n8890 & ~n8895;
  assign n10261 = n10259 & ~n10260;
  assign n10262 = ~n8893 & n10261;
  assign n10263 = ~n8893 & ~n10260;
  assign n10264 = ~n10259 & ~n10263;
  assign n10265 = ~n10262 & ~n10264;
  assign n10266 = ~n10252 & ~n10265;
  assign n10267 = n10259 & ~n10263;
  assign n10268 = ~n10259 & ~n10260;
  assign n10269 = ~n8893 & n10268;
  assign n10270 = ~n10267 & ~n10269;
  assign n10271 = pi273 & ~n10270;
  assign n10272 = pi130 & n10271;
  assign n10273 = ~n10266 & ~n10272;
  assign n10274 = ~n8901 & n8920;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 = ~n8904 & n10275;
  assign n10277 = ~n8904 & ~n10274;
  assign n10278 = n10273 & ~n10277;
  assign n10279 = ~n10276 & ~n10278;
  assign n10280 = ~n8921 & ~n10248;
  assign n10281 = ~n10247 & n10280;
  assign n10282 = ~n8938 & ~n10281;
  assign n10283 = ~n10279 & ~n10282;
  assign n10284 = ~n10251 & n10283;
  assign n10285 = ~n10251 & ~n10282;
  assign n10286 = n10279 & ~n10285;
  assign n10287 = ~n10284 & ~n10286;
  assign n10288 = ~n10246 & ~n10287;
  assign n10289 = n10279 & ~n10282;
  assign n10290 = ~n10251 & n10289;
  assign n10291 = ~n10279 & ~n10285;
  assign n10292 = ~n10290 & ~n10291;
  assign n10293 = pi272 & ~n10292;
  assign n10294 = pi131 & n10293;
  assign n10295 = ~n10288 & ~n10294;
  assign n10296 = n8942 & ~n8953;
  assign n10297 = ~n8942 & n8953;
  assign n10298 = ~n8944 & ~n10297;
  assign n10299 = ~n10296 & ~n10298;
  assign n10300 = n10295 & n10299;
  assign n10301 = ~n10295 & ~n10299;
  assign n10302 = ~n10300 & ~n10301;
  assign n10303 = pi133 & pi270;
  assign n10304 = pi132 & pi271;
  assign n10305 = n10303 & n10304;
  assign n10306 = ~n10303 & ~n10304;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n10302 & ~n10307;
  assign n10309 = ~n10295 & n10299;
  assign n10310 = n10295 & ~n10299;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = pi270 & ~n10304;
  assign n10313 = pi133 & n10312;
  assign n10314 = pi271 & ~n10303;
  assign n10315 = pi132 & n10314;
  assign n10316 = ~n10313 & ~n10315;
  assign n10317 = ~n10311 & ~n10316;
  assign n10318 = ~n10308 & ~n10317;
  assign n10319 = ~n8974 & ~n8978;
  assign n10320 = ~n8979 & ~n10319;
  assign n10321 = n10318 & n10320;
  assign n10322 = ~n10318 & ~n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = pi134 & pi269;
  assign n10325 = n8958 & ~n8971;
  assign n10326 = ~n8967 & n10325;
  assign n10327 = ~n8958 & ~n8974;
  assign n10328 = ~n10326 & ~n10327;
  assign n10329 = ~n8876 & ~n10328;
  assign n10330 = ~n8958 & ~n8971;
  assign n10331 = ~n8967 & n10330;
  assign n10332 = n8958 & ~n8974;
  assign n10333 = ~n10331 & ~n10332;
  assign n10334 = pi269 & ~n10333;
  assign n10335 = pi133 & n10334;
  assign n10336 = ~n10329 & ~n10335;
  assign n10337 = ~n8990 & ~n10336;
  assign n10338 = n8990 & n10336;
  assign n10339 = n8968 & ~n10338;
  assign n10340 = ~n10337 & ~n10339;
  assign n10341 = n10324 & ~n10340;
  assign n10342 = ~n8968 & ~n10337;
  assign n10343 = ~n10338 & ~n10342;
  assign n10344 = ~n10324 & ~n10343;
  assign n10345 = ~n10341 & ~n10344;
  assign n10346 = ~n10323 & ~n10345;
  assign n10347 = n10318 & ~n10320;
  assign n10348 = ~n10318 & n10320;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = ~n10324 & ~n10340;
  assign n10351 = n10324 & ~n10343;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = ~n10349 & ~n10352;
  assign n10354 = ~n10346 & ~n10353;
  assign n10355 = ~n8993 & ~n8994;
  assign n10356 = n8993 & n8994;
  assign n10357 = ~n8999 & ~n10356;
  assign n10358 = ~n10355 & ~n10357;
  assign n10359 = ~n10354 & n10358;
  assign n10360 = n10354 & ~n10358;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = pi136 & pi267;
  assign n10363 = pi135 & pi268;
  assign n10364 = n10362 & n10363;
  assign n10365 = ~n10362 & ~n10363;
  assign n10366 = ~n10364 & ~n10365;
  assign n10367 = ~n10361 & ~n10366;
  assign n10368 = n10354 & n10358;
  assign n10369 = ~n10354 & ~n10358;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = pi267 & ~n10363;
  assign n10372 = pi136 & n10371;
  assign n10373 = pi268 & ~n10362;
  assign n10374 = pi135 & n10373;
  assign n10375 = ~n10372 & ~n10374;
  assign n10376 = ~n10370 & ~n10375;
  assign n10377 = ~n10367 & ~n10376;
  assign n10378 = ~n9026 & ~n9030;
  assign n10379 = ~n9031 & ~n10378;
  assign n10380 = n10377 & n10379;
  assign n10381 = ~n10377 & ~n10379;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = pi137 & pi266;
  assign n10384 = n9010 & ~n9023;
  assign n10385 = ~n9019 & n10384;
  assign n10386 = ~n9010 & ~n9026;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n8875 & ~n10387;
  assign n10389 = ~n9010 & ~n9023;
  assign n10390 = ~n9019 & n10389;
  assign n10391 = n9010 & ~n9026;
  assign n10392 = ~n10390 & ~n10391;
  assign n10393 = pi266 & ~n10392;
  assign n10394 = pi136 & n10393;
  assign n10395 = ~n10388 & ~n10394;
  assign n10396 = ~n9042 & ~n10395;
  assign n10397 = n9042 & n10395;
  assign n10398 = n9020 & ~n10397;
  assign n10399 = ~n10396 & ~n10398;
  assign n10400 = n10383 & ~n10399;
  assign n10401 = ~n9020 & ~n10396;
  assign n10402 = ~n10397 & ~n10401;
  assign n10403 = ~n10383 & ~n10402;
  assign n10404 = ~n10400 & ~n10403;
  assign n10405 = ~n10382 & ~n10404;
  assign n10406 = n10377 & ~n10379;
  assign n10407 = ~n10377 & n10379;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = ~n10383 & ~n10399;
  assign n10410 = n10383 & ~n10402;
  assign n10411 = ~n10409 & ~n10410;
  assign n10412 = ~n10408 & ~n10411;
  assign n10413 = ~n10405 & ~n10412;
  assign n10414 = ~n9046 & ~n9057;
  assign n10415 = n9046 & n9057;
  assign n10416 = ~n9051 & ~n10415;
  assign n10417 = ~n10414 & ~n10416;
  assign n10418 = ~n10413 & n10417;
  assign n10419 = n10413 & ~n10417;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = pi139 & pi264;
  assign n10422 = pi138 & pi265;
  assign n10423 = n10421 & n10422;
  assign n10424 = ~n10421 & ~n10422;
  assign n10425 = ~n10423 & ~n10424;
  assign n10426 = ~n10420 & ~n10425;
  assign n10427 = n10413 & n10417;
  assign n10428 = ~n10413 & ~n10417;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = pi264 & ~n10422;
  assign n10431 = pi139 & n10430;
  assign n10432 = pi265 & ~n10421;
  assign n10433 = pi138 & n10432;
  assign n10434 = ~n10431 & ~n10433;
  assign n10435 = ~n10429 & ~n10434;
  assign n10436 = ~n10426 & ~n10435;
  assign n10437 = ~n9075 & ~n9082;
  assign n10438 = ~n9070 & n10437;
  assign n10439 = ~n9083 & ~n10438;
  assign n10440 = n10436 & n10439;
  assign n10441 = ~n10436 & ~n10439;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = pi140 & pi263;
  assign n10444 = ~n9062 & ~n9075;
  assign n10445 = ~n9070 & n10444;
  assign n10446 = n9062 & ~n9078;
  assign n10447 = ~n10445 & ~n10446;
  assign n10448 = ~n8874 & ~n10447;
  assign n10449 = n9062 & ~n9075;
  assign n10450 = ~n9070 & n10449;
  assign n10451 = ~n9062 & ~n9078;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = pi263 & ~n10452;
  assign n10454 = pi139 & n10453;
  assign n10455 = ~n10448 & ~n10454;
  assign n10456 = n9094 & n10455;
  assign n10457 = ~n9094 & ~n10455;
  assign n10458 = n9071 & ~n10457;
  assign n10459 = ~n10456 & ~n10458;
  assign n10460 = n10443 & ~n10459;
  assign n10461 = ~n9071 & ~n10456;
  assign n10462 = ~n10457 & ~n10461;
  assign n10463 = ~n10443 & ~n10462;
  assign n10464 = ~n10460 & ~n10463;
  assign n10465 = ~n10442 & ~n10464;
  assign n10466 = n10436 & ~n10439;
  assign n10467 = ~n10436 & n10439;
  assign n10468 = ~n10466 & ~n10467;
  assign n10469 = ~n10443 & ~n10459;
  assign n10470 = n10443 & ~n10462;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = ~n10468 & ~n10471;
  assign n10473 = ~n10465 & ~n10472;
  assign n10474 = ~n9101 & ~n9112;
  assign n10475 = n9101 & n9112;
  assign n10476 = ~n9103 & ~n10475;
  assign n10477 = ~n9100 & n10476;
  assign n10478 = ~n10474 & ~n10477;
  assign n10479 = ~n10473 & n10478;
  assign n10480 = n10473 & ~n10478;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = pi142 & pi261;
  assign n10483 = pi141 & pi262;
  assign n10484 = n10482 & n10483;
  assign n10485 = ~n10482 & ~n10483;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = ~n10481 & ~n10486;
  assign n10488 = n10473 & n10478;
  assign n10489 = ~n10473 & ~n10478;
  assign n10490 = ~n10488 & ~n10489;
  assign n10491 = pi261 & ~n10483;
  assign n10492 = pi142 & n10491;
  assign n10493 = pi262 & ~n10482;
  assign n10494 = pi141 & n10493;
  assign n10495 = ~n10492 & ~n10494;
  assign n10496 = ~n10490 & ~n10495;
  assign n10497 = ~n10487 & ~n10496;
  assign n10498 = ~n10245 & n10497;
  assign n10499 = n10245 & ~n10497;
  assign n10500 = ~n10498 & ~n10499;
  assign n10501 = ~n9144 & ~n9147;
  assign n10502 = ~n9133 & n10501;
  assign n10503 = ~n9145 & n9147;
  assign n10504 = ~n10502 & ~n10503;
  assign n10505 = ~n9161 & ~n10504;
  assign n10506 = ~n9144 & n9147;
  assign n10507 = ~n9133 & n10506;
  assign n10508 = ~n9145 & ~n9147;
  assign n10509 = ~n10507 & ~n10508;
  assign n10510 = ~n9127 & ~n10509;
  assign n10511 = ~n10505 & ~n10510;
  assign n10512 = n9146 & ~n10511;
  assign n10513 = pi144 & pi259;
  assign n10514 = n10512 & n10513;
  assign n10515 = ~n10512 & ~n10513;
  assign n10516 = ~n10514 & ~n10515;
  assign n10517 = ~n10500 & ~n10516;
  assign n10518 = n10245 & n10497;
  assign n10519 = ~n10245 & ~n10497;
  assign n10520 = ~n10518 & ~n10519;
  assign n10521 = ~n10512 & n10513;
  assign n10522 = n10512 & ~n10513;
  assign n10523 = ~n10521 & ~n10522;
  assign n10524 = ~n10520 & ~n10523;
  assign n10525 = ~n10517 & ~n10524;
  assign n10526 = ~n10244 & ~n10525;
  assign n10527 = n10235 & n10241;
  assign n10528 = ~n10235 & ~n10241;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = ~n10516 & ~n10520;
  assign n10531 = ~n10500 & ~n10523;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = ~n10529 & ~n10532;
  assign n10534 = ~n10526 & ~n10533;
  assign n10535 = ~n8513 & ~n10218;
  assign n10536 = ~n10219 & ~n10535;
  assign n10537 = n10534 & ~n10536;
  assign n10538 = ~n10534 & n10536;
  assign n10539 = ~n10537 & ~n10538;
  assign n10540 = ~n10231 & ~n10539;
  assign n10541 = n10534 & n10536;
  assign n10542 = ~n10534 & ~n10536;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = n9167 & n10228;
  assign n10545 = ~n9167 & ~n10228;
  assign n10546 = ~n10544 & ~n10545;
  assign n10547 = ~n10543 & ~n10546;
  assign n10548 = pi322 & ~n10547;
  assign n10549 = ~n10540 & n10548;
  assign n10550 = ~n10227 & ~n10549;
  assign n10551 = pi322 & ~n10226;
  assign n10552 = ~n10231 & ~n10543;
  assign n10553 = ~n10539 & ~n10546;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = n10551 & ~n10554;
  assign n10556 = pi323 & n10555;
  assign n10557 = ~n10550 & ~n10556;
  assign n10558 = pi325 & n9205;
  assign n10559 = ~n7601 & ~n9187;
  assign n10560 = n7601 & ~n9180;
  assign n10561 = ~n10559 & ~n10560;
  assign n10562 = pi324 & n10561;
  assign n10563 = n10558 & n10562;
  assign n10564 = ~n10558 & ~n10562;
  assign n10565 = ~n10563 & ~n10564;
  assign n10566 = ~n10557 & ~n10565;
  assign n10567 = ~n10558 & n10562;
  assign n10568 = n10558 & ~n10562;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = ~n10556 & ~n10569;
  assign n10571 = ~n10550 & n10570;
  assign n10572 = ~n10566 & ~n10571;
  assign n10573 = ~n10215 & ~n10572;
  assign n10574 = ~n10204 & ~n10212;
  assign n10575 = n10204 & n10212;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = ~n10557 & ~n10569;
  assign n10578 = ~n10556 & ~n10565;
  assign n10579 = ~n10550 & n10578;
  assign n10580 = ~n10577 & ~n10579;
  assign n10581 = ~n10576 & ~n10580;
  assign n10582 = ~n10573 & ~n10581;
  assign n10583 = n9202 & ~n9241;
  assign n10584 = ~n9206 & ~n10209;
  assign n10585 = n8860 & ~n9201;
  assign n10586 = ~n8860 & ~n9200;
  assign n10587 = ~n9192 & n10586;
  assign n10588 = ~n10585 & ~n10587;
  assign n10589 = n9205 & ~n10588;
  assign n10590 = pi324 & n10589;
  assign n10591 = ~n10584 & ~n10590;
  assign n10592 = n8868 & ~n10591;
  assign n10593 = ~n8868 & n10591;
  assign n10594 = ~n10592 & ~n10593;
  assign n10595 = ~n9202 & n9241;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10583 & ~n10596;
  assign n10598 = n10582 & n10597;
  assign n10599 = ~n10582 & ~n10597;
  assign n10600 = ~n10598 & ~n10599;
  assign n10601 = pi327 & n5973;
  assign n10602 = pi326 & n6556;
  assign n10603 = n10601 & n10602;
  assign n10604 = ~n10601 & ~n10602;
  assign n10605 = ~n10603 & ~n10604;
  assign n10606 = ~n10600 & ~n10605;
  assign n10607 = ~n10582 & n10597;
  assign n10608 = n10582 & ~n10597;
  assign n10609 = ~n10607 & ~n10608;
  assign n10610 = ~n10601 & n10602;
  assign n10611 = n10601 & ~n10602;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = ~n10609 & ~n10612;
  assign n10614 = ~n10606 & ~n10613;
  assign n10615 = ~n10202 & ~n10614;
  assign n10616 = n10179 & ~n10199;
  assign n10617 = ~n10179 & n10199;
  assign n10618 = ~n10616 & ~n10617;
  assign n10619 = ~n10605 & ~n10609;
  assign n10620 = ~n10600 & ~n10612;
  assign n10621 = ~n10619 & ~n10620;
  assign n10622 = ~n10618 & ~n10621;
  assign n10623 = ~n10615 & ~n10622;
  assign n10624 = ~n10175 & n10623;
  assign n10625 = n10175 & ~n10623;
  assign n10626 = ~n10624 & ~n10625;
  assign n10627 = n5732 & ~n10626;
  assign n10628 = pi328 & n10627;
  assign n10629 = pi328 & n5732;
  assign n10630 = n10175 & n10623;
  assign n10631 = ~n10175 & ~n10623;
  assign n10632 = ~n10630 & ~n10631;
  assign n10633 = ~n10629 & ~n10632;
  assign n10634 = ~n10628 & ~n10633;
  assign n10635 = ~n10174 & ~n10634;
  assign n10636 = n10159 & ~n10171;
  assign n10637 = ~n10159 & n10171;
  assign n10638 = ~n10636 & ~n10637;
  assign n10639 = n5732 & ~n10632;
  assign n10640 = pi328 & n10639;
  assign n10641 = ~n10626 & ~n10629;
  assign n10642 = ~n10640 & ~n10641;
  assign n10643 = ~n10638 & ~n10642;
  assign n10644 = ~n10635 & ~n10643;
  assign n10645 = ~n9305 & n9309;
  assign n10646 = ~n9288 & ~n9316;
  assign n10647 = n9288 & n9316;
  assign n10648 = ~n10646 & ~n10647;
  assign n10649 = n9305 & ~n9309;
  assign n10650 = ~n10648 & ~n10649;
  assign n10651 = ~n10645 & ~n10650;
  assign n10652 = n10644 & n10651;
  assign n10653 = ~n10644 & ~n10651;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = pi331 & n4596;
  assign n10656 = ~n9288 & n9311;
  assign n10657 = n9288 & ~n9311;
  assign n10658 = ~n4596 & ~n10657;
  assign n10659 = ~n10656 & ~n10658;
  assign n10660 = n5257 & ~n10659;
  assign n10661 = ~n5257 & ~n10656;
  assign n10662 = n4596 & n10661;
  assign n10663 = ~n10660 & ~n10662;
  assign n10664 = pi330 & ~n10663;
  assign n10665 = pi330 & n5257;
  assign n10666 = n9288 & ~n10665;
  assign n10667 = ~n9311 & n10666;
  assign n10668 = ~n10664 & ~n10667;
  assign n10669 = ~n10655 & n10668;
  assign n10670 = n10655 & ~n10668;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = pi332 & n2887;
  assign n10673 = ~n9319 & ~n9335;
  assign n10674 = ~n9342 & n10673;
  assign n10675 = ~n9333 & ~n9335;
  assign n10676 = ~n9308 & n10675;
  assign n10677 = ~n9334 & ~n10676;
  assign n10678 = ~n10674 & n10677;
  assign n10679 = n10672 & ~n10678;
  assign n10680 = ~n10672 & n10678;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = ~n10671 & ~n10681;
  assign n10683 = n10655 & n10668;
  assign n10684 = ~n10655 & ~n10668;
  assign n10685 = ~n10683 & ~n10684;
  assign n10686 = ~n10672 & ~n10678;
  assign n10687 = n10672 & n10678;
  assign n10688 = ~n10686 & ~n10687;
  assign n10689 = ~n10685 & ~n10688;
  assign n10690 = ~n10682 & ~n10689;
  assign n10691 = ~n10654 & ~n10690;
  assign n10692 = n10644 & ~n10651;
  assign n10693 = ~n10644 & n10651;
  assign n10694 = ~n10692 & ~n10693;
  assign n10695 = ~n10681 & ~n10685;
  assign n10696 = ~n10671 & ~n10688;
  assign n10697 = ~n10695 & ~n10696;
  assign n10698 = ~n10694 & ~n10697;
  assign n10699 = ~n10691 & ~n10698;
  assign n10700 = ~n10154 & n10699;
  assign n10701 = n10154 & ~n10699;
  assign n10702 = ~n10700 & ~n10701;
  assign n10703 = pi335 & n1729;
  assign n10704 = pi334 & n2091;
  assign n10705 = n1729 & ~n8798;
  assign n10706 = pi333 & n10705;
  assign n10707 = ~n8166 & ~n8789;
  assign n10708 = ~n9353 & ~n10707;
  assign n10709 = ~n10706 & n10708;
  assign n10710 = ~n9358 & ~n10709;
  assign n10711 = ~n9354 & n10710;
  assign n10712 = ~n10704 & ~n10711;
  assign n10713 = n8810 & n10712;
  assign n10714 = n9354 & ~n10710;
  assign n10715 = n10704 & ~n10714;
  assign n10716 = ~n8810 & n10715;
  assign n10717 = ~n10713 & ~n10716;
  assign n10718 = ~n10133 & ~n10717;
  assign n10719 = n8810 & n10715;
  assign n10720 = ~n8810 & n10712;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = ~n10142 & ~n10721;
  assign n10723 = ~n10704 & ~n10710;
  assign n10724 = n9354 & n10723;
  assign n10725 = n10704 & n10710;
  assign n10726 = ~n9354 & n10725;
  assign n10727 = ~n10724 & ~n10726;
  assign n10728 = ~n10722 & n10727;
  assign n10729 = ~n10718 & n10728;
  assign n10730 = n10703 & ~n10729;
  assign n10731 = ~n10703 & n10729;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 = ~n10702 & ~n10732;
  assign n10734 = n10154 & n10699;
  assign n10735 = ~n10154 & ~n10699;
  assign n10736 = ~n10734 & ~n10735;
  assign n10737 = ~n10703 & ~n10729;
  assign n10738 = n10703 & n10729;
  assign n10739 = ~n10737 & ~n10738;
  assign n10740 = ~n10736 & ~n10739;
  assign n10741 = ~n10733 & ~n10740;
  assign n10742 = ~n10153 & ~n10741;
  assign n10743 = ~n10130 & n10150;
  assign n10744 = n10130 & ~n10150;
  assign n10745 = ~n10743 & ~n10744;
  assign n10746 = ~n10732 & ~n10736;
  assign n10747 = ~n10702 & ~n10739;
  assign n10748 = ~n10746 & ~n10747;
  assign n10749 = ~n10745 & ~n10748;
  assign n10750 = ~n10742 & ~n10749;
  assign n10751 = ~n1154 & n8732;
  assign n10752 = pi337 & n10751;
  assign n10753 = ~n8732 & ~n9414;
  assign n10754 = ~n9395 & ~n9410;
  assign n10755 = ~n9404 & n10754;
  assign n10756 = n9395 & ~n9411;
  assign n10757 = ~n10755 & ~n10756;
  assign n10758 = ~n10753 & ~n10757;
  assign n10759 = ~n10752 & ~n10758;
  assign n10760 = n10750 & ~n10759;
  assign n10761 = ~n10750 & n10759;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = n9395 & ~n9410;
  assign n10764 = ~n9404 & ~n10763;
  assign n10765 = n1442 & n10764;
  assign n10766 = pi336 & n10765;
  assign n10767 = pi336 & n1442;
  assign n10768 = ~n10764 & ~n10767;
  assign n10769 = ~n10766 & ~n10768;
  assign n10770 = pi337 & ~n1256;
  assign n10771 = n10769 & ~n10770;
  assign n10772 = ~n1256 & ~n10769;
  assign n10773 = pi337 & n10772;
  assign n10774 = ~n10771 & ~n10773;
  assign n10775 = ~n10762 & ~n10774;
  assign n10776 = ~n10750 & ~n10759;
  assign n10777 = n10750 & n10759;
  assign n10778 = ~n10776 & ~n10777;
  assign n10779 = ~n10769 & ~n10770;
  assign n10780 = ~n1256 & n10769;
  assign n10781 = pi337 & n10780;
  assign n10782 = ~n10779 & ~n10781;
  assign n10783 = ~n10778 & ~n10782;
  assign n10784 = ~n10775 & ~n10783;
  assign n10785 = n10126 & ~n10784;
  assign n10786 = ~n10126 & n10784;
  assign n10787 = ~n10785 & ~n10786;
  assign n10788 = pi258 & ~n10787;
  assign n10789 = pi128 & n10788;
  assign n10790 = pi339 & n10789;
  assign n10791 = pi339 & n1156;
  assign n10792 = ~n10785 & ~n10791;
  assign n10793 = ~n10786 & n10792;
  assign n10794 = ~n10790 & ~n10793;
  assign n10795 = ~pi274 & ~n8782;
  assign n10796 = pi274 & n8782;
  assign n10797 = n9426 & ~n9436;
  assign n10798 = pi338 & ~n9426;
  assign n10799 = n1156 & n10798;
  assign n10800 = ~n10797 & ~n10799;
  assign n10801 = ~n10796 & ~n10800;
  assign n10802 = ~n10795 & ~n10801;
  assign n10803 = ~pi275 & ~n10802;
  assign n10804 = pi275 & n10802;
  assign n10805 = ~n10803 & ~n10804;
  assign n10806 = ~n10794 & ~n10805;
  assign n10807 = pi275 & ~n10802;
  assign n10808 = ~pi275 & n10802;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = ~n10793 & ~n10809;
  assign n10811 = ~n10790 & n10810;
  assign n10812 = ~n10806 & ~n10811;
  assign n10813 = ~n9441 & ~n9762;
  assign n10814 = ~n9440 & n9762;
  assign n10815 = ~n9439 & n10814;
  assign n10816 = ~n9758 & ~n10815;
  assign n10817 = ~n10813 & ~n10816;
  assign n10818 = n10812 & ~n10817;
  assign n10819 = ~n10812 & n10817;
  assign n10820 = ~n10818 & ~n10819;
  assign n10821 = ~n10120 & ~n10820;
  assign n10822 = n10812 & n10817;
  assign n10823 = ~n10812 & ~n10817;
  assign n10824 = ~n10822 & ~n10823;
  assign n10825 = n10120 & ~n10824;
  assign n10826 = ~n10821 & ~n10825;
  assign n10827 = ~n831 & ~n10826;
  assign n10828 = ~n9772 & ~n10827;
  assign n10829 = pi161 & ~n10828;
  assign n10830 = pi081 & ~pi161;
  assign n10831 = ~n10829 & ~n10830;
  assign po210 = ~pi160 & ~n10831;
  assign n10833 = pi276 & n831;
  assign n10834 = pi304 & ~n1568;
  assign n10835 = n10075 & n10094;
  assign n10836 = ~n10075 & ~n10094;
  assign n10837 = ~n10835 & ~n10836;
  assign n10838 = n10077 & ~n10095;
  assign n10839 = ~n10837 & ~n10838;
  assign n10840 = n1515 & ~n10077;
  assign n10841 = pi306 & n10840;
  assign n10842 = ~n10839 & ~n10841;
  assign n10843 = ~n10075 & ~n10091;
  assign n10844 = ~n9461 & n9733;
  assign n10845 = ~n9456 & ~n10844;
  assign n10846 = ~n10086 & ~n10845;
  assign n10847 = n10075 & n10091;
  assign n10848 = ~n10846 & ~n10847;
  assign n10849 = ~n10843 & ~n10848;
  assign n10850 = pi309 & n2183;
  assign n10851 = ~n10054 & ~n10061;
  assign n10852 = ~n10062 & ~n10851;
  assign n10853 = ~n10850 & ~n10852;
  assign n10854 = ~n10057 & ~n10062;
  assign n10855 = ~n10061 & ~n10854;
  assign n10856 = n10850 & ~n10855;
  assign n10857 = ~n10853 & ~n10856;
  assign n10858 = n9688 & n10014;
  assign n10859 = n9683 & n10858;
  assign n10860 = ~n9690 & ~n10030;
  assign n10861 = n1840 & n10860;
  assign n10862 = ~n9689 & ~n10014;
  assign n10863 = n2183 & ~n10862;
  assign n10864 = ~n10861 & ~n10863;
  assign n10865 = pi310 & ~n10864;
  assign n10866 = ~n10859 & ~n10865;
  assign n10867 = ~n9997 & ~n9998;
  assign n10868 = n9997 & n9998;
  assign n10869 = ~n10003 & ~n10868;
  assign n10870 = ~n10867 & ~n10869;
  assign n10871 = pi313 & n4086;
  assign n10872 = ~n9976 & ~n9983;
  assign n10873 = ~n9984 & ~n10872;
  assign n10874 = ~n10871 & ~n10873;
  assign n10875 = ~n9979 & ~n9984;
  assign n10876 = ~n9983 & ~n10875;
  assign n10877 = n10871 & ~n10876;
  assign n10878 = ~n10874 & ~n10877;
  assign n10879 = ~n9943 & ~n9944;
  assign n10880 = n9943 & n9944;
  assign n10881 = ~n9617 & ~n10880;
  assign n10882 = ~n9611 & n10881;
  assign n10883 = ~n10879 & ~n10882;
  assign n10884 = ~n9867 & n9872;
  assign n10885 = ~n9866 & ~n9872;
  assign n10886 = ~n9864 & n10885;
  assign n10887 = ~n10884 & ~n10886;
  assign n10888 = ~n9896 & ~n10887;
  assign n10889 = pi142 & pi144;
  assign n10890 = pi143 & n9788;
  assign n10891 = ~n10889 & ~n10890;
  assign n10892 = pi141 & ~n10891;
  assign n10893 = pi143 & pi145;
  assign n10894 = ~n9506 & ~n10893;
  assign n10895 = pi142 & ~n10894;
  assign n10896 = ~pi143 & ~pi145;
  assign n10897 = pi144 & ~n10896;
  assign n10898 = ~n10895 & ~n10897;
  assign n10899 = ~n10892 & n10898;
  assign n10900 = pi146 & n10899;
  assign n10901 = ~pi146 & ~n10899;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = pi145 & ~n10902;
  assign n10904 = pi146 & ~n10899;
  assign n10905 = ~pi146 & n10899;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = ~pi145 & ~n10906;
  assign n10908 = ~n10903 & ~n10907;
  assign n10909 = pi321 & n10908;
  assign n10910 = ~n9816 & n9822;
  assign n10911 = n9517 & ~n10910;
  assign n10912 = pi320 & n10911;
  assign n10913 = n9815 & ~n9822;
  assign n10914 = pi321 & n10913;
  assign n10915 = ~n10912 & ~n10914;
  assign n10916 = pi320 & n9815;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = n9815 & n10915;
  assign n10919 = pi320 & n10918;
  assign n10920 = ~n10917 & ~n10919;
  assign n10921 = ~n10909 & ~n10920;
  assign n10922 = n10915 & ~n10916;
  assign n10923 = n9815 & ~n10915;
  assign n10924 = pi320 & n10923;
  assign n10925 = ~n10922 & ~n10924;
  assign n10926 = n10908 & ~n10925;
  assign n10927 = pi321 & n10926;
  assign n10928 = ~n10921 & ~n10927;
  assign n10929 = pi319 & n9517;
  assign n10930 = n10928 & n10929;
  assign n10931 = ~n10928 & ~n10929;
  assign n10932 = ~n10930 & ~n10931;
  assign n10933 = ~n9835 & ~n9843;
  assign n10934 = n9835 & n9843;
  assign n10935 = n7874 & ~n10934;
  assign n10936 = pi319 & n10935;
  assign n10937 = ~n10933 & ~n10936;
  assign n10938 = n10932 & n10937;
  assign n10939 = ~n10932 & ~n10937;
  assign n10940 = ~n10938 & ~n10939;
  assign n10941 = n7874 & ~n10940;
  assign n10942 = pi318 & n10941;
  assign n10943 = pi318 & n7874;
  assign n10944 = ~n10932 & n10937;
  assign n10945 = n10932 & ~n10937;
  assign n10946 = ~n10944 & ~n10945;
  assign n10947 = ~n10943 & ~n10946;
  assign n10948 = ~n10942 & ~n10947;
  assign n10949 = n9849 & ~n9859;
  assign n10950 = ~n9849 & n9859;
  assign n10951 = ~n9852 & ~n10950;
  assign n10952 = ~n10949 & ~n10951;
  assign n10953 = n10948 & ~n10952;
  assign n10954 = ~n10948 & n10952;
  assign n10955 = ~n10953 & ~n10954;
  assign n10956 = pi317 & n7044;
  assign n10957 = ~n9866 & n9872;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = ~n9864 & n10958;
  assign n10960 = ~n9864 & ~n10957;
  assign n10961 = n10956 & ~n10960;
  assign n10962 = ~n10959 & ~n10961;
  assign n10963 = ~n10955 & ~n10962;
  assign n10964 = n10948 & n10952;
  assign n10965 = ~n10948 & ~n10952;
  assign n10966 = ~n10964 & ~n10965;
  assign n10967 = n10956 & ~n10957;
  assign n10968 = ~n9864 & n10967;
  assign n10969 = ~n10956 & ~n10960;
  assign n10970 = ~n10968 & ~n10969;
  assign n10971 = ~n10966 & ~n10970;
  assign n10972 = ~n10963 & ~n10971;
  assign n10973 = ~pi316 & ~n10972;
  assign n10974 = ~n6777 & ~n10972;
  assign n10975 = n6777 & n10972;
  assign n10976 = pi316 & n10975;
  assign n10977 = ~n10974 & ~n10976;
  assign n10978 = ~n5463 & ~n10977;
  assign n10979 = ~n10973 & ~n10978;
  assign n10980 = ~n10888 & ~n10979;
  assign n10981 = n9896 & n10972;
  assign n10982 = n10887 & n10981;
  assign n10983 = ~n9896 & ~n10972;
  assign n10984 = ~n10887 & n10983;
  assign n10985 = ~n10982 & ~n10984;
  assign n10986 = pi316 & ~n10985;
  assign n10987 = n9896 & ~n10887;
  assign n10988 = ~n9896 & n10887;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = ~n10972 & ~n10989;
  assign n10991 = n5463 & n10990;
  assign n10992 = ~n10986 & ~n10991;
  assign n10993 = n6777 & ~n10992;
  assign n10994 = n9896 & ~n10972;
  assign n10995 = n10887 & n10994;
  assign n10996 = n9896 & n10887;
  assign n10997 = n5463 & ~n10996;
  assign n10998 = pi316 & n10997;
  assign n10999 = ~n10888 & ~n10998;
  assign n11000 = n10972 & ~n10999;
  assign n11001 = ~n10995 & ~n11000;
  assign n11002 = ~n6777 & ~n11001;
  assign n11003 = ~pi316 & ~n10887;
  assign n11004 = ~n9896 & n10972;
  assign n11005 = n11003 & n11004;
  assign n11006 = ~n11002 & ~n11005;
  assign n11007 = ~n10993 & n11006;
  assign n11008 = ~n10980 & n11007;
  assign n11009 = n9902 & ~n9905;
  assign n11010 = ~n9606 & ~n9937;
  assign n11011 = n9606 & n9937;
  assign n11012 = n9584 & ~n11011;
  assign n11013 = ~n11010 & ~n11012;
  assign n11014 = ~n9902 & n9905;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = ~n11009 & ~n11015;
  assign n11017 = n11008 & n11016;
  assign n11018 = ~n11008 & ~n11016;
  assign n11019 = ~n11017 & ~n11018;
  assign n11020 = n5463 & ~n11019;
  assign n11021 = pi315 & n11020;
  assign n11022 = pi315 & n5463;
  assign n11023 = ~n11008 & n11016;
  assign n11024 = n11008 & ~n11016;
  assign n11025 = ~n11023 & ~n11024;
  assign n11026 = ~n11022 & ~n11025;
  assign n11027 = ~n11021 & ~n11026;
  assign n11028 = n4772 & ~n11027;
  assign n11029 = pi314 & n11028;
  assign n11030 = pi314 & n4772;
  assign n11031 = ~n11026 & ~n11030;
  assign n11032 = ~n11021 & n11031;
  assign n11033 = ~n11029 & ~n11032;
  assign n11034 = ~n10883 & ~n11033;
  assign n11035 = n10883 & ~n11032;
  assign n11036 = ~n11029 & n11035;
  assign n11037 = ~n11034 & ~n11036;
  assign n11038 = n10878 & ~n11037;
  assign n11039 = ~n10878 & n11037;
  assign n11040 = ~n11038 & ~n11039;
  assign n11041 = pi312 & n3552;
  assign n11042 = ~n3012 & ~n3552;
  assign n11043 = pi313 & ~n11042;
  assign n11044 = n9959 & ~n11043;
  assign n11045 = ~n3012 & n3552;
  assign n11046 = pi313 & ~n9959;
  assign n11047 = n11045 & n11046;
  assign n11048 = ~n11044 & ~n11047;
  assign n11049 = ~n9973 & ~n11048;
  assign n11050 = ~n3552 & n9959;
  assign n11051 = ~n9961 & ~n11050;
  assign n11052 = ~n9619 & ~n11051;
  assign n11053 = n9972 & n11052;
  assign n11054 = n3012 & ~n3552;
  assign n11055 = ~n9959 & n11054;
  assign n11056 = ~n3012 & ~n9619;
  assign n11057 = n3552 & ~n11056;
  assign n11058 = n9959 & n11057;
  assign n11059 = ~n11055 & ~n11058;
  assign n11060 = pi313 & ~n11059;
  assign n11061 = n9619 & n9983;
  assign n11062 = ~n11060 & ~n11061;
  assign n11063 = ~n9972 & ~n11062;
  assign n11064 = ~n3552 & ~n9959;
  assign n11065 = n3552 & n9959;
  assign n11066 = ~n11064 & ~n11065;
  assign n11067 = n3012 & ~n11066;
  assign n11068 = pi313 & n11067;
  assign n11069 = n9619 & n11068;
  assign n11070 = ~n11063 & ~n11069;
  assign n11071 = ~n11053 & n11070;
  assign n11072 = ~n11049 & n11071;
  assign n11073 = ~n9994 & ~n11072;
  assign n11074 = n9994 & n11072;
  assign n11075 = n9963 & ~n11074;
  assign n11076 = ~n11073 & ~n11075;
  assign n11077 = n11041 & ~n11076;
  assign n11078 = ~n9963 & ~n11073;
  assign n11079 = ~n11074 & ~n11078;
  assign n11080 = ~n11041 & ~n11079;
  assign n11081 = ~n11077 & ~n11080;
  assign n11082 = ~n11040 & ~n11081;
  assign n11083 = n10878 & n11037;
  assign n11084 = ~n10878 & ~n11037;
  assign n11085 = ~n11083 & ~n11084;
  assign n11086 = ~n11041 & ~n11076;
  assign n11087 = n11041 & ~n11079;
  assign n11088 = ~n11086 & ~n11087;
  assign n11089 = ~n11085 & ~n11088;
  assign n11090 = ~n11082 & ~n11089;
  assign n11091 = n10870 & n11090;
  assign n11092 = ~n10870 & ~n11090;
  assign n11093 = ~n11091 & ~n11092;
  assign n11094 = n3012 & ~n11093;
  assign n11095 = pi311 & n11094;
  assign n11096 = pi311 & n3012;
  assign n11097 = ~n10870 & n11090;
  assign n11098 = n10870 & ~n11090;
  assign n11099 = ~n11097 & ~n11098;
  assign n11100 = ~n11096 & ~n11099;
  assign n11101 = ~n11095 & ~n11100;
  assign n11102 = n2574 & ~n11101;
  assign n11103 = pi310 & n11102;
  assign n11104 = pi310 & n2574;
  assign n11105 = ~n11100 & ~n11104;
  assign n11106 = ~n11095 & n11105;
  assign n11107 = ~n11103 & ~n11106;
  assign n11108 = ~n10866 & ~n11107;
  assign n11109 = n10866 & ~n11106;
  assign n11110 = ~n11103 & n11109;
  assign n11111 = ~n11108 & ~n11110;
  assign n11112 = n10857 & n11111;
  assign n11113 = ~n10857 & ~n11111;
  assign n11114 = ~n11112 & ~n11113;
  assign n11115 = pi308 & n1840;
  assign n11116 = pi309 & ~n6883;
  assign n11117 = n10046 & ~n11116;
  assign n11118 = pi309 & ~n10046;
  assign n11119 = n6886 & n11118;
  assign n11120 = ~n11117 & ~n11119;
  assign n11121 = ~n10051 & ~n11120;
  assign n11122 = ~n1840 & n10046;
  assign n11123 = ~n10062 & ~n11122;
  assign n11124 = n9699 & ~n11123;
  assign n11125 = n9466 & n11124;
  assign n11126 = n6897 & ~n10046;
  assign n11127 = ~n1533 & n9699;
  assign n11128 = n1840 & ~n11127;
  assign n11129 = n10046 & n11128;
  assign n11130 = ~n11126 & ~n11129;
  assign n11131 = pi309 & ~n11130;
  assign n11132 = ~n9699 & n10047;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~n9466 & ~n11133;
  assign n11135 = ~n1840 & ~n10046;
  assign n11136 = n1840 & n10046;
  assign n11137 = ~n11135 & ~n11136;
  assign n11138 = n1533 & ~n11137;
  assign n11139 = pi309 & n11138;
  assign n11140 = ~n9699 & n11139;
  assign n11141 = ~n11134 & ~n11140;
  assign n11142 = ~n11125 & n11141;
  assign n11143 = ~n11121 & n11142;
  assign n11144 = n10072 & n11143;
  assign n11145 = ~n10072 & ~n11143;
  assign n11146 = n10050 & ~n11145;
  assign n11147 = ~n11144 & ~n11146;
  assign n11148 = n11115 & ~n11147;
  assign n11149 = ~n10050 & ~n11144;
  assign n11150 = ~n11145 & ~n11149;
  assign n11151 = ~n11115 & ~n11150;
  assign n11152 = ~n11148 & ~n11151;
  assign n11153 = ~n11114 & ~n11152;
  assign n11154 = n10857 & ~n11111;
  assign n11155 = ~n10857 & n11111;
  assign n11156 = ~n11154 & ~n11155;
  assign n11157 = ~n11115 & ~n11147;
  assign n11158 = n11115 & ~n11150;
  assign n11159 = ~n11157 & ~n11158;
  assign n11160 = ~n11156 & ~n11159;
  assign n11161 = ~n11153 & ~n11160;
  assign n11162 = n10849 & n11161;
  assign n11163 = ~n10849 & ~n11161;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = n1533 & ~n11164;
  assign n11166 = pi307 & n11165;
  assign n11167 = pi307 & n1533;
  assign n11168 = ~n10849 & n11161;
  assign n11169 = n10849 & ~n11161;
  assign n11170 = ~n11168 & ~n11169;
  assign n11171 = ~n11167 & ~n11170;
  assign n11172 = ~n11166 & ~n11171;
  assign n11173 = n1553 & ~n11172;
  assign n11174 = pi306 & n11173;
  assign n11175 = pi306 & n1553;
  assign n11176 = ~n11171 & ~n11175;
  assign n11177 = ~n11166 & n11176;
  assign n11178 = ~n11174 & ~n11177;
  assign n11179 = n10842 & ~n11178;
  assign n11180 = ~n10842 & ~n11177;
  assign n11181 = ~n11174 & n11180;
  assign n11182 = ~n11179 & ~n11181;
  assign n11183 = n10834 & ~n11182;
  assign n11184 = ~n10834 & n11182;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = pi304 & ~n10118;
  assign n11187 = pi128 & n11186;
  assign n11188 = ~pi130 & n10109;
  assign n11189 = n1335 & n11188;
  assign n11190 = ~pi129 & n9777;
  assign n11191 = pi129 & ~n9777;
  assign n11192 = n10109 & ~n11191;
  assign n11193 = pi128 & n11192;
  assign n11194 = ~n11190 & ~n11193;
  assign n11195 = pi130 & ~n11194;
  assign n11196 = ~n11189 & ~n11195;
  assign n11197 = pi305 & ~n11196;
  assign n11198 = n9777 & n10109;
  assign n11199 = ~pi130 & ~n11198;
  assign n11200 = pi128 & n11199;
  assign n11201 = ~pi128 & pi130;
  assign n11202 = pi305 & ~n11201;
  assign n11203 = ~n10109 & ~n11202;
  assign n11204 = ~n11200 & ~n11203;
  assign n11205 = pi129 & ~n11204;
  assign n11206 = pi128 & n10109;
  assign n11207 = ~pi130 & ~n11206;
  assign n11208 = ~pi129 & n11207;
  assign n11209 = pi305 & ~n11208;
  assign n11210 = ~n9777 & ~n11209;
  assign n11211 = ~n11205 & ~n11210;
  assign n11212 = ~n11197 & n11211;
  assign n11213 = n11187 & ~n11212;
  assign n11214 = ~n11187 & n11212;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = ~n11185 & ~n11215;
  assign n11217 = n10834 & n11182;
  assign n11218 = ~n10834 & ~n11182;
  assign n11219 = ~n11217 & ~n11218;
  assign n11220 = n11187 & n11212;
  assign n11221 = ~n11187 & ~n11212;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = ~n11219 & ~n11222;
  assign n11224 = ~n11216 & ~n11223;
  assign n11225 = n10794 & ~n10802;
  assign n11226 = ~n10794 & n10802;
  assign n11227 = ~pi275 & ~n11226;
  assign n11228 = ~n11225 & ~n11227;
  assign n11229 = ~n1154 & n10784;
  assign n11230 = n1154 & ~n10784;
  assign n11231 = n9426 & ~n11230;
  assign n11232 = n1156 & n11231;
  assign n11233 = ~n11229 & ~n11232;
  assign n11234 = n1256 & ~n11233;
  assign n11235 = ~n10121 & ~n11229;
  assign n11236 = ~n11230 & ~n11235;
  assign n11237 = ~n1256 & ~n11236;
  assign n11238 = ~n11234 & ~n11237;
  assign n11239 = pi338 & ~n11238;
  assign n11240 = ~n10130 & n10699;
  assign n11241 = n10130 & ~n10699;
  assign n11242 = ~n11240 & ~n11241;
  assign n11243 = n10150 & n10703;
  assign n11244 = n10154 & ~n10729;
  assign n11245 = ~n10154 & n10729;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = ~n11243 & ~n11246;
  assign n11248 = ~n11242 & n11247;
  assign n11249 = ~n10130 & ~n10699;
  assign n11250 = n10130 & n10699;
  assign n11251 = ~n11249 & ~n11250;
  assign n11252 = ~n10154 & ~n10729;
  assign n11253 = n10154 & n10729;
  assign n11254 = ~n11252 & ~n11253;
  assign n11255 = ~n11243 & ~n11254;
  assign n11256 = ~n11251 & n11255;
  assign n11257 = ~n10150 & ~n10703;
  assign n11258 = ~n11256 & ~n11257;
  assign n11259 = ~n11248 & n11258;
  assign n11260 = n10750 & n10769;
  assign n11261 = ~n10750 & ~n10769;
  assign n11262 = ~n11260 & ~n11261;
  assign n11263 = n10759 & ~n10770;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = ~n1256 & ~n10759;
  assign n11266 = pi337 & n11265;
  assign n11267 = ~n11264 & ~n11266;
  assign n11268 = n11259 & n11267;
  assign n11269 = ~n11259 & ~n11267;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 = pi335 & n2091;
  assign n11272 = ~n10171 & ~n10175;
  assign n11273 = n10171 & n10175;
  assign n11274 = ~n10159 & n10623;
  assign n11275 = n10159 & ~n10623;
  assign n11276 = ~n11274 & ~n11275;
  assign n11277 = n5732 & ~n11276;
  assign n11278 = pi328 & n11277;
  assign n11279 = ~n10159 & ~n10623;
  assign n11280 = n10159 & n10623;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = ~n10629 & ~n11281;
  assign n11283 = ~n11278 & ~n11282;
  assign n11284 = ~n11273 & ~n11283;
  assign n11285 = ~n11272 & ~n11284;
  assign n11286 = ~n10651 & n10655;
  assign n11287 = n10651 & ~n10655;
  assign n11288 = n4596 & ~n10656;
  assign n11289 = ~n10657 & ~n11288;
  assign n11290 = n5257 & ~n11289;
  assign n11291 = pi330 & n11290;
  assign n11292 = ~n5257 & ~n11288;
  assign n11293 = pi330 & ~n11292;
  assign n11294 = ~n10657 & ~n11293;
  assign n11295 = ~n11291 & ~n11294;
  assign n11296 = n10644 & ~n11295;
  assign n11297 = ~n10644 & n11295;
  assign n11298 = ~n11296 & ~n11297;
  assign n11299 = ~n11287 & ~n11298;
  assign n11300 = ~n11286 & ~n11299;
  assign n11301 = n11285 & n11300;
  assign n11302 = ~n11285 & ~n11300;
  assign n11303 = ~n11301 & ~n11302;
  assign n11304 = n10644 & ~n11294;
  assign n11305 = ~n11291 & ~n11304;
  assign n11306 = n5714 & n11305;
  assign n11307 = pi330 & n11306;
  assign n11308 = pi330 & n5714;
  assign n11309 = ~n11305 & ~n11308;
  assign n11310 = ~n11307 & ~n11309;
  assign n11311 = ~n10179 & ~n10597;
  assign n11312 = n10179 & n10597;
  assign n11313 = ~n11311 & ~n11312;
  assign n11314 = n10199 & n10601;
  assign n11315 = ~n10582 & n10602;
  assign n11316 = n10582 & ~n10602;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = ~n11314 & ~n11317;
  assign n11319 = ~n11313 & n11318;
  assign n11320 = ~n10179 & n10597;
  assign n11321 = n10179 & ~n10597;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = n10582 & n10602;
  assign n11324 = ~n10582 & ~n10602;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = ~n11314 & ~n11325;
  assign n11327 = ~n11322 & n11326;
  assign n11328 = ~n10199 & ~n10601;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~n11319 & n11329;
  assign n11331 = n5732 & ~n11280;
  assign n11332 = pi328 & n11331;
  assign n11333 = ~n11279 & ~n11332;
  assign n11334 = n11330 & ~n11333;
  assign n11335 = ~n11330 & n11333;
  assign n11336 = ~n11334 & ~n11335;
  assign n11337 = pi327 & n6556;
  assign n11338 = n10558 & ~n10597;
  assign n11339 = ~n10204 & ~n10557;
  assign n11340 = n10204 & ~n10556;
  assign n11341 = ~n10550 & n11340;
  assign n11342 = ~n11339 & ~n11341;
  assign n11343 = ~n10562 & ~n11342;
  assign n11344 = n10204 & ~n10557;
  assign n11345 = ~n10204 & ~n10556;
  assign n11346 = ~n10550 & n11345;
  assign n11347 = ~n11344 & ~n11346;
  assign n11348 = n10561 & ~n11347;
  assign n11349 = pi324 & n11348;
  assign n11350 = ~n11343 & ~n11349;
  assign n11351 = n10212 & ~n11350;
  assign n11352 = ~n10212 & n11350;
  assign n11353 = ~n11351 & ~n11352;
  assign n11354 = ~n10558 & n10597;
  assign n11355 = ~n11353 & ~n11354;
  assign n11356 = ~n11338 & ~n11355;
  assign n11357 = ~n10179 & n10602;
  assign n11358 = n10179 & ~n10602;
  assign n11359 = ~n10609 & ~n11358;
  assign n11360 = ~n11357 & ~n11359;
  assign n11361 = n11356 & ~n11360;
  assign n11362 = ~n11356 & n11360;
  assign n11363 = ~n11361 & ~n11362;
  assign n11364 = ~n8513 & ~n10224;
  assign n11365 = n8513 & ~n10220;
  assign n11366 = ~n11364 & ~n11365;
  assign n11367 = pi324 & n11366;
  assign n11368 = ~n10204 & ~n10550;
  assign n11369 = ~n10556 & ~n11368;
  assign n11370 = ~n11367 & ~n11369;
  assign n11371 = n11367 & n11369;
  assign n11372 = ~n11370 & ~n11371;
  assign n11373 = ~n10228 & n10534;
  assign n11374 = n10228 & ~n10534;
  assign n11375 = ~n11373 & ~n11374;
  assign n11376 = n10536 & ~n11375;
  assign n11377 = ~n10536 & n11375;
  assign n11378 = ~n11376 & ~n11377;
  assign n11379 = ~n9167 & ~n11378;
  assign n11380 = ~n10536 & ~n11375;
  assign n11381 = n10536 & n11375;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = n9167 & ~n11382;
  assign n11384 = ~n11379 & ~n11383;
  assign n11385 = pi323 & n11384;
  assign n11386 = n10241 & n10245;
  assign n11387 = ~n10241 & ~n10245;
  assign n11388 = pi262 & ~n10490;
  assign n11389 = pi141 & n11388;
  assign n11390 = ~n10481 & ~n10483;
  assign n11391 = ~n11389 & ~n11390;
  assign n11392 = pi261 & ~n11391;
  assign n11393 = pi142 & n11392;
  assign n11394 = ~n10482 & ~n11390;
  assign n11395 = ~n11389 & n11394;
  assign n11396 = ~n11393 & ~n11395;
  assign n11397 = n10235 & n11396;
  assign n11398 = ~n10235 & ~n11396;
  assign n11399 = ~n11397 & ~n11398;
  assign n11400 = ~n11387 & ~n11399;
  assign n11401 = ~n11386 & ~n11400;
  assign n11402 = ~n10500 & ~n10515;
  assign n11403 = ~n10529 & n11402;
  assign n11404 = ~n10515 & ~n10520;
  assign n11405 = ~n10244 & n11404;
  assign n11406 = ~n10514 & ~n11405;
  assign n11407 = ~n11403 & n11406;
  assign n11408 = ~n11401 & ~n11407;
  assign n11409 = n11401 & n11407;
  assign n11410 = ~n11408 & ~n11409;
  assign n11411 = pi143 & pi261;
  assign n11412 = pi139 & pi265;
  assign n11413 = pi136 & pi268;
  assign n11414 = pi133 & pi271;
  assign n11415 = pi130 & pi274;
  assign n11416 = pi128 & pi276;
  assign n11417 = pi275 & ~n11416;
  assign n11418 = pi129 & n11417;
  assign n11419 = pi129 & pi275;
  assign n11420 = pi276 & ~n11419;
  assign n11421 = pi128 & n11420;
  assign n11422 = ~n11418 & ~n11421;
  assign n11423 = ~n10253 & ~n10256;
  assign n11424 = n10253 & n10256;
  assign n11425 = ~n8246 & ~n8249;
  assign n11426 = n8246 & n8249;
  assign n11427 = n7371 & ~n8906;
  assign n11428 = ~n8907 & ~n11427;
  assign n11429 = ~n11426 & ~n11428;
  assign n11430 = ~n11425 & ~n11429;
  assign n11431 = ~n8895 & ~n11430;
  assign n11432 = ~n8893 & ~n11431;
  assign n11433 = ~n11424 & ~n11432;
  assign n11434 = ~n11423 & ~n11433;
  assign n11435 = ~n11422 & ~n11434;
  assign n11436 = ~n11423 & ~n11431;
  assign n11437 = ~n8893 & n11436;
  assign n11438 = ~n11424 & ~n11437;
  assign n11439 = n11422 & ~n11438;
  assign n11440 = ~n11435 & ~n11439;
  assign n11441 = n11415 & ~n11440;
  assign n11442 = n11422 & ~n11434;
  assign n11443 = ~n11422 & ~n11438;
  assign n11444 = ~n11442 & ~n11443;
  assign n11445 = ~n11415 & ~n11444;
  assign n11446 = ~n11441 & ~n11445;
  assign n11447 = n10252 & n10270;
  assign n11448 = ~n10252 & ~n10270;
  assign n11449 = ~n10274 & ~n11448;
  assign n11450 = ~n8904 & n11449;
  assign n11451 = ~n11447 & ~n11450;
  assign n11452 = pi131 & pi273;
  assign n11453 = ~n11451 & ~n11452;
  assign n11454 = pi273 & n11451;
  assign n11455 = pi131 & n11454;
  assign n11456 = ~n11453 & ~n11455;
  assign n11457 = ~n11446 & ~n11456;
  assign n11458 = n11451 & ~n11452;
  assign n11459 = pi273 & ~n11451;
  assign n11460 = pi131 & n11459;
  assign n11461 = ~n11458 & ~n11460;
  assign n11462 = ~n11445 & ~n11461;
  assign n11463 = ~n11441 & n11462;
  assign n11464 = ~n11457 & ~n11463;
  assign n11465 = ~n10246 & ~n10279;
  assign n11466 = ~n10285 & ~n11465;
  assign n11467 = pi272 & n10279;
  assign n11468 = pi131 & n11467;
  assign n11469 = ~n11466 & ~n11468;
  assign n11470 = n11464 & n11469;
  assign n11471 = ~n11464 & ~n11469;
  assign n11472 = ~n11470 & ~n11471;
  assign n11473 = pi132 & pi272;
  assign n11474 = n10304 & ~n10309;
  assign n11475 = ~n10310 & ~n11474;
  assign n11476 = n11473 & ~n11475;
  assign n11477 = ~n10304 & ~n10310;
  assign n11478 = ~n10309 & ~n11477;
  assign n11479 = ~n11473 & ~n11478;
  assign n11480 = ~n11476 & ~n11479;
  assign n11481 = ~n11472 & ~n11480;
  assign n11482 = n11464 & ~n11469;
  assign n11483 = ~n11464 & n11469;
  assign n11484 = ~n11482 & ~n11483;
  assign n11485 = ~n11473 & ~n11475;
  assign n11486 = n11473 & ~n11478;
  assign n11487 = ~n11485 & ~n11486;
  assign n11488 = ~n11484 & ~n11487;
  assign n11489 = ~n11481 & ~n11488;
  assign n11490 = ~n11414 & n11489;
  assign n11491 = n11414 & ~n11489;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = pi271 & ~n10311;
  assign n11494 = pi132 & n11493;
  assign n11495 = ~n10302 & ~n10304;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = pi270 & ~n11496;
  assign n11498 = pi133 & n11497;
  assign n11499 = pi134 & pi270;
  assign n11500 = ~n10303 & ~n11495;
  assign n11501 = ~n11494 & n11500;
  assign n11502 = ~n10320 & ~n11501;
  assign n11503 = ~n11499 & ~n11502;
  assign n11504 = ~n11498 & n11503;
  assign n11505 = ~n11498 & ~n11502;
  assign n11506 = n11499 & ~n11505;
  assign n11507 = ~n11504 & ~n11506;
  assign n11508 = ~n11492 & ~n11507;
  assign n11509 = ~n11414 & ~n11489;
  assign n11510 = n11414 & n11489;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = n11499 & ~n11502;
  assign n11513 = ~n11498 & n11512;
  assign n11514 = ~n11499 & ~n11505;
  assign n11515 = ~n11513 & ~n11514;
  assign n11516 = ~n11511 & ~n11515;
  assign n11517 = ~n11508 & ~n11516;
  assign n11518 = n10324 & ~n10349;
  assign n11519 = ~n10324 & n10349;
  assign n11520 = ~n10340 & ~n11519;
  assign n11521 = ~n11518 & ~n11520;
  assign n11522 = n11517 & n11521;
  assign n11523 = ~n11517 & ~n11521;
  assign n11524 = ~n11522 & ~n11523;
  assign n11525 = pi135 & pi269;
  assign n11526 = n10363 & ~n10369;
  assign n11527 = ~n10368 & ~n11526;
  assign n11528 = n11525 & ~n11527;
  assign n11529 = ~n10363 & ~n10368;
  assign n11530 = ~n10369 & ~n11529;
  assign n11531 = ~n11525 & ~n11530;
  assign n11532 = ~n11528 & ~n11531;
  assign n11533 = ~n11524 & ~n11532;
  assign n11534 = n11517 & ~n11521;
  assign n11535 = ~n11517 & n11521;
  assign n11536 = ~n11534 & ~n11535;
  assign n11537 = ~n11525 & ~n11527;
  assign n11538 = n11525 & ~n11530;
  assign n11539 = ~n11537 & ~n11538;
  assign n11540 = ~n11536 & ~n11539;
  assign n11541 = ~n11533 & ~n11540;
  assign n11542 = ~n11413 & n11541;
  assign n11543 = n11413 & ~n11541;
  assign n11544 = ~n11542 & ~n11543;
  assign n11545 = pi268 & ~n10370;
  assign n11546 = pi135 & n11545;
  assign n11547 = ~n10361 & ~n10363;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = pi267 & ~n11548;
  assign n11550 = pi136 & n11549;
  assign n11551 = pi137 & pi267;
  assign n11552 = ~n10362 & ~n11547;
  assign n11553 = ~n11546 & n11552;
  assign n11554 = ~n10379 & ~n11553;
  assign n11555 = ~n11551 & ~n11554;
  assign n11556 = ~n11550 & n11555;
  assign n11557 = ~n11550 & ~n11554;
  assign n11558 = n11551 & ~n11557;
  assign n11559 = ~n11556 & ~n11558;
  assign n11560 = ~n11544 & ~n11559;
  assign n11561 = ~n11413 & ~n11541;
  assign n11562 = n11413 & n11541;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = n11551 & ~n11554;
  assign n11565 = ~n11550 & n11564;
  assign n11566 = ~n11551 & ~n11557;
  assign n11567 = ~n11565 & ~n11566;
  assign n11568 = ~n11563 & ~n11567;
  assign n11569 = ~n11560 & ~n11568;
  assign n11570 = n10383 & ~n10408;
  assign n11571 = ~n10383 & n10408;
  assign n11572 = ~n10399 & ~n11571;
  assign n11573 = ~n11570 & ~n11572;
  assign n11574 = n11569 & ~n11573;
  assign n11575 = ~n11569 & n11573;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = pi138 & pi266;
  assign n11578 = n10422 & ~n10428;
  assign n11579 = ~n10427 & ~n11578;
  assign n11580 = n11577 & ~n11579;
  assign n11581 = ~n10422 & ~n10427;
  assign n11582 = ~n10428 & ~n11581;
  assign n11583 = ~n11577 & ~n11582;
  assign n11584 = ~n11580 & ~n11583;
  assign n11585 = ~n11576 & ~n11584;
  assign n11586 = n11569 & n11573;
  assign n11587 = ~n11569 & ~n11573;
  assign n11588 = ~n11586 & ~n11587;
  assign n11589 = ~n11577 & ~n11579;
  assign n11590 = n11577 & ~n11582;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = ~n11588 & ~n11591;
  assign n11593 = ~n11585 & ~n11592;
  assign n11594 = ~n11412 & ~n11593;
  assign n11595 = n11412 & n11593;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = pi265 & ~n10429;
  assign n11598 = pi138 & n11597;
  assign n11599 = ~n10420 & ~n10422;
  assign n11600 = ~n10421 & ~n11599;
  assign n11601 = ~n11598 & n11600;
  assign n11602 = pi140 & pi264;
  assign n11603 = ~n11598 & ~n11599;
  assign n11604 = pi264 & ~n11603;
  assign n11605 = pi139 & n11604;
  assign n11606 = n10439 & ~n11605;
  assign n11607 = n11602 & ~n11606;
  assign n11608 = ~n11601 & n11607;
  assign n11609 = ~n11601 & ~n11606;
  assign n11610 = ~n11602 & ~n11609;
  assign n11611 = ~n11608 & ~n11610;
  assign n11612 = ~n11596 & ~n11611;
  assign n11613 = ~n11412 & n11593;
  assign n11614 = n11412 & ~n11593;
  assign n11615 = ~n11613 & ~n11614;
  assign n11616 = ~n11602 & ~n11606;
  assign n11617 = ~n11601 & n11616;
  assign n11618 = n11602 & ~n11609;
  assign n11619 = ~n11617 & ~n11618;
  assign n11620 = ~n11615 & ~n11619;
  assign n11621 = ~n11612 & ~n11620;
  assign n11622 = ~n10442 & ~n10443;
  assign n11623 = n10442 & n10443;
  assign n11624 = ~n10462 & ~n11623;
  assign n11625 = ~n11622 & ~n11624;
  assign n11626 = n11621 & ~n11625;
  assign n11627 = ~n11621 & n11625;
  assign n11628 = ~n11626 & ~n11627;
  assign n11629 = pi263 & ~n11628;
  assign n11630 = pi141 & n11629;
  assign n11631 = pi141 & pi263;
  assign n11632 = ~n11621 & ~n11625;
  assign n11633 = n11621 & n11625;
  assign n11634 = ~n11632 & ~n11633;
  assign n11635 = ~n11631 & ~n11634;
  assign n11636 = ~n11630 & ~n11635;
  assign n11637 = n10478 & n10483;
  assign n11638 = ~n10478 & ~n10483;
  assign n11639 = n10473 & ~n11638;
  assign n11640 = ~n11637 & ~n11639;
  assign n11641 = n11636 & n11640;
  assign n11642 = ~n11636 & ~n11640;
  assign n11643 = ~n11641 & ~n11642;
  assign n11644 = pi142 & pi262;
  assign n11645 = n10235 & ~n11393;
  assign n11646 = n11644 & ~n11645;
  assign n11647 = ~n11395 & n11646;
  assign n11648 = ~n11395 & ~n11645;
  assign n11649 = ~n11644 & ~n11648;
  assign n11650 = ~n11647 & ~n11649;
  assign n11651 = ~n11643 & ~n11650;
  assign n11652 = n11636 & ~n11640;
  assign n11653 = ~n11636 & n11640;
  assign n11654 = ~n11652 & ~n11653;
  assign n11655 = ~n11644 & ~n11645;
  assign n11656 = ~n11395 & n11655;
  assign n11657 = n11644 & ~n11648;
  assign n11658 = ~n11656 & ~n11657;
  assign n11659 = ~n11654 & ~n11658;
  assign n11660 = ~n11651 & ~n11659;
  assign n11661 = ~n11411 & n11660;
  assign n11662 = n11411 & ~n11660;
  assign n11663 = ~n11661 & ~n11662;
  assign n11664 = pi260 & ~n11663;
  assign n11665 = pi144 & n11664;
  assign n11666 = pi144 & pi260;
  assign n11667 = n11411 & n11660;
  assign n11668 = ~n11411 & ~n11660;
  assign n11669 = ~n11667 & ~n11668;
  assign n11670 = ~n11666 & ~n11669;
  assign n11671 = ~n11665 & ~n11670;
  assign n11672 = ~n11410 & ~n11671;
  assign n11673 = ~n11401 & n11407;
  assign n11674 = n11401 & ~n11407;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = pi260 & ~n11669;
  assign n11677 = pi144 & n11676;
  assign n11678 = ~n11663 & ~n11666;
  assign n11679 = ~n11677 & ~n11678;
  assign n11680 = ~n11675 & ~n11679;
  assign n11681 = ~n11672 & ~n11680;
  assign n11682 = ~n9167 & ~n10536;
  assign n11683 = n9167 & n10536;
  assign n11684 = ~n11375 & ~n11683;
  assign n11685 = ~n11682 & ~n11684;
  assign n11686 = n11681 & n11685;
  assign n11687 = ~n11681 & ~n11685;
  assign n11688 = ~n11686 & ~n11687;
  assign n11689 = ~n10228 & ~n10534;
  assign n11690 = pi146 & pi258;
  assign n11691 = pi145 & pi259;
  assign n11692 = ~n11690 & ~n11691;
  assign n11693 = n11690 & n11691;
  assign n11694 = ~n11692 & ~n11693;
  assign n11695 = ~n11689 & ~n11694;
  assign n11696 = n11690 & ~n11691;
  assign n11697 = ~n11690 & n11691;
  assign n11698 = ~n11696 & ~n11697;
  assign n11699 = ~n10534 & ~n11698;
  assign n11700 = ~n10228 & n11699;
  assign n11701 = ~n11695 & ~n11700;
  assign n11702 = ~n11688 & ~n11701;
  assign n11703 = n11681 & ~n11685;
  assign n11704 = ~n11681 & n11685;
  assign n11705 = ~n11703 & ~n11704;
  assign n11706 = ~n11689 & ~n11698;
  assign n11707 = ~n10534 & ~n11694;
  assign n11708 = ~n10228 & n11707;
  assign n11709 = ~n11706 & ~n11708;
  assign n11710 = ~n11705 & ~n11709;
  assign n11711 = ~n11702 & ~n11710;
  assign n11712 = pi322 & n11711;
  assign n11713 = ~n11385 & ~n11712;
  assign n11714 = n11384 & n11711;
  assign n11715 = n1445 & n11714;
  assign n11716 = ~n11713 & ~n11715;
  assign n11717 = ~n11372 & ~n11716;
  assign n11718 = ~n11367 & n11369;
  assign n11719 = n11367 & ~n11369;
  assign n11720 = ~n11718 & ~n11719;
  assign n11721 = ~n11385 & n11711;
  assign n11722 = pi322 & n11721;
  assign n11723 = n11384 & ~n11712;
  assign n11724 = pi323 & n11723;
  assign n11725 = ~n11722 & ~n11724;
  assign n11726 = ~n11720 & ~n11725;
  assign n11727 = ~n11717 & ~n11726;
  assign n11728 = ~n10212 & n10562;
  assign n11729 = n10212 & ~n10562;
  assign n11730 = ~n11342 & ~n11729;
  assign n11731 = ~n11728 & ~n11730;
  assign n11732 = n11727 & ~n11731;
  assign n11733 = ~n11727 & n11731;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = pi326 & n9205;
  assign n11736 = pi325 & n10561;
  assign n11737 = n11735 & n11736;
  assign n11738 = ~n11735 & ~n11736;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = ~n11734 & ~n11739;
  assign n11741 = ~n11727 & ~n11731;
  assign n11742 = n11727 & n11731;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = ~n11735 & n11736;
  assign n11745 = n11735 & ~n11736;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = ~n11743 & ~n11746;
  assign n11748 = ~n11740 & ~n11747;
  assign n11749 = ~n11363 & ~n11748;
  assign n11750 = n11356 & n11360;
  assign n11751 = ~n11356 & ~n11360;
  assign n11752 = ~n11750 & ~n11751;
  assign n11753 = ~n11739 & ~n11743;
  assign n11754 = ~n11734 & ~n11746;
  assign n11755 = ~n11753 & ~n11754;
  assign n11756 = ~n11752 & ~n11755;
  assign n11757 = ~n11749 & ~n11756;
  assign n11758 = ~n11337 & n11757;
  assign n11759 = n11337 & ~n11757;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = pi329 & n5732;
  assign n11762 = pi328 & n5973;
  assign n11763 = n11761 & n11762;
  assign n11764 = ~n11761 & ~n11762;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = ~n11760 & ~n11765;
  assign n11767 = n11337 & n11757;
  assign n11768 = ~n11337 & ~n11757;
  assign n11769 = ~n11767 & ~n11768;
  assign n11770 = ~n11761 & n11762;
  assign n11771 = n11761 & ~n11762;
  assign n11772 = ~n11770 & ~n11771;
  assign n11773 = ~n11769 & ~n11772;
  assign n11774 = ~n11766 & ~n11773;
  assign n11775 = ~n11336 & ~n11774;
  assign n11776 = n11330 & n11333;
  assign n11777 = ~n11330 & ~n11333;
  assign n11778 = ~n11776 & ~n11777;
  assign n11779 = ~n11765 & ~n11769;
  assign n11780 = ~n11760 & ~n11772;
  assign n11781 = ~n11779 & ~n11780;
  assign n11782 = ~n11778 & ~n11781;
  assign n11783 = ~n11775 & ~n11782;
  assign n11784 = n11310 & n11783;
  assign n11785 = ~n11310 & ~n11783;
  assign n11786 = ~n11784 & ~n11785;
  assign n11787 = n5257 & ~n11786;
  assign n11788 = pi331 & n11787;
  assign n11789 = pi331 & n5257;
  assign n11790 = ~n11310 & n11783;
  assign n11791 = n11310 & ~n11783;
  assign n11792 = ~n11790 & ~n11791;
  assign n11793 = ~n11789 & ~n11792;
  assign n11794 = ~n11788 & ~n11793;
  assign n11795 = ~n11303 & ~n11794;
  assign n11796 = n11285 & ~n11300;
  assign n11797 = ~n11285 & n11300;
  assign n11798 = ~n11796 & ~n11797;
  assign n11799 = n5257 & ~n11792;
  assign n11800 = pi331 & n11799;
  assign n11801 = ~n11786 & ~n11789;
  assign n11802 = ~n11800 & ~n11801;
  assign n11803 = ~n11798 & ~n11802;
  assign n11804 = ~n11795 & ~n11803;
  assign n11805 = ~n10130 & n10154;
  assign n11806 = n10130 & ~n10154;
  assign n11807 = n10699 & ~n11806;
  assign n11808 = ~n11805 & ~n11807;
  assign n11809 = n11804 & n11808;
  assign n11810 = ~n11804 & ~n11808;
  assign n11811 = ~n11809 & ~n11810;
  assign n11812 = pi333 & n2887;
  assign n11813 = ~n10671 & ~n10687;
  assign n11814 = ~n10694 & n11813;
  assign n11815 = ~n10685 & ~n10687;
  assign n11816 = ~n10654 & n11815;
  assign n11817 = ~n10686 & ~n11816;
  assign n11818 = ~n11814 & n11817;
  assign n11819 = pi332 & n4596;
  assign n11820 = n11818 & ~n11819;
  assign n11821 = n4596 & ~n11818;
  assign n11822 = pi332 & n11821;
  assign n11823 = ~n11820 & ~n11822;
  assign n11824 = ~n11812 & n11823;
  assign n11825 = n11812 & ~n11823;
  assign n11826 = ~n11824 & ~n11825;
  assign n11827 = pi334 & n2464;
  assign n11828 = n10154 & ~n11242;
  assign n11829 = ~n10154 & ~n11251;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = n8810 & ~n10133;
  assign n11832 = ~n8810 & ~n10142;
  assign n11833 = ~n11831 & ~n11832;
  assign n11834 = ~n10711 & ~n11833;
  assign n11835 = ~n10714 & ~n11834;
  assign n11836 = ~n10704 & n11835;
  assign n11837 = ~n11830 & ~n11836;
  assign n11838 = n10704 & ~n11835;
  assign n11839 = ~n11837 & ~n11838;
  assign n11840 = n11827 & n11839;
  assign n11841 = ~n11827 & ~n11839;
  assign n11842 = ~n11840 & ~n11841;
  assign n11843 = ~n11826 & ~n11842;
  assign n11844 = n11812 & n11823;
  assign n11845 = ~n11812 & ~n11823;
  assign n11846 = ~n11844 & ~n11845;
  assign n11847 = ~n11827 & n11839;
  assign n11848 = n11827 & ~n11839;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = ~n11846 & ~n11849;
  assign n11851 = ~n11843 & ~n11850;
  assign n11852 = ~n11811 & ~n11851;
  assign n11853 = n11804 & ~n11808;
  assign n11854 = ~n11804 & n11808;
  assign n11855 = ~n11853 & ~n11854;
  assign n11856 = ~n11842 & ~n11846;
  assign n11857 = ~n11826 & ~n11849;
  assign n11858 = ~n11856 & ~n11857;
  assign n11859 = ~n11855 & ~n11858;
  assign n11860 = ~n11852 & ~n11859;
  assign n11861 = ~n11271 & n11860;
  assign n11862 = n11271 & ~n11860;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = pi337 & n1442;
  assign n11865 = ~n10750 & n10764;
  assign n11866 = n10750 & ~n10764;
  assign n11867 = ~n1442 & ~n11866;
  assign n11868 = ~n11865 & ~n11867;
  assign n11869 = n1729 & ~n11868;
  assign n11870 = ~n1729 & ~n11865;
  assign n11871 = n1442 & n11870;
  assign n11872 = ~n11869 & ~n11871;
  assign n11873 = pi336 & ~n11872;
  assign n11874 = pi336 & n1729;
  assign n11875 = n10750 & ~n11874;
  assign n11876 = ~n10764 & n11875;
  assign n11877 = ~n11873 & ~n11876;
  assign n11878 = n11864 & ~n11877;
  assign n11879 = ~n11864 & n11877;
  assign n11880 = ~n11878 & ~n11879;
  assign n11881 = ~n11863 & ~n11880;
  assign n11882 = n11271 & n11860;
  assign n11883 = ~n11271 & ~n11860;
  assign n11884 = ~n11882 & ~n11883;
  assign n11885 = ~n11864 & ~n11877;
  assign n11886 = n11864 & n11877;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11884 & ~n11887;
  assign n11889 = ~n11881 & ~n11888;
  assign n11890 = ~n11270 & ~n11889;
  assign n11891 = n11259 & ~n11267;
  assign n11892 = ~n11259 & n11267;
  assign n11893 = ~n11891 & ~n11892;
  assign n11894 = ~n11880 & ~n11884;
  assign n11895 = ~n11863 & ~n11887;
  assign n11896 = ~n11894 & ~n11895;
  assign n11897 = ~n11893 & ~n11896;
  assign n11898 = ~n11890 & ~n11897;
  assign n11899 = n11239 & n11898;
  assign n11900 = ~n11239 & ~n11898;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = pi339 & ~n1154;
  assign n11903 = n10790 & n11902;
  assign n11904 = ~n10790 & ~n11902;
  assign n11905 = ~n11903 & ~n11904;
  assign n11906 = n1156 & ~n11905;
  assign n11907 = pi340 & n11906;
  assign n11908 = pi340 & n1156;
  assign n11909 = ~n10790 & n11902;
  assign n11910 = n10790 & ~n11902;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n11908 & ~n11911;
  assign n11913 = ~n11907 & ~n11912;
  assign n11914 = ~n11901 & ~n11913;
  assign n11915 = ~n11239 & n11898;
  assign n11916 = n11239 & ~n11898;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = n1156 & ~n11911;
  assign n11919 = pi340 & n11918;
  assign n11920 = ~n11905 & ~n11908;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = ~n11917 & ~n11921;
  assign n11923 = ~n11914 & ~n11922;
  assign n11924 = ~n11228 & ~n11923;
  assign n11925 = n11228 & n11923;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = pi276 & ~n11926;
  assign n11928 = ~n11228 & n11923;
  assign n11929 = n11228 & ~n11923;
  assign n11930 = ~n11928 & ~n11929;
  assign n11931 = ~pi276 & ~n11930;
  assign n11932 = ~n11927 & ~n11931;
  assign n11933 = n11224 & n11932;
  assign n11934 = ~n11224 & ~n11932;
  assign n11935 = ~n11933 & ~n11934;
  assign n11936 = pi303 & ~n11935;
  assign n11937 = pi128 & n11936;
  assign n11938 = pi128 & pi303;
  assign n11939 = ~n11224 & n11932;
  assign n11940 = n11224 & ~n11932;
  assign n11941 = ~n11939 & ~n11940;
  assign n11942 = ~n11938 & ~n11941;
  assign n11943 = ~n11937 & ~n11942;
  assign n11944 = n10120 & ~n10822;
  assign n11945 = ~n10823 & ~n11944;
  assign n11946 = n11943 & ~n11945;
  assign n11947 = ~n11943 & n11945;
  assign n11948 = ~n11946 & ~n11947;
  assign n11949 = ~n831 & ~n11948;
  assign n11950 = ~n10833 & ~n11949;
  assign n11951 = pi161 & ~n11950;
  assign n11952 = pi082 & ~pi161;
  assign n11953 = ~n11951 & ~n11952;
  assign po211 = ~pi160 & ~n11953;
  assign n11955 = pi083 & ~pi161;
  assign n11956 = pi305 & n1553;
  assign n11957 = ~n1533 & ~n11161;
  assign n11958 = n1533 & n11161;
  assign n11959 = ~n10849 & ~n11958;
  assign n11960 = ~n11957 & ~n11959;
  assign n11961 = n1840 & ~n11960;
  assign n11962 = ~n1840 & ~n11163;
  assign n11963 = n1533 & n11962;
  assign n11964 = ~n11961 & ~n11963;
  assign n11965 = pi307 & ~n11964;
  assign n11966 = pi307 & n1840;
  assign n11967 = n11161 & ~n11966;
  assign n11968 = n10849 & n11967;
  assign n11969 = ~n11965 & ~n11968;
  assign n11970 = pi309 & n2574;
  assign n11971 = ~n3012 & ~n11090;
  assign n11972 = n3012 & n11090;
  assign n11973 = ~n10870 & ~n11972;
  assign n11974 = ~n11971 & ~n11973;
  assign n11975 = n3552 & ~n11974;
  assign n11976 = ~n3552 & ~n11092;
  assign n11977 = n3012 & n11976;
  assign n11978 = ~n11975 & ~n11977;
  assign n11979 = pi311 & ~n11978;
  assign n11980 = pi311 & n3552;
  assign n11981 = n11090 & ~n11980;
  assign n11982 = n10870 & n11981;
  assign n11983 = ~n11979 & ~n11982;
  assign n11984 = pi313 & n4772;
  assign n11985 = ~n10928 & ~n10937;
  assign n11986 = ~pi147 & n10899;
  assign n11987 = pi147 & ~n10899;
  assign n11988 = ~pi146 & n11987;
  assign n11989 = ~n11986 & ~n11988;
  assign n11990 = pi145 & ~n11989;
  assign n11991 = ~pi147 & ~n10899;
  assign n11992 = pi147 & n10899;
  assign n11993 = pi146 & n11992;
  assign n11994 = ~n11991 & ~n11993;
  assign n11995 = ~pi145 & ~n11994;
  assign n11996 = ~pi147 & ~n10906;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 = ~n11990 & n11997;
  assign n11999 = pi321 & n11998;
  assign n12000 = ~n10909 & n10915;
  assign n12001 = n9815 & ~n12000;
  assign n12002 = pi320 & n12001;
  assign n12003 = n10908 & ~n10915;
  assign n12004 = pi321 & n12003;
  assign n12005 = ~n12002 & ~n12004;
  assign n12006 = pi320 & n10908;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = n10908 & n12005;
  assign n12009 = pi320 & n12008;
  assign n12010 = ~n12007 & ~n12009;
  assign n12011 = ~n11999 & ~n12010;
  assign n12012 = n12005 & ~n12006;
  assign n12013 = n10908 & ~n12005;
  assign n12014 = pi320 & n12013;
  assign n12015 = ~n12012 & ~n12014;
  assign n12016 = n11998 & ~n12015;
  assign n12017 = pi321 & n12016;
  assign n12018 = ~n12011 & ~n12017;
  assign n12019 = pi319 & n9815;
  assign n12020 = n12018 & n12019;
  assign n12021 = ~n12018 & ~n12019;
  assign n12022 = ~n12020 & ~n12021;
  assign n12023 = ~n9517 & ~n12022;
  assign n12024 = ~pi318 & ~n12022;
  assign n12025 = n9517 & n12022;
  assign n12026 = pi318 & n12025;
  assign n12027 = ~n12024 & ~n12026;
  assign n12028 = ~pi319 & ~n12027;
  assign n12029 = ~n12023 & ~n12028;
  assign n12030 = ~n11985 & ~n12029;
  assign n12031 = n9517 & n10928;
  assign n12032 = n10937 & n12022;
  assign n12033 = n12031 & n12032;
  assign n12034 = n9517 & n11985;
  assign n12035 = ~n10928 & n10937;
  assign n12036 = n10928 & ~n10937;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = pi319 & ~n12037;
  assign n12039 = ~n12034 & ~n12038;
  assign n12040 = ~n12022 & ~n12039;
  assign n12041 = ~n12033 & ~n12040;
  assign n12042 = pi318 & ~n12041;
  assign n12043 = ~n10937 & n12022;
  assign n12044 = ~n9517 & ~n10928;
  assign n12045 = n12043 & n12044;
  assign n12046 = n10937 & ~n12022;
  assign n12047 = n10928 & n12046;
  assign n12048 = n10928 & n10937;
  assign n12049 = n9517 & ~n12048;
  assign n12050 = pi319 & n12049;
  assign n12051 = ~n11985 & ~n12050;
  assign n12052 = n12022 & ~n12051;
  assign n12053 = ~n12047 & ~n12052;
  assign n12054 = ~pi318 & ~n12053;
  assign n12055 = ~n12045 & ~n12054;
  assign n12056 = ~n12042 & n12055;
  assign n12057 = ~n12030 & n12056;
  assign n12058 = n10943 & ~n10946;
  assign n12059 = ~n9852 & ~n9859;
  assign n12060 = n9852 & n9859;
  assign n12061 = n9849 & ~n12060;
  assign n12062 = ~n12059 & ~n12061;
  assign n12063 = ~n10943 & n10946;
  assign n12064 = ~n12062 & ~n12063;
  assign n12065 = ~n12058 & ~n12064;
  assign n12066 = n12057 & ~n12065;
  assign n12067 = ~n12057 & n12065;
  assign n12068 = ~n12066 & ~n12067;
  assign n12069 = ~n10956 & ~n10966;
  assign n12070 = n10956 & n10966;
  assign n12071 = ~n10957 & ~n12070;
  assign n12072 = ~n9864 & n12071;
  assign n12073 = ~n12069 & ~n12072;
  assign n12074 = n12068 & n12073;
  assign n12075 = ~n12068 & ~n12073;
  assign n12076 = ~n12074 & ~n12075;
  assign n12077 = pi317 & n7874;
  assign n12078 = pi316 & n7044;
  assign n12079 = ~n12077 & ~n12078;
  assign n12080 = n12077 & n12078;
  assign n12081 = ~n12079 & ~n12080;
  assign n12082 = ~n12076 & ~n12081;
  assign n12083 = ~n12068 & n12073;
  assign n12084 = n12068 & ~n12073;
  assign n12085 = ~n12083 & ~n12084;
  assign n12086 = n7874 & ~n12078;
  assign n12087 = pi317 & n12086;
  assign n12088 = n7044 & ~n12077;
  assign n12089 = pi316 & n12088;
  assign n12090 = ~n12087 & ~n12089;
  assign n12091 = ~n12085 & ~n12090;
  assign n12092 = ~n12082 & ~n12091;
  assign n12093 = ~n6777 & n10972;
  assign n12094 = ~n10996 & ~n12093;
  assign n12095 = n5463 & n12094;
  assign n12096 = ~n10888 & n10972;
  assign n12097 = n6777 & ~n12096;
  assign n12098 = ~n12095 & ~n12097;
  assign n12099 = pi316 & ~n12098;
  assign n12100 = ~n10984 & ~n12099;
  assign n12101 = n12092 & n12100;
  assign n12102 = ~n12092 & ~n12100;
  assign n12103 = ~n12101 & ~n12102;
  assign n12104 = n6777 & ~n12103;
  assign n12105 = pi315 & n12104;
  assign n12106 = pi315 & n6777;
  assign n12107 = ~n12092 & n12100;
  assign n12108 = n12092 & ~n12100;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = ~n12106 & ~n12109;
  assign n12111 = ~n12105 & ~n12110;
  assign n12112 = ~n11016 & n11022;
  assign n12113 = n11016 & ~n11022;
  assign n12114 = ~n11008 & ~n12113;
  assign n12115 = ~n12112 & ~n12114;
  assign n12116 = n12111 & n12115;
  assign n12117 = ~n12111 & ~n12115;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = pi314 & n5463;
  assign n12120 = ~n11035 & ~n12119;
  assign n12121 = ~n11029 & n12120;
  assign n12122 = ~n11029 & ~n11035;
  assign n12123 = n12119 & ~n12122;
  assign n12124 = ~n12121 & ~n12123;
  assign n12125 = ~n12118 & ~n12124;
  assign n12126 = n12111 & ~n12115;
  assign n12127 = ~n12111 & n12115;
  assign n12128 = ~n12126 & ~n12127;
  assign n12129 = ~n11035 & n12119;
  assign n12130 = ~n11029 & n12129;
  assign n12131 = ~n12119 & ~n12122;
  assign n12132 = ~n12130 & ~n12131;
  assign n12133 = ~n12128 & ~n12132;
  assign n12134 = ~n12125 & ~n12133;
  assign n12135 = ~n11984 & n12134;
  assign n12136 = n11984 & ~n12134;
  assign n12137 = ~n12135 & ~n12136;
  assign n12138 = pi312 & n4086;
  assign n12139 = n9619 & ~n9983;
  assign n12140 = n3012 & ~n11064;
  assign n12141 = pi313 & n12140;
  assign n12142 = ~n12139 & ~n12141;
  assign n12143 = ~n9972 & ~n12142;
  assign n12144 = n9619 & n12140;
  assign n12145 = ~n11065 & ~n12144;
  assign n12146 = pi313 & ~n12145;
  assign n12147 = ~n12143 & ~n12146;
  assign n12148 = n11037 & ~n12147;
  assign n12149 = ~n11037 & n12147;
  assign n12150 = n10871 & ~n12149;
  assign n12151 = ~n12148 & ~n12150;
  assign n12152 = n12138 & ~n12151;
  assign n12153 = ~n10871 & ~n12148;
  assign n12154 = ~n12149 & ~n12153;
  assign n12155 = ~n12138 & ~n12154;
  assign n12156 = ~n12152 & ~n12155;
  assign n12157 = ~n12137 & ~n12156;
  assign n12158 = ~n11984 & ~n12134;
  assign n12159 = n11984 & n12134;
  assign n12160 = ~n12158 & ~n12159;
  assign n12161 = ~n12138 & ~n12151;
  assign n12162 = n12138 & ~n12154;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n12160 & ~n12163;
  assign n12165 = ~n12157 & ~n12164;
  assign n12166 = n11041 & ~n11085;
  assign n12167 = ~n11041 & n11085;
  assign n12168 = ~n11076 & ~n12167;
  assign n12169 = ~n12166 & ~n12168;
  assign n12170 = ~n12165 & ~n12169;
  assign n12171 = n12165 & n12169;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = n11983 & n12172;
  assign n12174 = ~n11983 & ~n12172;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = pi310 & n3012;
  assign n12177 = ~n10866 & ~n11106;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = ~n11103 & n12178;
  assign n12180 = ~n11103 & ~n12177;
  assign n12181 = n12176 & ~n12180;
  assign n12182 = ~n12179 & ~n12181;
  assign n12183 = ~n12175 & ~n12182;
  assign n12184 = n11983 & ~n12172;
  assign n12185 = ~n11983 & n12172;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = n12176 & ~n12177;
  assign n12188 = ~n11103 & n12187;
  assign n12189 = ~n12176 & ~n12180;
  assign n12190 = ~n12188 & ~n12189;
  assign n12191 = ~n12186 & ~n12190;
  assign n12192 = ~n12183 & ~n12191;
  assign n12193 = ~n11970 & ~n12192;
  assign n12194 = n11970 & n12192;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = pi308 & n2183;
  assign n12197 = n1533 & ~n11122;
  assign n12198 = pi309 & n12197;
  assign n12199 = ~n9699 & ~n10061;
  assign n12200 = ~n12198 & ~n12199;
  assign n12201 = ~n9466 & ~n12200;
  assign n12202 = n1840 & ~n10046;
  assign n12203 = ~n9699 & n12197;
  assign n12204 = ~n12202 & ~n12203;
  assign n12205 = pi309 & ~n12204;
  assign n12206 = ~n12201 & ~n12205;
  assign n12207 = ~n11111 & ~n12206;
  assign n12208 = n11111 & n12206;
  assign n12209 = n10850 & ~n12208;
  assign n12210 = ~n12207 & ~n12209;
  assign n12211 = n12196 & ~n12210;
  assign n12212 = ~n10850 & ~n12207;
  assign n12213 = ~n12208 & ~n12212;
  assign n12214 = ~n12196 & ~n12213;
  assign n12215 = ~n12211 & ~n12214;
  assign n12216 = ~n12195 & ~n12215;
  assign n12217 = ~n11970 & n12192;
  assign n12218 = n11970 & ~n12192;
  assign n12219 = ~n12217 & ~n12218;
  assign n12220 = ~n12196 & ~n12210;
  assign n12221 = n12196 & ~n12213;
  assign n12222 = ~n12220 & ~n12221;
  assign n12223 = ~n12219 & ~n12222;
  assign n12224 = ~n12216 & ~n12223;
  assign n12225 = ~n11114 & ~n11115;
  assign n12226 = n11114 & n11115;
  assign n12227 = ~n11150 & ~n12226;
  assign n12228 = ~n12225 & ~n12227;
  assign n12229 = n12224 & ~n12228;
  assign n12230 = ~n12224 & n12228;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = n11969 & ~n12231;
  assign n12233 = ~n11969 & n12231;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = pi306 & n1533;
  assign n12236 = n10842 & ~n11174;
  assign n12237 = n12235 & ~n12236;
  assign n12238 = ~n11177 & n12237;
  assign n12239 = ~n11177 & ~n12236;
  assign n12240 = ~n12235 & ~n12239;
  assign n12241 = ~n12238 & ~n12240;
  assign n12242 = ~n12234 & ~n12241;
  assign n12243 = n11969 & n12231;
  assign n12244 = ~n11969 & ~n12231;
  assign n12245 = ~n12243 & ~n12244;
  assign n12246 = ~n12235 & ~n12236;
  assign n12247 = ~n11177 & n12246;
  assign n12248 = n12235 & ~n12239;
  assign n12249 = ~n12247 & ~n12248;
  assign n12250 = ~n12245 & ~n12249;
  assign n12251 = ~n12242 & ~n12250;
  assign n12252 = ~n11956 & n12251;
  assign n12253 = n11956 & ~n12251;
  assign n12254 = ~n12252 & ~n12253;
  assign n12255 = pi304 & n1515;
  assign n12256 = n11182 & n11211;
  assign n12257 = ~n12255 & ~n12256;
  assign n12258 = ~n11197 & n12257;
  assign n12259 = ~n11197 & ~n12256;
  assign n12260 = n12255 & ~n12259;
  assign n12261 = ~n12258 & ~n12260;
  assign n12262 = ~n12254 & ~n12261;
  assign n12263 = ~n11956 & ~n12251;
  assign n12264 = n11956 & n12251;
  assign n12265 = ~n12263 & ~n12264;
  assign n12266 = n12255 & ~n12256;
  assign n12267 = ~n11197 & n12266;
  assign n12268 = ~n12255 & ~n12259;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = ~n12265 & ~n12269;
  assign n12271 = ~n12262 & ~n12270;
  assign n12272 = n10834 & n11187;
  assign n12273 = ~n10834 & ~n11187;
  assign n12274 = n11182 & ~n11212;
  assign n12275 = ~n11182 & n11212;
  assign n12276 = ~n12274 & ~n12275;
  assign n12277 = ~n12273 & ~n12276;
  assign n12278 = ~n12272 & ~n12277;
  assign n12279 = ~n12271 & ~n12278;
  assign n12280 = n12271 & n12278;
  assign n12281 = ~n12279 & ~n12280;
  assign n12282 = pi130 & pi305;
  assign n12283 = ~pi129 & ~n12282;
  assign n12284 = pi128 & ~pi130;
  assign n12285 = pi305 & ~n12284;
  assign n12286 = ~n1514 & n12285;
  assign n12287 = n10109 & ~n12286;
  assign n12288 = ~n12283 & ~n12287;
  assign n12289 = n9777 & ~n12288;
  assign n12290 = ~pi129 & n11188;
  assign n12291 = pi130 & ~n10109;
  assign n12292 = pi129 & n12291;
  assign n12293 = ~n12290 & ~n12292;
  assign n12294 = pi128 & ~n12293;
  assign n12295 = ~n9777 & n10109;
  assign n12296 = pi130 & n12295;
  assign n12297 = ~pi130 & ~n10109;
  assign n12298 = pi129 & n12297;
  assign n12299 = ~n12296 & ~n12298;
  assign n12300 = ~pi128 & ~n12299;
  assign n12301 = pi129 & n10109;
  assign n12302 = ~pi129 & ~n10109;
  assign n12303 = ~n12301 & ~n12302;
  assign n12304 = ~n9777 & ~n12303;
  assign n12305 = pi130 & n12304;
  assign n12306 = ~n12300 & ~n12305;
  assign n12307 = ~n12294 & n12306;
  assign n12308 = pi305 & ~n12307;
  assign n12309 = ~n12289 & ~n12308;
  assign n12310 = n11182 & n12309;
  assign n12311 = ~n11182 & ~n12309;
  assign n12312 = ~n12310 & ~n12311;
  assign n12313 = ~n12272 & ~n12273;
  assign n12314 = ~n12312 & ~n12313;
  assign n12315 = ~n11182 & n12309;
  assign n12316 = n11182 & ~n12309;
  assign n12317 = ~n12315 & ~n12316;
  assign n12318 = ~n10834 & n11187;
  assign n12319 = n10834 & ~n11187;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = ~n12317 & ~n12320;
  assign n12322 = ~n12314 & ~n12321;
  assign n12323 = pi303 & ~n12322;
  assign n12324 = pi128 & n12323;
  assign n12325 = pi129 & n12324;
  assign n12326 = pi303 & ~n1568;
  assign n12327 = ~n12324 & n12326;
  assign n12328 = ~n12325 & ~n12327;
  assign n12329 = ~n12281 & ~n12328;
  assign n12330 = n12271 & ~n12278;
  assign n12331 = ~n12271 & n12278;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = ~pi129 & n12324;
  assign n12334 = ~n12324 & ~n12326;
  assign n12335 = ~n12333 & ~n12334;
  assign n12336 = ~n12332 & ~n12335;
  assign n12337 = ~n12329 & ~n12336;
  assign n12338 = ~n11932 & ~n11945;
  assign n12339 = n11932 & n11945;
  assign n12340 = ~n11224 & ~n11938;
  assign n12341 = pi303 & n11224;
  assign n12342 = pi128 & n12341;
  assign n12343 = ~n12340 & ~n12342;
  assign n12344 = ~n12339 & ~n12343;
  assign n12345 = ~n12338 & ~n12344;
  assign n12346 = ~n12337 & n12345;
  assign n12347 = n12337 & ~n12345;
  assign n12348 = ~n12346 & ~n12347;
  assign n12349 = ~pi276 & ~n11925;
  assign n12350 = ~n11924 & ~n12349;
  assign n12351 = pi340 & ~n1154;
  assign n12352 = ~n11901 & ~n11905;
  assign n12353 = pi128 & pi340;
  assign n12354 = pi258 & n12353;
  assign n12355 = ~n11911 & ~n11917;
  assign n12356 = n12354 & ~n12355;
  assign n12357 = ~n12352 & n12356;
  assign n12358 = ~n12351 & ~n12357;
  assign n12359 = pi339 & n10790;
  assign n12360 = ~pi339 & ~n10790;
  assign n12361 = ~n12359 & ~n12360;
  assign n12362 = ~n11917 & ~n12361;
  assign n12363 = pi339 & ~n10790;
  assign n12364 = ~pi339 & n10790;
  assign n12365 = ~n12363 & ~n12364;
  assign n12366 = ~n11901 & ~n12365;
  assign n12367 = ~n12362 & ~n12366;
  assign n12368 = n12354 & ~n12367;
  assign n12369 = ~n1154 & n12368;
  assign n12370 = ~n12358 & ~n12369;
  assign n12371 = n11259 & n11271;
  assign n12372 = ~n11259 & ~n11271;
  assign n12373 = n11860 & ~n12372;
  assign n12374 = ~n12371 & ~n12373;
  assign n12375 = ~n11259 & n11860;
  assign n12376 = n11259 & ~n11860;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = n11271 & ~n11877;
  assign n12379 = ~n11271 & n11877;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = n11267 & ~n11864;
  assign n12382 = ~n12380 & ~n12381;
  assign n12383 = ~n12377 & n12382;
  assign n12384 = ~n11267 & n11864;
  assign n12385 = ~n11259 & ~n11860;
  assign n12386 = n11259 & n11860;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = ~n11271 & ~n11877;
  assign n12389 = n11271 & n11877;
  assign n12390 = ~n12388 & ~n12389;
  assign n12391 = ~n12381 & ~n12390;
  assign n12392 = ~n12387 & n12391;
  assign n12393 = ~n12384 & ~n12392;
  assign n12394 = ~n12383 & n12393;
  assign n12395 = ~n12374 & n12394;
  assign n12396 = n12374 & ~n12394;
  assign n12397 = ~n12395 & ~n12396;
  assign n12398 = pi335 & n2464;
  assign n12399 = n11285 & n11761;
  assign n12400 = n5973 & ~n11760;
  assign n12401 = pi328 & n12400;
  assign n12402 = ~n11762 & ~n11769;
  assign n12403 = ~n12401 & ~n12402;
  assign n12404 = ~n11336 & ~n12403;
  assign n12405 = n5973 & ~n11769;
  assign n12406 = pi328 & n12405;
  assign n12407 = ~n11760 & ~n11762;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = ~n11778 & ~n12408;
  assign n12410 = ~n12404 & ~n12409;
  assign n12411 = ~n11285 & ~n11761;
  assign n12412 = n12410 & ~n12411;
  assign n12413 = ~n12399 & ~n12412;
  assign n12414 = ~n11285 & n11783;
  assign n12415 = n11285 & ~n11783;
  assign n12416 = ~n12414 & ~n12415;
  assign n12417 = ~n11310 & ~n12416;
  assign n12418 = n11285 & n11783;
  assign n12419 = ~n11285 & ~n11783;
  assign n12420 = ~n12418 & ~n12419;
  assign n12421 = n11310 & ~n12420;
  assign n12422 = ~n12417 & ~n12421;
  assign n12423 = n11300 & ~n11789;
  assign n12424 = ~n12422 & ~n12423;
  assign n12425 = n5257 & ~n11300;
  assign n12426 = pi331 & n12425;
  assign n12427 = ~n12424 & ~n12426;
  assign n12428 = ~n12413 & n12427;
  assign n12429 = n12413 & ~n12427;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = ~pi330 & ~n11305;
  assign n12432 = n11305 & ~n11308;
  assign n12433 = ~n5732 & ~n12432;
  assign n12434 = ~n12431 & ~n12433;
  assign n12435 = ~n12420 & ~n12434;
  assign n12436 = ~n5732 & ~n11305;
  assign n12437 = n5714 & n12436;
  assign n12438 = ~n5714 & n11305;
  assign n12439 = n5714 & ~n11305;
  assign n12440 = ~n12416 & ~n12439;
  assign n12441 = ~n12438 & ~n12440;
  assign n12442 = n5732 & ~n12441;
  assign n12443 = ~n12437 & ~n12442;
  assign n12444 = pi330 & ~n12443;
  assign n12445 = ~n12435 & ~n12444;
  assign n12446 = n11330 & n11337;
  assign n12447 = ~n11330 & ~n11337;
  assign n12448 = n11757 & ~n12447;
  assign n12449 = ~n12446 & ~n12448;
  assign n12450 = ~n11333 & n11762;
  assign n12451 = ~n11330 & ~n11757;
  assign n12452 = n11330 & n11757;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = n11337 & ~n12453;
  assign n12455 = n11330 & ~n11757;
  assign n12456 = ~n11330 & n11757;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~n11337 & ~n12457;
  assign n12459 = ~n12454 & ~n12458;
  assign n12460 = n11333 & ~n11762;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~n12450 & ~n12461;
  assign n12463 = ~n12449 & ~n12462;
  assign n12464 = n12449 & n12462;
  assign n12465 = ~n12463 & ~n12464;
  assign n12466 = pi327 & n9205;
  assign n12467 = ~n11356 & n11736;
  assign n12468 = n11356 & ~n11736;
  assign n12469 = ~n11734 & ~n12468;
  assign n12470 = ~n12467 & ~n12469;
  assign n12471 = ~n11356 & n11731;
  assign n12472 = n11356 & ~n11731;
  assign n12473 = ~n12471 & ~n12472;
  assign n12474 = ~n11727 & n11736;
  assign n12475 = n11727 & ~n11736;
  assign n12476 = ~n12474 & ~n12475;
  assign n12477 = n11360 & ~n11735;
  assign n12478 = ~n12476 & ~n12477;
  assign n12479 = ~n12473 & n12478;
  assign n12480 = ~n11360 & n11735;
  assign n12481 = ~n11356 & ~n11731;
  assign n12482 = n11356 & n11731;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = n11727 & n11736;
  assign n12485 = ~n11727 & ~n11736;
  assign n12486 = ~n12484 & ~n12485;
  assign n12487 = ~n12477 & ~n12486;
  assign n12488 = ~n12483 & n12487;
  assign n12489 = ~n12480 & ~n12488;
  assign n12490 = ~n12479 & n12489;
  assign n12491 = n12470 & ~n12490;
  assign n12492 = ~n12470 & n12490;
  assign n12493 = ~n12491 & ~n12492;
  assign n12494 = pi324 & n11384;
  assign n12495 = ~n11369 & n11384;
  assign n12496 = pi323 & n12495;
  assign n12497 = n11369 & ~n11385;
  assign n12498 = n11711 & ~n12497;
  assign n12499 = pi322 & n12498;
  assign n12500 = ~n12496 & ~n12499;
  assign n12501 = ~n12494 & ~n12500;
  assign n12502 = n12494 & n12500;
  assign n12503 = ~n12501 & ~n12502;
  assign n12504 = pi323 & n11711;
  assign n12505 = pi259 & n11681;
  assign n12506 = ~pi259 & ~n11681;
  assign n12507 = pi258 & ~n12506;
  assign n12508 = n10534 & n12507;
  assign n12509 = ~n12505 & ~n12508;
  assign n12510 = pi145 & ~n12509;
  assign n12511 = ~n11681 & ~n11691;
  assign n12512 = n11681 & n11691;
  assign n12513 = ~n12511 & ~n12512;
  assign n12514 = n10534 & n11690;
  assign n12515 = n10228 & n12514;
  assign n12516 = ~n11685 & ~n11689;
  assign n12517 = ~n11690 & ~n12516;
  assign n12518 = ~n12515 & ~n12517;
  assign n12519 = ~n12513 & ~n12518;
  assign n12520 = ~n10534 & n11685;
  assign n12521 = ~n10228 & n12520;
  assign n12522 = ~n11681 & n11691;
  assign n12523 = n11681 & ~n11691;
  assign n12524 = ~n12522 & ~n12523;
  assign n12525 = n10534 & ~n11690;
  assign n12526 = n10228 & n12525;
  assign n12527 = n11690 & ~n12516;
  assign n12528 = ~n12526 & ~n12527;
  assign n12529 = ~n12524 & ~n12528;
  assign n12530 = ~n12521 & ~n12529;
  assign n12531 = ~n12519 & n12530;
  assign n12532 = n12510 & n12531;
  assign n12533 = ~n12510 & ~n12531;
  assign n12534 = ~n12532 & ~n12533;
  assign n12535 = ~n10534 & n11681;
  assign n12536 = pi259 & n12535;
  assign n12537 = n10534 & ~n11681;
  assign n12538 = pi258 & n12537;
  assign n12539 = ~n12536 & ~n12538;
  assign n12540 = pi145 & ~n12539;
  assign n12541 = pi259 & ~n11681;
  assign n12542 = ~pi259 & n11681;
  assign n12543 = pi258 & n12542;
  assign n12544 = ~n12541 & ~n12543;
  assign n12545 = ~pi145 & ~n12544;
  assign n12546 = n1147 & n12535;
  assign n12547 = ~n1146 & ~n12546;
  assign n12548 = ~n12545 & n12547;
  assign n12549 = ~n12540 & n12548;
  assign n12550 = pi146 & ~n12549;
  assign n12551 = pi131 & pi274;
  assign n12552 = ~n11445 & n11451;
  assign n12553 = ~n11441 & n12552;
  assign n12554 = ~n11446 & ~n11451;
  assign n12555 = ~n12553 & ~n12554;
  assign n12556 = pi273 & ~n12555;
  assign n12557 = pi131 & n12556;
  assign n12558 = n11416 & n11419;
  assign n12559 = ~n11416 & ~n11419;
  assign n12560 = ~n11438 & ~n12559;
  assign n12561 = ~n12558 & ~n12560;
  assign n12562 = pi128 & pi277;
  assign n12563 = pi276 & ~n12562;
  assign n12564 = pi129 & n12563;
  assign n12565 = pi129 & pi276;
  assign n12566 = pi277 & ~n12565;
  assign n12567 = pi128 & n12566;
  assign n12568 = ~n12564 & ~n12567;
  assign n12569 = ~n12561 & n12568;
  assign n12570 = n12561 & ~n12568;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = pi275 & ~n12571;
  assign n12573 = pi130 & n12572;
  assign n12574 = pi130 & pi275;
  assign n12575 = ~n12570 & ~n12574;
  assign n12576 = ~n12569 & n12575;
  assign n12577 = ~n12573 & ~n12576;
  assign n12578 = ~n11441 & n11451;
  assign n12579 = ~n11445 & ~n12578;
  assign n12580 = ~n12577 & ~n12579;
  assign n12581 = ~n12576 & ~n12578;
  assign n12582 = ~n12573 & n12581;
  assign n12583 = ~n11445 & n12582;
  assign n12584 = ~n12580 & ~n12583;
  assign n12585 = ~n11452 & ~n12553;
  assign n12586 = ~n12554 & n12585;
  assign n12587 = ~n11469 & ~n12586;
  assign n12588 = ~n12584 & ~n12587;
  assign n12589 = ~n12557 & n12588;
  assign n12590 = ~n12557 & ~n12587;
  assign n12591 = n12584 & ~n12590;
  assign n12592 = ~n12589 & ~n12591;
  assign n12593 = ~n12551 & ~n12592;
  assign n12594 = n12584 & ~n12587;
  assign n12595 = ~n12557 & n12594;
  assign n12596 = ~n12584 & ~n12590;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = pi274 & ~n12597;
  assign n12599 = pi131 & n12598;
  assign n12600 = ~n12593 & ~n12599;
  assign n12601 = n11473 & ~n11484;
  assign n12602 = ~n11473 & n11484;
  assign n12603 = ~n11475 & ~n12602;
  assign n12604 = ~n12601 & ~n12603;
  assign n12605 = n12600 & n12604;
  assign n12606 = ~n12600 & ~n12604;
  assign n12607 = ~n12605 & ~n12606;
  assign n12608 = pi133 & pi272;
  assign n12609 = pi132 & pi273;
  assign n12610 = n12608 & n12609;
  assign n12611 = ~n12608 & ~n12609;
  assign n12612 = ~n12610 & ~n12611;
  assign n12613 = ~n12607 & ~n12612;
  assign n12614 = ~n12600 & n12604;
  assign n12615 = n12600 & ~n12604;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = pi272 & ~n12609;
  assign n12618 = pi133 & n12617;
  assign n12619 = pi273 & ~n12608;
  assign n12620 = pi132 & n12619;
  assign n12621 = ~n12618 & ~n12620;
  assign n12622 = ~n12616 & ~n12621;
  assign n12623 = ~n12613 & ~n12622;
  assign n12624 = ~n11505 & ~n11509;
  assign n12625 = ~n11510 & ~n12624;
  assign n12626 = n12623 & n12625;
  assign n12627 = ~n12623 & ~n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = pi134 & pi271;
  assign n12630 = n11489 & ~n11502;
  assign n12631 = ~n11498 & n12630;
  assign n12632 = ~n11489 & ~n11505;
  assign n12633 = ~n12631 & ~n12632;
  assign n12634 = ~n11414 & ~n12633;
  assign n12635 = ~n11489 & ~n11502;
  assign n12636 = ~n11498 & n12635;
  assign n12637 = n11489 & ~n11505;
  assign n12638 = ~n12636 & ~n12637;
  assign n12639 = pi271 & ~n12638;
  assign n12640 = pi133 & n12639;
  assign n12641 = ~n12634 & ~n12640;
  assign n12642 = ~n11521 & ~n12641;
  assign n12643 = n11521 & n12641;
  assign n12644 = n11499 & ~n12643;
  assign n12645 = ~n12642 & ~n12644;
  assign n12646 = n12629 & ~n12645;
  assign n12647 = ~n11499 & ~n12642;
  assign n12648 = ~n12643 & ~n12647;
  assign n12649 = ~n12629 & ~n12648;
  assign n12650 = ~n12646 & ~n12649;
  assign n12651 = ~n12628 & ~n12650;
  assign n12652 = n12623 & ~n12625;
  assign n12653 = ~n12623 & n12625;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = ~n12629 & ~n12645;
  assign n12656 = n12629 & ~n12648;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12654 & ~n12657;
  assign n12659 = ~n12651 & ~n12658;
  assign n12660 = ~n11524 & ~n11525;
  assign n12661 = n11524 & n11525;
  assign n12662 = ~n11530 & ~n12661;
  assign n12663 = ~n12660 & ~n12662;
  assign n12664 = ~n12659 & n12663;
  assign n12665 = n12659 & ~n12663;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = pi136 & pi269;
  assign n12668 = pi135 & pi270;
  assign n12669 = n12667 & n12668;
  assign n12670 = ~n12667 & ~n12668;
  assign n12671 = ~n12669 & ~n12670;
  assign n12672 = ~n12666 & ~n12671;
  assign n12673 = n12659 & n12663;
  assign n12674 = ~n12659 & ~n12663;
  assign n12675 = ~n12673 & ~n12674;
  assign n12676 = pi269 & ~n12668;
  assign n12677 = pi136 & n12676;
  assign n12678 = pi270 & ~n12667;
  assign n12679 = pi135 & n12678;
  assign n12680 = ~n12677 & ~n12679;
  assign n12681 = ~n12675 & ~n12680;
  assign n12682 = ~n12672 & ~n12681;
  assign n12683 = ~n11557 & ~n11561;
  assign n12684 = ~n11562 & ~n12683;
  assign n12685 = n12682 & n12684;
  assign n12686 = ~n12682 & ~n12684;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = pi137 & pi268;
  assign n12689 = n11541 & ~n11554;
  assign n12690 = ~n11550 & n12689;
  assign n12691 = ~n11541 & ~n11557;
  assign n12692 = ~n12690 & ~n12691;
  assign n12693 = ~n11413 & ~n12692;
  assign n12694 = ~n11541 & ~n11554;
  assign n12695 = ~n11550 & n12694;
  assign n12696 = n11541 & ~n11557;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = pi268 & ~n12697;
  assign n12699 = pi136 & n12698;
  assign n12700 = ~n12693 & ~n12699;
  assign n12701 = ~n11573 & ~n12700;
  assign n12702 = n11573 & n12700;
  assign n12703 = n11551 & ~n12702;
  assign n12704 = ~n12701 & ~n12703;
  assign n12705 = n12688 & ~n12704;
  assign n12706 = ~n11551 & ~n12701;
  assign n12707 = ~n12702 & ~n12706;
  assign n12708 = ~n12688 & ~n12707;
  assign n12709 = ~n12705 & ~n12708;
  assign n12710 = ~n12687 & ~n12709;
  assign n12711 = n12682 & ~n12684;
  assign n12712 = ~n12682 & n12684;
  assign n12713 = ~n12711 & ~n12712;
  assign n12714 = ~n12688 & ~n12704;
  assign n12715 = n12688 & ~n12707;
  assign n12716 = ~n12714 & ~n12715;
  assign n12717 = ~n12713 & ~n12716;
  assign n12718 = ~n12710 & ~n12717;
  assign n12719 = ~n11577 & ~n11588;
  assign n12720 = n11577 & n11588;
  assign n12721 = ~n11582 & ~n12720;
  assign n12722 = ~n12719 & ~n12721;
  assign n12723 = ~n12718 & n12722;
  assign n12724 = n12718 & ~n12722;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = pi139 & pi266;
  assign n12727 = pi138 & pi267;
  assign n12728 = n12726 & n12727;
  assign n12729 = ~n12726 & ~n12727;
  assign n12730 = ~n12728 & ~n12729;
  assign n12731 = ~n12725 & ~n12730;
  assign n12732 = n12718 & n12722;
  assign n12733 = ~n12718 & ~n12722;
  assign n12734 = ~n12732 & ~n12733;
  assign n12735 = pi266 & ~n12727;
  assign n12736 = pi139 & n12735;
  assign n12737 = pi267 & ~n12726;
  assign n12738 = pi138 & n12737;
  assign n12739 = ~n12736 & ~n12738;
  assign n12740 = ~n12734 & ~n12739;
  assign n12741 = ~n12731 & ~n12740;
  assign n12742 = ~n11606 & ~n11613;
  assign n12743 = ~n11601 & n12742;
  assign n12744 = ~n11614 & ~n12743;
  assign n12745 = n12741 & n12744;
  assign n12746 = ~n12741 & ~n12744;
  assign n12747 = ~n12745 & ~n12746;
  assign n12748 = pi140 & pi265;
  assign n12749 = ~n11593 & ~n11606;
  assign n12750 = ~n11601 & n12749;
  assign n12751 = n11593 & ~n11609;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = ~n11412 & ~n12752;
  assign n12754 = n11593 & ~n11606;
  assign n12755 = ~n11601 & n12754;
  assign n12756 = ~n11593 & ~n11609;
  assign n12757 = ~n12755 & ~n12756;
  assign n12758 = pi265 & ~n12757;
  assign n12759 = pi139 & n12758;
  assign n12760 = ~n12753 & ~n12759;
  assign n12761 = n11625 & n12760;
  assign n12762 = ~n11625 & ~n12760;
  assign n12763 = n11602 & ~n12762;
  assign n12764 = ~n12761 & ~n12763;
  assign n12765 = n12748 & ~n12764;
  assign n12766 = ~n11602 & ~n12761;
  assign n12767 = ~n12762 & ~n12766;
  assign n12768 = ~n12748 & ~n12767;
  assign n12769 = ~n12765 & ~n12768;
  assign n12770 = ~n12747 & ~n12769;
  assign n12771 = n12741 & ~n12744;
  assign n12772 = ~n12741 & n12744;
  assign n12773 = ~n12771 & ~n12772;
  assign n12774 = ~n12748 & ~n12764;
  assign n12775 = n12748 & ~n12767;
  assign n12776 = ~n12774 & ~n12775;
  assign n12777 = ~n12773 & ~n12776;
  assign n12778 = ~n12770 & ~n12777;
  assign n12779 = ~n11628 & ~n11631;
  assign n12780 = ~n10483 & ~n10488;
  assign n12781 = ~n10489 & ~n12780;
  assign n12782 = n11628 & n11631;
  assign n12783 = ~n12781 & ~n12782;
  assign n12784 = ~n12779 & ~n12783;
  assign n12785 = ~n12778 & n12784;
  assign n12786 = n12778 & ~n12784;
  assign n12787 = ~n12785 & ~n12786;
  assign n12788 = pi142 & pi263;
  assign n12789 = pi141 & pi264;
  assign n12790 = n12788 & n12789;
  assign n12791 = ~n12788 & ~n12789;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = ~n12787 & ~n12792;
  assign n12794 = n12778 & n12784;
  assign n12795 = ~n12778 & ~n12784;
  assign n12796 = ~n12794 & ~n12795;
  assign n12797 = pi263 & ~n12789;
  assign n12798 = pi142 & n12797;
  assign n12799 = pi264 & ~n12788;
  assign n12800 = pi141 & n12799;
  assign n12801 = ~n12798 & ~n12800;
  assign n12802 = ~n12796 & ~n12801;
  assign n12803 = ~n12793 & ~n12802;
  assign n12804 = n11644 & ~n11654;
  assign n12805 = ~n11644 & n11654;
  assign n12806 = ~n11645 & ~n12805;
  assign n12807 = ~n11395 & n12806;
  assign n12808 = ~n12804 & ~n12807;
  assign n12809 = n12803 & ~n12808;
  assign n12810 = ~n12803 & n12808;
  assign n12811 = ~n12809 & ~n12810;
  assign n12812 = pi143 & pi262;
  assign n12813 = ~n11401 & n11660;
  assign n12814 = n11401 & ~n11660;
  assign n12815 = n11411 & ~n12814;
  assign n12816 = ~n12813 & ~n12815;
  assign n12817 = n12812 & ~n12816;
  assign n12818 = ~n11411 & ~n12813;
  assign n12819 = ~n12814 & ~n12818;
  assign n12820 = ~n12812 & ~n12819;
  assign n12821 = ~n12817 & ~n12820;
  assign n12822 = ~n12811 & ~n12821;
  assign n12823 = n12803 & n12808;
  assign n12824 = ~n12803 & ~n12808;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = ~n12812 & ~n12816;
  assign n12827 = n12812 & ~n12819;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = ~n12825 & ~n12828;
  assign n12830 = ~n12822 & ~n12829;
  assign n12831 = n11401 & n11660;
  assign n12832 = ~n11401 & ~n11660;
  assign n12833 = ~n12831 & ~n12832;
  assign n12834 = ~n11411 & ~n12833;
  assign n12835 = ~n12813 & ~n12814;
  assign n12836 = n11411 & ~n12835;
  assign n12837 = ~n12834 & ~n12836;
  assign n12838 = n11407 & ~n11666;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = pi260 & ~n11407;
  assign n12841 = pi144 & n12840;
  assign n12842 = ~n12839 & ~n12841;
  assign n12843 = ~n12830 & n12842;
  assign n12844 = n12830 & ~n12842;
  assign n12845 = ~n12843 & ~n12844;
  assign n12846 = pi145 & pi260;
  assign n12847 = pi144 & pi261;
  assign n12848 = n12846 & n12847;
  assign n12849 = ~n12846 & ~n12847;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = ~n12845 & ~n12850;
  assign n12852 = n12830 & n12842;
  assign n12853 = ~n12830 & ~n12842;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = pi260 & ~n12847;
  assign n12856 = pi145 & n12855;
  assign n12857 = pi261 & ~n12846;
  assign n12858 = pi144 & n12857;
  assign n12859 = ~n12856 & ~n12858;
  assign n12860 = ~n12854 & ~n12859;
  assign n12861 = ~n12851 & ~n12860;
  assign n12862 = ~n12550 & n12861;
  assign n12863 = n12550 & ~n12861;
  assign n12864 = ~n12862 & ~n12863;
  assign n12865 = ~pi146 & ~pi259;
  assign n12866 = pi146 & pi259;
  assign n12867 = n10228 & n12866;
  assign n12868 = ~n12865 & ~n12867;
  assign n12869 = ~n10534 & ~n12868;
  assign n12870 = ~pi145 & ~n11690;
  assign n12871 = ~n6503 & ~n12870;
  assign n12872 = pi146 & ~pi259;
  assign n12873 = pi145 & n12872;
  assign n12874 = ~pi146 & pi259;
  assign n12875 = pi258 & n12874;
  assign n12876 = ~n12873 & ~n12875;
  assign n12877 = n10534 & ~n12876;
  assign n12878 = n12871 & ~n12877;
  assign n12879 = ~n12869 & n12878;
  assign n12880 = n11681 & ~n12879;
  assign n12881 = pi258 & n12872;
  assign n12882 = pi145 & n12874;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = ~n10534 & ~n12883;
  assign n12885 = ~pi145 & pi146;
  assign n12886 = pi145 & n12865;
  assign n12887 = ~n12866 & ~n12886;
  assign n12888 = n10534 & ~n12887;
  assign n12889 = ~n12885 & ~n12888;
  assign n12890 = pi258 & ~n12889;
  assign n12891 = pi145 & n1146;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = ~n12884 & n12892;
  assign n12894 = ~n11681 & ~n12893;
  assign n12895 = ~n12880 & ~n12894;
  assign n12896 = pi147 & pi258;
  assign n12897 = ~n12895 & n12896;
  assign n12898 = n12895 & ~n12896;
  assign n12899 = ~n12897 & ~n12898;
  assign n12900 = ~n12864 & ~n12899;
  assign n12901 = n12550 & n12861;
  assign n12902 = ~n12550 & ~n12861;
  assign n12903 = ~n12901 & ~n12902;
  assign n12904 = n12895 & n12896;
  assign n12905 = ~n12895 & ~n12896;
  assign n12906 = ~n12904 & ~n12905;
  assign n12907 = ~n12903 & ~n12906;
  assign n12908 = ~n12900 & ~n12907;
  assign n12909 = ~n12534 & ~n12908;
  assign n12910 = n12510 & ~n12531;
  assign n12911 = ~n12510 & n12531;
  assign n12912 = ~n12910 & ~n12911;
  assign n12913 = ~n12899 & ~n12903;
  assign n12914 = ~n12864 & ~n12906;
  assign n12915 = ~n12913 & ~n12914;
  assign n12916 = ~n12912 & ~n12915;
  assign n12917 = ~n12909 & ~n12916;
  assign n12918 = pi322 & n12917;
  assign n12919 = ~n12504 & ~n12918;
  assign n12920 = n11711 & n12917;
  assign n12921 = n1445 & n12920;
  assign n12922 = ~n12919 & ~n12921;
  assign n12923 = ~n12503 & ~n12922;
  assign n12924 = ~n12494 & n12500;
  assign n12925 = n12494 & ~n12500;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = ~n12504 & n12917;
  assign n12928 = pi322 & n12927;
  assign n12929 = n11711 & ~n12918;
  assign n12930 = pi323 & n12929;
  assign n12931 = ~n12928 & ~n12930;
  assign n12932 = ~n12926 & ~n12931;
  assign n12933 = ~n12923 & ~n12932;
  assign n12934 = n11367 & ~n11731;
  assign n12935 = ~n11369 & ~n11712;
  assign n12936 = n11369 & n11711;
  assign n12937 = pi322 & n12936;
  assign n12938 = ~n12935 & ~n12937;
  assign n12939 = ~n11385 & ~n12938;
  assign n12940 = n11369 & ~n11712;
  assign n12941 = ~n11369 & n11711;
  assign n12942 = pi322 & n12941;
  assign n12943 = ~n12940 & ~n12942;
  assign n12944 = n11384 & ~n12943;
  assign n12945 = pi323 & n12944;
  assign n12946 = ~n12939 & ~n12945;
  assign n12947 = ~n11367 & n11731;
  assign n12948 = ~n12946 & ~n12947;
  assign n12949 = ~n12934 & ~n12948;
  assign n12950 = n12933 & ~n12949;
  assign n12951 = ~n12933 & n12949;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = pi326 & n10561;
  assign n12954 = pi325 & n11366;
  assign n12955 = n12953 & n12954;
  assign n12956 = ~n12953 & ~n12954;
  assign n12957 = ~n12955 & ~n12956;
  assign n12958 = ~n12952 & ~n12957;
  assign n12959 = ~n12933 & ~n12949;
  assign n12960 = n12933 & n12949;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = ~n12953 & n12954;
  assign n12963 = n12953 & ~n12954;
  assign n12964 = ~n12962 & ~n12963;
  assign n12965 = ~n12961 & ~n12964;
  assign n12966 = ~n12958 & ~n12965;
  assign n12967 = ~n12493 & ~n12966;
  assign n12968 = n12470 & n12490;
  assign n12969 = ~n12470 & ~n12490;
  assign n12970 = ~n12968 & ~n12969;
  assign n12971 = ~n12957 & ~n12961;
  assign n12972 = ~n12952 & ~n12964;
  assign n12973 = ~n12971 & ~n12972;
  assign n12974 = ~n12970 & ~n12973;
  assign n12975 = ~n12967 & ~n12974;
  assign n12976 = ~n12466 & n12975;
  assign n12977 = n12466 & ~n12975;
  assign n12978 = ~n12976 & ~n12977;
  assign n12979 = pi329 & n5973;
  assign n12980 = pi328 & n6556;
  assign n12981 = n12979 & n12980;
  assign n12982 = ~n12979 & ~n12980;
  assign n12983 = ~n12981 & ~n12982;
  assign n12984 = ~n12978 & ~n12983;
  assign n12985 = n12466 & n12975;
  assign n12986 = ~n12466 & ~n12975;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~n12979 & n12980;
  assign n12989 = n12979 & ~n12980;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = ~n12987 & ~n12990;
  assign n12992 = ~n12984 & ~n12991;
  assign n12993 = ~n12465 & ~n12992;
  assign n12994 = ~n12449 & n12462;
  assign n12995 = n12449 & ~n12462;
  assign n12996 = ~n12994 & ~n12995;
  assign n12997 = ~n12983 & ~n12987;
  assign n12998 = ~n12978 & ~n12990;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = ~n12996 & ~n12999;
  assign n13001 = ~n12993 & ~n13000;
  assign n13002 = n12445 & n13001;
  assign n13003 = ~n12445 & ~n13001;
  assign n13004 = ~n13002 & ~n13003;
  assign n13005 = n5714 & ~n13004;
  assign n13006 = pi331 & n13005;
  assign n13007 = pi331 & n5714;
  assign n13008 = ~n12445 & n13001;
  assign n13009 = n12445 & ~n13001;
  assign n13010 = ~n13008 & ~n13009;
  assign n13011 = ~n13007 & ~n13010;
  assign n13012 = ~n13006 & ~n13011;
  assign n13013 = ~n12430 & ~n13012;
  assign n13014 = ~n12413 & ~n12427;
  assign n13015 = n12413 & n12427;
  assign n13016 = ~n13014 & ~n13015;
  assign n13017 = n5714 & ~n13010;
  assign n13018 = pi331 & n13017;
  assign n13019 = ~n13004 & ~n13007;
  assign n13020 = ~n13018 & ~n13019;
  assign n13021 = ~n13016 & ~n13020;
  assign n13022 = ~n13013 & ~n13021;
  assign n13023 = ~n11808 & n11812;
  assign n13024 = ~n11804 & ~n11823;
  assign n13025 = n11804 & n11823;
  assign n13026 = ~n13024 & ~n13025;
  assign n13027 = n11808 & ~n11812;
  assign n13028 = ~n13026 & ~n13027;
  assign n13029 = ~n13023 & ~n13028;
  assign n13030 = n13022 & n13029;
  assign n13031 = ~n13022 & ~n13029;
  assign n13032 = ~n13030 & ~n13031;
  assign n13033 = pi333 & n4596;
  assign n13034 = ~n11804 & ~n11818;
  assign n13035 = n11804 & n11818;
  assign n13036 = ~n4596 & ~n13035;
  assign n13037 = ~n13034 & ~n13036;
  assign n13038 = n5257 & ~n13037;
  assign n13039 = ~n5257 & ~n13034;
  assign n13040 = n4596 & n13039;
  assign n13041 = ~n13038 & ~n13040;
  assign n13042 = pi332 & ~n13041;
  assign n13043 = pi332 & n5257;
  assign n13044 = n11804 & ~n13043;
  assign n13045 = n11818 & n13044;
  assign n13046 = ~n13042 & ~n13045;
  assign n13047 = ~n13033 & n13046;
  assign n13048 = n13033 & ~n13046;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = pi334 & n2887;
  assign n13051 = ~n11826 & ~n11848;
  assign n13052 = ~n11855 & n13051;
  assign n13053 = ~n11846 & ~n11848;
  assign n13054 = ~n11811 & n13053;
  assign n13055 = ~n11847 & ~n13054;
  assign n13056 = ~n13052 & n13055;
  assign n13057 = n13050 & ~n13056;
  assign n13058 = ~n13050 & n13056;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = ~n13049 & ~n13059;
  assign n13061 = n13033 & n13046;
  assign n13062 = ~n13033 & ~n13046;
  assign n13063 = ~n13061 & ~n13062;
  assign n13064 = ~n13050 & ~n13056;
  assign n13065 = n13050 & n13056;
  assign n13066 = ~n13064 & ~n13065;
  assign n13067 = ~n13063 & ~n13066;
  assign n13068 = ~n13060 & ~n13067;
  assign n13069 = ~n13032 & ~n13068;
  assign n13070 = n13022 & ~n13029;
  assign n13071 = ~n13022 & n13029;
  assign n13072 = ~n13070 & ~n13071;
  assign n13073 = ~n13059 & ~n13063;
  assign n13074 = ~n13049 & ~n13066;
  assign n13075 = ~n13073 & ~n13074;
  assign n13076 = ~n13072 & ~n13075;
  assign n13077 = ~n13069 & ~n13076;
  assign n13078 = ~n12398 & n13077;
  assign n13079 = n12398 & ~n13077;
  assign n13080 = ~n13078 & ~n13079;
  assign n13081 = pi337 & n1729;
  assign n13082 = n1442 & ~n11865;
  assign n13083 = ~n1729 & ~n13082;
  assign n13084 = pi336 & ~n13083;
  assign n13085 = ~n11866 & ~n13084;
  assign n13086 = pi336 & n2091;
  assign n13087 = n11271 & ~n13086;
  assign n13088 = ~n13085 & n13087;
  assign n13089 = ~n11866 & ~n13082;
  assign n13090 = n1729 & ~n13089;
  assign n13091 = pi336 & n13090;
  assign n13092 = ~n11271 & n13086;
  assign n13093 = ~n13091 & n13092;
  assign n13094 = ~n13088 & ~n13093;
  assign n13095 = ~n12387 & ~n13094;
  assign n13096 = n11271 & n13086;
  assign n13097 = ~n13091 & n13096;
  assign n13098 = ~n11271 & ~n13086;
  assign n13099 = ~n13085 & n13098;
  assign n13100 = ~n13097 & ~n13099;
  assign n13101 = ~n12377 & ~n13100;
  assign n13102 = ~n13086 & n13091;
  assign n13103 = n13085 & n13086;
  assign n13104 = ~n13091 & n13103;
  assign n13105 = ~n13102 & ~n13104;
  assign n13106 = ~n13101 & n13105;
  assign n13107 = ~n13095 & n13106;
  assign n13108 = n13081 & ~n13107;
  assign n13109 = ~n13081 & n13107;
  assign n13110 = ~n13108 & ~n13109;
  assign n13111 = ~n13080 & ~n13110;
  assign n13112 = n12398 & n13077;
  assign n13113 = ~n12398 & ~n13077;
  assign n13114 = ~n13112 & ~n13113;
  assign n13115 = ~n13081 & ~n13107;
  assign n13116 = n13081 & n13107;
  assign n13117 = ~n13115 & ~n13116;
  assign n13118 = ~n13114 & ~n13117;
  assign n13119 = ~n13111 & ~n13118;
  assign n13120 = ~n12397 & ~n13119;
  assign n13121 = ~n12374 & ~n12394;
  assign n13122 = n12374 & n12394;
  assign n13123 = ~n13121 & ~n13122;
  assign n13124 = ~n13110 & ~n13114;
  assign n13125 = ~n13080 & ~n13117;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = ~n13123 & ~n13126;
  assign n13128 = ~n13120 & ~n13127;
  assign n13129 = ~n1256 & ~n11233;
  assign n13130 = pi338 & n13129;
  assign n13131 = n1256 & ~n11229;
  assign n13132 = ~n11232 & n13131;
  assign n13133 = pi338 & ~n13132;
  assign n13134 = ~n13130 & n13133;
  assign n13135 = n11898 & ~n13134;
  assign n13136 = ~n11898 & n13134;
  assign n13137 = ~n13135 & ~n13136;
  assign n13138 = ~n11904 & ~n13137;
  assign n13139 = ~n11903 & ~n13138;
  assign n13140 = ~n13128 & n13139;
  assign n13141 = n13128 & ~n13139;
  assign n13142 = ~n13140 & ~n13141;
  assign n13143 = n11898 & n13133;
  assign n13144 = ~n13130 & ~n13143;
  assign n13145 = n1442 & ~n13144;
  assign n13146 = pi338 & n13145;
  assign n13147 = pi338 & n1442;
  assign n13148 = ~n13143 & ~n13147;
  assign n13149 = ~n13130 & n13148;
  assign n13150 = ~n13146 & ~n13149;
  assign n13151 = ~n1256 & ~n13150;
  assign n13152 = pi339 & n13151;
  assign n13153 = pi339 & ~n1256;
  assign n13154 = ~n13149 & ~n13153;
  assign n13155 = ~n13146 & n13154;
  assign n13156 = ~n13152 & ~n13155;
  assign n13157 = ~n13142 & ~n13156;
  assign n13158 = n13128 & n13139;
  assign n13159 = ~n13128 & ~n13139;
  assign n13160 = ~n13158 & ~n13159;
  assign n13161 = n13150 & n13153;
  assign n13162 = ~n13150 & ~n13153;
  assign n13163 = ~n13161 & ~n13162;
  assign n13164 = ~n13160 & ~n13163;
  assign n13165 = ~n13157 & ~n13164;
  assign n13166 = pi341 & n1156;
  assign n13167 = ~n13165 & ~n13166;
  assign n13168 = pi341 & n13165;
  assign n13169 = n1156 & n13168;
  assign n13170 = ~n13167 & ~n13169;
  assign n13171 = ~n12370 & ~n13170;
  assign n13172 = pi341 & ~n13165;
  assign n13173 = n1156 & n13172;
  assign n13174 = n13165 & ~n13166;
  assign n13175 = ~n13173 & ~n13174;
  assign n13176 = ~n12369 & ~n13175;
  assign n13177 = ~n12358 & n13176;
  assign n13178 = ~n13171 & ~n13177;
  assign n13179 = ~n12350 & ~n13178;
  assign n13180 = n12350 & n13178;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = pi277 & ~n13181;
  assign n13183 = ~n12350 & n13178;
  assign n13184 = n12350 & ~n13178;
  assign n13185 = ~n13183 & ~n13184;
  assign n13186 = ~pi277 & ~n13185;
  assign n13187 = ~n13182 & ~n13186;
  assign n13188 = pi128 & pi302;
  assign n13189 = ~n13187 & n13188;
  assign n13190 = n13187 & ~n13188;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n12348 & ~n13191;
  assign n13193 = ~n12337 & ~n12345;
  assign n13194 = n12337 & n12345;
  assign n13195 = ~n13193 & ~n13194;
  assign n13196 = ~n13187 & ~n13188;
  assign n13197 = n13187 & n13188;
  assign n13198 = ~n13196 & ~n13197;
  assign n13199 = ~n13195 & ~n13198;
  assign n13200 = ~n13192 & ~n13199;
  assign n13201 = ~n831 & ~n13200;
  assign n13202 = ~pi277 & n831;
  assign n13203 = ~n13201 & ~n13202;
  assign n13204 = pi161 & n13203;
  assign n13205 = ~n11955 & ~n13204;
  assign po212 = ~pi160 & ~n13205;
  assign n13207 = pi278 & n831;
  assign n13208 = ~pi277 & ~n13180;
  assign n13209 = ~n13179 & ~n13208;
  assign n13210 = n1442 & n13144;
  assign n13211 = pi338 & n13210;
  assign n13212 = ~n13144 & ~n13147;
  assign n13213 = ~n13211 & ~n13212;
  assign n13214 = ~n13153 & n13213;
  assign n13215 = n13153 & ~n13213;
  assign n13216 = ~n13214 & ~n13215;
  assign n13217 = ~n13160 & ~n13216;
  assign n13218 = n13153 & n13213;
  assign n13219 = ~n13153 & ~n13213;
  assign n13220 = ~n13218 & ~n13219;
  assign n13221 = ~n13142 & ~n13220;
  assign n13222 = ~n12369 & ~n13221;
  assign n13223 = ~n13217 & n13222;
  assign n13224 = ~n12358 & ~n13223;
  assign n13225 = pi340 & ~n1256;
  assign n13226 = n13224 & ~n13225;
  assign n13227 = ~n1256 & ~n13224;
  assign n13228 = pi340 & n13227;
  assign n13229 = ~n13226 & ~n13228;
  assign n13230 = ~n12374 & n12398;
  assign n13231 = n12374 & ~n12398;
  assign n13232 = n13077 & ~n13231;
  assign n13233 = ~n13230 & ~n13232;
  assign n13234 = n12374 & n13077;
  assign n13235 = ~n12374 & ~n13077;
  assign n13236 = ~n13234 & ~n13235;
  assign n13237 = n12398 & ~n13107;
  assign n13238 = ~n12398 & n13107;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = n12394 & ~n13081;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = ~n13236 & n13241;
  assign n13243 = ~n12394 & n13081;
  assign n13244 = n12374 & ~n13077;
  assign n13245 = ~n12374 & n13077;
  assign n13246 = ~n13244 & ~n13245;
  assign n13247 = ~n12398 & ~n13107;
  assign n13248 = n12398 & n13107;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = ~n13240 & ~n13249;
  assign n13251 = ~n13246 & n13250;
  assign n13252 = ~n13243 & ~n13251;
  assign n13253 = ~n13242 & n13252;
  assign n13254 = ~n13233 & n13253;
  assign n13255 = n13233 & ~n13253;
  assign n13256 = ~n13254 & ~n13255;
  assign n13257 = pi335 & n2887;
  assign n13258 = ~n12449 & ~n12975;
  assign n13259 = n12449 & n12975;
  assign n13260 = ~n13258 & ~n13259;
  assign n13261 = ~n12466 & ~n12980;
  assign n13262 = n12466 & n12980;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = ~n13260 & ~n13263;
  assign n13265 = n12449 & ~n12975;
  assign n13266 = ~n12449 & n12975;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = n6556 & ~n12466;
  assign n13269 = pi328 & n13268;
  assign n13270 = n9205 & ~n12980;
  assign n13271 = pi327 & n13270;
  assign n13272 = ~n13269 & ~n13271;
  assign n13273 = ~n13267 & ~n13272;
  assign n13274 = ~n13264 & ~n13273;
  assign n13275 = ~n12462 & n13274;
  assign n13276 = n12462 & ~n13274;
  assign n13277 = ~n13275 & ~n13276;
  assign n13278 = n12413 & ~n12979;
  assign n13279 = ~n13277 & ~n13278;
  assign n13280 = ~n12413 & n12979;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = n12413 & n13001;
  assign n13283 = ~n12413 & ~n13001;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = ~n12445 & ~n13284;
  assign n13286 = ~n12413 & n13001;
  assign n13287 = n12413 & ~n13001;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = n12445 & ~n13288;
  assign n13290 = ~n13285 & ~n13289;
  assign n13291 = n12427 & ~n13007;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = n5714 & ~n12427;
  assign n13294 = pi331 & n13293;
  assign n13295 = ~n13292 & ~n13294;
  assign n13296 = ~n13281 & n13295;
  assign n13297 = n13281 & ~n13295;
  assign n13298 = ~n13296 & ~n13297;
  assign n13299 = pi329 & n6556;
  assign n13300 = ~n12449 & n12466;
  assign n13301 = n12449 & ~n12466;
  assign n13302 = n12975 & ~n13301;
  assign n13303 = ~n13300 & ~n13302;
  assign n13304 = ~n12462 & n12980;
  assign n13305 = n12466 & ~n13267;
  assign n13306 = ~n12466 & ~n13260;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = n12462 & ~n12980;
  assign n13309 = ~n13307 & ~n13308;
  assign n13310 = ~n13304 & ~n13309;
  assign n13311 = ~n13303 & ~n13310;
  assign n13312 = n13303 & n13310;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = n12494 & ~n12949;
  assign n13315 = ~n12500 & ~n12918;
  assign n13316 = n12500 & n12917;
  assign n13317 = pi322 & n13316;
  assign n13318 = ~n13315 & ~n13317;
  assign n13319 = ~n12504 & ~n13318;
  assign n13320 = n12500 & ~n12918;
  assign n13321 = ~n12500 & n12917;
  assign n13322 = pi322 & n13321;
  assign n13323 = ~n13320 & ~n13322;
  assign n13324 = n11711 & ~n13323;
  assign n13325 = pi323 & n13324;
  assign n13326 = ~n13319 & ~n13325;
  assign n13327 = ~n12494 & n12949;
  assign n13328 = ~n13326 & ~n13327;
  assign n13329 = ~n13314 & ~n13328;
  assign n13330 = ~n12470 & n12954;
  assign n13331 = n12470 & ~n12954;
  assign n13332 = ~n12952 & ~n13331;
  assign n13333 = ~n13330 & ~n13332;
  assign n13334 = ~n13329 & n13333;
  assign n13335 = n13329 & ~n13333;
  assign n13336 = ~n13334 & ~n13335;
  assign n13337 = pi324 & n11711;
  assign n13338 = pi323 & n12917;
  assign n13339 = n11711 & ~n12500;
  assign n13340 = pi323 & n13339;
  assign n13341 = n12500 & ~n12504;
  assign n13342 = n12917 & ~n13341;
  assign n13343 = pi322 & n13342;
  assign n13344 = ~n13340 & ~n13343;
  assign n13345 = pi146 & pi260;
  assign n13346 = pi145 & n12537;
  assign n13347 = pi145 & n10534;
  assign n13348 = n11681 & ~n13347;
  assign n13349 = ~n13346 & ~n13348;
  assign n13350 = pi258 & ~n13349;
  assign n13351 = ~pi259 & ~n13350;
  assign n13352 = pi146 & ~n13351;
  assign n13353 = ~n12522 & ~n12542;
  assign n13354 = ~n10534 & ~n13353;
  assign n13355 = ~pi145 & n11681;
  assign n13356 = pi145 & ~pi259;
  assign n13357 = ~n11681 & n13356;
  assign n13358 = ~n12505 & ~n13357;
  assign n13359 = n10534 & ~n13358;
  assign n13360 = ~n13355 & ~n13359;
  assign n13361 = ~n13354 & n13360;
  assign n13362 = pi146 & ~n13361;
  assign n13363 = pi258 & n13362;
  assign n13364 = pi259 & n13363;
  assign n13365 = ~n12510 & n12861;
  assign n13366 = n12510 & ~n12861;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = ~n13364 & ~n13367;
  assign n13369 = n13352 & ~n13368;
  assign n13370 = n13345 & ~n13369;
  assign n13371 = ~n12510 & ~n12861;
  assign n13372 = n12510 & n12861;
  assign n13373 = ~n13371 & ~n13372;
  assign n13374 = ~n13364 & n13373;
  assign n13375 = ~n13345 & ~n13374;
  assign n13376 = n13352 & n13375;
  assign n13377 = ~n13370 & ~n13376;
  assign n13378 = pi142 & pi264;
  assign n13379 = pi139 & pi267;
  assign n13380 = pi136 & pi270;
  assign n13381 = pi134 & pi272;
  assign n13382 = pi273 & ~n12616;
  assign n13383 = pi132 & n13382;
  assign n13384 = ~n12607 & ~n12609;
  assign n13385 = ~n13383 & ~n13384;
  assign n13386 = pi272 & ~n13385;
  assign n13387 = pi133 & n13386;
  assign n13388 = pi132 & pi274;
  assign n13389 = pi131 & pi275;
  assign n13390 = ~n12561 & n12562;
  assign n13391 = pi128 & pi278;
  assign n13392 = pi277 & ~n13391;
  assign n13393 = pi129 & n13392;
  assign n13394 = pi129 & pi277;
  assign n13395 = pi278 & ~n13394;
  assign n13396 = pi128 & n13395;
  assign n13397 = ~n13393 & ~n13396;
  assign n13398 = ~pi276 & ~n13397;
  assign n13399 = ~pi130 & ~n13397;
  assign n13400 = pi276 & n13397;
  assign n13401 = pi130 & n13400;
  assign n13402 = ~n13399 & ~n13401;
  assign n13403 = ~pi129 & ~n13402;
  assign n13404 = ~n13398 & ~n13403;
  assign n13405 = ~n13390 & ~n13404;
  assign n13406 = n12561 & n12562;
  assign n13407 = ~n12561 & ~n12562;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = pi129 & ~n13408;
  assign n13410 = pi276 & n13390;
  assign n13411 = ~n13409 & ~n13410;
  assign n13412 = ~n13397 & ~n13411;
  assign n13413 = pi276 & n12561;
  assign n13414 = ~n12562 & n13397;
  assign n13415 = n13413 & n13414;
  assign n13416 = ~n13412 & ~n13415;
  assign n13417 = pi130 & ~n13416;
  assign n13418 = ~n12562 & ~n13397;
  assign n13419 = n12561 & n13418;
  assign n13420 = n12561 & ~n12562;
  assign n13421 = pi276 & ~n13420;
  assign n13422 = pi129 & n13421;
  assign n13423 = ~n13390 & ~n13422;
  assign n13424 = n13397 & ~n13423;
  assign n13425 = ~n13419 & ~n13424;
  assign n13426 = ~pi130 & ~n13425;
  assign n13427 = n12562 & n13397;
  assign n13428 = ~pi276 & ~n12561;
  assign n13429 = n13427 & n13428;
  assign n13430 = ~n13426 & ~n13429;
  assign n13431 = ~n13417 & n13430;
  assign n13432 = ~n13405 & n13431;
  assign n13433 = ~n13389 & ~n13432;
  assign n13434 = n13389 & n13432;
  assign n13435 = ~n13433 & ~n13434;
  assign n13436 = ~n10277 & ~n11447;
  assign n13437 = ~n11448 & ~n13436;
  assign n13438 = ~n11441 & ~n13437;
  assign n13439 = ~n11445 & ~n13438;
  assign n13440 = ~n12573 & ~n13439;
  assign n13441 = ~n12576 & ~n13440;
  assign n13442 = ~n13435 & ~n13441;
  assign n13443 = ~n13389 & n13432;
  assign n13444 = n13389 & ~n13432;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = ~n13440 & ~n13445;
  assign n13447 = ~n12576 & n13446;
  assign n13448 = ~n13442 & ~n13447;
  assign n13449 = n12551 & n12584;
  assign n13450 = ~n12551 & ~n12584;
  assign n13451 = ~n12590 & ~n13450;
  assign n13452 = ~n13449 & ~n13451;
  assign n13453 = ~n13448 & ~n13452;
  assign n13454 = ~n12587 & ~n13449;
  assign n13455 = ~n12557 & n13454;
  assign n13456 = ~n13450 & ~n13455;
  assign n13457 = n13448 & ~n13456;
  assign n13458 = ~n13453 & ~n13457;
  assign n13459 = ~n13388 & n13458;
  assign n13460 = n13388 & ~n13458;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = pi133 & pi273;
  assign n13463 = n12609 & ~n12614;
  assign n13464 = ~n12615 & ~n13463;
  assign n13465 = n13462 & ~n13464;
  assign n13466 = ~n12609 & ~n12615;
  assign n13467 = ~n12614 & ~n13466;
  assign n13468 = ~n13462 & ~n13467;
  assign n13469 = ~n13465 & ~n13468;
  assign n13470 = ~n13461 & ~n13469;
  assign n13471 = ~n13388 & ~n13458;
  assign n13472 = n13388 & n13458;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = ~n13462 & ~n13464;
  assign n13475 = n13462 & ~n13467;
  assign n13476 = ~n13474 & ~n13475;
  assign n13477 = ~n13473 & ~n13476;
  assign n13478 = ~n13470 & ~n13477;
  assign n13479 = ~n12608 & ~n13384;
  assign n13480 = ~n13383 & n13479;
  assign n13481 = ~n12625 & ~n13480;
  assign n13482 = ~n13478 & ~n13481;
  assign n13483 = ~n13387 & n13482;
  assign n13484 = ~n13387 & ~n13481;
  assign n13485 = n13478 & ~n13484;
  assign n13486 = ~n13483 & ~n13485;
  assign n13487 = ~n13381 & ~n13486;
  assign n13488 = n13478 & ~n13481;
  assign n13489 = ~n13387 & n13488;
  assign n13490 = ~n13478 & ~n13484;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = pi272 & ~n13491;
  assign n13493 = pi134 & n13492;
  assign n13494 = ~n13487 & ~n13493;
  assign n13495 = n12629 & ~n12654;
  assign n13496 = ~n12629 & n12654;
  assign n13497 = ~n12645 & ~n13496;
  assign n13498 = ~n13495 & ~n13497;
  assign n13499 = n13494 & n13498;
  assign n13500 = ~n13494 & ~n13498;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = pi135 & pi271;
  assign n13503 = n12668 & ~n12674;
  assign n13504 = ~n12673 & ~n13503;
  assign n13505 = n13502 & ~n13504;
  assign n13506 = ~n12668 & ~n12673;
  assign n13507 = ~n12674 & ~n13506;
  assign n13508 = ~n13502 & ~n13507;
  assign n13509 = ~n13505 & ~n13508;
  assign n13510 = ~n13501 & ~n13509;
  assign n13511 = n13494 & ~n13498;
  assign n13512 = ~n13494 & n13498;
  assign n13513 = ~n13511 & ~n13512;
  assign n13514 = ~n13502 & ~n13504;
  assign n13515 = n13502 & ~n13507;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = ~n13513 & ~n13516;
  assign n13518 = ~n13510 & ~n13517;
  assign n13519 = ~n13380 & n13518;
  assign n13520 = n13380 & ~n13518;
  assign n13521 = ~n13519 & ~n13520;
  assign n13522 = pi270 & ~n12675;
  assign n13523 = pi135 & n13522;
  assign n13524 = ~n12666 & ~n12668;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = pi269 & ~n13525;
  assign n13527 = pi136 & n13526;
  assign n13528 = pi137 & pi269;
  assign n13529 = ~n12667 & ~n13524;
  assign n13530 = ~n13523 & n13529;
  assign n13531 = ~n12684 & ~n13530;
  assign n13532 = ~n13528 & ~n13531;
  assign n13533 = ~n13527 & n13532;
  assign n13534 = ~n13527 & ~n13531;
  assign n13535 = n13528 & ~n13534;
  assign n13536 = ~n13533 & ~n13535;
  assign n13537 = ~n13521 & ~n13536;
  assign n13538 = ~n13380 & ~n13518;
  assign n13539 = n13380 & n13518;
  assign n13540 = ~n13538 & ~n13539;
  assign n13541 = n13528 & ~n13531;
  assign n13542 = ~n13527 & n13541;
  assign n13543 = ~n13528 & ~n13534;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = ~n13540 & ~n13544;
  assign n13546 = ~n13537 & ~n13545;
  assign n13547 = n12688 & ~n12713;
  assign n13548 = ~n12688 & n12713;
  assign n13549 = ~n12704 & ~n13548;
  assign n13550 = ~n13547 & ~n13549;
  assign n13551 = n13546 & ~n13550;
  assign n13552 = ~n13546 & n13550;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = pi138 & pi268;
  assign n13555 = n12727 & ~n12733;
  assign n13556 = ~n12732 & ~n13555;
  assign n13557 = n13554 & ~n13556;
  assign n13558 = ~n12727 & ~n12732;
  assign n13559 = ~n12733 & ~n13558;
  assign n13560 = ~n13554 & ~n13559;
  assign n13561 = ~n13557 & ~n13560;
  assign n13562 = ~n13553 & ~n13561;
  assign n13563 = n13546 & n13550;
  assign n13564 = ~n13546 & ~n13550;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = ~n13554 & ~n13556;
  assign n13567 = n13554 & ~n13559;
  assign n13568 = ~n13566 & ~n13567;
  assign n13569 = ~n13565 & ~n13568;
  assign n13570 = ~n13562 & ~n13569;
  assign n13571 = ~n13379 & ~n13570;
  assign n13572 = n13379 & n13570;
  assign n13573 = ~n13571 & ~n13572;
  assign n13574 = pi267 & ~n12734;
  assign n13575 = pi138 & n13574;
  assign n13576 = ~n12725 & ~n12727;
  assign n13577 = ~n12726 & ~n13576;
  assign n13578 = ~n13575 & n13577;
  assign n13579 = pi140 & pi266;
  assign n13580 = ~n13575 & ~n13576;
  assign n13581 = pi266 & ~n13580;
  assign n13582 = pi139 & n13581;
  assign n13583 = n12744 & ~n13582;
  assign n13584 = n13579 & ~n13583;
  assign n13585 = ~n13578 & n13584;
  assign n13586 = ~n13578 & ~n13583;
  assign n13587 = ~n13579 & ~n13586;
  assign n13588 = ~n13585 & ~n13587;
  assign n13589 = ~n13573 & ~n13588;
  assign n13590 = ~n13379 & n13570;
  assign n13591 = n13379 & ~n13570;
  assign n13592 = ~n13590 & ~n13591;
  assign n13593 = ~n13579 & ~n13583;
  assign n13594 = ~n13578 & n13593;
  assign n13595 = n13579 & ~n13586;
  assign n13596 = ~n13594 & ~n13595;
  assign n13597 = ~n13592 & ~n13596;
  assign n13598 = ~n13589 & ~n13597;
  assign n13599 = ~n12747 & ~n12748;
  assign n13600 = n12747 & n12748;
  assign n13601 = ~n12767 & ~n13600;
  assign n13602 = ~n13599 & ~n13601;
  assign n13603 = n13598 & n13602;
  assign n13604 = ~n13598 & ~n13602;
  assign n13605 = ~n13603 & ~n13604;
  assign n13606 = pi141 & pi265;
  assign n13607 = n12789 & ~n12795;
  assign n13608 = ~n12794 & ~n13607;
  assign n13609 = n13606 & ~n13608;
  assign n13610 = ~n12789 & ~n12794;
  assign n13611 = ~n12795 & ~n13610;
  assign n13612 = ~n13606 & ~n13611;
  assign n13613 = ~n13609 & ~n13612;
  assign n13614 = ~n13605 & ~n13613;
  assign n13615 = n13598 & ~n13602;
  assign n13616 = ~n13598 & n13602;
  assign n13617 = ~n13615 & ~n13616;
  assign n13618 = ~n13606 & ~n13608;
  assign n13619 = n13606 & ~n13611;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = ~n13617 & ~n13620;
  assign n13622 = ~n13614 & ~n13621;
  assign n13623 = ~n13378 & ~n13622;
  assign n13624 = n13378 & n13622;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = pi264 & ~n12796;
  assign n13627 = pi141 & n13626;
  assign n13628 = ~n12787 & ~n12789;
  assign n13629 = ~n12788 & ~n13628;
  assign n13630 = ~n13627 & n13629;
  assign n13631 = pi143 & pi263;
  assign n13632 = ~n13627 & ~n13628;
  assign n13633 = pi263 & ~n13632;
  assign n13634 = pi142 & n13633;
  assign n13635 = n12808 & ~n13634;
  assign n13636 = n13631 & ~n13635;
  assign n13637 = ~n13630 & n13636;
  assign n13638 = ~n13630 & ~n13635;
  assign n13639 = ~n13631 & ~n13638;
  assign n13640 = ~n13637 & ~n13639;
  assign n13641 = ~n13625 & ~n13640;
  assign n13642 = ~n13378 & n13622;
  assign n13643 = n13378 & ~n13622;
  assign n13644 = ~n13642 & ~n13643;
  assign n13645 = ~n13631 & ~n13635;
  assign n13646 = ~n13630 & n13645;
  assign n13647 = n13631 & ~n13638;
  assign n13648 = ~n13646 & ~n13647;
  assign n13649 = ~n13644 & ~n13648;
  assign n13650 = ~n13641 & ~n13649;
  assign n13651 = ~n12812 & ~n12825;
  assign n13652 = n12812 & n12825;
  assign n13653 = ~n12819 & ~n13652;
  assign n13654 = ~n13651 & ~n13653;
  assign n13655 = n13650 & ~n13654;
  assign n13656 = ~n13650 & n13654;
  assign n13657 = ~n13655 & ~n13656;
  assign n13658 = pi262 & ~n13657;
  assign n13659 = pi144 & n13658;
  assign n13660 = pi144 & pi262;
  assign n13661 = ~n13650 & ~n13654;
  assign n13662 = n13650 & n13654;
  assign n13663 = ~n13661 & ~n13662;
  assign n13664 = ~n13660 & ~n13663;
  assign n13665 = ~n13659 & ~n13664;
  assign n13666 = ~n12842 & n12847;
  assign n13667 = n12842 & ~n12847;
  assign n13668 = ~n12830 & ~n13667;
  assign n13669 = ~n13666 & ~n13668;
  assign n13670 = n13665 & n13669;
  assign n13671 = ~n13665 & ~n13669;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = pi261 & ~n12854;
  assign n13674 = pi144 & n13673;
  assign n13675 = ~n12845 & ~n12847;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = pi260 & ~n13676;
  assign n13678 = pi145 & n13677;
  assign n13679 = pi145 & pi261;
  assign n13680 = ~n12846 & ~n13675;
  assign n13681 = ~n13674 & n13680;
  assign n13682 = n12510 & ~n13681;
  assign n13683 = ~n13679 & ~n13682;
  assign n13684 = ~n13678 & n13683;
  assign n13685 = ~n13678 & ~n13682;
  assign n13686 = n13679 & ~n13685;
  assign n13687 = ~n13684 & ~n13686;
  assign n13688 = ~n13672 & ~n13687;
  assign n13689 = n13665 & ~n13669;
  assign n13690 = ~n13665 & n13669;
  assign n13691 = ~n13689 & ~n13690;
  assign n13692 = n13679 & ~n13682;
  assign n13693 = ~n13678 & n13692;
  assign n13694 = ~n13679 & ~n13685;
  assign n13695 = ~n13693 & ~n13694;
  assign n13696 = ~n13691 & ~n13695;
  assign n13697 = ~n13688 & ~n13696;
  assign n13698 = n13377 & n13697;
  assign n13699 = ~n13377 & ~n13697;
  assign n13700 = ~n13698 & ~n13699;
  assign n13701 = pi148 & pi258;
  assign n13702 = pi147 & pi259;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = n13701 & n13702;
  assign n13705 = ~n13703 & ~n13704;
  assign n13706 = ~n13678 & ~n13681;
  assign n13707 = ~n12510 & n12550;
  assign n13708 = n12510 & ~n12550;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = ~n13706 & ~n13709;
  assign n13711 = ~n12510 & ~n12550;
  assign n13712 = n12510 & n12550;
  assign n13713 = ~n13711 & ~n13712;
  assign n13714 = ~n13681 & ~n13713;
  assign n13715 = ~n13678 & n13714;
  assign n13716 = ~n13710 & ~n13715;
  assign n13717 = pi258 & ~n13716;
  assign n13718 = pi147 & n13717;
  assign n13719 = pi258 & ~n13706;
  assign n13720 = pi147 & n13719;
  assign n13721 = ~n12896 & ~n13681;
  assign n13722 = ~n13678 & n13721;
  assign n13723 = ~n13720 & ~n13722;
  assign n13724 = ~n13713 & ~n13723;
  assign n13725 = n12896 & n13706;
  assign n13726 = ~n12896 & ~n13706;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = ~n13709 & ~n13727;
  assign n13729 = ~n13724 & ~n13728;
  assign n13730 = n13718 & ~n13729;
  assign n13731 = ~n13718 & n13729;
  assign n13732 = ~n13730 & ~n13731;
  assign n13733 = ~n13705 & ~n13732;
  assign n13734 = n13701 & ~n13702;
  assign n13735 = ~n13701 & n13702;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = ~n13718 & ~n13729;
  assign n13738 = n13718 & n13729;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = ~n13736 & ~n13739;
  assign n13741 = ~n13733 & ~n13740;
  assign n13742 = ~n13700 & ~n13741;
  assign n13743 = n13377 & ~n13697;
  assign n13744 = ~n13377 & n13697;
  assign n13745 = ~n13743 & ~n13744;
  assign n13746 = ~n13732 & ~n13736;
  assign n13747 = ~n13705 & ~n13739;
  assign n13748 = ~n13746 & ~n13747;
  assign n13749 = ~n13745 & ~n13748;
  assign n13750 = ~n13742 & ~n13749;
  assign n13751 = n12531 & ~n13729;
  assign n13752 = ~n12531 & n13729;
  assign n13753 = ~n12895 & ~n13752;
  assign n13754 = ~n13751 & ~n13753;
  assign n13755 = n13750 & ~n13754;
  assign n13756 = ~n13750 & n13754;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = n13344 & ~n13757;
  assign n13759 = pi322 & n13758;
  assign n13760 = ~n13750 & ~n13754;
  assign n13761 = n13750 & n13754;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = pi322 & n13762;
  assign n13764 = ~n13344 & ~n13763;
  assign n13765 = ~n13759 & ~n13764;
  assign n13766 = ~n13338 & ~n13765;
  assign n13767 = ~n13344 & ~n13757;
  assign n13768 = pi322 & n13767;
  assign n13769 = n13344 & ~n13763;
  assign n13770 = ~n13768 & ~n13769;
  assign n13771 = n12917 & ~n13770;
  assign n13772 = pi323 & n13771;
  assign n13773 = ~n13766 & ~n13772;
  assign n13774 = ~n13337 & n13773;
  assign n13775 = n13337 & ~n13773;
  assign n13776 = ~n13774 & ~n13775;
  assign n13777 = pi326 & n11366;
  assign n13778 = pi325 & n11384;
  assign n13779 = n13777 & n13778;
  assign n13780 = ~n13777 & ~n13778;
  assign n13781 = ~n13779 & ~n13780;
  assign n13782 = ~n13776 & ~n13781;
  assign n13783 = n13337 & n13773;
  assign n13784 = ~n13337 & ~n13773;
  assign n13785 = ~n13783 & ~n13784;
  assign n13786 = ~n13777 & n13778;
  assign n13787 = n13777 & ~n13778;
  assign n13788 = ~n13786 & ~n13787;
  assign n13789 = ~n13785 & ~n13788;
  assign n13790 = ~n13782 & ~n13789;
  assign n13791 = ~n13336 & ~n13790;
  assign n13792 = ~n13329 & ~n13333;
  assign n13793 = n13329 & n13333;
  assign n13794 = ~n13792 & ~n13793;
  assign n13795 = ~n13781 & ~n13785;
  assign n13796 = ~n13776 & ~n13788;
  assign n13797 = ~n13795 & ~n13796;
  assign n13798 = ~n13794 & ~n13797;
  assign n13799 = ~n13791 & ~n13798;
  assign n13800 = ~n12470 & n12949;
  assign n13801 = n12470 & ~n12949;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~n12933 & n12954;
  assign n13804 = n12933 & ~n12954;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = n12490 & ~n12953;
  assign n13807 = ~n13805 & ~n13806;
  assign n13808 = ~n13802 & n13807;
  assign n13809 = ~n12490 & n12953;
  assign n13810 = ~n12470 & ~n12949;
  assign n13811 = n12470 & n12949;
  assign n13812 = ~n13810 & ~n13811;
  assign n13813 = n12933 & n12954;
  assign n13814 = ~n12933 & ~n12954;
  assign n13815 = ~n13813 & ~n13814;
  assign n13816 = ~n13806 & ~n13815;
  assign n13817 = ~n13812 & n13816;
  assign n13818 = ~n13809 & ~n13817;
  assign n13819 = ~n13808 & n13818;
  assign n13820 = n13799 & n13819;
  assign n13821 = ~n13799 & ~n13819;
  assign n13822 = ~n13820 & ~n13821;
  assign n13823 = pi328 & n9205;
  assign n13824 = pi327 & n10561;
  assign n13825 = n13823 & n13824;
  assign n13826 = ~n13823 & ~n13824;
  assign n13827 = ~n13825 & ~n13826;
  assign n13828 = ~n13822 & ~n13827;
  assign n13829 = ~n13799 & n13819;
  assign n13830 = n13799 & ~n13819;
  assign n13831 = ~n13829 & ~n13830;
  assign n13832 = ~n13823 & n13824;
  assign n13833 = n13823 & ~n13824;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = ~n13831 & ~n13834;
  assign n13836 = ~n13828 & ~n13835;
  assign n13837 = ~n13313 & ~n13836;
  assign n13838 = ~n13303 & n13310;
  assign n13839 = n13303 & ~n13310;
  assign n13840 = ~n13838 & ~n13839;
  assign n13841 = ~n13827 & ~n13831;
  assign n13842 = ~n13822 & ~n13834;
  assign n13843 = ~n13841 & ~n13842;
  assign n13844 = ~n13840 & ~n13843;
  assign n13845 = ~n13837 & ~n13844;
  assign n13846 = ~n13299 & n13845;
  assign n13847 = n13299 & ~n13845;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = pi331 & n5732;
  assign n13850 = pi330 & n12439;
  assign n13851 = ~n12420 & ~n12432;
  assign n13852 = ~n13850 & ~n13851;
  assign n13853 = ~pi330 & ~n13852;
  assign n13854 = pi330 & n5732;
  assign n13855 = n13852 & ~n13854;
  assign n13856 = ~n5973 & ~n13855;
  assign n13857 = ~n13853 & ~n13856;
  assign n13858 = ~n13288 & ~n13857;
  assign n13859 = ~n5973 & ~n13852;
  assign n13860 = n5732 & n13859;
  assign n13861 = ~n5732 & n13852;
  assign n13862 = n5732 & ~n13852;
  assign n13863 = ~n13284 & ~n13862;
  assign n13864 = ~n13861 & ~n13863;
  assign n13865 = n5973 & ~n13864;
  assign n13866 = ~n13860 & ~n13865;
  assign n13867 = pi330 & ~n13866;
  assign n13868 = ~n13858 & ~n13867;
  assign n13869 = n13849 & ~n13868;
  assign n13870 = ~n13849 & n13868;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13848 & ~n13871;
  assign n13873 = n13299 & n13845;
  assign n13874 = ~n13299 & ~n13845;
  assign n13875 = ~n13873 & ~n13874;
  assign n13876 = ~n13849 & ~n13868;
  assign n13877 = n13849 & n13868;
  assign n13878 = ~n13876 & ~n13877;
  assign n13879 = ~n13875 & ~n13878;
  assign n13880 = ~n13872 & ~n13879;
  assign n13881 = ~n13298 & ~n13880;
  assign n13882 = ~n13281 & ~n13295;
  assign n13883 = n13281 & n13295;
  assign n13884 = ~n13882 & ~n13883;
  assign n13885 = ~n13871 & ~n13875;
  assign n13886 = ~n13848 & ~n13878;
  assign n13887 = ~n13885 & ~n13886;
  assign n13888 = ~n13884 & ~n13887;
  assign n13889 = ~n13881 & ~n13888;
  assign n13890 = ~n13029 & n13033;
  assign n13891 = ~n13022 & ~n13046;
  assign n13892 = n13022 & n13046;
  assign n13893 = ~n13891 & ~n13892;
  assign n13894 = n13029 & ~n13033;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = ~n13890 & ~n13895;
  assign n13897 = n13889 & n13896;
  assign n13898 = ~n13889 & ~n13896;
  assign n13899 = ~n13897 & ~n13898;
  assign n13900 = pi333 & n5257;
  assign n13901 = n4596 & ~n13034;
  assign n13902 = pi332 & n13901;
  assign n13903 = ~n13035 & ~n13902;
  assign n13904 = ~n13022 & n13903;
  assign n13905 = n13022 & ~n13903;
  assign n13906 = ~n5257 & ~n13905;
  assign n13907 = ~n13904 & ~n13906;
  assign n13908 = n5714 & ~n13907;
  assign n13909 = ~n5714 & ~n13904;
  assign n13910 = n5257 & n13909;
  assign n13911 = ~n13908 & ~n13910;
  assign n13912 = pi332 & ~n13911;
  assign n13913 = pi332 & n5714;
  assign n13914 = n13022 & ~n13913;
  assign n13915 = ~n13903 & n13914;
  assign n13916 = ~n13912 & ~n13915;
  assign n13917 = ~n13900 & n13916;
  assign n13918 = n13900 & ~n13916;
  assign n13919 = ~n13917 & ~n13918;
  assign n13920 = pi334 & n4596;
  assign n13921 = ~n13049 & ~n13065;
  assign n13922 = ~n13072 & n13921;
  assign n13923 = ~n13063 & ~n13065;
  assign n13924 = ~n13032 & n13923;
  assign n13925 = ~n13064 & ~n13924;
  assign n13926 = ~n13922 & n13925;
  assign n13927 = n13920 & ~n13926;
  assign n13928 = ~n13920 & n13926;
  assign n13929 = ~n13927 & ~n13928;
  assign n13930 = ~n13919 & ~n13929;
  assign n13931 = n13900 & n13916;
  assign n13932 = ~n13900 & ~n13916;
  assign n13933 = ~n13931 & ~n13932;
  assign n13934 = ~n13920 & ~n13926;
  assign n13935 = n13920 & n13926;
  assign n13936 = ~n13934 & ~n13935;
  assign n13937 = ~n13933 & ~n13936;
  assign n13938 = ~n13930 & ~n13937;
  assign n13939 = ~n13899 & ~n13938;
  assign n13940 = n13889 & ~n13896;
  assign n13941 = ~n13889 & n13896;
  assign n13942 = ~n13940 & ~n13941;
  assign n13943 = ~n13929 & ~n13933;
  assign n13944 = ~n13919 & ~n13936;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = ~n13942 & ~n13945;
  assign n13947 = ~n13939 & ~n13946;
  assign n13948 = ~n13257 & n13947;
  assign n13949 = n13257 & ~n13947;
  assign n13950 = ~n13948 & ~n13949;
  assign n13951 = pi337 & n2091;
  assign n13952 = pi336 & n2464;
  assign n13953 = n2091 & ~n12377;
  assign n13954 = pi335 & n13953;
  assign n13955 = ~n11271 & ~n12387;
  assign n13956 = ~n13085 & ~n13955;
  assign n13957 = ~n13954 & n13956;
  assign n13958 = ~n13091 & ~n13957;
  assign n13959 = ~n13086 & n13958;
  assign n13960 = ~n13952 & ~n13959;
  assign n13961 = n12398 & n13960;
  assign n13962 = n13086 & ~n13958;
  assign n13963 = n13952 & ~n13962;
  assign n13964 = ~n12398 & n13963;
  assign n13965 = ~n13961 & ~n13964;
  assign n13966 = ~n13246 & ~n13965;
  assign n13967 = n12398 & n13963;
  assign n13968 = ~n12398 & n13960;
  assign n13969 = ~n13967 & ~n13968;
  assign n13970 = ~n13236 & ~n13969;
  assign n13971 = ~n13952 & ~n13958;
  assign n13972 = n13086 & n13971;
  assign n13973 = n13952 & n13958;
  assign n13974 = ~n13086 & n13973;
  assign n13975 = ~n13972 & ~n13974;
  assign n13976 = ~n13970 & n13975;
  assign n13977 = ~n13966 & n13976;
  assign n13978 = n13951 & ~n13977;
  assign n13979 = ~n13951 & n13977;
  assign n13980 = ~n13978 & ~n13979;
  assign n13981 = ~n13950 & ~n13980;
  assign n13982 = n13257 & n13947;
  assign n13983 = ~n13257 & ~n13947;
  assign n13984 = ~n13982 & ~n13983;
  assign n13985 = ~n13951 & ~n13977;
  assign n13986 = n13951 & n13977;
  assign n13987 = ~n13985 & ~n13986;
  assign n13988 = ~n13984 & ~n13987;
  assign n13989 = ~n13981 & ~n13988;
  assign n13990 = ~n13256 & ~n13989;
  assign n13991 = ~n13233 & ~n13253;
  assign n13992 = n13233 & n13253;
  assign n13993 = ~n13991 & ~n13992;
  assign n13994 = ~n13980 & ~n13984;
  assign n13995 = ~n13950 & ~n13987;
  assign n13996 = ~n13994 & ~n13995;
  assign n13997 = ~n13993 & ~n13996;
  assign n13998 = ~n13990 & ~n13997;
  assign n13999 = ~n13139 & n13153;
  assign n14000 = n13139 & ~n13153;
  assign n14001 = n13128 & ~n13150;
  assign n14002 = ~n13128 & n13150;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = ~n14000 & ~n14003;
  assign n14005 = ~n13999 & ~n14004;
  assign n14006 = n13998 & n14005;
  assign n14007 = ~n13998 & ~n14005;
  assign n14008 = ~n14006 & ~n14007;
  assign n14009 = pi339 & n1442;
  assign n14010 = n13128 & ~n13149;
  assign n14011 = ~n13146 & ~n14010;
  assign n14012 = ~n14009 & ~n14011;
  assign n14013 = n14009 & n14011;
  assign n14014 = ~n14012 & ~n14013;
  assign n14015 = n1729 & ~n14014;
  assign n14016 = pi338 & n14015;
  assign n14017 = pi338 & n1729;
  assign n14018 = n14009 & ~n14011;
  assign n14019 = ~n14009 & n14011;
  assign n14020 = ~n14018 & ~n14019;
  assign n14021 = ~n14017 & ~n14020;
  assign n14022 = ~n14016 & ~n14021;
  assign n14023 = ~n14008 & ~n14022;
  assign n14024 = n13998 & ~n14005;
  assign n14025 = ~n13998 & n14005;
  assign n14026 = ~n14024 & ~n14025;
  assign n14027 = n1729 & ~n14020;
  assign n14028 = pi338 & n14027;
  assign n14029 = ~n14014 & ~n14017;
  assign n14030 = ~n14028 & ~n14029;
  assign n14031 = ~n14026 & ~n14030;
  assign n14032 = ~n14023 & ~n14031;
  assign n14033 = n13229 & n14032;
  assign n14034 = ~n13229 & ~n14032;
  assign n14035 = ~n14033 & ~n14034;
  assign n14036 = ~n12369 & n13165;
  assign n14037 = ~n12358 & n14036;
  assign n14038 = ~n12370 & ~n13165;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = pi258 & ~n14039;
  assign n14041 = pi128 & n14040;
  assign n14042 = pi341 & n14041;
  assign n14043 = pi341 & ~n1154;
  assign n14044 = n14042 & n14043;
  assign n14045 = ~n14042 & ~n14043;
  assign n14046 = ~n14044 & ~n14045;
  assign n14047 = n1156 & ~n14046;
  assign n14048 = pi342 & n14047;
  assign n14049 = pi342 & n1156;
  assign n14050 = ~n14042 & n14043;
  assign n14051 = n14042 & ~n14043;
  assign n14052 = ~n14050 & ~n14051;
  assign n14053 = ~n14049 & ~n14052;
  assign n14054 = ~n14048 & ~n14053;
  assign n14055 = ~n14035 & ~n14054;
  assign n14056 = ~n13229 & n14032;
  assign n14057 = n13229 & ~n14032;
  assign n14058 = ~n14056 & ~n14057;
  assign n14059 = n1156 & ~n14052;
  assign n14060 = pi342 & n14059;
  assign n14061 = ~n14046 & ~n14049;
  assign n14062 = ~n14060 & ~n14061;
  assign n14063 = ~n14058 & ~n14062;
  assign n14064 = ~n14055 & ~n14063;
  assign n14065 = pi278 & ~n14064;
  assign n14066 = ~pi278 & n14064;
  assign n14067 = ~n14065 & ~n14066;
  assign n14068 = n13209 & ~n14067;
  assign n14069 = ~n13209 & n14067;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 = pi303 & n1515;
  assign n14072 = ~n12281 & ~n12333;
  assign n14073 = ~n12334 & ~n14072;
  assign n14074 = n14071 & ~n14073;
  assign n14075 = ~n12332 & ~n12334;
  assign n14076 = ~n12333 & ~n14075;
  assign n14077 = ~n14071 & ~n14076;
  assign n14078 = ~n14074 & ~n14077;
  assign n14079 = pi305 & n1533;
  assign n14080 = ~n12259 & ~n12263;
  assign n14081 = ~n12264 & ~n14080;
  assign n14082 = ~n14079 & ~n14081;
  assign n14083 = ~n12256 & ~n12264;
  assign n14084 = ~n11197 & n14083;
  assign n14085 = ~n12263 & ~n14084;
  assign n14086 = n14079 & ~n14085;
  assign n14087 = ~n14082 & ~n14086;
  assign n14088 = ~n11966 & ~n12231;
  assign n14089 = ~n11162 & ~n11167;
  assign n14090 = ~n11163 & ~n14089;
  assign n14091 = n11966 & n12231;
  assign n14092 = ~n14090 & ~n14091;
  assign n14093 = ~n14088 & ~n14092;
  assign n14094 = pi309 & n3012;
  assign n14095 = ~n12210 & ~n12217;
  assign n14096 = ~n12218 & ~n14095;
  assign n14097 = ~n14094 & ~n14096;
  assign n14098 = ~n12213 & ~n12218;
  assign n14099 = ~n12217 & ~n14098;
  assign n14100 = n14094 & ~n14099;
  assign n14101 = ~n14097 & ~n14100;
  assign n14102 = ~n11980 & ~n12172;
  assign n14103 = ~n11091 & ~n11096;
  assign n14104 = ~n11092 & ~n14103;
  assign n14105 = n11980 & n12172;
  assign n14106 = ~n14104 & ~n14105;
  assign n14107 = ~n14102 & ~n14106;
  assign n14108 = pi313 & n5463;
  assign n14109 = ~n12151 & ~n12158;
  assign n14110 = ~n12159 & ~n14109;
  assign n14111 = ~n14108 & ~n14110;
  assign n14112 = ~n12154 & ~n12159;
  assign n14113 = ~n12158 & ~n14112;
  assign n14114 = n14108 & ~n14113;
  assign n14115 = ~n14111 & ~n14114;
  assign n14116 = ~n12118 & ~n12119;
  assign n14117 = n12118 & n12119;
  assign n14118 = ~n11035 & ~n14117;
  assign n14119 = ~n11029 & n14118;
  assign n14120 = ~n14116 & ~n14119;
  assign n14121 = pi316 & n7874;
  assign n14122 = ~n10929 & n10937;
  assign n14123 = ~n10928 & ~n14122;
  assign n14124 = n10929 & ~n10937;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = n12022 & ~n14125;
  assign n14127 = ~n10929 & ~n11985;
  assign n14128 = ~n12048 & ~n14127;
  assign n14129 = ~n12022 & ~n14128;
  assign n14130 = ~n14126 & ~n14129;
  assign n14131 = ~n12065 & ~n14130;
  assign n14132 = ~pi148 & ~n10899;
  assign n14133 = pi147 & n14132;
  assign n14134 = ~pi147 & pi148;
  assign n14135 = pi146 & n14134;
  assign n14136 = ~n14133 & ~n14135;
  assign n14137 = pi145 & ~n14136;
  assign n14138 = pi147 & pi148;
  assign n14139 = ~pi146 & n14138;
  assign n14140 = ~pi148 & n10899;
  assign n14141 = ~pi147 & n14140;
  assign n14142 = ~n14139 & ~n14141;
  assign n14143 = ~pi145 & ~n14142;
  assign n14144 = pi147 & ~pi148;
  assign n14145 = pi148 & ~n10899;
  assign n14146 = ~pi147 & n14145;
  assign n14147 = ~n14144 & ~n14146;
  assign n14148 = pi146 & ~n14147;
  assign n14149 = ~pi147 & ~pi148;
  assign n14150 = pi148 & n10899;
  assign n14151 = pi147 & n14150;
  assign n14152 = ~n14149 & ~n14151;
  assign n14153 = ~pi146 & ~n14152;
  assign n14154 = ~n14148 & ~n14153;
  assign n14155 = ~n14143 & n14154;
  assign n14156 = ~n14137 & n14155;
  assign n14157 = pi321 & n14156;
  assign n14158 = ~n11999 & n12005;
  assign n14159 = n10908 & ~n14158;
  assign n14160 = pi320 & n14159;
  assign n14161 = n11998 & ~n12005;
  assign n14162 = pi321 & n14161;
  assign n14163 = ~n14160 & ~n14162;
  assign n14164 = pi320 & n11998;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = n11998 & n14163;
  assign n14167 = pi320 & n14166;
  assign n14168 = ~n14165 & ~n14167;
  assign n14169 = ~n14157 & ~n14168;
  assign n14170 = n14163 & ~n14164;
  assign n14171 = n11998 & ~n14163;
  assign n14172 = pi320 & n14171;
  assign n14173 = ~n14170 & ~n14172;
  assign n14174 = n14156 & ~n14173;
  assign n14175 = pi321 & n14174;
  assign n14176 = ~n14169 & ~n14175;
  assign n14177 = pi319 & n10908;
  assign n14178 = n14176 & n14177;
  assign n14179 = ~n14176 & ~n14177;
  assign n14180 = ~n14178 & ~n14179;
  assign n14181 = ~n12018 & n12019;
  assign n14182 = n12018 & ~n12019;
  assign n14183 = n10929 & ~n12048;
  assign n14184 = ~n11985 & ~n14183;
  assign n14185 = ~n14182 & ~n14184;
  assign n14186 = ~n14181 & ~n14185;
  assign n14187 = n14180 & ~n14186;
  assign n14188 = ~n14128 & ~n14181;
  assign n14189 = ~n14182 & ~n14188;
  assign n14190 = ~n14180 & ~n14189;
  assign n14191 = ~n14187 & ~n14190;
  assign n14192 = ~pi318 & ~n14191;
  assign n14193 = ~n9815 & ~n14191;
  assign n14194 = n9815 & n14191;
  assign n14195 = pi318 & n14194;
  assign n14196 = ~n14193 & ~n14195;
  assign n14197 = ~n9517 & ~n14196;
  assign n14198 = ~n14192 & ~n14197;
  assign n14199 = ~n14131 & ~n14198;
  assign n14200 = n12065 & n14191;
  assign n14201 = n14130 & n14200;
  assign n14202 = ~n12065 & ~n14191;
  assign n14203 = ~n14130 & n14202;
  assign n14204 = ~n14201 & ~n14203;
  assign n14205 = pi318 & ~n14204;
  assign n14206 = ~n12065 & n14130;
  assign n14207 = n12065 & ~n14130;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~n14191 & ~n14208;
  assign n14210 = n9517 & n14209;
  assign n14211 = ~n14205 & ~n14210;
  assign n14212 = n9815 & ~n14211;
  assign n14213 = n12065 & ~n14191;
  assign n14214 = n14130 & n14213;
  assign n14215 = n12065 & n14130;
  assign n14216 = n9517 & ~n14215;
  assign n14217 = pi318 & n14216;
  assign n14218 = ~n14131 & ~n14217;
  assign n14219 = n14191 & ~n14218;
  assign n14220 = ~n14214 & ~n14219;
  assign n14221 = ~n9815 & ~n14220;
  assign n14222 = ~pi318 & ~n14130;
  assign n14223 = ~n12065 & n14191;
  assign n14224 = n14222 & n14223;
  assign n14225 = ~n14221 & ~n14224;
  assign n14226 = ~n14212 & n14225;
  assign n14227 = ~n14199 & n14226;
  assign n14228 = ~pi317 & ~n14227;
  assign n14229 = ~n9517 & ~n14227;
  assign n14230 = n9517 & n14227;
  assign n14231 = pi317 & n14230;
  assign n14232 = ~n14229 & ~n14231;
  assign n14233 = ~n7874 & ~n14232;
  assign n14234 = ~n14228 & ~n14233;
  assign n14235 = ~n12083 & ~n14234;
  assign n14236 = ~n12073 & n14227;
  assign n14237 = n12068 & n14236;
  assign n14238 = n12073 & ~n14227;
  assign n14239 = ~n12068 & n14238;
  assign n14240 = ~n14237 & ~n14239;
  assign n14241 = pi317 & ~n14240;
  assign n14242 = ~n12076 & ~n14227;
  assign n14243 = n7874 & n14242;
  assign n14244 = ~n14241 & ~n14243;
  assign n14245 = n9517 & ~n14244;
  assign n14246 = ~n12073 & ~n14227;
  assign n14247 = n12068 & n14246;
  assign n14248 = n7874 & ~n12084;
  assign n14249 = pi317 & n14248;
  assign n14250 = ~n12083 & ~n14249;
  assign n14251 = n14227 & ~n14250;
  assign n14252 = ~n14247 & ~n14251;
  assign n14253 = ~n9517 & ~n14252;
  assign n14254 = ~pi317 & ~n12068;
  assign n14255 = n12073 & n14227;
  assign n14256 = n14254 & n14255;
  assign n14257 = ~n14253 & ~n14256;
  assign n14258 = ~n14245 & n14257;
  assign n14259 = ~n14235 & n14258;
  assign n14260 = ~n14121 & ~n14259;
  assign n14261 = n14121 & n14259;
  assign n14262 = ~n14260 & ~n14261;
  assign n14263 = pi315 & n7044;
  assign n14264 = n7874 & ~n12085;
  assign n14265 = pi317 & n14264;
  assign n14266 = ~n12076 & ~n12077;
  assign n14267 = ~n14265 & ~n14266;
  assign n14268 = ~n12100 & ~n14267;
  assign n14269 = n12100 & n14267;
  assign n14270 = n12078 & ~n14269;
  assign n14271 = ~n14268 & ~n14270;
  assign n14272 = n14263 & ~n14271;
  assign n14273 = ~n12078 & ~n14268;
  assign n14274 = ~n14269 & ~n14273;
  assign n14275 = ~n14263 & ~n14274;
  assign n14276 = ~n14272 & ~n14275;
  assign n14277 = ~n14262 & ~n14276;
  assign n14278 = ~n14121 & n14259;
  assign n14279 = n14121 & ~n14259;
  assign n14280 = ~n14278 & ~n14279;
  assign n14281 = ~n14263 & ~n14271;
  assign n14282 = n14263 & ~n14274;
  assign n14283 = ~n14281 & ~n14282;
  assign n14284 = ~n14280 & ~n14283;
  assign n14285 = ~n14277 & ~n14284;
  assign n14286 = n12106 & ~n12109;
  assign n14287 = ~n11017 & n11022;
  assign n14288 = ~n11018 & ~n14287;
  assign n14289 = ~n12106 & n12109;
  assign n14290 = ~n14288 & ~n14289;
  assign n14291 = ~n14286 & ~n14290;
  assign n14292 = ~n14285 & n14291;
  assign n14293 = n14285 & ~n14291;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = n6777 & ~n14294;
  assign n14296 = pi314 & n14295;
  assign n14297 = pi314 & n6777;
  assign n14298 = ~n14293 & ~n14297;
  assign n14299 = ~n14292 & n14298;
  assign n14300 = ~n14296 & ~n14299;
  assign n14301 = ~n14120 & ~n14300;
  assign n14302 = n14120 & ~n14299;
  assign n14303 = ~n14296 & n14302;
  assign n14304 = ~n14301 & ~n14303;
  assign n14305 = n14115 & ~n14304;
  assign n14306 = ~n14115 & n14304;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = pi312 & n4772;
  assign n14309 = pi313 & ~n9912;
  assign n14310 = n12134 & ~n14309;
  assign n14311 = pi313 & ~n12134;
  assign n14312 = n9909 & n14311;
  assign n14313 = ~n14310 & ~n14312;
  assign n14314 = ~n12148 & ~n14313;
  assign n14315 = ~n4772 & n12134;
  assign n14316 = ~n12136 & ~n14315;
  assign n14317 = ~n11037 & ~n14316;
  assign n14318 = n12147 & n14317;
  assign n14319 = n9924 & ~n12134;
  assign n14320 = ~n4086 & ~n11037;
  assign n14321 = n4772 & ~n14320;
  assign n14322 = n12134 & n14321;
  assign n14323 = ~n14319 & ~n14322;
  assign n14324 = pi313 & ~n14323;
  assign n14325 = n11037 & n12158;
  assign n14326 = ~n14324 & ~n14325;
  assign n14327 = ~n12147 & ~n14326;
  assign n14328 = ~n4772 & ~n12134;
  assign n14329 = n4772 & n12134;
  assign n14330 = ~n14328 & ~n14329;
  assign n14331 = n4086 & ~n14330;
  assign n14332 = pi313 & n14331;
  assign n14333 = n11037 & n14332;
  assign n14334 = ~n14327 & ~n14333;
  assign n14335 = ~n14318 & n14334;
  assign n14336 = ~n14314 & n14335;
  assign n14337 = ~n12169 & ~n14336;
  assign n14338 = n12169 & n14336;
  assign n14339 = n12138 & ~n14338;
  assign n14340 = ~n14337 & ~n14339;
  assign n14341 = n14308 & ~n14340;
  assign n14342 = ~n12138 & ~n14337;
  assign n14343 = ~n14338 & ~n14342;
  assign n14344 = ~n14308 & ~n14343;
  assign n14345 = ~n14341 & ~n14344;
  assign n14346 = ~n14307 & ~n14345;
  assign n14347 = n14115 & n14304;
  assign n14348 = ~n14115 & ~n14304;
  assign n14349 = ~n14347 & ~n14348;
  assign n14350 = ~n14308 & ~n14340;
  assign n14351 = n14308 & ~n14343;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = ~n14349 & ~n14352;
  assign n14354 = ~n14346 & ~n14353;
  assign n14355 = n14107 & ~n14354;
  assign n14356 = ~n14107 & n14354;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = n4086 & ~n14357;
  assign n14359 = pi311 & n14358;
  assign n14360 = pi311 & n4086;
  assign n14361 = ~n14107 & ~n14354;
  assign n14362 = n14107 & n14354;
  assign n14363 = ~n14361 & ~n14362;
  assign n14364 = ~n14360 & ~n14363;
  assign n14365 = ~n14359 & ~n14364;
  assign n14366 = ~n12176 & ~n12186;
  assign n14367 = n12176 & n12186;
  assign n14368 = ~n12177 & ~n14367;
  assign n14369 = ~n11103 & n14368;
  assign n14370 = ~n14366 & ~n14369;
  assign n14371 = n14365 & n14370;
  assign n14372 = ~n14365 & ~n14370;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = n3552 & ~n14373;
  assign n14375 = pi310 & n14374;
  assign n14376 = pi310 & n3552;
  assign n14377 = ~n14365 & n14370;
  assign n14378 = n14365 & ~n14370;
  assign n14379 = ~n14377 & ~n14378;
  assign n14380 = ~n14376 & ~n14379;
  assign n14381 = ~n14375 & ~n14380;
  assign n14382 = n14101 & n14381;
  assign n14383 = ~n14101 & ~n14381;
  assign n14384 = ~n14382 & ~n14383;
  assign n14385 = pi308 & n2574;
  assign n14386 = pi309 & ~n9624;
  assign n14387 = n12192 & ~n14386;
  assign n14388 = pi309 & ~n12192;
  assign n14389 = n9627 & n14388;
  assign n14390 = ~n14387 & ~n14389;
  assign n14391 = ~n12207 & ~n14390;
  assign n14392 = ~n2574 & n12192;
  assign n14393 = ~n12218 & ~n14392;
  assign n14394 = n11111 & ~n14393;
  assign n14395 = n12206 & n14394;
  assign n14396 = n9636 & ~n12192;
  assign n14397 = ~n2183 & n11111;
  assign n14398 = n2574 & ~n14397;
  assign n14399 = n12192 & n14398;
  assign n14400 = ~n14396 & ~n14399;
  assign n14401 = pi309 & ~n14400;
  assign n14402 = ~n11111 & n12193;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = ~n12206 & ~n14403;
  assign n14405 = ~n2574 & ~n12192;
  assign n14406 = n2574 & n12192;
  assign n14407 = ~n14405 & ~n14406;
  assign n14408 = n2183 & ~n14407;
  assign n14409 = pi309 & n14408;
  assign n14410 = ~n11111 & n14409;
  assign n14411 = ~n14404 & ~n14410;
  assign n14412 = ~n14395 & n14411;
  assign n14413 = ~n14391 & n14412;
  assign n14414 = n12228 & n14413;
  assign n14415 = ~n12228 & ~n14413;
  assign n14416 = n12196 & ~n14415;
  assign n14417 = ~n14414 & ~n14416;
  assign n14418 = n14385 & ~n14417;
  assign n14419 = ~n12196 & ~n14414;
  assign n14420 = ~n14415 & ~n14419;
  assign n14421 = ~n14385 & ~n14420;
  assign n14422 = ~n14418 & ~n14421;
  assign n14423 = ~n14384 & ~n14422;
  assign n14424 = n14101 & ~n14381;
  assign n14425 = ~n14101 & n14381;
  assign n14426 = ~n14424 & ~n14425;
  assign n14427 = ~n14385 & ~n14417;
  assign n14428 = n14385 & ~n14420;
  assign n14429 = ~n14427 & ~n14428;
  assign n14430 = ~n14426 & ~n14429;
  assign n14431 = ~n14423 & ~n14430;
  assign n14432 = ~n14093 & ~n14431;
  assign n14433 = n14093 & n14431;
  assign n14434 = ~n14432 & ~n14433;
  assign n14435 = n2183 & ~n14434;
  assign n14436 = pi307 & n14435;
  assign n14437 = pi307 & n2183;
  assign n14438 = n14093 & ~n14431;
  assign n14439 = ~n14093 & n14431;
  assign n14440 = ~n14438 & ~n14439;
  assign n14441 = ~n14437 & ~n14440;
  assign n14442 = ~n14436 & ~n14441;
  assign n14443 = n12235 & ~n12245;
  assign n14444 = ~n12235 & n12245;
  assign n14445 = ~n12236 & ~n14444;
  assign n14446 = ~n11177 & n14445;
  assign n14447 = ~n14443 & ~n14446;
  assign n14448 = ~n14442 & n14447;
  assign n14449 = n14442 & ~n14447;
  assign n14450 = ~n14448 & ~n14449;
  assign n14451 = n1840 & ~n14450;
  assign n14452 = pi306 & n14451;
  assign n14453 = pi306 & n1840;
  assign n14454 = n14442 & n14447;
  assign n14455 = ~n14442 & ~n14447;
  assign n14456 = ~n14454 & ~n14455;
  assign n14457 = ~n14453 & ~n14456;
  assign n14458 = ~n14452 & ~n14457;
  assign n14459 = n14087 & n14458;
  assign n14460 = ~n14087 & ~n14458;
  assign n14461 = ~n14459 & ~n14460;
  assign n14462 = pi304 & n1553;
  assign n14463 = ~n12251 & ~n12256;
  assign n14464 = ~n11197 & n14463;
  assign n14465 = n12251 & ~n12259;
  assign n14466 = ~n14464 & ~n14465;
  assign n14467 = ~n11956 & ~n14466;
  assign n14468 = n12251 & ~n12256;
  assign n14469 = ~n11197 & n14468;
  assign n14470 = ~n12251 & ~n12259;
  assign n14471 = ~n14469 & ~n14470;
  assign n14472 = n1553 & ~n14471;
  assign n14473 = pi305 & n14472;
  assign n14474 = ~n14467 & ~n14473;
  assign n14475 = ~n12278 & n14474;
  assign n14476 = n12278 & ~n14474;
  assign n14477 = n12255 & ~n14476;
  assign n14478 = ~n14475 & ~n14477;
  assign n14479 = n14462 & ~n14478;
  assign n14480 = ~n12255 & ~n14475;
  assign n14481 = ~n14476 & ~n14480;
  assign n14482 = ~n14462 & ~n14481;
  assign n14483 = ~n14479 & ~n14482;
  assign n14484 = ~n14461 & ~n14483;
  assign n14485 = n14087 & ~n14458;
  assign n14486 = ~n14087 & n14458;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = ~n14462 & ~n14478;
  assign n14489 = n14462 & ~n14481;
  assign n14490 = ~n14488 & ~n14489;
  assign n14491 = ~n14487 & ~n14490;
  assign n14492 = ~n14484 & ~n14491;
  assign n14493 = ~n14078 & n14492;
  assign n14494 = n14078 & ~n14492;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = pi302 & ~n1568;
  assign n14497 = ~n12337 & n14496;
  assign n14498 = n13188 & n14497;
  assign n14499 = ~n12337 & n13188;
  assign n14500 = ~n14496 & ~n14499;
  assign n14501 = ~n14498 & ~n14500;
  assign n14502 = ~n14495 & ~n14501;
  assign n14503 = ~n14078 & ~n14492;
  assign n14504 = n14078 & n14492;
  assign n14505 = ~n14503 & ~n14504;
  assign n14506 = n14496 & ~n14499;
  assign n14507 = ~n12337 & ~n14496;
  assign n14508 = n13188 & n14507;
  assign n14509 = ~n14506 & ~n14508;
  assign n14510 = ~n14505 & ~n14509;
  assign n14511 = ~n14502 & ~n14510;
  assign n14512 = pi301 & ~n14511;
  assign n14513 = pi128 & n14512;
  assign n14514 = pi128 & pi301;
  assign n14515 = n14511 & ~n14514;
  assign n14516 = ~n14513 & ~n14515;
  assign n14517 = ~n14070 & ~n14516;
  assign n14518 = ~n13209 & ~n14067;
  assign n14519 = n13209 & n14067;
  assign n14520 = ~n14518 & ~n14519;
  assign n14521 = ~n14511 & ~n14514;
  assign n14522 = pi301 & n14511;
  assign n14523 = pi128 & n14522;
  assign n14524 = ~n14521 & ~n14523;
  assign n14525 = ~n14520 & ~n14524;
  assign n14526 = ~n14517 & ~n14525;
  assign n14527 = ~n12345 & ~n13187;
  assign n14528 = n12345 & n13187;
  assign n14529 = n12337 & ~n13188;
  assign n14530 = ~n14499 & ~n14529;
  assign n14531 = ~n14528 & ~n14530;
  assign n14532 = ~n14527 & ~n14531;
  assign n14533 = n14526 & ~n14532;
  assign n14534 = ~n14526 & n14532;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~n831 & ~n14535;
  assign n14537 = ~n13207 & ~n14536;
  assign n14538 = pi161 & ~n14537;
  assign n14539 = pi084 & ~pi161;
  assign n14540 = ~n14538 & ~n14539;
  assign po213 = ~pi160 & ~n14540;
  assign n14542 = ~pi085 & ~pi161;
  assign n14543 = ~pi279 & n831;
  assign n14544 = n14496 & n14499;
  assign n14545 = ~n14500 & ~n14544;
  assign n14546 = ~n14495 & ~n14545;
  assign n14547 = ~n14496 & n14499;
  assign n14548 = ~n14506 & ~n14547;
  assign n14549 = ~n14505 & ~n14548;
  assign n14550 = ~n14546 & ~n14549;
  assign n14551 = pi301 & ~n14550;
  assign n14552 = pi128 & n14551;
  assign n14553 = ~pi128 & pi301;
  assign n14554 = ~n14552 & ~n14553;
  assign n14555 = pi129 & ~n14554;
  assign n14556 = pi301 & ~n14552;
  assign n14557 = n1567 & n14556;
  assign n14558 = ~n14555 & ~n14557;
  assign n14559 = ~n1515 & n14492;
  assign n14560 = n1515 & ~n14492;
  assign n14561 = n14076 & ~n14560;
  assign n14562 = ~n14559 & ~n14561;
  assign n14563 = n1553 & ~n14562;
  assign n14564 = n14076 & n14492;
  assign n14565 = ~n1553 & ~n14564;
  assign n14566 = n1515 & n14565;
  assign n14567 = ~n14563 & ~n14566;
  assign n14568 = pi303 & ~n14567;
  assign n14569 = pi303 & n1553;
  assign n14570 = ~n14492 & ~n14569;
  assign n14571 = ~n14076 & n14570;
  assign n14572 = ~n14568 & ~n14571;
  assign n14573 = pi302 & n1515;
  assign n14574 = n14572 & ~n14573;
  assign n14575 = n1515 & ~n14572;
  assign n14576 = pi302 & n14575;
  assign n14577 = ~n14574 & ~n14576;
  assign n14578 = pi305 & n1840;
  assign n14579 = pi309 & n3552;
  assign n14580 = pi313 & n6777;
  assign n14581 = ~n9815 & n14191;
  assign n14582 = ~n14215 & ~n14581;
  assign n14583 = n9517 & n14582;
  assign n14584 = ~n14131 & n14191;
  assign n14585 = n9815 & ~n14584;
  assign n14586 = ~n14583 & ~n14585;
  assign n14587 = pi318 & ~n14586;
  assign n14588 = ~n14203 & ~n14587;
  assign n14589 = pi148 & ~pi149;
  assign n14590 = pi146 & n14589;
  assign n14591 = pi149 & ~n10899;
  assign n14592 = n14144 & n14591;
  assign n14593 = ~n14590 & ~n14592;
  assign n14594 = pi145 & ~n14593;
  assign n14595 = pi149 & n10899;
  assign n14596 = n14134 & n14595;
  assign n14597 = ~pi148 & ~pi149;
  assign n14598 = ~pi146 & n14597;
  assign n14599 = ~n14596 & ~n14598;
  assign n14600 = ~pi145 & ~n14599;
  assign n14601 = ~pi148 & pi149;
  assign n14602 = pi147 & n14601;
  assign n14603 = ~pi149 & ~n10899;
  assign n14604 = pi148 & n14603;
  assign n14605 = ~n14602 & ~n14604;
  assign n14606 = pi146 & ~n14605;
  assign n14607 = pi148 & pi149;
  assign n14608 = ~pi147 & n14607;
  assign n14609 = ~pi149 & n10899;
  assign n14610 = ~pi148 & n14609;
  assign n14611 = ~n14608 & ~n14610;
  assign n14612 = ~pi146 & ~n14611;
  assign n14613 = ~n14138 & ~n14149;
  assign n14614 = ~pi149 & ~n14613;
  assign n14615 = ~n14612 & ~n14614;
  assign n14616 = ~n14606 & n14615;
  assign n14617 = ~n14600 & n14616;
  assign n14618 = ~n14594 & n14617;
  assign n14619 = pi321 & n14618;
  assign n14620 = ~n14157 & n14163;
  assign n14621 = n11998 & ~n14620;
  assign n14622 = pi320 & n14621;
  assign n14623 = n14156 & ~n14163;
  assign n14624 = pi321 & n14623;
  assign n14625 = ~n14622 & ~n14624;
  assign n14626 = pi320 & n14156;
  assign n14627 = ~n14625 & ~n14626;
  assign n14628 = n14156 & n14625;
  assign n14629 = pi320 & n14628;
  assign n14630 = ~n14627 & ~n14629;
  assign n14631 = ~n14619 & ~n14630;
  assign n14632 = n14625 & ~n14626;
  assign n14633 = n14156 & ~n14625;
  assign n14634 = pi320 & n14633;
  assign n14635 = ~n14632 & ~n14634;
  assign n14636 = n14618 & ~n14635;
  assign n14637 = pi321 & n14636;
  assign n14638 = ~n14631 & ~n14637;
  assign n14639 = pi319 & n11998;
  assign n14640 = n14638 & n14639;
  assign n14641 = ~n14638 & ~n14639;
  assign n14642 = ~n14640 & ~n14641;
  assign n14643 = ~n10937 & ~n14182;
  assign n14644 = ~n9815 & n12018;
  assign n14645 = n9517 & ~n14644;
  assign n14646 = pi319 & n14645;
  assign n14647 = ~n14643 & ~n14646;
  assign n14648 = ~n10928 & ~n14647;
  assign n14649 = n9815 & ~n12018;
  assign n14650 = ~n10937 & n14645;
  assign n14651 = ~n14649 & ~n14650;
  assign n14652 = pi319 & ~n14651;
  assign n14653 = ~n14648 & ~n14652;
  assign n14654 = ~n14176 & ~n14653;
  assign n14655 = n14176 & n14653;
  assign n14656 = pi319 & ~n14655;
  assign n14657 = ~n14654 & ~n14656;
  assign n14658 = n14642 & ~n14657;
  assign n14659 = ~pi319 & ~n14654;
  assign n14660 = ~n14655 & ~n14659;
  assign n14661 = ~n14642 & ~n14660;
  assign n14662 = ~n14658 & ~n14661;
  assign n14663 = n10908 & ~n14662;
  assign n14664 = pi318 & n14663;
  assign n14665 = n10908 & ~n14655;
  assign n14666 = pi319 & n14665;
  assign n14667 = ~n14654 & ~n14666;
  assign n14668 = ~n14642 & ~n14667;
  assign n14669 = n14642 & ~n14660;
  assign n14670 = ~n14668 & ~n14669;
  assign n14671 = ~pi318 & ~n14670;
  assign n14672 = ~n14642 & ~n14653;
  assign n14673 = ~n14176 & n14672;
  assign n14674 = n14642 & ~n14654;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = ~n10908 & ~n14675;
  assign n14677 = ~n14671 & ~n14676;
  assign n14678 = ~n14664 & n14677;
  assign n14679 = ~n14588 & ~n14678;
  assign n14680 = n14588 & n14678;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = n9815 & ~n14681;
  assign n14683 = pi317 & n14682;
  assign n14684 = pi317 & n9815;
  assign n14685 = ~n14680 & ~n14684;
  assign n14686 = ~n14679 & n14685;
  assign n14687 = ~n14683 & ~n14686;
  assign n14688 = ~n9517 & n14227;
  assign n14689 = ~n12084 & ~n14688;
  assign n14690 = n7874 & n14689;
  assign n14691 = ~n12083 & n14227;
  assign n14692 = n9517 & ~n14691;
  assign n14693 = ~n14690 & ~n14692;
  assign n14694 = pi317 & ~n14693;
  assign n14695 = ~n14239 & ~n14694;
  assign n14696 = pi316 & n9517;
  assign n14697 = ~n14695 & ~n14696;
  assign n14698 = n9517 & n14695;
  assign n14699 = pi316 & n14698;
  assign n14700 = ~n14697 & ~n14699;
  assign n14701 = ~n14687 & ~n14700;
  assign n14702 = n14695 & ~n14696;
  assign n14703 = n9517 & ~n14695;
  assign n14704 = pi316 & n14703;
  assign n14705 = ~n14702 & ~n14704;
  assign n14706 = ~n14686 & ~n14705;
  assign n14707 = ~n14683 & n14706;
  assign n14708 = ~n14701 & ~n14707;
  assign n14709 = ~n12100 & ~n14278;
  assign n14710 = ~n7874 & n14259;
  assign n14711 = n7044 & ~n14710;
  assign n14712 = pi316 & n14711;
  assign n14713 = ~n14709 & ~n14712;
  assign n14714 = ~n14267 & ~n14713;
  assign n14715 = n7874 & ~n14259;
  assign n14716 = ~n12100 & n14711;
  assign n14717 = ~n14715 & ~n14716;
  assign n14718 = pi316 & ~n14717;
  assign n14719 = ~n14714 & ~n14718;
  assign n14720 = n14708 & n14719;
  assign n14721 = ~n14708 & ~n14719;
  assign n14722 = ~n14720 & ~n14721;
  assign n14723 = n7874 & ~n14722;
  assign n14724 = pi315 & n14723;
  assign n14725 = pi315 & n7874;
  assign n14726 = ~n14708 & n14719;
  assign n14727 = n14708 & ~n14719;
  assign n14728 = ~n14726 & ~n14727;
  assign n14729 = ~n14725 & ~n14728;
  assign n14730 = ~n14724 & ~n14729;
  assign n14731 = n14263 & ~n14291;
  assign n14732 = ~n7044 & n7874;
  assign n14733 = pi316 & n14259;
  assign n14734 = n14732 & n14733;
  assign n14735 = ~n7044 & ~n7874;
  assign n14736 = pi316 & ~n14735;
  assign n14737 = ~n14259 & ~n14736;
  assign n14738 = ~n14734 & ~n14737;
  assign n14739 = ~n14268 & ~n14738;
  assign n14740 = ~n7874 & ~n14259;
  assign n14741 = ~n14261 & ~n14740;
  assign n14742 = n12100 & ~n14741;
  assign n14743 = n14267 & n14742;
  assign n14744 = ~n7044 & n12100;
  assign n14745 = n7874 & ~n14744;
  assign n14746 = ~n14259 & n14745;
  assign n14747 = n7044 & ~n7874;
  assign n14748 = n14259 & n14747;
  assign n14749 = ~n14746 & ~n14748;
  assign n14750 = pi316 & ~n14749;
  assign n14751 = ~n12100 & n14278;
  assign n14752 = ~n14750 & ~n14751;
  assign n14753 = ~n14267 & ~n14752;
  assign n14754 = ~n14710 & ~n14715;
  assign n14755 = n7044 & ~n14754;
  assign n14756 = pi316 & n14755;
  assign n14757 = ~n12100 & n14756;
  assign n14758 = ~n14753 & ~n14757;
  assign n14759 = ~n14743 & n14758;
  assign n14760 = ~n14739 & n14759;
  assign n14761 = ~n14263 & n14291;
  assign n14762 = ~n14760 & ~n14761;
  assign n14763 = ~n14731 & ~n14762;
  assign n14764 = n14730 & n14763;
  assign n14765 = ~n14730 & ~n14763;
  assign n14766 = ~n14764 & ~n14765;
  assign n14767 = pi314 & n7044;
  assign n14768 = ~n14302 & ~n14767;
  assign n14769 = ~n14296 & n14768;
  assign n14770 = ~n14296 & ~n14302;
  assign n14771 = n14767 & ~n14770;
  assign n14772 = ~n14769 & ~n14771;
  assign n14773 = ~n14766 & ~n14772;
  assign n14774 = n14730 & ~n14763;
  assign n14775 = ~n14730 & n14763;
  assign n14776 = ~n14774 & ~n14775;
  assign n14777 = ~n14302 & n14767;
  assign n14778 = ~n14296 & n14777;
  assign n14779 = ~n14767 & ~n14770;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = ~n14776 & ~n14780;
  assign n14782 = ~n14773 & ~n14781;
  assign n14783 = ~n14580 & n14782;
  assign n14784 = n14580 & ~n14782;
  assign n14785 = ~n14783 & ~n14784;
  assign n14786 = pi312 & n5463;
  assign n14787 = n11037 & ~n12158;
  assign n14788 = n4086 & ~n14328;
  assign n14789 = pi313 & n14788;
  assign n14790 = ~n14787 & ~n14789;
  assign n14791 = ~n12147 & ~n14790;
  assign n14792 = n11037 & n14788;
  assign n14793 = ~n14329 & ~n14792;
  assign n14794 = pi313 & ~n14793;
  assign n14795 = ~n14791 & ~n14794;
  assign n14796 = n14304 & ~n14795;
  assign n14797 = ~n14304 & n14795;
  assign n14798 = n14108 & ~n14797;
  assign n14799 = ~n14796 & ~n14798;
  assign n14800 = n14786 & ~n14799;
  assign n14801 = ~n14108 & ~n14796;
  assign n14802 = ~n14797 & ~n14801;
  assign n14803 = ~n14786 & ~n14802;
  assign n14804 = ~n14800 & ~n14803;
  assign n14805 = ~n14785 & ~n14804;
  assign n14806 = ~n14580 & ~n14782;
  assign n14807 = n14580 & n14782;
  assign n14808 = ~n14806 & ~n14807;
  assign n14809 = ~n14786 & ~n14799;
  assign n14810 = n14786 & ~n14802;
  assign n14811 = ~n14809 & ~n14810;
  assign n14812 = ~n14808 & ~n14811;
  assign n14813 = ~n14805 & ~n14812;
  assign n14814 = n14308 & ~n14349;
  assign n14815 = ~n14308 & n14349;
  assign n14816 = ~n14340 & ~n14815;
  assign n14817 = ~n14814 & ~n14816;
  assign n14818 = n14813 & n14817;
  assign n14819 = ~n14813 & ~n14817;
  assign n14820 = ~n14818 & ~n14819;
  assign n14821 = pi311 & n4772;
  assign n14822 = n14360 & ~n14361;
  assign n14823 = ~n14362 & ~n14822;
  assign n14824 = n14821 & ~n14823;
  assign n14825 = ~n14360 & ~n14362;
  assign n14826 = ~n14361 & ~n14825;
  assign n14827 = ~n14821 & ~n14826;
  assign n14828 = ~n14824 & ~n14827;
  assign n14829 = ~n14820 & ~n14828;
  assign n14830 = n14813 & ~n14817;
  assign n14831 = ~n14813 & n14817;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~n14821 & ~n14823;
  assign n14834 = n14821 & ~n14826;
  assign n14835 = ~n14833 & ~n14834;
  assign n14836 = ~n14832 & ~n14835;
  assign n14837 = ~n14829 & ~n14836;
  assign n14838 = ~pi310 & n14837;
  assign n14839 = ~n4086 & n14837;
  assign n14840 = n4086 & ~n14837;
  assign n14841 = pi310 & n14840;
  assign n14842 = ~n14839 & ~n14841;
  assign n14843 = ~n3552 & ~n14842;
  assign n14844 = ~n14838 & ~n14843;
  assign n14845 = ~n14371 & ~n14844;
  assign n14846 = n14370 & n14837;
  assign n14847 = n14365 & n14846;
  assign n14848 = ~n14370 & ~n14837;
  assign n14849 = ~n14365 & n14848;
  assign n14850 = ~n14847 & ~n14849;
  assign n14851 = pi310 & ~n14850;
  assign n14852 = ~n14379 & n14837;
  assign n14853 = n3552 & n14852;
  assign n14854 = ~n14851 & ~n14853;
  assign n14855 = n4086 & ~n14854;
  assign n14856 = n14370 & ~n14837;
  assign n14857 = ~pi310 & n14365;
  assign n14858 = n14856 & n14857;
  assign n14859 = ~n14370 & n14837;
  assign n14860 = ~n14365 & n14859;
  assign n14861 = n3552 & ~n14372;
  assign n14862 = pi310 & n14861;
  assign n14863 = ~n14371 & ~n14862;
  assign n14864 = ~n14837 & ~n14863;
  assign n14865 = ~n14860 & ~n14864;
  assign n14866 = ~n4086 & ~n14865;
  assign n14867 = ~n14858 & ~n14866;
  assign n14868 = ~n14855 & n14867;
  assign n14869 = ~n14845 & n14868;
  assign n14870 = ~n14579 & ~n14869;
  assign n14871 = n14579 & n14869;
  assign n14872 = ~n14870 & ~n14871;
  assign n14873 = pi308 & n3012;
  assign n14874 = n2183 & ~n14392;
  assign n14875 = pi309 & n14874;
  assign n14876 = ~n11111 & ~n12217;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = ~n12206 & ~n14877;
  assign n14879 = n2574 & ~n12192;
  assign n14880 = ~n11111 & n14874;
  assign n14881 = ~n14879 & ~n14880;
  assign n14882 = pi309 & ~n14881;
  assign n14883 = ~n14878 & ~n14882;
  assign n14884 = ~n14381 & ~n14883;
  assign n14885 = n14381 & n14883;
  assign n14886 = n14094 & ~n14885;
  assign n14887 = ~n14884 & ~n14886;
  assign n14888 = n14873 & ~n14887;
  assign n14889 = ~n14094 & ~n14884;
  assign n14890 = ~n14885 & ~n14889;
  assign n14891 = ~n14873 & ~n14890;
  assign n14892 = ~n14888 & ~n14891;
  assign n14893 = ~n14872 & ~n14892;
  assign n14894 = ~n14579 & n14869;
  assign n14895 = n14579 & ~n14869;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = ~n14873 & ~n14887;
  assign n14898 = n14873 & ~n14890;
  assign n14899 = ~n14897 & ~n14898;
  assign n14900 = ~n14896 & ~n14899;
  assign n14901 = ~n14893 & ~n14900;
  assign n14902 = ~n14384 & ~n14385;
  assign n14903 = n14384 & n14385;
  assign n14904 = ~n14420 & ~n14903;
  assign n14905 = ~n14902 & ~n14904;
  assign n14906 = n14901 & n14905;
  assign n14907 = ~n14901 & ~n14905;
  assign n14908 = ~n14906 & ~n14907;
  assign n14909 = pi307 & n2574;
  assign n14910 = ~n14432 & n14437;
  assign n14911 = ~n14433 & ~n14910;
  assign n14912 = n14909 & ~n14911;
  assign n14913 = ~n14433 & ~n14437;
  assign n14914 = ~n14432 & ~n14913;
  assign n14915 = ~n14909 & ~n14914;
  assign n14916 = ~n14912 & ~n14915;
  assign n14917 = ~n14908 & ~n14916;
  assign n14918 = n14901 & ~n14905;
  assign n14919 = ~n14901 & n14905;
  assign n14920 = ~n14918 & ~n14919;
  assign n14921 = ~n14909 & ~n14911;
  assign n14922 = n14909 & ~n14914;
  assign n14923 = ~n14921 & ~n14922;
  assign n14924 = ~n14920 & ~n14923;
  assign n14925 = ~n14917 & ~n14924;
  assign n14926 = ~pi306 & n14925;
  assign n14927 = ~n2183 & n14925;
  assign n14928 = n2183 & ~n14925;
  assign n14929 = pi306 & n14928;
  assign n14930 = ~n14927 & ~n14929;
  assign n14931 = ~n1840 & ~n14930;
  assign n14932 = ~n14926 & ~n14931;
  assign n14933 = ~n14455 & ~n14932;
  assign n14934 = ~n14447 & n14925;
  assign n14935 = ~n14442 & n14934;
  assign n14936 = n14447 & ~n14925;
  assign n14937 = n14442 & n14936;
  assign n14938 = ~n14935 & ~n14937;
  assign n14939 = pi306 & ~n14938;
  assign n14940 = ~n14450 & n14925;
  assign n14941 = n1840 & n14940;
  assign n14942 = ~n14939 & ~n14941;
  assign n14943 = n2183 & ~n14942;
  assign n14944 = ~pi306 & ~n14442;
  assign n14945 = ~n14447 & ~n14925;
  assign n14946 = n14944 & n14945;
  assign n14947 = n14447 & n14925;
  assign n14948 = n14442 & n14947;
  assign n14949 = n1840 & ~n14454;
  assign n14950 = pi306 & n14949;
  assign n14951 = ~n14455 & ~n14950;
  assign n14952 = ~n14925 & ~n14951;
  assign n14953 = ~n14948 & ~n14952;
  assign n14954 = ~n2183 & ~n14953;
  assign n14955 = ~n14946 & ~n14954;
  assign n14956 = ~n14943 & n14955;
  assign n14957 = ~n14933 & n14956;
  assign n14958 = ~n14578 & n14957;
  assign n14959 = n14578 & ~n14957;
  assign n14960 = ~n14958 & ~n14959;
  assign n14961 = pi304 & n1533;
  assign n14962 = ~n14081 & n14458;
  assign n14963 = n14081 & ~n14458;
  assign n14964 = n14079 & ~n14963;
  assign n14965 = ~n14962 & ~n14964;
  assign n14966 = n14961 & ~n14965;
  assign n14967 = ~n14079 & ~n14962;
  assign n14968 = ~n14963 & ~n14967;
  assign n14969 = ~n14961 & ~n14968;
  assign n14970 = ~n14966 & ~n14969;
  assign n14971 = ~n14960 & ~n14970;
  assign n14972 = ~n14578 & ~n14957;
  assign n14973 = n14578 & n14957;
  assign n14974 = ~n14972 & ~n14973;
  assign n14975 = ~n14961 & ~n14965;
  assign n14976 = n14961 & ~n14968;
  assign n14977 = ~n14975 & ~n14976;
  assign n14978 = ~n14974 & ~n14977;
  assign n14979 = ~n14971 & ~n14978;
  assign n14980 = ~n14462 & ~n14487;
  assign n14981 = n14462 & n14487;
  assign n14982 = ~n14481 & ~n14981;
  assign n14983 = ~n14980 & ~n14982;
  assign n14984 = ~n14979 & ~n14983;
  assign n14985 = n14979 & n14983;
  assign n14986 = ~n14984 & ~n14985;
  assign n14987 = ~n14495 & ~n14500;
  assign n14988 = ~n14498 & ~n14987;
  assign n14989 = ~n14986 & ~n14988;
  assign n14990 = n14986 & n14988;
  assign n14991 = ~n14989 & ~n14990;
  assign n14992 = ~n14577 & ~n14991;
  assign n14993 = n14986 & ~n14988;
  assign n14994 = ~n14986 & n14988;
  assign n14995 = ~n14993 & ~n14994;
  assign n14996 = ~n14572 & ~n14573;
  assign n14997 = n1515 & n14572;
  assign n14998 = pi302 & n14997;
  assign n14999 = ~n14996 & ~n14998;
  assign n15000 = ~n14995 & ~n14999;
  assign n15001 = ~n14992 & ~n15000;
  assign n15002 = ~n14558 & n15001;
  assign n15003 = n14558 & ~n15001;
  assign n15004 = ~n15002 & ~n15003;
  assign n15005 = pi300 & ~n15004;
  assign n15006 = pi128 & n15005;
  assign n15007 = pi128 & pi300;
  assign n15008 = n14558 & n15001;
  assign n15009 = ~n14558 & ~n15001;
  assign n15010 = ~n15008 & ~n15009;
  assign n15011 = ~n15007 & ~n15010;
  assign n15012 = ~n15006 & ~n15011;
  assign n15013 = ~n13209 & ~n14064;
  assign n15014 = n13209 & n14064;
  assign n15015 = ~pi278 & ~n15014;
  assign n15016 = ~n15013 & ~n15015;
  assign n15017 = ~n13233 & ~n13947;
  assign n15018 = n13233 & n13947;
  assign n15019 = ~n15017 & ~n15018;
  assign n15020 = n13257 & ~n13977;
  assign n15021 = ~n13257 & n13977;
  assign n15022 = ~n15020 & ~n15021;
  assign n15023 = n13253 & ~n13951;
  assign n15024 = ~n15022 & ~n15023;
  assign n15025 = ~n15019 & n15024;
  assign n15026 = ~n13253 & n13951;
  assign n15027 = ~n13233 & n13947;
  assign n15028 = n13233 & ~n13947;
  assign n15029 = ~n15027 & ~n15028;
  assign n15030 = ~n13257 & ~n13977;
  assign n15031 = n13257 & n13977;
  assign n15032 = ~n15030 & ~n15031;
  assign n15033 = ~n15023 & ~n15032;
  assign n15034 = ~n15029 & n15033;
  assign n15035 = ~n15026 & ~n15034;
  assign n15036 = ~n15025 & n15035;
  assign n15037 = n14005 & ~n14009;
  assign n15038 = ~n14005 & n14009;
  assign n15039 = ~n13998 & ~n14011;
  assign n15040 = n13998 & n14011;
  assign n15041 = ~n15039 & ~n15040;
  assign n15042 = n1729 & ~n15041;
  assign n15043 = pi338 & n15042;
  assign n15044 = ~n13998 & n14011;
  assign n15045 = n13998 & ~n14011;
  assign n15046 = ~n15044 & ~n15045;
  assign n15047 = ~n14017 & ~n15046;
  assign n15048 = ~n15043 & ~n15047;
  assign n15049 = ~n15038 & ~n15048;
  assign n15050 = ~n15037 & ~n15049;
  assign n15051 = n15036 & n15050;
  assign n15052 = ~n15036 & ~n15050;
  assign n15053 = ~n15051 & ~n15052;
  assign n15054 = pi337 & n2464;
  assign n15055 = n13281 & n13845;
  assign n15056 = ~n13281 & ~n13845;
  assign n15057 = ~n15055 & ~n15056;
  assign n15058 = n13299 & ~n13868;
  assign n15059 = ~n13299 & n13868;
  assign n15060 = ~n15058 & ~n15059;
  assign n15061 = n13295 & ~n13849;
  assign n15062 = ~n15060 & ~n15061;
  assign n15063 = ~n15057 & n15062;
  assign n15064 = ~n13295 & n13849;
  assign n15065 = n13281 & ~n13845;
  assign n15066 = ~n13281 & n13845;
  assign n15067 = ~n15065 & ~n15066;
  assign n15068 = ~n13299 & ~n13868;
  assign n15069 = n13299 & n13868;
  assign n15070 = ~n15068 & ~n15069;
  assign n15071 = ~n15061 & ~n15070;
  assign n15072 = ~n15067 & n15071;
  assign n15073 = ~n15064 & ~n15072;
  assign n15074 = ~n15063 & n15073;
  assign n15075 = ~n13896 & n13900;
  assign n15076 = ~n13889 & ~n13916;
  assign n15077 = n13889 & n13916;
  assign n15078 = ~n15076 & ~n15077;
  assign n15079 = n13896 & ~n13900;
  assign n15080 = ~n15078 & ~n15079;
  assign n15081 = ~n15075 & ~n15080;
  assign n15082 = n15074 & ~n15081;
  assign n15083 = ~n15074 & n15081;
  assign n15084 = ~n15082 & ~n15083;
  assign n15085 = pi331 & n5973;
  assign n15086 = n13303 & ~n13819;
  assign n15087 = ~n13303 & n13819;
  assign n15088 = ~n15086 & ~n15087;
  assign n15089 = ~n13799 & n13824;
  assign n15090 = n13799 & ~n13824;
  assign n15091 = ~n15089 & ~n15090;
  assign n15092 = n13310 & ~n13823;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = ~n15088 & n15093;
  assign n15095 = ~n13310 & n13823;
  assign n15096 = n13303 & n13819;
  assign n15097 = ~n13303 & ~n13819;
  assign n15098 = ~n15096 & ~n15097;
  assign n15099 = n13799 & n13824;
  assign n15100 = ~n13799 & ~n13824;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = ~n15092 & ~n15101;
  assign n15103 = ~n15098 & n15102;
  assign n15104 = ~n15095 & ~n15103;
  assign n15105 = ~n15094 & n15104;
  assign n15106 = ~n13281 & n13299;
  assign n15107 = n13281 & ~n13299;
  assign n15108 = n13845 & ~n15107;
  assign n15109 = ~n15106 & ~n15108;
  assign n15110 = n15105 & ~n15109;
  assign n15111 = ~n15105 & n15109;
  assign n15112 = ~n15110 & ~n15111;
  assign n15113 = pi328 & n10561;
  assign n15114 = n13777 & ~n13819;
  assign n15115 = n11384 & ~n13776;
  assign n15116 = pi325 & n15115;
  assign n15117 = ~n13778 & ~n13785;
  assign n15118 = ~n15116 & ~n15117;
  assign n15119 = ~n13794 & ~n15118;
  assign n15120 = n11384 & ~n13785;
  assign n15121 = pi325 & n15120;
  assign n15122 = ~n13776 & ~n13778;
  assign n15123 = ~n15121 & ~n15122;
  assign n15124 = ~n13336 & ~n15123;
  assign n15125 = ~n15119 & ~n15124;
  assign n15126 = ~n13777 & n13819;
  assign n15127 = ~n15125 & ~n15126;
  assign n15128 = ~n15114 & ~n15127;
  assign n15129 = n13303 & ~n13824;
  assign n15130 = ~n13831 & ~n15129;
  assign n15131 = ~n13303 & n13824;
  assign n15132 = ~n15130 & ~n15131;
  assign n15133 = n15128 & ~n15132;
  assign n15134 = ~n15128 & n15132;
  assign n15135 = ~n15133 & ~n15134;
  assign n15136 = n12917 & ~n13344;
  assign n15137 = pi323 & n15136;
  assign n15138 = ~n13338 & n13344;
  assign n15139 = n13762 & ~n15138;
  assign n15140 = pi322 & n15139;
  assign n15141 = ~n15137 & ~n15140;
  assign n15142 = ~n13329 & n13337;
  assign n15143 = n13329 & ~n13337;
  assign n15144 = ~n13773 & ~n15143;
  assign n15145 = ~n15142 & ~n15144;
  assign n15146 = ~n15141 & n15145;
  assign n15147 = n15141 & ~n15145;
  assign n15148 = ~n15146 & ~n15147;
  assign n15149 = pi323 & n13762;
  assign n15150 = n13702 & n13718;
  assign n15151 = ~n13702 & ~n13718;
  assign n15152 = ~n15150 & ~n15151;
  assign n15153 = pi258 & ~n15152;
  assign n15154 = pi148 & n15153;
  assign n15155 = n13702 & ~n13718;
  assign n15156 = ~n13702 & n13718;
  assign n15157 = ~n15155 & ~n15156;
  assign n15158 = ~n13701 & ~n15157;
  assign n15159 = ~n15154 & ~n15158;
  assign n15160 = ~n13745 & ~n15159;
  assign n15161 = pi258 & ~n15157;
  assign n15162 = pi148 & n15161;
  assign n15163 = ~n13701 & ~n15152;
  assign n15164 = ~n15162 & ~n15163;
  assign n15165 = ~n13700 & ~n15164;
  assign n15166 = ~n15160 & ~n15165;
  assign n15167 = ~n13432 & ~n13441;
  assign n15168 = n13432 & ~n13440;
  assign n15169 = ~n12576 & n15168;
  assign n15170 = ~n15167 & ~n15169;
  assign n15171 = n13389 & ~n15170;
  assign n15172 = n13432 & ~n13441;
  assign n15173 = ~n13432 & ~n13440;
  assign n15174 = ~n12576 & n15173;
  assign n15175 = ~n15172 & ~n15174;
  assign n15176 = ~n13389 & ~n15175;
  assign n15177 = ~n13452 & ~n15176;
  assign n15178 = ~n15171 & ~n15177;
  assign n15179 = pi129 & pi278;
  assign n15180 = pi128 & pi279;
  assign n15181 = ~n15179 & ~n15180;
  assign n15182 = pi278 & n1175;
  assign n15183 = pi279 & n15182;
  assign n15184 = ~n15181 & ~n15183;
  assign n15185 = pi129 & n13391;
  assign n15186 = ~n12562 & ~n12565;
  assign n15187 = ~n12561 & ~n15186;
  assign n15188 = n12562 & n12565;
  assign n15189 = ~n15187 & ~n15188;
  assign n15190 = ~pi129 & ~n13391;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = ~n15185 & ~n15191;
  assign n15193 = ~n15184 & ~n15192;
  assign n15194 = ~n15185 & n15189;
  assign n15195 = ~n15190 & ~n15194;
  assign n15196 = n15184 & ~n15195;
  assign n15197 = ~n15193 & ~n15196;
  assign n15198 = pi277 & ~n15197;
  assign n15199 = pi130 & n15198;
  assign n15200 = n13391 & ~n15189;
  assign n15201 = ~n13391 & n15189;
  assign n15202 = pi129 & ~n15201;
  assign n15203 = pi277 & n15202;
  assign n15204 = ~n15200 & ~n15203;
  assign n15205 = n15184 & ~n15204;
  assign n15206 = ~n15184 & ~n15195;
  assign n15207 = ~n15205 & ~n15206;
  assign n15208 = ~pi130 & ~n15207;
  assign n15209 = ~n15184 & ~n15200;
  assign n15210 = n13391 & n15184;
  assign n15211 = ~n15189 & n15210;
  assign n15212 = ~n15209 & ~n15211;
  assign n15213 = ~pi277 & ~n15212;
  assign n15214 = ~n15208 & ~n15213;
  assign n15215 = ~n13397 & ~n13423;
  assign n15216 = ~pi129 & ~n13390;
  assign n15217 = ~n13420 & ~n15216;
  assign n15218 = n13397 & ~n15217;
  assign n15219 = ~n15215 & ~n15218;
  assign n15220 = ~pi130 & ~n15219;
  assign n15221 = ~n13390 & n13397;
  assign n15222 = n12562 & ~n13397;
  assign n15223 = ~n12561 & n15222;
  assign n15224 = ~n15221 & ~n15223;
  assign n15225 = ~pi276 & ~n15224;
  assign n15226 = ~n15220 & ~n15225;
  assign n15227 = pi129 & ~n13420;
  assign n15228 = ~n13390 & ~n15227;
  assign n15229 = n13397 & ~n15228;
  assign n15230 = ~n13397 & ~n15217;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = pi276 & ~n15231;
  assign n15233 = pi130 & n15232;
  assign n15234 = ~n13441 & ~n15233;
  assign n15235 = n15226 & ~n15234;
  assign n15236 = n15214 & ~n15235;
  assign n15237 = ~n15199 & n15236;
  assign n15238 = ~n15199 & n15214;
  assign n15239 = n15235 & ~n15238;
  assign n15240 = ~n15237 & ~n15239;
  assign n15241 = pi276 & ~n15240;
  assign n15242 = pi131 & n15241;
  assign n15243 = pi131 & pi276;
  assign n15244 = ~n15237 & ~n15243;
  assign n15245 = ~n15239 & n15244;
  assign n15246 = ~n15242 & ~n15245;
  assign n15247 = ~n15178 & ~n15246;
  assign n15248 = n15178 & n15246;
  assign n15249 = ~n15247 & ~n15248;
  assign n15250 = pi275 & ~n15249;
  assign n15251 = pi132 & n15250;
  assign n15252 = pi132 & pi275;
  assign n15253 = ~n15248 & ~n15252;
  assign n15254 = ~n15247 & n15253;
  assign n15255 = ~n15251 & ~n15254;
  assign n15256 = pi274 & n13458;
  assign n15257 = ~pi274 & ~n13458;
  assign n15258 = pi273 & ~n15257;
  assign n15259 = ~n12604 & n15258;
  assign n15260 = ~n15256 & ~n15259;
  assign n15261 = pi132 & ~n15260;
  assign n15262 = ~n12604 & ~n13471;
  assign n15263 = pi132 & n15258;
  assign n15264 = ~n15262 & ~n15263;
  assign n15265 = n12600 & ~n15264;
  assign n15266 = ~n15261 & ~n15265;
  assign n15267 = pi133 & pi274;
  assign n15268 = ~n15266 & ~n15267;
  assign n15269 = pi274 & n15266;
  assign n15270 = pi133 & n15269;
  assign n15271 = ~n15268 & ~n15270;
  assign n15272 = ~n15255 & ~n15271;
  assign n15273 = pi274 & ~n15266;
  assign n15274 = pi133 & n15273;
  assign n15275 = n15266 & ~n15267;
  assign n15276 = ~n15274 & ~n15275;
  assign n15277 = ~n15254 & ~n15276;
  assign n15278 = ~n15251 & n15277;
  assign n15279 = ~n15272 & ~n15278;
  assign n15280 = ~pi273 & ~pi274;
  assign n15281 = pi132 & ~n15280;
  assign n15282 = ~n13458 & ~n15281;
  assign n15283 = ~pi273 & pi274;
  assign n15284 = pi132 & n13458;
  assign n15285 = n15283 & n15284;
  assign n15286 = ~n15282 & ~n15285;
  assign n15287 = ~n12615 & ~n15286;
  assign n15288 = ~n13472 & ~n15257;
  assign n15289 = n12604 & ~n15288;
  assign n15290 = ~n12600 & n15289;
  assign n15291 = pi274 & ~n13458;
  assign n15292 = ~pi274 & n13458;
  assign n15293 = ~n15291 & ~n15292;
  assign n15294 = pi273 & ~n15293;
  assign n15295 = pi132 & n15294;
  assign n15296 = ~n12604 & n15295;
  assign n15297 = ~pi273 & n12604;
  assign n15298 = pi274 & ~n15297;
  assign n15299 = ~n13458 & n15298;
  assign n15300 = pi273 & ~pi274;
  assign n15301 = n13458 & n15300;
  assign n15302 = ~n15299 & ~n15301;
  assign n15303 = pi132 & ~n15302;
  assign n15304 = ~n12604 & n13459;
  assign n15305 = ~n15303 & ~n15304;
  assign n15306 = n12600 & ~n15305;
  assign n15307 = ~n15296 & ~n15306;
  assign n15308 = ~n15290 & n15307;
  assign n15309 = ~n15287 & n15308;
  assign n15310 = n13462 & n15309;
  assign n15311 = ~n13462 & ~n15309;
  assign n15312 = ~n13484 & ~n15311;
  assign n15313 = ~n15310 & ~n15312;
  assign n15314 = n15279 & n15313;
  assign n15315 = ~n15279 & ~n15313;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = pi134 & pi273;
  assign n15318 = ~n13486 & ~n13498;
  assign n15319 = n13486 & n13498;
  assign n15320 = n13381 & ~n15319;
  assign n15321 = ~n15318 & ~n15320;
  assign n15322 = n15317 & ~n15321;
  assign n15323 = ~n13381 & ~n15318;
  assign n15324 = ~n15319 & ~n15323;
  assign n15325 = ~n15317 & ~n15324;
  assign n15326 = ~n15322 & ~n15325;
  assign n15327 = ~n15316 & ~n15326;
  assign n15328 = n15279 & ~n15313;
  assign n15329 = ~n15279 & n15313;
  assign n15330 = ~n15328 & ~n15329;
  assign n15331 = ~n15317 & ~n15321;
  assign n15332 = n15317 & ~n15324;
  assign n15333 = ~n15331 & ~n15332;
  assign n15334 = ~n15330 & ~n15333;
  assign n15335 = ~n15327 & ~n15334;
  assign n15336 = ~n13501 & ~n13502;
  assign n15337 = n13501 & n13502;
  assign n15338 = ~n13507 & ~n15337;
  assign n15339 = ~n15336 & ~n15338;
  assign n15340 = ~n15335 & n15339;
  assign n15341 = n15335 & ~n15339;
  assign n15342 = ~n15340 & ~n15341;
  assign n15343 = pi136 & pi271;
  assign n15344 = pi135 & pi272;
  assign n15345 = n15343 & n15344;
  assign n15346 = ~n15343 & ~n15344;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = ~n15342 & ~n15347;
  assign n15349 = n15335 & n15339;
  assign n15350 = ~n15335 & ~n15339;
  assign n15351 = ~n15349 & ~n15350;
  assign n15352 = pi271 & ~n15344;
  assign n15353 = pi136 & n15352;
  assign n15354 = pi272 & ~n15343;
  assign n15355 = pi135 & n15354;
  assign n15356 = ~n15353 & ~n15355;
  assign n15357 = ~n15351 & ~n15356;
  assign n15358 = ~n15348 & ~n15357;
  assign n15359 = ~n13534 & ~n13538;
  assign n15360 = ~n13539 & ~n15359;
  assign n15361 = n15358 & n15360;
  assign n15362 = ~n15358 & ~n15360;
  assign n15363 = ~n15361 & ~n15362;
  assign n15364 = pi137 & pi270;
  assign n15365 = n13518 & ~n13531;
  assign n15366 = ~n13527 & n15365;
  assign n15367 = ~n13518 & ~n13534;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = ~n13380 & ~n15368;
  assign n15370 = ~n13518 & ~n13531;
  assign n15371 = ~n13527 & n15370;
  assign n15372 = n13518 & ~n13534;
  assign n15373 = ~n15371 & ~n15372;
  assign n15374 = pi270 & ~n15373;
  assign n15375 = pi136 & n15374;
  assign n15376 = ~n15369 & ~n15375;
  assign n15377 = ~n13550 & ~n15376;
  assign n15378 = n13550 & n15376;
  assign n15379 = n13528 & ~n15378;
  assign n15380 = ~n15377 & ~n15379;
  assign n15381 = n15364 & ~n15380;
  assign n15382 = ~n13528 & ~n15377;
  assign n15383 = ~n15378 & ~n15382;
  assign n15384 = ~n15364 & ~n15383;
  assign n15385 = ~n15381 & ~n15384;
  assign n15386 = ~n15363 & ~n15385;
  assign n15387 = n15358 & ~n15360;
  assign n15388 = ~n15358 & n15360;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = ~n15364 & ~n15380;
  assign n15391 = n15364 & ~n15383;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = ~n15389 & ~n15392;
  assign n15394 = ~n15386 & ~n15393;
  assign n15395 = ~n13554 & ~n13565;
  assign n15396 = n13554 & n13565;
  assign n15397 = ~n13559 & ~n15396;
  assign n15398 = ~n15395 & ~n15397;
  assign n15399 = ~n15394 & n15398;
  assign n15400 = n15394 & ~n15398;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = pi139 & pi268;
  assign n15403 = pi138 & pi269;
  assign n15404 = n15402 & n15403;
  assign n15405 = ~n15402 & ~n15403;
  assign n15406 = ~n15404 & ~n15405;
  assign n15407 = ~n15401 & ~n15406;
  assign n15408 = n15394 & n15398;
  assign n15409 = ~n15394 & ~n15398;
  assign n15410 = ~n15408 & ~n15409;
  assign n15411 = pi268 & ~n15403;
  assign n15412 = pi139 & n15411;
  assign n15413 = pi269 & ~n15402;
  assign n15414 = pi138 & n15413;
  assign n15415 = ~n15412 & ~n15414;
  assign n15416 = ~n15410 & ~n15415;
  assign n15417 = ~n15407 & ~n15416;
  assign n15418 = ~n13583 & ~n13590;
  assign n15419 = ~n13578 & n15418;
  assign n15420 = ~n13591 & ~n15419;
  assign n15421 = n15417 & n15420;
  assign n15422 = ~n15417 & ~n15420;
  assign n15423 = ~n15421 & ~n15422;
  assign n15424 = pi140 & pi267;
  assign n15425 = ~n13570 & ~n13583;
  assign n15426 = ~n13578 & n15425;
  assign n15427 = n13570 & ~n13586;
  assign n15428 = ~n15426 & ~n15427;
  assign n15429 = ~n13379 & ~n15428;
  assign n15430 = n13570 & ~n13583;
  assign n15431 = ~n13578 & n15430;
  assign n15432 = ~n13570 & ~n13586;
  assign n15433 = ~n15431 & ~n15432;
  assign n15434 = pi267 & ~n15433;
  assign n15435 = pi139 & n15434;
  assign n15436 = ~n15429 & ~n15435;
  assign n15437 = n13602 & n15436;
  assign n15438 = ~n13602 & ~n15436;
  assign n15439 = n13579 & ~n15438;
  assign n15440 = ~n15437 & ~n15439;
  assign n15441 = n15424 & ~n15440;
  assign n15442 = ~n13579 & ~n15437;
  assign n15443 = ~n15438 & ~n15442;
  assign n15444 = ~n15424 & ~n15443;
  assign n15445 = ~n15441 & ~n15444;
  assign n15446 = ~n15423 & ~n15445;
  assign n15447 = n15417 & ~n15420;
  assign n15448 = ~n15417 & n15420;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = ~n15424 & ~n15440;
  assign n15451 = n15424 & ~n15443;
  assign n15452 = ~n15450 & ~n15451;
  assign n15453 = ~n15449 & ~n15452;
  assign n15454 = ~n15446 & ~n15453;
  assign n15455 = ~n13606 & ~n13617;
  assign n15456 = n13606 & n13617;
  assign n15457 = ~n13611 & ~n15456;
  assign n15458 = ~n15455 & ~n15457;
  assign n15459 = ~n15454 & n15458;
  assign n15460 = n15454 & ~n15458;
  assign n15461 = ~n15459 & ~n15460;
  assign n15462 = pi142 & pi265;
  assign n15463 = pi141 & pi266;
  assign n15464 = n15462 & n15463;
  assign n15465 = ~n15462 & ~n15463;
  assign n15466 = ~n15464 & ~n15465;
  assign n15467 = ~n15461 & ~n15466;
  assign n15468 = n15454 & n15458;
  assign n15469 = ~n15454 & ~n15458;
  assign n15470 = ~n15468 & ~n15469;
  assign n15471 = pi265 & ~n15463;
  assign n15472 = pi142 & n15471;
  assign n15473 = pi266 & ~n15462;
  assign n15474 = pi141 & n15473;
  assign n15475 = ~n15472 & ~n15474;
  assign n15476 = ~n15470 & ~n15475;
  assign n15477 = ~n15467 & ~n15476;
  assign n15478 = ~n13635 & ~n13642;
  assign n15479 = ~n13630 & n15478;
  assign n15480 = ~n13643 & ~n15479;
  assign n15481 = n15477 & ~n15480;
  assign n15482 = ~n15477 & n15480;
  assign n15483 = ~n15481 & ~n15482;
  assign n15484 = pi143 & pi264;
  assign n15485 = ~n13622 & ~n13635;
  assign n15486 = ~n13630 & n15485;
  assign n15487 = n13622 & ~n13638;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = ~n13378 & ~n15488;
  assign n15490 = n13622 & ~n13635;
  assign n15491 = ~n13630 & n15490;
  assign n15492 = ~n13622 & ~n13638;
  assign n15493 = ~n15491 & ~n15492;
  assign n15494 = pi264 & ~n15493;
  assign n15495 = pi142 & n15494;
  assign n15496 = ~n15489 & ~n15495;
  assign n15497 = n13654 & n15496;
  assign n15498 = ~n13654 & ~n15496;
  assign n15499 = n13631 & ~n15498;
  assign n15500 = ~n15497 & ~n15499;
  assign n15501 = n15484 & ~n15500;
  assign n15502 = ~n13631 & ~n15497;
  assign n15503 = ~n15498 & ~n15502;
  assign n15504 = ~n15484 & ~n15503;
  assign n15505 = ~n15501 & ~n15504;
  assign n15506 = ~n15483 & ~n15505;
  assign n15507 = n15477 & n15480;
  assign n15508 = ~n15477 & ~n15480;
  assign n15509 = ~n15507 & ~n15508;
  assign n15510 = ~n15484 & ~n15500;
  assign n15511 = n15484 & ~n15503;
  assign n15512 = ~n15510 & ~n15511;
  assign n15513 = ~n15509 & ~n15512;
  assign n15514 = ~n15506 & ~n15513;
  assign n15515 = n13660 & ~n13663;
  assign n15516 = n12847 & ~n12852;
  assign n15517 = ~n12853 & ~n15516;
  assign n15518 = ~n13660 & n13663;
  assign n15519 = ~n15517 & ~n15518;
  assign n15520 = ~n15515 & ~n15519;
  assign n15521 = ~n15514 & n15520;
  assign n15522 = n15514 & ~n15520;
  assign n15523 = ~n15521 & ~n15522;
  assign n15524 = pi145 & pi262;
  assign n15525 = pi144 & pi263;
  assign n15526 = n15524 & n15525;
  assign n15527 = ~n15524 & ~n15525;
  assign n15528 = ~n15526 & ~n15527;
  assign n15529 = ~n15523 & ~n15528;
  assign n15530 = n15514 & n15520;
  assign n15531 = ~n15514 & ~n15520;
  assign n15532 = ~n15530 & ~n15531;
  assign n15533 = pi262 & ~n15525;
  assign n15534 = pi145 & n15533;
  assign n15535 = pi263 & ~n15524;
  assign n15536 = pi144 & n15535;
  assign n15537 = ~n15534 & ~n15536;
  assign n15538 = ~n15532 & ~n15537;
  assign n15539 = ~n15529 & ~n15538;
  assign n15540 = ~n13672 & ~n13679;
  assign n15541 = n13672 & n13679;
  assign n15542 = ~n13682 & ~n15541;
  assign n15543 = ~n13678 & n15542;
  assign n15544 = ~n15540 & ~n15543;
  assign n15545 = n15539 & n15544;
  assign n15546 = ~n15539 & ~n15544;
  assign n15547 = ~n15545 & ~n15546;
  assign n15548 = pi146 & pi261;
  assign n15549 = n12510 & ~n13706;
  assign n15550 = ~n12510 & n13706;
  assign n15551 = ~n13364 & ~n15550;
  assign n15552 = ~n15549 & n15551;
  assign n15553 = n13352 & ~n15552;
  assign n15554 = n13697 & n15553;
  assign n15555 = ~n13697 & ~n15553;
  assign n15556 = n13345 & ~n15555;
  assign n15557 = ~n15554 & ~n15556;
  assign n15558 = n15548 & ~n15557;
  assign n15559 = ~n13345 & ~n15554;
  assign n15560 = ~n15555 & ~n15559;
  assign n15561 = ~n15548 & ~n15560;
  assign n15562 = ~n15558 & ~n15561;
  assign n15563 = ~n15547 & ~n15562;
  assign n15564 = n15539 & ~n15544;
  assign n15565 = ~n15539 & n15544;
  assign n15566 = ~n15564 & ~n15565;
  assign n15567 = ~n15548 & ~n15557;
  assign n15568 = n15548 & ~n15560;
  assign n15569 = ~n15567 & ~n15568;
  assign n15570 = ~n15566 & ~n15569;
  assign n15571 = ~n15563 & ~n15570;
  assign n15572 = ~n13700 & ~n15151;
  assign n15573 = ~n15150 & ~n15572;
  assign n15574 = n15571 & ~n15573;
  assign n15575 = ~n15571 & n15573;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = pi148 & pi259;
  assign n15578 = ~n13745 & ~n15152;
  assign n15579 = ~n13700 & ~n15157;
  assign n15580 = n13701 & ~n15579;
  assign n15581 = ~n15578 & n15580;
  assign n15582 = ~n15577 & ~n15581;
  assign n15583 = pi147 & n13718;
  assign n15584 = ~pi147 & ~n13718;
  assign n15585 = ~n15583 & ~n15584;
  assign n15586 = ~n13700 & ~n15585;
  assign n15587 = pi147 & ~n13718;
  assign n15588 = ~pi147 & n13718;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = ~n13745 & ~n15589;
  assign n15591 = ~n15586 & ~n15590;
  assign n15592 = n13701 & ~n15591;
  assign n15593 = pi259 & n15592;
  assign n15594 = ~n15582 & ~n15593;
  assign n15595 = pi149 & pi258;
  assign n15596 = pi147 & pi260;
  assign n15597 = ~n15595 & ~n15596;
  assign n15598 = n15595 & n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = ~n15594 & ~n15599;
  assign n15601 = ~n15595 & n15596;
  assign n15602 = n15595 & ~n15596;
  assign n15603 = ~n15601 & ~n15602;
  assign n15604 = ~n15593 & ~n15603;
  assign n15605 = ~n15582 & n15604;
  assign n15606 = ~n15600 & ~n15605;
  assign n15607 = ~n15576 & ~n15606;
  assign n15608 = n15571 & n15573;
  assign n15609 = ~n15571 & ~n15573;
  assign n15610 = ~n15608 & ~n15609;
  assign n15611 = ~n15594 & ~n15603;
  assign n15612 = ~n15593 & ~n15599;
  assign n15613 = ~n15582 & n15612;
  assign n15614 = ~n15611 & ~n15613;
  assign n15615 = ~n15610 & ~n15614;
  assign n15616 = ~n15607 & ~n15615;
  assign n15617 = ~n13754 & ~n15166;
  assign n15618 = n13754 & n15166;
  assign n15619 = ~n13729 & ~n15618;
  assign n15620 = ~n15617 & ~n15619;
  assign n15621 = n15616 & n15620;
  assign n15622 = ~n15616 & ~n15620;
  assign n15623 = ~n15621 & ~n15622;
  assign n15624 = ~n15166 & ~n15623;
  assign n15625 = n15616 & ~n15620;
  assign n15626 = ~n15616 & n15620;
  assign n15627 = ~n15625 & ~n15626;
  assign n15628 = n15166 & ~n15627;
  assign n15629 = ~n15624 & ~n15628;
  assign n15630 = pi322 & ~n15629;
  assign n15631 = ~n15149 & ~n15630;
  assign n15632 = n13762 & ~n15629;
  assign n15633 = pi323 & n15632;
  assign n15634 = pi322 & n15633;
  assign n15635 = ~n15631 & ~n15634;
  assign n15636 = pi325 & n11711;
  assign n15637 = pi324 & n12917;
  assign n15638 = n15636 & n15637;
  assign n15639 = ~n15636 & ~n15637;
  assign n15640 = ~n15638 & ~n15639;
  assign n15641 = ~n15635 & ~n15640;
  assign n15642 = ~n15636 & n15637;
  assign n15643 = n15636 & ~n15637;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = ~n15634 & ~n15644;
  assign n15646 = ~n15631 & n15645;
  assign n15647 = ~n15641 & ~n15646;
  assign n15648 = ~n15148 & ~n15647;
  assign n15649 = ~n15141 & ~n15145;
  assign n15650 = n15141 & n15145;
  assign n15651 = ~n15649 & ~n15650;
  assign n15652 = ~n15635 & ~n15644;
  assign n15653 = ~n15634 & ~n15640;
  assign n15654 = ~n15631 & n15653;
  assign n15655 = ~n15652 & ~n15654;
  assign n15656 = ~n15651 & ~n15655;
  assign n15657 = ~n15648 & ~n15656;
  assign n15658 = ~n13333 & n13778;
  assign n15659 = ~n13329 & ~n13773;
  assign n15660 = n13329 & n13773;
  assign n15661 = ~n15659 & ~n15660;
  assign n15662 = n13337 & ~n15661;
  assign n15663 = n13329 & ~n13773;
  assign n15664 = ~n13329 & n13773;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = ~n13337 & ~n15665;
  assign n15667 = ~n15662 & ~n15666;
  assign n15668 = n13333 & ~n13778;
  assign n15669 = ~n15667 & ~n15668;
  assign n15670 = ~n15658 & ~n15669;
  assign n15671 = n15657 & n15670;
  assign n15672 = ~n15657 & ~n15670;
  assign n15673 = ~n15671 & ~n15672;
  assign n15674 = pi327 & n11366;
  assign n15675 = pi326 & n11384;
  assign n15676 = n15674 & n15675;
  assign n15677 = ~n15674 & ~n15675;
  assign n15678 = ~n15676 & ~n15677;
  assign n15679 = ~n15673 & ~n15678;
  assign n15680 = ~n15657 & n15670;
  assign n15681 = n15657 & ~n15670;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = ~n15674 & n15675;
  assign n15684 = n15674 & ~n15675;
  assign n15685 = ~n15683 & ~n15684;
  assign n15686 = ~n15682 & ~n15685;
  assign n15687 = ~n15679 & ~n15686;
  assign n15688 = ~n15135 & ~n15687;
  assign n15689 = n15128 & n15132;
  assign n15690 = ~n15128 & ~n15132;
  assign n15691 = ~n15689 & ~n15690;
  assign n15692 = ~n15678 & ~n15682;
  assign n15693 = ~n15673 & ~n15685;
  assign n15694 = ~n15692 & ~n15693;
  assign n15695 = ~n15691 & ~n15694;
  assign n15696 = ~n15688 & ~n15695;
  assign n15697 = ~n15113 & n15696;
  assign n15698 = n15113 & ~n15696;
  assign n15699 = ~n15697 & ~n15698;
  assign n15700 = pi330 & n6556;
  assign n15701 = pi330 & n5973;
  assign n15702 = pi330 & n13862;
  assign n15703 = ~n13288 & ~n13855;
  assign n15704 = ~n15702 & ~n15703;
  assign n15705 = ~n15701 & n15704;
  assign n15706 = ~n15700 & ~n15705;
  assign n15707 = n13299 & n15706;
  assign n15708 = n15701 & ~n15704;
  assign n15709 = n15700 & ~n15708;
  assign n15710 = ~n13299 & n15709;
  assign n15711 = ~n15707 & ~n15710;
  assign n15712 = ~n15067 & ~n15711;
  assign n15713 = n13299 & n15709;
  assign n15714 = ~n13299 & n15706;
  assign n15715 = ~n15713 & ~n15714;
  assign n15716 = ~n15057 & ~n15715;
  assign n15717 = ~n15700 & ~n15704;
  assign n15718 = n15701 & n15717;
  assign n15719 = n15700 & n15704;
  assign n15720 = ~n15701 & n15719;
  assign n15721 = ~n15718 & ~n15720;
  assign n15722 = ~n15716 & n15721;
  assign n15723 = ~n15712 & n15722;
  assign n15724 = pi329 & n9205;
  assign n15725 = ~n15723 & n15724;
  assign n15726 = n15723 & ~n15724;
  assign n15727 = ~n15725 & ~n15726;
  assign n15728 = ~n15699 & ~n15727;
  assign n15729 = n15113 & n15696;
  assign n15730 = ~n15113 & ~n15696;
  assign n15731 = ~n15729 & ~n15730;
  assign n15732 = n15723 & n15724;
  assign n15733 = ~n15723 & ~n15724;
  assign n15734 = ~n15732 & ~n15733;
  assign n15735 = ~n15731 & ~n15734;
  assign n15736 = ~n15728 & ~n15735;
  assign n15737 = ~n15112 & ~n15736;
  assign n15738 = n15105 & n15109;
  assign n15739 = ~n15105 & ~n15109;
  assign n15740 = ~n15738 & ~n15739;
  assign n15741 = ~n15727 & ~n15731;
  assign n15742 = ~n15699 & ~n15734;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = ~n15740 & ~n15743;
  assign n15745 = ~n15737 & ~n15744;
  assign n15746 = ~n15085 & n15745;
  assign n15747 = n15085 & ~n15745;
  assign n15748 = ~n15746 & ~n15747;
  assign n15749 = pi333 & n5714;
  assign n15750 = n5257 & ~n13904;
  assign n15751 = pi332 & n15750;
  assign n15752 = ~n13905 & ~n15751;
  assign n15753 = ~n13889 & n15752;
  assign n15754 = n13889 & ~n15752;
  assign n15755 = ~n5714 & ~n15754;
  assign n15756 = ~n15753 & ~n15755;
  assign n15757 = n5732 & ~n15756;
  assign n15758 = ~n5732 & ~n15753;
  assign n15759 = n5714 & n15758;
  assign n15760 = ~n15757 & ~n15759;
  assign n15761 = pi332 & ~n15760;
  assign n15762 = pi332 & n5732;
  assign n15763 = n13889 & ~n15762;
  assign n15764 = ~n15752 & n15763;
  assign n15765 = ~n15761 & ~n15764;
  assign n15766 = n15749 & ~n15765;
  assign n15767 = ~n15749 & n15765;
  assign n15768 = ~n15766 & ~n15767;
  assign n15769 = ~n15748 & ~n15768;
  assign n15770 = n15085 & n15745;
  assign n15771 = ~n15085 & ~n15745;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = ~n15749 & ~n15765;
  assign n15774 = n15749 & n15765;
  assign n15775 = ~n15773 & ~n15774;
  assign n15776 = ~n15772 & ~n15775;
  assign n15777 = ~n15769 & ~n15776;
  assign n15778 = ~n15084 & ~n15777;
  assign n15779 = n15074 & n15081;
  assign n15780 = ~n15074 & ~n15081;
  assign n15781 = ~n15779 & ~n15780;
  assign n15782 = ~n15768 & ~n15772;
  assign n15783 = ~n15748 & ~n15775;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = ~n15781 & ~n15784;
  assign n15786 = ~n15778 & ~n15785;
  assign n15787 = ~n13233 & n13257;
  assign n15788 = n13233 & ~n13257;
  assign n15789 = n13947 & ~n15788;
  assign n15790 = ~n15787 & ~n15789;
  assign n15791 = n15786 & n15790;
  assign n15792 = ~n15786 & ~n15790;
  assign n15793 = ~n15791 & ~n15792;
  assign n15794 = pi335 & n4596;
  assign n15795 = ~n13919 & ~n13935;
  assign n15796 = ~n13942 & n15795;
  assign n15797 = ~n13933 & ~n13935;
  assign n15798 = ~n13899 & n15797;
  assign n15799 = ~n13934 & ~n15798;
  assign n15800 = ~n15796 & n15799;
  assign n15801 = pi334 & n5257;
  assign n15802 = n15800 & ~n15801;
  assign n15803 = n5257 & ~n15800;
  assign n15804 = pi334 & n15803;
  assign n15805 = ~n15802 & ~n15804;
  assign n15806 = ~n15794 & n15805;
  assign n15807 = n15794 & ~n15805;
  assign n15808 = ~n15806 & ~n15807;
  assign n15809 = pi336 & n2887;
  assign n15810 = n13257 & ~n15029;
  assign n15811 = ~n13257 & ~n15019;
  assign n15812 = ~n15810 & ~n15811;
  assign n15813 = n12398 & ~n13246;
  assign n15814 = ~n12398 & ~n13236;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = ~n13959 & ~n15815;
  assign n15817 = ~n13962 & ~n15816;
  assign n15818 = ~n13952 & n15817;
  assign n15819 = ~n15812 & ~n15818;
  assign n15820 = n13952 & ~n15817;
  assign n15821 = ~n15819 & ~n15820;
  assign n15822 = n15809 & n15821;
  assign n15823 = ~n15809 & ~n15821;
  assign n15824 = ~n15822 & ~n15823;
  assign n15825 = ~n15808 & ~n15824;
  assign n15826 = n15794 & n15805;
  assign n15827 = ~n15794 & ~n15805;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = ~n15809 & n15821;
  assign n15830 = n15809 & ~n15821;
  assign n15831 = ~n15829 & ~n15830;
  assign n15832 = ~n15828 & ~n15831;
  assign n15833 = ~n15825 & ~n15832;
  assign n15834 = ~n15793 & ~n15833;
  assign n15835 = n15786 & ~n15790;
  assign n15836 = ~n15786 & n15790;
  assign n15837 = ~n15835 & ~n15836;
  assign n15838 = ~n15824 & ~n15828;
  assign n15839 = ~n15808 & ~n15831;
  assign n15840 = ~n15838 & ~n15839;
  assign n15841 = ~n15837 & ~n15840;
  assign n15842 = ~n15834 & ~n15841;
  assign n15843 = ~n15054 & n15842;
  assign n15844 = n15054 & ~n15842;
  assign n15845 = ~n15843 & ~n15844;
  assign n15846 = pi339 & n1729;
  assign n15847 = ~n1729 & ~n15045;
  assign n15848 = ~n15044 & ~n15847;
  assign n15849 = n2091 & ~n15848;
  assign n15850 = ~n2091 & ~n15044;
  assign n15851 = n1729 & n15850;
  assign n15852 = ~n15849 & ~n15851;
  assign n15853 = pi338 & ~n15852;
  assign n15854 = pi338 & n2091;
  assign n15855 = n13998 & ~n15854;
  assign n15856 = ~n14011 & n15855;
  assign n15857 = ~n15853 & ~n15856;
  assign n15858 = n15846 & ~n15857;
  assign n15859 = ~n15846 & n15857;
  assign n15860 = ~n15858 & ~n15859;
  assign n15861 = ~n15845 & ~n15860;
  assign n15862 = n15054 & n15842;
  assign n15863 = ~n15054 & ~n15842;
  assign n15864 = ~n15862 & ~n15863;
  assign n15865 = ~n15846 & ~n15857;
  assign n15866 = n15846 & n15857;
  assign n15867 = ~n15865 & ~n15866;
  assign n15868 = ~n15864 & ~n15867;
  assign n15869 = ~n15861 & ~n15868;
  assign n15870 = ~n15053 & ~n15869;
  assign n15871 = n15036 & ~n15050;
  assign n15872 = ~n15036 & n15050;
  assign n15873 = ~n15871 & ~n15872;
  assign n15874 = ~n15860 & ~n15864;
  assign n15875 = ~n15845 & ~n15867;
  assign n15876 = ~n15874 & ~n15875;
  assign n15877 = ~n15873 & ~n15876;
  assign n15878 = ~n15870 & ~n15877;
  assign n15879 = ~n14045 & ~n14058;
  assign n15880 = ~n14044 & ~n15879;
  assign n15881 = ~n15878 & n15880;
  assign n15882 = n15878 & ~n15880;
  assign n15883 = ~n15881 & ~n15882;
  assign n15884 = n13224 & ~n14032;
  assign n15885 = ~n13224 & n14032;
  assign n15886 = ~n1256 & ~n15885;
  assign n15887 = ~n15884 & ~n15886;
  assign n15888 = n1442 & ~n15887;
  assign n15889 = pi340 & n15888;
  assign n15890 = ~n1442 & ~n15886;
  assign n15891 = pi340 & ~n15890;
  assign n15892 = ~n15884 & ~n15891;
  assign n15893 = ~n15889 & ~n15892;
  assign n15894 = ~n1256 & ~n15893;
  assign n15895 = pi341 & n15894;
  assign n15896 = pi341 & ~n1256;
  assign n15897 = ~n15892 & ~n15896;
  assign n15898 = ~n15889 & n15897;
  assign n15899 = ~n15895 & ~n15898;
  assign n15900 = ~n15883 & ~n15899;
  assign n15901 = n15878 & n15880;
  assign n15902 = ~n15878 & ~n15880;
  assign n15903 = ~n15901 & ~n15902;
  assign n15904 = n15893 & n15896;
  assign n15905 = ~n15893 & ~n15896;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = ~n15903 & ~n15906;
  assign n15908 = ~n15900 & ~n15907;
  assign n15909 = pi342 & ~n1154;
  assign n15910 = ~n14035 & ~n14046;
  assign n15911 = pi128 & pi342;
  assign n15912 = pi258 & n15911;
  assign n15913 = ~n14052 & ~n14058;
  assign n15914 = n15912 & ~n15913;
  assign n15915 = ~n15910 & n15914;
  assign n15916 = ~n15909 & ~n15915;
  assign n15917 = pi341 & n14042;
  assign n15918 = ~pi341 & ~n14042;
  assign n15919 = ~n15917 & ~n15918;
  assign n15920 = ~n14058 & ~n15919;
  assign n15921 = pi341 & ~n14042;
  assign n15922 = ~pi341 & n14042;
  assign n15923 = ~n15921 & ~n15922;
  assign n15924 = ~n14035 & ~n15923;
  assign n15925 = ~n15920 & ~n15924;
  assign n15926 = n15912 & ~n15925;
  assign n15927 = ~n1154 & n15926;
  assign n15928 = ~n15916 & ~n15927;
  assign n15929 = n15908 & ~n15928;
  assign n15930 = ~n15908 & ~n15927;
  assign n15931 = ~n15916 & n15930;
  assign n15932 = ~n15929 & ~n15931;
  assign n15933 = pi279 & n15932;
  assign n15934 = ~pi279 & ~n15932;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = pi258 & ~n15935;
  assign n15937 = pi128 & n15936;
  assign n15938 = pi343 & n15937;
  assign n15939 = pi279 & ~n15932;
  assign n15940 = ~pi279 & n15932;
  assign n15941 = ~n15939 & ~n15940;
  assign n15942 = pi343 & n1156;
  assign n15943 = ~n15941 & ~n15942;
  assign n15944 = ~n15938 & ~n15943;
  assign n15945 = ~n15016 & ~n15944;
  assign n15946 = n15016 & n15944;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = ~n15012 & ~n15947;
  assign n15949 = ~n15016 & n15944;
  assign n15950 = n15016 & ~n15944;
  assign n15951 = ~n15949 & ~n15950;
  assign n15952 = n15012 & ~n15951;
  assign n15953 = ~n15948 & ~n15952;
  assign n15954 = ~n14520 & ~n14532;
  assign n15955 = ~n14519 & n14532;
  assign n15956 = ~n14518 & n15955;
  assign n15957 = ~n14516 & ~n15956;
  assign n15958 = ~n15954 & ~n15957;
  assign n15959 = n15953 & n15958;
  assign n15960 = ~n15953 & ~n15958;
  assign n15961 = ~n15959 & ~n15960;
  assign n15962 = ~n831 & ~n15961;
  assign n15963 = ~n14543 & ~n15962;
  assign n15964 = pi161 & ~n15963;
  assign n15965 = ~n14542 & ~n15964;
  assign po214 = ~pi160 & n15965;
  assign n15967 = pi086 & ~pi161;
  assign n15968 = n1256 & ~n15884;
  assign n15969 = ~n15885 & ~n15968;
  assign n15970 = n1442 & ~n15969;
  assign n15971 = ~n1442 & ~n15885;
  assign n15972 = ~n1256 & n15971;
  assign n15973 = ~n15970 & ~n15972;
  assign n15974 = pi340 & ~n15973;
  assign n15975 = pi340 & n1442;
  assign n15976 = ~n14032 & ~n15975;
  assign n15977 = n13224 & n15976;
  assign n15978 = ~n15974 & ~n15977;
  assign n15979 = ~n15896 & n15978;
  assign n15980 = n15896 & ~n15978;
  assign n15981 = ~n15979 & ~n15980;
  assign n15982 = ~n15883 & ~n15981;
  assign n15983 = n15896 & n15978;
  assign n15984 = ~n15896 & ~n15978;
  assign n15985 = ~n15983 & ~n15984;
  assign n15986 = ~n15903 & ~n15985;
  assign n15987 = ~n15927 & ~n15986;
  assign n15988 = ~n15982 & n15987;
  assign n15989 = ~n15916 & ~n15988;
  assign n15990 = pi342 & ~n1256;
  assign n15991 = n15989 & ~n15990;
  assign n15992 = ~n1256 & ~n15989;
  assign n15993 = pi342 & n15992;
  assign n15994 = ~n15991 & ~n15993;
  assign n15995 = ~n15036 & ~n15842;
  assign n15996 = n15036 & n15842;
  assign n15997 = ~n15995 & ~n15996;
  assign n15998 = n15050 & n15846;
  assign n15999 = n15054 & ~n15857;
  assign n16000 = ~n15054 & n15857;
  assign n16001 = ~n15999 & ~n16000;
  assign n16002 = ~n15998 & ~n16001;
  assign n16003 = ~n15997 & n16002;
  assign n16004 = ~n15036 & n15842;
  assign n16005 = n15036 & ~n15842;
  assign n16006 = ~n16004 & ~n16005;
  assign n16007 = ~n15054 & ~n15857;
  assign n16008 = n15054 & n15857;
  assign n16009 = ~n16007 & ~n16008;
  assign n16010 = ~n15998 & ~n16009;
  assign n16011 = ~n16006 & n16010;
  assign n16012 = ~n15050 & ~n15846;
  assign n16013 = ~n16011 & ~n16012;
  assign n16014 = ~n16003 & n16013;
  assign n16015 = ~n15880 & n15896;
  assign n16016 = n15880 & ~n15896;
  assign n16017 = n15878 & n15893;
  assign n16018 = ~n15878 & ~n15893;
  assign n16019 = ~n16017 & ~n16018;
  assign n16020 = ~n16016 & ~n16019;
  assign n16021 = ~n16015 & ~n16020;
  assign n16022 = n16014 & n16021;
  assign n16023 = ~n16014 & ~n16021;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = ~n15878 & ~n15892;
  assign n16026 = ~n15889 & ~n16025;
  assign n16027 = n1729 & n16026;
  assign n16028 = pi340 & n16027;
  assign n16029 = pi340 & n1729;
  assign n16030 = ~n16026 & ~n16029;
  assign n16031 = ~n16028 & ~n16030;
  assign n16032 = ~n15074 & ~n15745;
  assign n16033 = n15074 & n15745;
  assign n16034 = ~n16032 & ~n16033;
  assign n16035 = ~n15081 & n15749;
  assign n16036 = n15085 & ~n15765;
  assign n16037 = ~n15085 & n15765;
  assign n16038 = ~n16036 & ~n16037;
  assign n16039 = ~n16035 & ~n16038;
  assign n16040 = ~n16034 & n16039;
  assign n16041 = ~n15074 & n15745;
  assign n16042 = n15074 & ~n15745;
  assign n16043 = ~n16041 & ~n16042;
  assign n16044 = ~n15085 & ~n15765;
  assign n16045 = n15085 & n15765;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = ~n16035 & ~n16046;
  assign n16048 = ~n16043 & n16047;
  assign n16049 = n15081 & ~n15749;
  assign n16050 = ~n16048 & ~n16049;
  assign n16051 = ~n16040 & n16050;
  assign n16052 = ~n15786 & n15805;
  assign n16053 = n15786 & ~n15805;
  assign n16054 = ~n16052 & ~n16053;
  assign n16055 = n15790 & ~n15794;
  assign n16056 = ~n16054 & ~n16055;
  assign n16057 = ~n15790 & n15794;
  assign n16058 = ~n16056 & ~n16057;
  assign n16059 = n16051 & n16058;
  assign n16060 = ~n16051 & ~n16058;
  assign n16061 = ~n16059 & ~n16060;
  assign n16062 = n15786 & ~n15800;
  assign n16063 = ~n15786 & n15800;
  assign n16064 = ~n5257 & ~n16063;
  assign n16065 = ~n16062 & ~n16064;
  assign n16066 = n5714 & ~n16065;
  assign n16067 = ~n5714 & ~n16062;
  assign n16068 = n5257 & n16067;
  assign n16069 = ~n16066 & ~n16068;
  assign n16070 = pi334 & ~n16069;
  assign n16071 = pi334 & n5714;
  assign n16072 = ~n15786 & ~n16071;
  assign n16073 = n15800 & n16072;
  assign n16074 = ~n16070 & ~n16073;
  assign n16075 = ~n15105 & n15113;
  assign n16076 = n15105 & ~n15113;
  assign n16077 = ~n15696 & ~n16076;
  assign n16078 = ~n16075 & ~n16077;
  assign n16079 = ~n15109 & n15724;
  assign n16080 = ~n15105 & ~n15696;
  assign n16081 = n15105 & n15696;
  assign n16082 = ~n16080 & ~n16081;
  assign n16083 = n15113 & ~n16082;
  assign n16084 = n15105 & ~n15696;
  assign n16085 = ~n15105 & n15696;
  assign n16086 = ~n16084 & ~n16085;
  assign n16087 = ~n15113 & ~n16086;
  assign n16088 = ~n16083 & ~n16087;
  assign n16089 = n15109 & ~n15724;
  assign n16090 = ~n16088 & ~n16089;
  assign n16091 = ~n16079 & ~n16090;
  assign n16092 = n16078 & ~n16091;
  assign n16093 = ~n16078 & n16091;
  assign n16094 = ~n16092 & ~n16093;
  assign n16095 = pi329 & n10561;
  assign n16096 = ~n15128 & n15675;
  assign n16097 = n15128 & ~n15675;
  assign n16098 = ~n15682 & ~n16097;
  assign n16099 = ~n16096 & ~n16098;
  assign n16100 = ~n15128 & ~n15670;
  assign n16101 = n15128 & n15670;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = ~n15132 & n15674;
  assign n16104 = ~n15657 & n15675;
  assign n16105 = n15657 & ~n15675;
  assign n16106 = ~n16104 & ~n16105;
  assign n16107 = ~n16103 & ~n16106;
  assign n16108 = ~n16102 & n16107;
  assign n16109 = ~n15128 & n15670;
  assign n16110 = n15128 & ~n15670;
  assign n16111 = ~n16109 & ~n16110;
  assign n16112 = n15657 & n15675;
  assign n16113 = ~n15657 & ~n15675;
  assign n16114 = ~n16112 & ~n16113;
  assign n16115 = ~n16103 & ~n16114;
  assign n16116 = ~n16111 & n16115;
  assign n16117 = n15132 & ~n15674;
  assign n16118 = ~n16116 & ~n16117;
  assign n16119 = ~n16108 & n16118;
  assign n16120 = n16099 & n16119;
  assign n16121 = ~n16099 & ~n16119;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = ~n15141 & ~n15631;
  assign n16124 = ~n15634 & ~n16123;
  assign n16125 = ~n15145 & n15637;
  assign n16126 = ~n15141 & ~n15635;
  assign n16127 = n15141 & ~n15634;
  assign n16128 = ~n15631 & n16127;
  assign n16129 = ~n16126 & ~n16128;
  assign n16130 = n15145 & ~n15637;
  assign n16131 = ~n16129 & ~n16130;
  assign n16132 = ~n16125 & ~n16131;
  assign n16133 = ~n16124 & n16132;
  assign n16134 = n16124 & ~n16132;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = pi145 & pi263;
  assign n16137 = pi142 & pi266;
  assign n16138 = pi139 & pi269;
  assign n16139 = pi136 & pi272;
  assign n16140 = ~n15255 & n15266;
  assign n16141 = ~n15254 & ~n15266;
  assign n16142 = ~n15251 & n16141;
  assign n16143 = ~n16140 & ~n16142;
  assign n16144 = ~n15313 & n16143;
  assign n16145 = pi132 & pi276;
  assign n16146 = ~n13391 & ~n13394;
  assign n16147 = n13391 & n13394;
  assign n16148 = n12561 & ~n15188;
  assign n16149 = ~n15186 & ~n16148;
  assign n16150 = ~n16147 & ~n16149;
  assign n16151 = ~n16146 & ~n16150;
  assign n16152 = ~n15183 & ~n16151;
  assign n16153 = ~n15181 & ~n16152;
  assign n16154 = pi128 & pi280;
  assign n16155 = pi279 & ~n16154;
  assign n16156 = pi129 & n16155;
  assign n16157 = pi129 & pi279;
  assign n16158 = pi280 & ~n16157;
  assign n16159 = pi128 & n16158;
  assign n16160 = ~n16156 & ~n16159;
  assign n16161 = pi130 & pi278;
  assign n16162 = ~n16160 & ~n16161;
  assign n16163 = pi278 & n16160;
  assign n16164 = pi130 & n16163;
  assign n16165 = ~n16162 & ~n16164;
  assign n16166 = ~n16153 & ~n16165;
  assign n16167 = n16160 & ~n16161;
  assign n16168 = pi278 & ~n16160;
  assign n16169 = pi130 & n16168;
  assign n16170 = ~n16167 & ~n16169;
  assign n16171 = ~n16152 & ~n16170;
  assign n16172 = ~n15181 & n16171;
  assign n16173 = ~n16166 & ~n16172;
  assign n16174 = ~n15199 & ~n15235;
  assign n16175 = n16173 & ~n16174;
  assign n16176 = n15214 & n16175;
  assign n16177 = n15214 & ~n16174;
  assign n16178 = ~n16173 & ~n16177;
  assign n16179 = ~n16176 & ~n16178;
  assign n16180 = pi277 & ~n16179;
  assign n16181 = pi131 & n16180;
  assign n16182 = pi131 & pi277;
  assign n16183 = ~n16178 & ~n16182;
  assign n16184 = ~n16176 & n16183;
  assign n16185 = ~n16181 & ~n16184;
  assign n16186 = ~n15178 & ~n15245;
  assign n16187 = ~n16185 & ~n16186;
  assign n16188 = ~n15242 & n16187;
  assign n16189 = ~n15242 & ~n16186;
  assign n16190 = ~n16184 & ~n16189;
  assign n16191 = ~n16181 & n16190;
  assign n16192 = ~n16188 & ~n16191;
  assign n16193 = ~n16145 & n16192;
  assign n16194 = n16145 & ~n16192;
  assign n16195 = ~n16193 & ~n16194;
  assign n16196 = pi133 & pi275;
  assign n16197 = ~n15251 & n15266;
  assign n16198 = n16196 & ~n16197;
  assign n16199 = ~n15254 & n16198;
  assign n16200 = ~n15254 & ~n16197;
  assign n16201 = ~n16196 & ~n16200;
  assign n16202 = ~n16199 & ~n16201;
  assign n16203 = ~n16195 & ~n16202;
  assign n16204 = ~n16145 & ~n16192;
  assign n16205 = n16145 & n16192;
  assign n16206 = ~n16204 & ~n16205;
  assign n16207 = ~n16196 & ~n16197;
  assign n16208 = ~n15254 & n16207;
  assign n16209 = n16196 & ~n16200;
  assign n16210 = ~n16208 & ~n16209;
  assign n16211 = ~n16206 & ~n16210;
  assign n16212 = ~n16203 & ~n16211;
  assign n16213 = ~pi274 & ~n16212;
  assign n16214 = ~pi134 & ~n16212;
  assign n16215 = pi274 & n16212;
  assign n16216 = pi134 & n16215;
  assign n16217 = ~n16214 & ~n16216;
  assign n16218 = ~pi133 & ~n16217;
  assign n16219 = ~n16213 & ~n16218;
  assign n16220 = ~n16144 & ~n16219;
  assign n16221 = n15313 & n16212;
  assign n16222 = pi274 & ~n16143;
  assign n16223 = n16221 & n16222;
  assign n16224 = n15313 & n16143;
  assign n16225 = ~n15313 & ~n16143;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = pi133 & ~n16226;
  assign n16228 = pi274 & n16144;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = ~n16212 & ~n16229;
  assign n16231 = ~n16223 & ~n16230;
  assign n16232 = pi134 & ~n16231;
  assign n16233 = ~pi274 & n16143;
  assign n16234 = ~n15313 & n16212;
  assign n16235 = n16233 & n16234;
  assign n16236 = n15313 & ~n16212;
  assign n16237 = ~n16143 & n16236;
  assign n16238 = n15313 & ~n16143;
  assign n16239 = pi274 & ~n16238;
  assign n16240 = pi133 & n16239;
  assign n16241 = ~n16144 & ~n16240;
  assign n16242 = n16212 & ~n16241;
  assign n16243 = ~n16237 & ~n16242;
  assign n16244 = ~pi134 & ~n16243;
  assign n16245 = ~n16235 & ~n16244;
  assign n16246 = ~n16232 & n16245;
  assign n16247 = ~n16220 & n16246;
  assign n16248 = n15317 & ~n15330;
  assign n16249 = ~n15317 & n15330;
  assign n16250 = ~n15321 & ~n16249;
  assign n16251 = ~n16248 & ~n16250;
  assign n16252 = n16247 & n16251;
  assign n16253 = ~n16247 & ~n16251;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = pi135 & pi273;
  assign n16256 = n15344 & ~n15350;
  assign n16257 = ~n15349 & ~n16256;
  assign n16258 = n16255 & ~n16257;
  assign n16259 = ~n15344 & ~n15349;
  assign n16260 = ~n15350 & ~n16259;
  assign n16261 = ~n16255 & ~n16260;
  assign n16262 = ~n16258 & ~n16261;
  assign n16263 = ~n16254 & ~n16262;
  assign n16264 = n16247 & ~n16251;
  assign n16265 = ~n16247 & n16251;
  assign n16266 = ~n16264 & ~n16265;
  assign n16267 = ~n16255 & ~n16257;
  assign n16268 = n16255 & ~n16260;
  assign n16269 = ~n16267 & ~n16268;
  assign n16270 = ~n16266 & ~n16269;
  assign n16271 = ~n16263 & ~n16270;
  assign n16272 = ~n16139 & n16271;
  assign n16273 = n16139 & ~n16271;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = pi272 & ~n15351;
  assign n16276 = pi135 & n16275;
  assign n16277 = ~n15342 & ~n15344;
  assign n16278 = ~n16276 & ~n16277;
  assign n16279 = pi271 & ~n16278;
  assign n16280 = pi136 & n16279;
  assign n16281 = pi137 & pi271;
  assign n16282 = ~n15343 & ~n16277;
  assign n16283 = ~n16276 & n16282;
  assign n16284 = ~n15360 & ~n16283;
  assign n16285 = ~n16281 & ~n16284;
  assign n16286 = ~n16280 & n16285;
  assign n16287 = ~n16280 & ~n16284;
  assign n16288 = n16281 & ~n16287;
  assign n16289 = ~n16286 & ~n16288;
  assign n16290 = ~n16274 & ~n16289;
  assign n16291 = ~n16139 & ~n16271;
  assign n16292 = n16139 & n16271;
  assign n16293 = ~n16291 & ~n16292;
  assign n16294 = n16281 & ~n16284;
  assign n16295 = ~n16280 & n16294;
  assign n16296 = ~n16281 & ~n16287;
  assign n16297 = ~n16295 & ~n16296;
  assign n16298 = ~n16293 & ~n16297;
  assign n16299 = ~n16290 & ~n16298;
  assign n16300 = n15364 & ~n15389;
  assign n16301 = ~n15364 & n15389;
  assign n16302 = ~n15380 & ~n16301;
  assign n16303 = ~n16300 & ~n16302;
  assign n16304 = n16299 & ~n16303;
  assign n16305 = ~n16299 & n16303;
  assign n16306 = ~n16304 & ~n16305;
  assign n16307 = pi138 & pi270;
  assign n16308 = n15403 & ~n15409;
  assign n16309 = ~n15408 & ~n16308;
  assign n16310 = n16307 & ~n16309;
  assign n16311 = ~n15403 & ~n15408;
  assign n16312 = ~n15409 & ~n16311;
  assign n16313 = ~n16307 & ~n16312;
  assign n16314 = ~n16310 & ~n16313;
  assign n16315 = ~n16306 & ~n16314;
  assign n16316 = n16299 & n16303;
  assign n16317 = ~n16299 & ~n16303;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = ~n16307 & ~n16309;
  assign n16320 = n16307 & ~n16312;
  assign n16321 = ~n16319 & ~n16320;
  assign n16322 = ~n16318 & ~n16321;
  assign n16323 = ~n16315 & ~n16322;
  assign n16324 = ~n16138 & ~n16323;
  assign n16325 = n16138 & n16323;
  assign n16326 = ~n16324 & ~n16325;
  assign n16327 = pi269 & ~n15410;
  assign n16328 = pi138 & n16327;
  assign n16329 = ~n15401 & ~n15403;
  assign n16330 = ~n15402 & ~n16329;
  assign n16331 = ~n16328 & n16330;
  assign n16332 = pi140 & pi268;
  assign n16333 = ~n16328 & ~n16329;
  assign n16334 = pi268 & ~n16333;
  assign n16335 = pi139 & n16334;
  assign n16336 = n15420 & ~n16335;
  assign n16337 = n16332 & ~n16336;
  assign n16338 = ~n16331 & n16337;
  assign n16339 = ~n16331 & ~n16336;
  assign n16340 = ~n16332 & ~n16339;
  assign n16341 = ~n16338 & ~n16340;
  assign n16342 = ~n16326 & ~n16341;
  assign n16343 = ~n16138 & n16323;
  assign n16344 = n16138 & ~n16323;
  assign n16345 = ~n16343 & ~n16344;
  assign n16346 = ~n16332 & ~n16336;
  assign n16347 = ~n16331 & n16346;
  assign n16348 = n16332 & ~n16339;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = ~n16345 & ~n16349;
  assign n16351 = ~n16342 & ~n16350;
  assign n16352 = ~n15423 & ~n15424;
  assign n16353 = n15423 & n15424;
  assign n16354 = ~n15443 & ~n16353;
  assign n16355 = ~n16352 & ~n16354;
  assign n16356 = n16351 & n16355;
  assign n16357 = ~n16351 & ~n16355;
  assign n16358 = ~n16356 & ~n16357;
  assign n16359 = pi141 & pi267;
  assign n16360 = n15463 & ~n15469;
  assign n16361 = ~n15468 & ~n16360;
  assign n16362 = n16359 & ~n16361;
  assign n16363 = ~n15463 & ~n15468;
  assign n16364 = ~n15469 & ~n16363;
  assign n16365 = ~n16359 & ~n16364;
  assign n16366 = ~n16362 & ~n16365;
  assign n16367 = ~n16358 & ~n16366;
  assign n16368 = n16351 & ~n16355;
  assign n16369 = ~n16351 & n16355;
  assign n16370 = ~n16368 & ~n16369;
  assign n16371 = ~n16359 & ~n16361;
  assign n16372 = n16359 & ~n16364;
  assign n16373 = ~n16371 & ~n16372;
  assign n16374 = ~n16370 & ~n16373;
  assign n16375 = ~n16367 & ~n16374;
  assign n16376 = ~n16137 & ~n16375;
  assign n16377 = n16137 & n16375;
  assign n16378 = ~n16376 & ~n16377;
  assign n16379 = pi266 & ~n15470;
  assign n16380 = pi141 & n16379;
  assign n16381 = ~n15461 & ~n15463;
  assign n16382 = ~n15462 & ~n16381;
  assign n16383 = ~n16380 & n16382;
  assign n16384 = pi143 & pi265;
  assign n16385 = ~n16380 & ~n16381;
  assign n16386 = pi265 & ~n16385;
  assign n16387 = pi142 & n16386;
  assign n16388 = n15480 & ~n16387;
  assign n16389 = n16384 & ~n16388;
  assign n16390 = ~n16383 & n16389;
  assign n16391 = ~n16383 & ~n16388;
  assign n16392 = ~n16384 & ~n16391;
  assign n16393 = ~n16390 & ~n16392;
  assign n16394 = ~n16378 & ~n16393;
  assign n16395 = ~n16137 & n16375;
  assign n16396 = n16137 & ~n16375;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = ~n16384 & ~n16388;
  assign n16399 = ~n16383 & n16398;
  assign n16400 = n16384 & ~n16391;
  assign n16401 = ~n16399 & ~n16400;
  assign n16402 = ~n16397 & ~n16401;
  assign n16403 = ~n16394 & ~n16402;
  assign n16404 = ~n15484 & ~n15509;
  assign n16405 = n15484 & n15509;
  assign n16406 = ~n15503 & ~n16405;
  assign n16407 = ~n16404 & ~n16406;
  assign n16408 = n16403 & ~n16407;
  assign n16409 = ~n16403 & n16407;
  assign n16410 = ~n16408 & ~n16409;
  assign n16411 = pi144 & pi264;
  assign n16412 = n15525 & ~n15530;
  assign n16413 = ~n15531 & ~n16412;
  assign n16414 = n16411 & ~n16413;
  assign n16415 = ~n15525 & ~n15531;
  assign n16416 = ~n15530 & ~n16415;
  assign n16417 = ~n16411 & ~n16416;
  assign n16418 = ~n16414 & ~n16417;
  assign n16419 = ~n16410 & ~n16418;
  assign n16420 = n16403 & n16407;
  assign n16421 = ~n16403 & ~n16407;
  assign n16422 = ~n16420 & ~n16421;
  assign n16423 = ~n16411 & ~n16413;
  assign n16424 = n16411 & ~n16416;
  assign n16425 = ~n16423 & ~n16424;
  assign n16426 = ~n16422 & ~n16425;
  assign n16427 = ~n16419 & ~n16426;
  assign n16428 = ~n16136 & n16427;
  assign n16429 = n16136 & ~n16427;
  assign n16430 = ~n16428 & ~n16429;
  assign n16431 = pi263 & ~n15532;
  assign n16432 = pi144 & n16431;
  assign n16433 = ~n15523 & ~n15525;
  assign n16434 = ~n16432 & ~n16433;
  assign n16435 = pi262 & ~n16434;
  assign n16436 = pi145 & n16435;
  assign n16437 = pi146 & pi262;
  assign n16438 = ~n15524 & ~n16433;
  assign n16439 = ~n16432 & n16438;
  assign n16440 = n15544 & ~n16439;
  assign n16441 = ~n16437 & ~n16440;
  assign n16442 = ~n16436 & n16441;
  assign n16443 = ~n16436 & ~n16440;
  assign n16444 = n16437 & ~n16443;
  assign n16445 = ~n16442 & ~n16444;
  assign n16446 = ~n16430 & ~n16445;
  assign n16447 = ~n16136 & ~n16427;
  assign n16448 = n16136 & n16427;
  assign n16449 = ~n16447 & ~n16448;
  assign n16450 = n16437 & ~n16440;
  assign n16451 = ~n16436 & n16450;
  assign n16452 = ~n16437 & ~n16443;
  assign n16453 = ~n16451 & ~n16452;
  assign n16454 = ~n16449 & ~n16453;
  assign n16455 = ~n16446 & ~n16454;
  assign n16456 = ~n15548 & ~n15566;
  assign n16457 = n15548 & n15566;
  assign n16458 = ~n15560 & ~n16457;
  assign n16459 = ~n16456 & ~n16458;
  assign n16460 = n16455 & ~n16459;
  assign n16461 = ~n16455 & n16459;
  assign n16462 = ~n16460 & ~n16461;
  assign n16463 = pi147 & pi261;
  assign n16464 = n15596 & ~n15608;
  assign n16465 = ~n15609 & ~n16464;
  assign n16466 = n16463 & ~n16465;
  assign n16467 = ~n15596 & ~n15609;
  assign n16468 = ~n15608 & ~n16467;
  assign n16469 = ~n16463 & ~n16468;
  assign n16470 = ~n16466 & ~n16469;
  assign n16471 = ~n16462 & ~n16470;
  assign n16472 = n16455 & n16459;
  assign n16473 = ~n16455 & ~n16459;
  assign n16474 = ~n16472 & ~n16473;
  assign n16475 = ~n16463 & ~n16465;
  assign n16476 = n16463 & ~n16468;
  assign n16477 = ~n16475 & ~n16476;
  assign n16478 = ~n16474 & ~n16477;
  assign n16479 = ~n16471 & ~n16478;
  assign n16480 = pi260 & ~n15610;
  assign n16481 = pi147 & n16480;
  assign n16482 = ~n15576 & ~n15596;
  assign n16483 = ~n15593 & ~n16482;
  assign n16484 = ~n16481 & n16483;
  assign n16485 = ~n15582 & ~n16484;
  assign n16486 = n16479 & ~n16485;
  assign n16487 = ~n16479 & n16485;
  assign n16488 = ~n16486 & ~n16487;
  assign n16489 = pi149 & pi259;
  assign n16490 = pi148 & pi260;
  assign n16491 = ~n16489 & ~n16490;
  assign n16492 = n16489 & n16490;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = ~n15593 & ~n15596;
  assign n16495 = ~n15582 & n16494;
  assign n16496 = ~n15594 & n15596;
  assign n16497 = ~n16495 & ~n16496;
  assign n16498 = ~n15610 & ~n16497;
  assign n16499 = ~n15593 & n15596;
  assign n16500 = ~n15582 & n16499;
  assign n16501 = ~n15594 & ~n15596;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n15576 & ~n16502;
  assign n16504 = ~n16498 & ~n16503;
  assign n16505 = n15595 & ~n16504;
  assign n16506 = pi150 & pi258;
  assign n16507 = n16505 & n16506;
  assign n16508 = ~n16505 & ~n16506;
  assign n16509 = ~n16507 & ~n16508;
  assign n16510 = ~n16493 & ~n16509;
  assign n16511 = n16489 & ~n16490;
  assign n16512 = ~n16489 & n16490;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = ~n16505 & n16506;
  assign n16515 = n16505 & ~n16506;
  assign n16516 = ~n16514 & ~n16515;
  assign n16517 = ~n16513 & ~n16516;
  assign n16518 = ~n16510 & ~n16517;
  assign n16519 = ~n16488 & ~n16518;
  assign n16520 = n16479 & n16485;
  assign n16521 = ~n16479 & ~n16485;
  assign n16522 = ~n16520 & ~n16521;
  assign n16523 = ~n16509 & ~n16513;
  assign n16524 = ~n16493 & ~n16516;
  assign n16525 = ~n16523 & ~n16524;
  assign n16526 = ~n16522 & ~n16525;
  assign n16527 = ~n16519 & ~n16526;
  assign n16528 = n15620 & ~n16527;
  assign n16529 = ~n15620 & n16527;
  assign n16530 = n15616 & n16529;
  assign n16531 = ~n16528 & ~n16530;
  assign n16532 = ~n15166 & ~n16531;
  assign n16533 = ~n15620 & ~n16527;
  assign n16534 = n15620 & n16527;
  assign n16535 = ~n15616 & n16534;
  assign n16536 = ~n16533 & ~n16535;
  assign n16537 = n15166 & ~n16536;
  assign n16538 = ~n15623 & ~n16527;
  assign n16539 = ~n16537 & ~n16538;
  assign n16540 = ~n16532 & n16539;
  assign n16541 = pi322 & ~n16540;
  assign n16542 = pi323 & ~n15629;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = n15166 & n15625;
  assign n16545 = ~n15624 & ~n16544;
  assign n16546 = ~n16527 & ~n16545;
  assign n16547 = n15166 & ~n15616;
  assign n16548 = n16534 & n16547;
  assign n16549 = ~n16546 & ~n16548;
  assign n16550 = pi323 & ~n16549;
  assign n16551 = pi322 & n16550;
  assign n16552 = ~n16543 & ~n16551;
  assign n16553 = pi325 & n12917;
  assign n16554 = pi324 & n13762;
  assign n16555 = n16553 & n16554;
  assign n16556 = ~n16553 & ~n16554;
  assign n16557 = ~n16555 & ~n16556;
  assign n16558 = ~n16552 & ~n16557;
  assign n16559 = ~n16553 & n16554;
  assign n16560 = n16553 & ~n16554;
  assign n16561 = ~n16559 & ~n16560;
  assign n16562 = ~n16551 & ~n16561;
  assign n16563 = ~n16543 & n16562;
  assign n16564 = ~n16558 & ~n16563;
  assign n16565 = ~n16135 & ~n16564;
  assign n16566 = ~n16124 & ~n16132;
  assign n16567 = n16124 & n16132;
  assign n16568 = ~n16566 & ~n16567;
  assign n16569 = ~n16552 & ~n16561;
  assign n16570 = ~n16551 & ~n16557;
  assign n16571 = ~n16543 & n16570;
  assign n16572 = ~n16569 & ~n16571;
  assign n16573 = ~n16568 & ~n16572;
  assign n16574 = ~n16565 & ~n16573;
  assign n16575 = n15636 & ~n15670;
  assign n16576 = ~n15145 & ~n16129;
  assign n16577 = n15145 & n16129;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = n15637 & ~n16578;
  assign n16580 = n15145 & ~n16129;
  assign n16581 = ~n15145 & n16129;
  assign n16582 = ~n16580 & ~n16581;
  assign n16583 = ~n15637 & ~n16582;
  assign n16584 = ~n16579 & ~n16583;
  assign n16585 = ~n15636 & n15670;
  assign n16586 = ~n16584 & ~n16585;
  assign n16587 = ~n16575 & ~n16586;
  assign n16588 = n16574 & n16587;
  assign n16589 = ~n16574 & ~n16587;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = pi327 & n11384;
  assign n16592 = pi326 & n11711;
  assign n16593 = n16591 & n16592;
  assign n16594 = ~n16591 & ~n16592;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = ~n16590 & ~n16595;
  assign n16597 = ~n16574 & n16587;
  assign n16598 = n16574 & ~n16587;
  assign n16599 = ~n16597 & ~n16598;
  assign n16600 = ~n16591 & n16592;
  assign n16601 = n16591 & ~n16592;
  assign n16602 = ~n16600 & ~n16601;
  assign n16603 = ~n16599 & ~n16602;
  assign n16604 = ~n16596 & ~n16603;
  assign n16605 = ~n16122 & ~n16604;
  assign n16606 = n16099 & ~n16119;
  assign n16607 = ~n16099 & n16119;
  assign n16608 = ~n16606 & ~n16607;
  assign n16609 = ~n16595 & ~n16599;
  assign n16610 = ~n16590 & ~n16602;
  assign n16611 = ~n16609 & ~n16610;
  assign n16612 = ~n16608 & ~n16611;
  assign n16613 = ~n16605 & ~n16612;
  assign n16614 = ~n16095 & n16613;
  assign n16615 = n16095 & ~n16613;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = n11366 & ~n16616;
  assign n16618 = pi328 & n16617;
  assign n16619 = pi328 & n11366;
  assign n16620 = n16095 & n16613;
  assign n16621 = ~n16095 & ~n16613;
  assign n16622 = ~n16620 & ~n16621;
  assign n16623 = ~n16619 & ~n16622;
  assign n16624 = ~n16618 & ~n16623;
  assign n16625 = ~n16094 & ~n16624;
  assign n16626 = n16078 & n16091;
  assign n16627 = ~n16078 & ~n16091;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = n11366 & ~n16622;
  assign n16630 = pi328 & n16629;
  assign n16631 = ~n16616 & ~n16619;
  assign n16632 = ~n16630 & ~n16631;
  assign n16633 = ~n16628 & ~n16632;
  assign n16634 = ~n16625 & ~n16633;
  assign n16635 = ~n15074 & n15085;
  assign n16636 = n15074 & ~n15085;
  assign n16637 = ~n15745 & ~n16636;
  assign n16638 = ~n16635 & ~n16637;
  assign n16639 = n16634 & n16638;
  assign n16640 = ~n16634 & ~n16638;
  assign n16641 = ~n16639 & ~n16640;
  assign n16642 = pi331 & n6556;
  assign n16643 = n13299 & ~n15067;
  assign n16644 = ~n13299 & ~n15057;
  assign n16645 = ~n16643 & ~n16644;
  assign n16646 = ~n15705 & ~n16645;
  assign n16647 = ~n15708 & ~n16646;
  assign n16648 = n9205 & ~n15699;
  assign n16649 = pi329 & n16648;
  assign n16650 = ~n15724 & ~n15731;
  assign n16651 = ~n16649 & ~n16650;
  assign n16652 = ~n15112 & ~n16651;
  assign n16653 = n9205 & ~n15731;
  assign n16654 = pi329 & n16653;
  assign n16655 = ~n15699 & ~n15724;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = ~n15740 & ~n16656;
  assign n16658 = ~n16652 & ~n16657;
  assign n16659 = n16647 & ~n16658;
  assign n16660 = ~n16647 & n16658;
  assign n16661 = ~n6556 & ~n16660;
  assign n16662 = ~n16659 & ~n16661;
  assign n16663 = n9205 & ~n16662;
  assign n16664 = ~n9205 & ~n16659;
  assign n16665 = n6556 & n16664;
  assign n16666 = ~n16663 & ~n16665;
  assign n16667 = pi330 & ~n16666;
  assign n16668 = pi330 & n9205;
  assign n16669 = n16658 & ~n16668;
  assign n16670 = ~n16647 & n16669;
  assign n16671 = ~n16667 & ~n16670;
  assign n16672 = ~n16642 & n16671;
  assign n16673 = n16642 & ~n16671;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = pi333 & n5732;
  assign n16676 = n5714 & ~n15753;
  assign n16677 = ~n5732 & ~n16676;
  assign n16678 = pi332 & ~n16677;
  assign n16679 = ~n15754 & ~n16678;
  assign n16680 = pi332 & n5973;
  assign n16681 = n15085 & ~n16680;
  assign n16682 = ~n16679 & n16681;
  assign n16683 = ~n15754 & ~n16676;
  assign n16684 = n5732 & ~n16683;
  assign n16685 = pi332 & n16684;
  assign n16686 = ~n15085 & n16680;
  assign n16687 = ~n16685 & n16686;
  assign n16688 = ~n16682 & ~n16687;
  assign n16689 = ~n16034 & ~n16688;
  assign n16690 = n15085 & n16680;
  assign n16691 = ~n16685 & n16690;
  assign n16692 = ~n15085 & ~n16680;
  assign n16693 = ~n16679 & n16692;
  assign n16694 = ~n16691 & ~n16693;
  assign n16695 = ~n16043 & ~n16694;
  assign n16696 = ~n16680 & n16685;
  assign n16697 = n16679 & n16680;
  assign n16698 = ~n16685 & n16697;
  assign n16699 = ~n16696 & ~n16698;
  assign n16700 = ~n16695 & n16699;
  assign n16701 = ~n16689 & n16700;
  assign n16702 = n16675 & ~n16701;
  assign n16703 = ~n16675 & n16701;
  assign n16704 = ~n16702 & ~n16703;
  assign n16705 = ~n16674 & ~n16704;
  assign n16706 = n16642 & n16671;
  assign n16707 = ~n16642 & ~n16671;
  assign n16708 = ~n16706 & ~n16707;
  assign n16709 = ~n16675 & ~n16701;
  assign n16710 = n16675 & n16701;
  assign n16711 = ~n16709 & ~n16710;
  assign n16712 = ~n16708 & ~n16711;
  assign n16713 = ~n16705 & ~n16712;
  assign n16714 = ~n16641 & ~n16713;
  assign n16715 = n16634 & ~n16638;
  assign n16716 = ~n16634 & n16638;
  assign n16717 = ~n16715 & ~n16716;
  assign n16718 = ~n16704 & ~n16708;
  assign n16719 = ~n16674 & ~n16711;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = ~n16717 & ~n16720;
  assign n16722 = ~n16714 & ~n16721;
  assign n16723 = n16074 & n16722;
  assign n16724 = ~n16074 & ~n16722;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = n5257 & ~n16725;
  assign n16727 = pi335 & n16726;
  assign n16728 = pi335 & n5257;
  assign n16729 = ~n16074 & n16722;
  assign n16730 = n16074 & ~n16722;
  assign n16731 = ~n16729 & ~n16730;
  assign n16732 = ~n16728 & ~n16731;
  assign n16733 = ~n16727 & ~n16732;
  assign n16734 = ~n16061 & ~n16733;
  assign n16735 = n16051 & ~n16058;
  assign n16736 = ~n16051 & n16058;
  assign n16737 = ~n16735 & ~n16736;
  assign n16738 = n5257 & ~n16731;
  assign n16739 = pi335 & n16738;
  assign n16740 = ~n16725 & ~n16728;
  assign n16741 = ~n16739 & ~n16740;
  assign n16742 = ~n16737 & ~n16741;
  assign n16743 = ~n16734 & ~n16742;
  assign n16744 = ~n15036 & n15054;
  assign n16745 = n15036 & ~n15054;
  assign n16746 = ~n15842 & ~n16745;
  assign n16747 = ~n16744 & ~n16746;
  assign n16748 = n16743 & n16747;
  assign n16749 = ~n16743 & ~n16747;
  assign n16750 = ~n16748 & ~n16749;
  assign n16751 = pi337 & n2887;
  assign n16752 = ~n15808 & ~n15830;
  assign n16753 = ~n15793 & n16752;
  assign n16754 = ~n15828 & ~n15830;
  assign n16755 = ~n15837 & n16754;
  assign n16756 = ~n15829 & ~n16755;
  assign n16757 = ~n16753 & n16756;
  assign n16758 = pi336 & n4596;
  assign n16759 = n16757 & ~n16758;
  assign n16760 = n4596 & ~n16757;
  assign n16761 = pi336 & n16760;
  assign n16762 = ~n16759 & ~n16761;
  assign n16763 = ~n16751 & n16762;
  assign n16764 = n16751 & ~n16762;
  assign n16765 = ~n16763 & ~n16764;
  assign n16766 = pi339 & n2091;
  assign n16767 = n1729 & ~n15044;
  assign n16768 = ~n2091 & ~n16767;
  assign n16769 = pi338 & ~n16768;
  assign n16770 = ~n15045 & ~n16769;
  assign n16771 = pi338 & n2464;
  assign n16772 = n15054 & ~n16771;
  assign n16773 = ~n16770 & n16772;
  assign n16774 = ~n15045 & ~n16767;
  assign n16775 = n2091 & ~n16774;
  assign n16776 = pi338 & n16775;
  assign n16777 = ~n15054 & n16771;
  assign n16778 = ~n16776 & n16777;
  assign n16779 = ~n16773 & ~n16778;
  assign n16780 = ~n15997 & ~n16779;
  assign n16781 = n15054 & n16771;
  assign n16782 = ~n16776 & n16781;
  assign n16783 = ~n15054 & ~n16771;
  assign n16784 = ~n16770 & n16783;
  assign n16785 = ~n16782 & ~n16784;
  assign n16786 = ~n16006 & ~n16785;
  assign n16787 = ~n16771 & n16776;
  assign n16788 = n16770 & n16771;
  assign n16789 = ~n16776 & n16788;
  assign n16790 = ~n16787 & ~n16789;
  assign n16791 = ~n16786 & n16790;
  assign n16792 = ~n16780 & n16791;
  assign n16793 = n16766 & ~n16792;
  assign n16794 = ~n16766 & n16792;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~n16765 & ~n16795;
  assign n16797 = n16751 & n16762;
  assign n16798 = ~n16751 & ~n16762;
  assign n16799 = ~n16797 & ~n16798;
  assign n16800 = ~n16766 & ~n16792;
  assign n16801 = n16766 & n16792;
  assign n16802 = ~n16800 & ~n16801;
  assign n16803 = ~n16799 & ~n16802;
  assign n16804 = ~n16796 & ~n16803;
  assign n16805 = ~n16750 & ~n16804;
  assign n16806 = n16743 & ~n16747;
  assign n16807 = ~n16743 & n16747;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = ~n16795 & ~n16799;
  assign n16810 = ~n16765 & ~n16802;
  assign n16811 = ~n16809 & ~n16810;
  assign n16812 = ~n16808 & ~n16811;
  assign n16813 = ~n16805 & ~n16812;
  assign n16814 = n16031 & n16813;
  assign n16815 = ~n16031 & ~n16813;
  assign n16816 = ~n16814 & ~n16815;
  assign n16817 = n1442 & ~n16816;
  assign n16818 = pi341 & n16817;
  assign n16819 = pi341 & n1442;
  assign n16820 = ~n16031 & n16813;
  assign n16821 = n16031 & ~n16813;
  assign n16822 = ~n16820 & ~n16821;
  assign n16823 = ~n16819 & ~n16822;
  assign n16824 = ~n16818 & ~n16823;
  assign n16825 = ~n16024 & ~n16824;
  assign n16826 = n16014 & ~n16021;
  assign n16827 = ~n16014 & n16021;
  assign n16828 = ~n16826 & ~n16827;
  assign n16829 = n1442 & ~n16822;
  assign n16830 = pi341 & n16829;
  assign n16831 = ~n16816 & ~n16819;
  assign n16832 = ~n16830 & ~n16831;
  assign n16833 = ~n16828 & ~n16832;
  assign n16834 = ~n16825 & ~n16833;
  assign n16835 = n15994 & ~n16834;
  assign n16836 = ~n15994 & n16834;
  assign n16837 = ~n16835 & ~n16836;
  assign n16838 = pi258 & ~n15932;
  assign n16839 = pi128 & n16838;
  assign n16840 = pi343 & n16839;
  assign n16841 = pi343 & ~n1154;
  assign n16842 = ~n16840 & ~n16841;
  assign n16843 = n16840 & n16841;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = n1156 & ~n16844;
  assign n16846 = pi344 & n16845;
  assign n16847 = pi344 & n1156;
  assign n16848 = n16840 & ~n16841;
  assign n16849 = ~n16840 & n16841;
  assign n16850 = ~n16848 & ~n16849;
  assign n16851 = ~n16847 & ~n16850;
  assign n16852 = ~n16846 & ~n16851;
  assign n16853 = ~n16837 & ~n16852;
  assign n16854 = n15994 & n16834;
  assign n16855 = ~n15994 & ~n16834;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = n1156 & ~n16850;
  assign n16858 = pi344 & n16857;
  assign n16859 = ~n16844 & ~n16847;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = ~n16856 & ~n16860;
  assign n16862 = ~n16853 & ~n16861;
  assign n16863 = n15012 & ~n15958;
  assign n16864 = ~n15012 & n15958;
  assign n16865 = ~n15947 & ~n16864;
  assign n16866 = ~n16863 & ~n16865;
  assign n16867 = n16862 & n16866;
  assign n16868 = ~n16862 & ~n16866;
  assign n16869 = ~n16867 & ~n16868;
  assign n16870 = pi130 & pi301;
  assign n16871 = ~pi129 & ~n16870;
  assign n16872 = pi301 & ~n12284;
  assign n16873 = ~n1514 & n16872;
  assign n16874 = n15001 & ~n16873;
  assign n16875 = ~n16871 & ~n16874;
  assign n16876 = n14552 & ~n16875;
  assign n16877 = ~pi130 & n15001;
  assign n16878 = ~pi129 & n16877;
  assign n16879 = pi130 & ~n15001;
  assign n16880 = pi129 & n16879;
  assign n16881 = ~n16878 & ~n16880;
  assign n16882 = pi128 & ~n16881;
  assign n16883 = ~n14552 & n15001;
  assign n16884 = pi130 & n16883;
  assign n16885 = ~pi130 & ~n15001;
  assign n16886 = pi129 & n16885;
  assign n16887 = ~n16884 & ~n16886;
  assign n16888 = ~pi128 & ~n16887;
  assign n16889 = pi129 & n15001;
  assign n16890 = ~pi129 & ~n15001;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = ~n14552 & ~n16891;
  assign n16893 = pi130 & n16892;
  assign n16894 = ~n16888 & ~n16893;
  assign n16895 = ~n16882 & n16894;
  assign n16896 = pi301 & ~n16895;
  assign n16897 = ~n16876 & ~n16896;
  assign n16898 = n1515 & ~n14988;
  assign n16899 = pi302 & n16898;
  assign n16900 = ~n14572 & n14986;
  assign n16901 = n14572 & ~n14986;
  assign n16902 = ~n16900 & ~n16901;
  assign n16903 = ~n14573 & n14988;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = ~n16899 & ~n16904;
  assign n16906 = n14979 & ~n14983;
  assign n16907 = ~n14979 & n14983;
  assign n16908 = ~n16906 & ~n16907;
  assign n16909 = ~n14569 & ~n16908;
  assign n16910 = ~n14076 & ~n14492;
  assign n16911 = ~n14071 & ~n16910;
  assign n16912 = ~n14564 & ~n16911;
  assign n16913 = n14569 & n16908;
  assign n16914 = ~n16912 & ~n16913;
  assign n16915 = ~n16909 & ~n16914;
  assign n16916 = pi305 & n2183;
  assign n16917 = ~n14965 & ~n14972;
  assign n16918 = ~n14973 & ~n16917;
  assign n16919 = ~n16916 & ~n16918;
  assign n16920 = ~n14968 & ~n14973;
  assign n16921 = ~n14972 & ~n16920;
  assign n16922 = n16916 & ~n16921;
  assign n16923 = ~n16919 & ~n16922;
  assign n16924 = ~n14442 & n14945;
  assign n16925 = ~n14454 & ~n14927;
  assign n16926 = n1840 & n16925;
  assign n16927 = ~n14455 & n14925;
  assign n16928 = n2183 & ~n16927;
  assign n16929 = ~n16926 & ~n16928;
  assign n16930 = pi306 & ~n16929;
  assign n16931 = ~n16924 & ~n16930;
  assign n16932 = ~n14909 & ~n14920;
  assign n16933 = n14909 & n14920;
  assign n16934 = ~n14914 & ~n16933;
  assign n16935 = ~n16932 & ~n16934;
  assign n16936 = pi309 & n4086;
  assign n16937 = ~n14887 & ~n14894;
  assign n16938 = ~n14895 & ~n16937;
  assign n16939 = ~n16936 & ~n16938;
  assign n16940 = ~n14890 & ~n14895;
  assign n16941 = ~n14894 & ~n16940;
  assign n16942 = n16936 & ~n16941;
  assign n16943 = ~n16939 & ~n16942;
  assign n16944 = ~n14820 & ~n14821;
  assign n16945 = n14820 & n14821;
  assign n16946 = ~n14826 & ~n16945;
  assign n16947 = ~n16944 & ~n16946;
  assign n16948 = pi313 & n7044;
  assign n16949 = ~n14799 & ~n14806;
  assign n16950 = ~n14807 & ~n16949;
  assign n16951 = ~n16948 & ~n16950;
  assign n16952 = ~n14802 & ~n14807;
  assign n16953 = ~n14806 & ~n16952;
  assign n16954 = n16948 & ~n16953;
  assign n16955 = ~n16951 & ~n16954;
  assign n16956 = ~n14766 & ~n14767;
  assign n16957 = n14766 & n14767;
  assign n16958 = ~n14302 & ~n16957;
  assign n16959 = ~n14296 & n16958;
  assign n16960 = ~n16956 & ~n16959;
  assign n16961 = ~n14687 & ~n14695;
  assign n16962 = ~n14686 & n14695;
  assign n16963 = ~n14683 & n16962;
  assign n16964 = ~n16961 & ~n16963;
  assign n16965 = ~n14719 & ~n16964;
  assign n16966 = pi146 & pi148;
  assign n16967 = pi147 & n14591;
  assign n16968 = ~n16966 & ~n16967;
  assign n16969 = pi145 & ~n16968;
  assign n16970 = pi147 & pi149;
  assign n16971 = ~n14145 & ~n16970;
  assign n16972 = pi146 & ~n16971;
  assign n16973 = ~pi147 & ~pi149;
  assign n16974 = pi148 & ~n16973;
  assign n16975 = ~n16972 & ~n16974;
  assign n16976 = ~n16969 & n16975;
  assign n16977 = pi150 & n16976;
  assign n16978 = ~pi150 & ~n16976;
  assign n16979 = ~n16977 & ~n16978;
  assign n16980 = pi149 & ~n16979;
  assign n16981 = pi150 & ~n16976;
  assign n16982 = ~pi150 & n16976;
  assign n16983 = ~n16981 & ~n16982;
  assign n16984 = ~pi149 & ~n16983;
  assign n16985 = ~n16980 & ~n16984;
  assign n16986 = pi321 & n16985;
  assign n16987 = ~n14619 & n14625;
  assign n16988 = n14156 & ~n16987;
  assign n16989 = pi320 & n16988;
  assign n16990 = n14618 & ~n14625;
  assign n16991 = pi321 & n16990;
  assign n16992 = ~n16989 & ~n16991;
  assign n16993 = pi320 & n14618;
  assign n16994 = ~n16992 & ~n16993;
  assign n16995 = n14618 & n16992;
  assign n16996 = pi320 & n16995;
  assign n16997 = ~n16994 & ~n16996;
  assign n16998 = ~n16986 & ~n16997;
  assign n16999 = n16992 & ~n16993;
  assign n17000 = n14618 & ~n16992;
  assign n17001 = pi320 & n17000;
  assign n17002 = ~n16999 & ~n17001;
  assign n17003 = n16985 & ~n17002;
  assign n17004 = pi321 & n17003;
  assign n17005 = ~n16998 & ~n17004;
  assign n17006 = pi319 & n14156;
  assign n17007 = ~n17005 & n17006;
  assign n17008 = n17005 & ~n17006;
  assign n17009 = ~n17007 & ~n17008;
  assign n17010 = n14638 & ~n14639;
  assign n17011 = ~n14653 & ~n17010;
  assign n17012 = ~n11998 & n14638;
  assign n17013 = n10908 & ~n17012;
  assign n17014 = pi319 & n17013;
  assign n17015 = ~n17011 & ~n17014;
  assign n17016 = ~n14176 & ~n17015;
  assign n17017 = n11998 & ~n14638;
  assign n17018 = ~n14653 & n17013;
  assign n17019 = ~n17017 & ~n17018;
  assign n17020 = pi319 & ~n17019;
  assign n17021 = ~n17016 & ~n17020;
  assign n17022 = pi318 & n11998;
  assign n17023 = n17021 & n17022;
  assign n17024 = ~n17021 & ~n17022;
  assign n17025 = ~n17023 & ~n17024;
  assign n17026 = ~n17009 & ~n17025;
  assign n17027 = ~n17021 & n17022;
  assign n17028 = n17021 & ~n17022;
  assign n17029 = ~n17027 & ~n17028;
  assign n17030 = ~n17008 & ~n17029;
  assign n17031 = ~n17007 & n17030;
  assign n17032 = ~n17026 & ~n17031;
  assign n17033 = n14588 & ~n14664;
  assign n17034 = n14677 & ~n17033;
  assign n17035 = n17032 & n17034;
  assign n17036 = ~n17032 & ~n17034;
  assign n17037 = ~n17035 & ~n17036;
  assign n17038 = pi317 & n10908;
  assign n17039 = ~n14686 & ~n14695;
  assign n17040 = ~n17038 & ~n17039;
  assign n17041 = ~n14683 & n17040;
  assign n17042 = ~n14683 & ~n17039;
  assign n17043 = n17038 & ~n17042;
  assign n17044 = ~n17041 & ~n17043;
  assign n17045 = ~n17037 & ~n17044;
  assign n17046 = n17032 & ~n17034;
  assign n17047 = ~n17032 & n17034;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = n17038 & ~n17039;
  assign n17050 = ~n14683 & n17049;
  assign n17051 = ~n17038 & ~n17042;
  assign n17052 = ~n17050 & ~n17051;
  assign n17053 = ~n17048 & ~n17052;
  assign n17054 = ~n17045 & ~n17053;
  assign n17055 = ~pi316 & ~n17054;
  assign n17056 = ~n9815 & ~n17054;
  assign n17057 = n9815 & n17054;
  assign n17058 = pi316 & n17057;
  assign n17059 = ~n17056 & ~n17058;
  assign n17060 = ~n9517 & ~n17059;
  assign n17061 = ~n17055 & ~n17060;
  assign n17062 = ~n16965 & ~n17061;
  assign n17063 = n14719 & n17054;
  assign n17064 = n16964 & n17063;
  assign n17065 = ~n14719 & ~n17054;
  assign n17066 = ~n16964 & n17065;
  assign n17067 = ~n17064 & ~n17066;
  assign n17068 = pi316 & ~n17067;
  assign n17069 = n14719 & ~n16964;
  assign n17070 = ~n14719 & n16964;
  assign n17071 = ~n17069 & ~n17070;
  assign n17072 = ~n17054 & ~n17071;
  assign n17073 = n9517 & n17072;
  assign n17074 = ~n17068 & ~n17073;
  assign n17075 = n9815 & ~n17074;
  assign n17076 = n14719 & ~n17054;
  assign n17077 = n16964 & n17076;
  assign n17078 = n14719 & n16964;
  assign n17079 = n9517 & ~n17078;
  assign n17080 = pi316 & n17079;
  assign n17081 = ~n16965 & ~n17080;
  assign n17082 = n17054 & ~n17081;
  assign n17083 = ~n17077 & ~n17082;
  assign n17084 = ~n9815 & ~n17083;
  assign n17085 = ~pi316 & ~n16964;
  assign n17086 = ~n14719 & n17054;
  assign n17087 = n17085 & n17086;
  assign n17088 = ~n17084 & ~n17087;
  assign n17089 = ~n17075 & n17088;
  assign n17090 = ~n17062 & n17089;
  assign n17091 = n14725 & ~n14728;
  assign n17092 = ~n14291 & ~n14760;
  assign n17093 = n14291 & n14760;
  assign n17094 = n14263 & ~n17093;
  assign n17095 = ~n17092 & ~n17094;
  assign n17096 = ~n14725 & n14728;
  assign n17097 = ~n17095 & ~n17096;
  assign n17098 = ~n17091 & ~n17097;
  assign n17099 = n17090 & n17098;
  assign n17100 = ~n17090 & ~n17098;
  assign n17101 = ~n17099 & ~n17100;
  assign n17102 = n9517 & ~n17101;
  assign n17103 = pi315 & n17102;
  assign n17104 = pi315 & n9517;
  assign n17105 = ~n17090 & n17098;
  assign n17106 = n17090 & ~n17098;
  assign n17107 = ~n17105 & ~n17106;
  assign n17108 = ~n17104 & ~n17107;
  assign n17109 = ~n17103 & ~n17108;
  assign n17110 = n7874 & ~n17109;
  assign n17111 = pi314 & n17110;
  assign n17112 = pi314 & n7874;
  assign n17113 = ~n17108 & ~n17112;
  assign n17114 = ~n17103 & n17113;
  assign n17115 = ~n17111 & ~n17114;
  assign n17116 = ~n16960 & ~n17115;
  assign n17117 = n16960 & ~n17114;
  assign n17118 = ~n17111 & n17117;
  assign n17119 = ~n17116 & ~n17118;
  assign n17120 = n16955 & ~n17119;
  assign n17121 = ~n16955 & n17119;
  assign n17122 = ~n17120 & ~n17121;
  assign n17123 = pi312 & n6777;
  assign n17124 = ~n5463 & ~n6777;
  assign n17125 = pi313 & ~n17124;
  assign n17126 = n14782 & ~n17125;
  assign n17127 = ~n5463 & n6777;
  assign n17128 = pi313 & ~n14782;
  assign n17129 = n17127 & n17128;
  assign n17130 = ~n17126 & ~n17129;
  assign n17131 = ~n14796 & ~n17130;
  assign n17132 = ~n6777 & n14782;
  assign n17133 = ~n14784 & ~n17132;
  assign n17134 = ~n14304 & ~n17133;
  assign n17135 = n14795 & n17134;
  assign n17136 = n5463 & ~n6777;
  assign n17137 = ~n14782 & n17136;
  assign n17138 = ~n5463 & ~n14304;
  assign n17139 = n6777 & ~n17138;
  assign n17140 = n14782 & n17139;
  assign n17141 = ~n17137 & ~n17140;
  assign n17142 = pi313 & ~n17141;
  assign n17143 = n14304 & n14806;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = ~n14795 & ~n17144;
  assign n17146 = ~n6777 & ~n14782;
  assign n17147 = n6777 & n14782;
  assign n17148 = ~n17146 & ~n17147;
  assign n17149 = n5463 & ~n17148;
  assign n17150 = pi313 & n17149;
  assign n17151 = n14304 & n17150;
  assign n17152 = ~n17145 & ~n17151;
  assign n17153 = ~n17135 & n17152;
  assign n17154 = ~n17131 & n17153;
  assign n17155 = ~n14817 & ~n17154;
  assign n17156 = n14817 & n17154;
  assign n17157 = n14786 & ~n17156;
  assign n17158 = ~n17155 & ~n17157;
  assign n17159 = n17123 & ~n17158;
  assign n17160 = ~n14786 & ~n17155;
  assign n17161 = ~n17156 & ~n17160;
  assign n17162 = ~n17123 & ~n17161;
  assign n17163 = ~n17159 & ~n17162;
  assign n17164 = ~n17122 & ~n17163;
  assign n17165 = n16955 & n17119;
  assign n17166 = ~n16955 & ~n17119;
  assign n17167 = ~n17165 & ~n17166;
  assign n17168 = ~n17123 & ~n17158;
  assign n17169 = n17123 & ~n17161;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = ~n17167 & ~n17170;
  assign n17172 = ~n17164 & ~n17171;
  assign n17173 = n16947 & ~n17172;
  assign n17174 = ~n16947 & n17172;
  assign n17175 = ~n17173 & ~n17174;
  assign n17176 = n5463 & ~n17175;
  assign n17177 = pi311 & n17176;
  assign n17178 = pi311 & n5463;
  assign n17179 = ~n16947 & ~n17172;
  assign n17180 = n16947 & n17172;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = ~n17178 & ~n17181;
  assign n17183 = ~n17177 & ~n17182;
  assign n17184 = ~n4086 & ~n14837;
  assign n17185 = ~n14372 & ~n17184;
  assign n17186 = n3552 & n17185;
  assign n17187 = ~n14371 & ~n14837;
  assign n17188 = n4086 & ~n17187;
  assign n17189 = ~n17186 & ~n17188;
  assign n17190 = pi310 & ~n17189;
  assign n17191 = ~n14847 & ~n17190;
  assign n17192 = n17183 & ~n17191;
  assign n17193 = ~n17183 & n17191;
  assign n17194 = ~n17192 & ~n17193;
  assign n17195 = n4772 & ~n17194;
  assign n17196 = pi310 & n17195;
  assign n17197 = pi310 & n4772;
  assign n17198 = ~n17183 & ~n17191;
  assign n17199 = n17183 & n17191;
  assign n17200 = ~n17198 & ~n17199;
  assign n17201 = ~n17197 & ~n17200;
  assign n17202 = ~n17196 & ~n17201;
  assign n17203 = n16943 & n17202;
  assign n17204 = ~n16943 & ~n17202;
  assign n17205 = ~n17203 & ~n17204;
  assign n17206 = pi308 & n3552;
  assign n17207 = pi309 & ~n11042;
  assign n17208 = n14869 & ~n17207;
  assign n17209 = pi309 & ~n14869;
  assign n17210 = n11045 & n17209;
  assign n17211 = ~n17208 & ~n17210;
  assign n17212 = ~n14884 & ~n17211;
  assign n17213 = ~n3552 & n14869;
  assign n17214 = ~n14895 & ~n17213;
  assign n17215 = n14381 & ~n17214;
  assign n17216 = n14883 & n17215;
  assign n17217 = n11054 & ~n14869;
  assign n17218 = ~n3012 & n14381;
  assign n17219 = n3552 & ~n17218;
  assign n17220 = n14869 & n17219;
  assign n17221 = ~n17217 & ~n17220;
  assign n17222 = pi309 & ~n17221;
  assign n17223 = ~n14381 & n14870;
  assign n17224 = ~n17222 & ~n17223;
  assign n17225 = ~n14883 & ~n17224;
  assign n17226 = ~n3552 & ~n14869;
  assign n17227 = n3552 & n14869;
  assign n17228 = ~n17226 & ~n17227;
  assign n17229 = n3012 & ~n17228;
  assign n17230 = pi309 & n17229;
  assign n17231 = ~n14381 & n17230;
  assign n17232 = ~n17225 & ~n17231;
  assign n17233 = ~n17216 & n17232;
  assign n17234 = ~n17212 & n17233;
  assign n17235 = n14905 & n17234;
  assign n17236 = ~n14905 & ~n17234;
  assign n17237 = n14873 & ~n17236;
  assign n17238 = ~n17235 & ~n17237;
  assign n17239 = n17206 & ~n17238;
  assign n17240 = ~n14873 & ~n17235;
  assign n17241 = ~n17236 & ~n17240;
  assign n17242 = ~n17206 & ~n17241;
  assign n17243 = ~n17239 & ~n17242;
  assign n17244 = ~n17205 & ~n17243;
  assign n17245 = n16943 & ~n17202;
  assign n17246 = ~n16943 & n17202;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = ~n17206 & ~n17238;
  assign n17249 = n17206 & ~n17241;
  assign n17250 = ~n17248 & ~n17249;
  assign n17251 = ~n17247 & ~n17250;
  assign n17252 = ~n17244 & ~n17251;
  assign n17253 = n16935 & n17252;
  assign n17254 = ~n16935 & ~n17252;
  assign n17255 = ~n17253 & ~n17254;
  assign n17256 = n3012 & ~n17255;
  assign n17257 = pi307 & n17256;
  assign n17258 = pi307 & n3012;
  assign n17259 = ~n16935 & n17252;
  assign n17260 = n16935 & ~n17252;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = ~n17258 & ~n17261;
  assign n17263 = ~n17257 & ~n17262;
  assign n17264 = n2574 & ~n17263;
  assign n17265 = pi306 & n17264;
  assign n17266 = pi306 & n2574;
  assign n17267 = ~n17262 & ~n17266;
  assign n17268 = ~n17257 & n17267;
  assign n17269 = ~n17265 & ~n17268;
  assign n17270 = n16931 & ~n17269;
  assign n17271 = ~n16931 & ~n17268;
  assign n17272 = ~n17265 & n17271;
  assign n17273 = ~n17270 & ~n17272;
  assign n17274 = n16923 & n17273;
  assign n17275 = ~n16923 & ~n17273;
  assign n17276 = ~n17274 & ~n17275;
  assign n17277 = pi304 & n1840;
  assign n17278 = pi305 & n14957;
  assign n17279 = n6886 & n17278;
  assign n17280 = pi305 & ~n6883;
  assign n17281 = ~n14957 & ~n17280;
  assign n17282 = ~n17279 & ~n17281;
  assign n17283 = ~n14962 & ~n17282;
  assign n17284 = ~n1840 & ~n14957;
  assign n17285 = ~n14973 & ~n17284;
  assign n17286 = ~n14458 & ~n17285;
  assign n17287 = n14081 & n17286;
  assign n17288 = n1840 & ~n14957;
  assign n17289 = ~n1840 & n14957;
  assign n17290 = ~n17288 & ~n17289;
  assign n17291 = n1533 & ~n17290;
  assign n17292 = pi305 & n17291;
  assign n17293 = n14458 & n17292;
  assign n17294 = ~n1533 & ~n14458;
  assign n17295 = n1840 & ~n17294;
  assign n17296 = ~n14957 & n17295;
  assign n17297 = n6897 & n14957;
  assign n17298 = ~n17296 & ~n17297;
  assign n17299 = pi305 & ~n17298;
  assign n17300 = n14458 & n14958;
  assign n17301 = ~n17299 & ~n17300;
  assign n17302 = ~n14081 & ~n17301;
  assign n17303 = ~n17293 & ~n17302;
  assign n17304 = ~n17287 & n17303;
  assign n17305 = ~n17283 & n17304;
  assign n17306 = n14983 & n17305;
  assign n17307 = ~n14983 & ~n17305;
  assign n17308 = n14961 & ~n17307;
  assign n17309 = ~n17306 & ~n17308;
  assign n17310 = n17277 & ~n17309;
  assign n17311 = ~n14961 & ~n17306;
  assign n17312 = ~n17307 & ~n17311;
  assign n17313 = ~n17277 & ~n17312;
  assign n17314 = ~n17310 & ~n17313;
  assign n17315 = ~n17276 & ~n17314;
  assign n17316 = n16923 & ~n17273;
  assign n17317 = ~n16923 & n17273;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = ~n17277 & ~n17309;
  assign n17320 = n17277 & ~n17312;
  assign n17321 = ~n17319 & ~n17320;
  assign n17322 = ~n17318 & ~n17321;
  assign n17323 = ~n17315 & ~n17322;
  assign n17324 = ~n16915 & n17323;
  assign n17325 = n16915 & ~n17323;
  assign n17326 = ~n17324 & ~n17325;
  assign n17327 = n1533 & ~n17326;
  assign n17328 = pi303 & n17327;
  assign n17329 = pi303 & n1533;
  assign n17330 = n16915 & n17323;
  assign n17331 = ~n16915 & ~n17323;
  assign n17332 = ~n17330 & ~n17331;
  assign n17333 = ~n17329 & ~n17332;
  assign n17334 = ~n17328 & ~n17333;
  assign n17335 = n1553 & ~n17334;
  assign n17336 = pi302 & n17335;
  assign n17337 = pi302 & n1553;
  assign n17338 = ~n17333 & ~n17337;
  assign n17339 = ~n17328 & n17338;
  assign n17340 = ~n17336 & ~n17339;
  assign n17341 = n16905 & ~n17340;
  assign n17342 = ~n16905 & ~n17339;
  assign n17343 = ~n17336 & n17342;
  assign n17344 = ~n17341 & ~n17343;
  assign n17345 = n16897 & ~n17344;
  assign n17346 = ~n16897 & n17344;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = pi300 & ~n15010;
  assign n17349 = pi128 & n17348;
  assign n17350 = pi300 & ~n1568;
  assign n17351 = ~n17349 & ~n17350;
  assign n17352 = n17349 & n17350;
  assign n17353 = ~n17351 & ~n17352;
  assign n17354 = pi299 & ~n17353;
  assign n17355 = pi128 & n17354;
  assign n17356 = pi128 & pi299;
  assign n17357 = n17349 & ~n17350;
  assign n17358 = ~n17349 & n17350;
  assign n17359 = ~n17357 & ~n17358;
  assign n17360 = ~n17356 & ~n17359;
  assign n17361 = ~n17355 & ~n17360;
  assign n17362 = ~n17347 & ~n17361;
  assign n17363 = n16897 & n17344;
  assign n17364 = ~n16897 & ~n17344;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = pi299 & ~n17359;
  assign n17367 = pi128 & n17366;
  assign n17368 = ~n17353 & ~n17356;
  assign n17369 = ~n17367 & ~n17368;
  assign n17370 = ~n17365 & ~n17369;
  assign n17371 = ~n17362 & ~n17370;
  assign n17372 = ~pi279 & ~n15016;
  assign n17373 = pi279 & n15016;
  assign n17374 = ~n15932 & ~n15942;
  assign n17375 = pi343 & n15932;
  assign n17376 = n1156 & n17375;
  assign n17377 = ~n17374 & ~n17376;
  assign n17378 = ~n17373 & ~n17377;
  assign n17379 = ~n17372 & ~n17378;
  assign n17380 = n17371 & n17379;
  assign n17381 = ~n17371 & ~n17379;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = pi280 & ~n17382;
  assign n17384 = ~n17371 & n17379;
  assign n17385 = n17371 & ~n17379;
  assign n17386 = ~n17384 & ~n17385;
  assign n17387 = ~pi280 & ~n17386;
  assign n17388 = ~n17383 & ~n17387;
  assign n17389 = ~n16869 & ~n17388;
  assign n17390 = n16862 & ~n16866;
  assign n17391 = ~n16862 & n16866;
  assign n17392 = ~n17390 & ~n17391;
  assign n17393 = pi280 & ~n17386;
  assign n17394 = ~pi280 & ~n17382;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = ~n17392 & ~n17395;
  assign n17397 = ~n17389 & ~n17396;
  assign n17398 = ~n831 & ~n17397;
  assign n17399 = ~pi280 & n831;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = pi161 & n17400;
  assign n17402 = ~n15967 & ~n17401;
  assign po215 = ~pi160 & ~n17402;
  assign n17404 = ~pi087 & ~pi161;
  assign n17405 = ~pi281 & n831;
  assign n17406 = pi301 & n1553;
  assign n17407 = ~n1533 & n17323;
  assign n17408 = n1533 & ~n17323;
  assign n17409 = ~n16915 & ~n17408;
  assign n17410 = ~n17407 & ~n17409;
  assign n17411 = n1840 & ~n17410;
  assign n17412 = ~n1840 & ~n17324;
  assign n17413 = n1533 & n17412;
  assign n17414 = ~n17411 & ~n17413;
  assign n17415 = pi303 & ~n17414;
  assign n17416 = pi303 & n1840;
  assign n17417 = ~n17323 & ~n17416;
  assign n17418 = n16915 & n17417;
  assign n17419 = ~n17415 & ~n17418;
  assign n17420 = pi305 & n2574;
  assign n17421 = ~n3012 & ~n17252;
  assign n17422 = n3012 & n17252;
  assign n17423 = ~n16935 & ~n17422;
  assign n17424 = ~n17421 & ~n17423;
  assign n17425 = n3552 & ~n17424;
  assign n17426 = ~n3552 & ~n17254;
  assign n17427 = n3012 & n17426;
  assign n17428 = ~n17425 & ~n17427;
  assign n17429 = pi307 & ~n17428;
  assign n17430 = pi307 & n3552;
  assign n17431 = n17252 & ~n17430;
  assign n17432 = n16935 & n17431;
  assign n17433 = ~n17429 & ~n17432;
  assign n17434 = pi309 & n4772;
  assign n17435 = pi313 & n7874;
  assign n17436 = ~n14638 & n14639;
  assign n17437 = n14177 & ~n14655;
  assign n17438 = ~n14654 & ~n17437;
  assign n17439 = ~n17010 & ~n17438;
  assign n17440 = ~n17436 & ~n17439;
  assign n17441 = ~n17008 & ~n17440;
  assign n17442 = ~n17007 & ~n17441;
  assign n17443 = ~pi151 & n16976;
  assign n17444 = pi151 & ~n16976;
  assign n17445 = ~pi150 & n17444;
  assign n17446 = ~n17443 & ~n17445;
  assign n17447 = pi149 & ~n17446;
  assign n17448 = ~pi151 & ~n16976;
  assign n17449 = pi151 & n16976;
  assign n17450 = pi150 & n17449;
  assign n17451 = ~n17448 & ~n17450;
  assign n17452 = ~pi149 & ~n17451;
  assign n17453 = ~pi151 & ~n16983;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = ~n17447 & n17454;
  assign n17456 = pi321 & n17455;
  assign n17457 = ~n16986 & n16992;
  assign n17458 = n14618 & ~n17457;
  assign n17459 = pi320 & n17458;
  assign n17460 = n16985 & ~n16992;
  assign n17461 = pi321 & n17460;
  assign n17462 = ~n17459 & ~n17461;
  assign n17463 = pi320 & n16985;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = n16985 & n17462;
  assign n17466 = pi320 & n17465;
  assign n17467 = ~n17464 & ~n17466;
  assign n17468 = ~n17456 & ~n17467;
  assign n17469 = n17462 & ~n17463;
  assign n17470 = n16985 & ~n17462;
  assign n17471 = pi320 & n17470;
  assign n17472 = ~n17469 & ~n17471;
  assign n17473 = n17455 & ~n17472;
  assign n17474 = pi321 & n17473;
  assign n17475 = ~n17468 & ~n17474;
  assign n17476 = pi319 & n14618;
  assign n17477 = ~n17475 & n17476;
  assign n17478 = n17475 & ~n17476;
  assign n17479 = ~n17477 & ~n17478;
  assign n17480 = ~n17442 & ~n17479;
  assign n17481 = n17442 & n17479;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = n14156 & ~n17482;
  assign n17484 = pi318 & n17483;
  assign n17485 = pi318 & n14156;
  assign n17486 = ~n17481 & ~n17485;
  assign n17487 = ~n17480 & n17486;
  assign n17488 = ~n17009 & ~n17021;
  assign n17489 = n17009 & n17021;
  assign n17490 = ~n17488 & ~n17489;
  assign n17491 = n17022 & ~n17490;
  assign n17492 = ~n17022 & n17490;
  assign n17493 = ~n17033 & ~n17492;
  assign n17494 = n14677 & n17493;
  assign n17495 = ~n17491 & ~n17494;
  assign n17496 = ~n17487 & n17495;
  assign n17497 = ~n17484 & n17496;
  assign n17498 = ~n17484 & ~n17487;
  assign n17499 = ~n17495 & ~n17498;
  assign n17500 = ~n17497 & ~n17499;
  assign n17501 = n11998 & ~n17500;
  assign n17502 = pi317 & n17501;
  assign n17503 = pi317 & n11998;
  assign n17504 = ~n17497 & ~n17503;
  assign n17505 = ~n17499 & n17504;
  assign n17506 = ~n17502 & ~n17505;
  assign n17507 = ~n17038 & ~n17048;
  assign n17508 = n17038 & n17048;
  assign n17509 = ~n17039 & ~n17508;
  assign n17510 = ~n14683 & n17509;
  assign n17511 = ~n17507 & ~n17510;
  assign n17512 = pi316 & n10908;
  assign n17513 = n17511 & ~n17512;
  assign n17514 = n10908 & ~n17511;
  assign n17515 = pi316 & n17514;
  assign n17516 = ~n17513 & ~n17515;
  assign n17517 = ~n17506 & ~n17516;
  assign n17518 = ~n17511 & ~n17512;
  assign n17519 = n10908 & n17511;
  assign n17520 = pi316 & n17519;
  assign n17521 = ~n17518 & ~n17520;
  assign n17522 = ~n17505 & ~n17521;
  assign n17523 = ~n17502 & n17522;
  assign n17524 = ~n17517 & ~n17523;
  assign n17525 = ~n9815 & n17054;
  assign n17526 = ~n17078 & ~n17525;
  assign n17527 = n9517 & n17526;
  assign n17528 = ~n16965 & n17054;
  assign n17529 = n9815 & ~n17528;
  assign n17530 = ~n17527 & ~n17529;
  assign n17531 = pi316 & ~n17530;
  assign n17532 = ~n17066 & ~n17531;
  assign n17533 = n17524 & n17532;
  assign n17534 = ~n17524 & ~n17532;
  assign n17535 = ~n17533 & ~n17534;
  assign n17536 = n9815 & ~n17535;
  assign n17537 = pi315 & n17536;
  assign n17538 = pi315 & n9815;
  assign n17539 = ~n17524 & n17532;
  assign n17540 = n17524 & ~n17532;
  assign n17541 = ~n17539 & ~n17540;
  assign n17542 = ~n17538 & ~n17541;
  assign n17543 = ~n17537 & ~n17542;
  assign n17544 = ~n17098 & n17104;
  assign n17545 = n17098 & ~n17104;
  assign n17546 = ~n17090 & ~n17545;
  assign n17547 = ~n17544 & ~n17546;
  assign n17548 = n17543 & n17547;
  assign n17549 = ~n17543 & ~n17547;
  assign n17550 = ~n17548 & ~n17549;
  assign n17551 = pi314 & n9517;
  assign n17552 = ~n17117 & ~n17551;
  assign n17553 = ~n17111 & n17552;
  assign n17554 = ~n17111 & ~n17117;
  assign n17555 = n17551 & ~n17554;
  assign n17556 = ~n17553 & ~n17555;
  assign n17557 = ~n17550 & ~n17556;
  assign n17558 = n17543 & ~n17547;
  assign n17559 = ~n17543 & n17547;
  assign n17560 = ~n17558 & ~n17559;
  assign n17561 = ~n17117 & n17551;
  assign n17562 = ~n17111 & n17561;
  assign n17563 = ~n17551 & ~n17554;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = ~n17560 & ~n17564;
  assign n17566 = ~n17557 & ~n17565;
  assign n17567 = ~n17435 & n17566;
  assign n17568 = n17435 & ~n17566;
  assign n17569 = ~n17567 & ~n17568;
  assign n17570 = pi312 & n7044;
  assign n17571 = n14304 & ~n14806;
  assign n17572 = n5463 & ~n17146;
  assign n17573 = pi313 & n17572;
  assign n17574 = ~n17571 & ~n17573;
  assign n17575 = ~n14795 & ~n17574;
  assign n17576 = n14304 & n17572;
  assign n17577 = ~n17147 & ~n17576;
  assign n17578 = pi313 & ~n17577;
  assign n17579 = ~n17575 & ~n17578;
  assign n17580 = n17119 & ~n17579;
  assign n17581 = ~n17119 & n17579;
  assign n17582 = n16948 & ~n17581;
  assign n17583 = ~n17580 & ~n17582;
  assign n17584 = n17570 & ~n17583;
  assign n17585 = ~n16948 & ~n17580;
  assign n17586 = ~n17581 & ~n17585;
  assign n17587 = ~n17570 & ~n17586;
  assign n17588 = ~n17584 & ~n17587;
  assign n17589 = ~n17569 & ~n17588;
  assign n17590 = ~n17435 & ~n17566;
  assign n17591 = n17435 & n17566;
  assign n17592 = ~n17590 & ~n17591;
  assign n17593 = ~n17570 & ~n17583;
  assign n17594 = n17570 & ~n17586;
  assign n17595 = ~n17593 & ~n17594;
  assign n17596 = ~n17592 & ~n17595;
  assign n17597 = ~n17589 & ~n17596;
  assign n17598 = n17123 & ~n17167;
  assign n17599 = ~n17123 & n17167;
  assign n17600 = ~n17158 & ~n17599;
  assign n17601 = ~n17598 & ~n17600;
  assign n17602 = n17597 & n17601;
  assign n17603 = ~n17597 & ~n17601;
  assign n17604 = ~n17602 & ~n17603;
  assign n17605 = pi311 & n6777;
  assign n17606 = n17178 & ~n17179;
  assign n17607 = ~n17180 & ~n17606;
  assign n17608 = n17605 & ~n17607;
  assign n17609 = ~n17178 & ~n17180;
  assign n17610 = ~n17179 & ~n17609;
  assign n17611 = ~n17605 & ~n17610;
  assign n17612 = ~n17608 & ~n17611;
  assign n17613 = ~n17604 & ~n17612;
  assign n17614 = n17597 & ~n17601;
  assign n17615 = ~n17597 & n17601;
  assign n17616 = ~n17614 & ~n17615;
  assign n17617 = ~n17605 & ~n17607;
  assign n17618 = n17605 & ~n17610;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = ~n17616 & ~n17619;
  assign n17621 = ~n17613 & ~n17620;
  assign n17622 = ~pi310 & n17621;
  assign n17623 = ~n5463 & n17621;
  assign n17624 = n5463 & ~n17621;
  assign n17625 = pi310 & n17624;
  assign n17626 = ~n17623 & ~n17625;
  assign n17627 = ~n4772 & ~n17626;
  assign n17628 = ~n17622 & ~n17627;
  assign n17629 = ~n17192 & ~n17628;
  assign n17630 = ~n17191 & n17621;
  assign n17631 = n17183 & n17630;
  assign n17632 = n17191 & ~n17621;
  assign n17633 = ~n17183 & n17632;
  assign n17634 = ~n17631 & ~n17633;
  assign n17635 = pi310 & ~n17634;
  assign n17636 = ~n17200 & n17621;
  assign n17637 = n4772 & n17636;
  assign n17638 = ~n17635 & ~n17637;
  assign n17639 = n5463 & ~n17638;
  assign n17640 = ~n17191 & ~n17621;
  assign n17641 = ~pi310 & n17183;
  assign n17642 = n17640 & n17641;
  assign n17643 = n17191 & n17621;
  assign n17644 = ~n17183 & n17643;
  assign n17645 = n4772 & ~n17193;
  assign n17646 = pi310 & n17645;
  assign n17647 = ~n17192 & ~n17646;
  assign n17648 = ~n17621 & ~n17647;
  assign n17649 = ~n17644 & ~n17648;
  assign n17650 = ~n5463 & ~n17649;
  assign n17651 = ~n17642 & ~n17650;
  assign n17652 = ~n17639 & n17651;
  assign n17653 = ~n17629 & n17652;
  assign n17654 = ~n17434 & ~n17653;
  assign n17655 = n17434 & n17653;
  assign n17656 = ~n17654 & ~n17655;
  assign n17657 = pi308 & n4086;
  assign n17658 = n3012 & ~n17213;
  assign n17659 = pi309 & n17658;
  assign n17660 = ~n14381 & ~n14894;
  assign n17661 = ~n17659 & ~n17660;
  assign n17662 = ~n14883 & ~n17661;
  assign n17663 = n3552 & ~n14869;
  assign n17664 = ~n14381 & n17658;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = pi309 & ~n17665;
  assign n17667 = ~n17662 & ~n17666;
  assign n17668 = ~n17202 & ~n17667;
  assign n17669 = n17202 & n17667;
  assign n17670 = n16936 & ~n17669;
  assign n17671 = ~n17668 & ~n17670;
  assign n17672 = n17657 & ~n17671;
  assign n17673 = ~n16936 & ~n17668;
  assign n17674 = ~n17669 & ~n17673;
  assign n17675 = ~n17657 & ~n17674;
  assign n17676 = ~n17672 & ~n17675;
  assign n17677 = ~n17656 & ~n17676;
  assign n17678 = ~n17434 & n17653;
  assign n17679 = n17434 & ~n17653;
  assign n17680 = ~n17678 & ~n17679;
  assign n17681 = ~n17657 & ~n17671;
  assign n17682 = n17657 & ~n17674;
  assign n17683 = ~n17681 & ~n17682;
  assign n17684 = ~n17680 & ~n17683;
  assign n17685 = ~n17677 & ~n17684;
  assign n17686 = ~n17205 & ~n17206;
  assign n17687 = n17205 & n17206;
  assign n17688 = ~n17241 & ~n17687;
  assign n17689 = ~n17686 & ~n17688;
  assign n17690 = n17685 & ~n17689;
  assign n17691 = ~n17685 & n17689;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 = n17433 & ~n17692;
  assign n17694 = ~n17433 & n17692;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = pi306 & n3012;
  assign n17697 = n16931 & ~n17265;
  assign n17698 = n17696 & ~n17697;
  assign n17699 = ~n17268 & n17698;
  assign n17700 = ~n17268 & ~n17697;
  assign n17701 = ~n17696 & ~n17700;
  assign n17702 = ~n17699 & ~n17701;
  assign n17703 = ~n17695 & ~n17702;
  assign n17704 = n17433 & n17692;
  assign n17705 = ~n17433 & ~n17692;
  assign n17706 = ~n17704 & ~n17705;
  assign n17707 = ~n17696 & ~n17697;
  assign n17708 = ~n17268 & n17707;
  assign n17709 = n17696 & ~n17700;
  assign n17710 = ~n17708 & ~n17709;
  assign n17711 = ~n17706 & ~n17710;
  assign n17712 = ~n17703 & ~n17711;
  assign n17713 = ~n17420 & n17712;
  assign n17714 = n17420 & ~n17712;
  assign n17715 = ~n17713 & ~n17714;
  assign n17716 = pi304 & n2183;
  assign n17717 = n14458 & ~n14972;
  assign n17718 = n1533 & ~n17284;
  assign n17719 = pi305 & n17718;
  assign n17720 = ~n17717 & ~n17719;
  assign n17721 = ~n14081 & ~n17720;
  assign n17722 = n1840 & n14957;
  assign n17723 = n14458 & n17718;
  assign n17724 = ~n17722 & ~n17723;
  assign n17725 = pi305 & ~n17724;
  assign n17726 = ~n17721 & ~n17725;
  assign n17727 = n17273 & ~n17726;
  assign n17728 = ~n17273 & n17726;
  assign n17729 = n16916 & ~n17728;
  assign n17730 = ~n17727 & ~n17729;
  assign n17731 = n17716 & ~n17730;
  assign n17732 = ~n16916 & ~n17727;
  assign n17733 = ~n17728 & ~n17732;
  assign n17734 = ~n17716 & ~n17733;
  assign n17735 = ~n17731 & ~n17734;
  assign n17736 = ~n17715 & ~n17735;
  assign n17737 = ~n17420 & ~n17712;
  assign n17738 = n17420 & n17712;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = ~n17716 & ~n17730;
  assign n17741 = n17716 & ~n17733;
  assign n17742 = ~n17740 & ~n17741;
  assign n17743 = ~n17739 & ~n17742;
  assign n17744 = ~n17736 & ~n17743;
  assign n17745 = ~n17277 & ~n17318;
  assign n17746 = n17277 & n17318;
  assign n17747 = ~n17312 & ~n17746;
  assign n17748 = ~n17745 & ~n17747;
  assign n17749 = ~n17744 & ~n17748;
  assign n17750 = n17744 & n17748;
  assign n17751 = ~n17749 & ~n17750;
  assign n17752 = n17419 & n17751;
  assign n17753 = ~n17419 & ~n17751;
  assign n17754 = ~n17752 & ~n17753;
  assign n17755 = pi302 & n1533;
  assign n17756 = ~n17342 & ~n17755;
  assign n17757 = ~n17336 & n17756;
  assign n17758 = ~n17336 & ~n17342;
  assign n17759 = n17755 & ~n17758;
  assign n17760 = ~n17757 & ~n17759;
  assign n17761 = ~n17754 & ~n17760;
  assign n17762 = n17419 & ~n17751;
  assign n17763 = ~n17419 & n17751;
  assign n17764 = ~n17762 & ~n17763;
  assign n17765 = ~n17342 & n17755;
  assign n17766 = ~n17336 & n17765;
  assign n17767 = ~n17755 & ~n17758;
  assign n17768 = ~n17766 & ~n17767;
  assign n17769 = ~n17764 & ~n17768;
  assign n17770 = ~n17761 & ~n17769;
  assign n17771 = ~n17406 & n17770;
  assign n17772 = n17406 & ~n17770;
  assign n17773 = ~n17771 & ~n17772;
  assign n17774 = n1335 & n16877;
  assign n17775 = ~pi129 & n14552;
  assign n17776 = pi129 & ~n14552;
  assign n17777 = n15001 & ~n17776;
  assign n17778 = pi128 & n17777;
  assign n17779 = ~n17775 & ~n17778;
  assign n17780 = pi130 & ~n17779;
  assign n17781 = ~n17774 & ~n17780;
  assign n17782 = pi301 & ~n17781;
  assign n17783 = pi300 & n1515;
  assign n17784 = n14552 & n15001;
  assign n17785 = ~pi130 & ~n17784;
  assign n17786 = pi128 & n17785;
  assign n17787 = pi301 & ~n11201;
  assign n17788 = ~n15001 & ~n17787;
  assign n17789 = ~n17786 & ~n17788;
  assign n17790 = pi129 & ~n17789;
  assign n17791 = pi128 & n15001;
  assign n17792 = ~pi130 & ~n17791;
  assign n17793 = ~pi129 & n17792;
  assign n17794 = pi301 & ~n17793;
  assign n17795 = ~n14552 & ~n17794;
  assign n17796 = ~n17790 & ~n17795;
  assign n17797 = n17344 & n17796;
  assign n17798 = ~n17783 & ~n17797;
  assign n17799 = ~n17782 & n17798;
  assign n17800 = ~n17782 & ~n17797;
  assign n17801 = n17783 & ~n17800;
  assign n17802 = ~n17799 & ~n17801;
  assign n17803 = ~n17773 & ~n17802;
  assign n17804 = ~n17406 & ~n17770;
  assign n17805 = n17406 & n17770;
  assign n17806 = ~n17804 & ~n17805;
  assign n17807 = n17783 & ~n17797;
  assign n17808 = ~n17782 & n17807;
  assign n17809 = ~n17783 & ~n17800;
  assign n17810 = ~n17808 & ~n17809;
  assign n17811 = ~n17806 & ~n17810;
  assign n17812 = ~n17803 & ~n17811;
  assign n17813 = ~n17782 & n17796;
  assign n17814 = n17344 & ~n17813;
  assign n17815 = ~n17344 & n17813;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = ~n17351 & ~n17816;
  assign n17818 = ~n17352 & ~n17817;
  assign n17819 = ~n17812 & ~n17818;
  assign n17820 = n17812 & n17818;
  assign n17821 = ~n17819 & ~n17820;
  assign n17822 = ~n17353 & ~n17365;
  assign n17823 = ~n17347 & ~n17359;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = pi299 & ~n17824;
  assign n17826 = pi128 & n17825;
  assign n17827 = pi129 & n17826;
  assign n17828 = pi299 & ~n1568;
  assign n17829 = ~n17826 & n17828;
  assign n17830 = ~n17827 & ~n17829;
  assign n17831 = ~n17821 & ~n17830;
  assign n17832 = n17812 & ~n17818;
  assign n17833 = ~n17812 & n17818;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = ~pi129 & n17826;
  assign n17836 = ~n17826 & ~n17828;
  assign n17837 = ~n17835 & ~n17836;
  assign n17838 = ~n17834 & ~n17837;
  assign n17839 = ~n17831 & ~n17838;
  assign n17840 = ~n16844 & ~n16856;
  assign n17841 = ~n16837 & ~n16850;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = n1156 & ~n17842;
  assign n17844 = pi344 & n17843;
  assign n17845 = n1154 & n17844;
  assign n17846 = ~n1154 & ~n17844;
  assign n17847 = pi344 & n17846;
  assign n17848 = ~n17845 & ~n17847;
  assign n17849 = n16014 & n16766;
  assign n17850 = ~n16762 & ~n16792;
  assign n17851 = n16762 & n16792;
  assign n17852 = ~n17850 & ~n17851;
  assign n17853 = n2887 & ~n17852;
  assign n17854 = pi337 & n17853;
  assign n17855 = ~n16762 & n16792;
  assign n17856 = n16762 & ~n16792;
  assign n17857 = ~n17855 & ~n17856;
  assign n17858 = ~n16751 & ~n17857;
  assign n17859 = ~n17854 & ~n17858;
  assign n17860 = ~n16750 & ~n17859;
  assign n17861 = n2887 & ~n17857;
  assign n17862 = pi337 & n17861;
  assign n17863 = ~n16751 & ~n17852;
  assign n17864 = ~n17862 & ~n17863;
  assign n17865 = ~n16808 & ~n17864;
  assign n17866 = ~n17860 & ~n17865;
  assign n17867 = ~n16014 & ~n16766;
  assign n17868 = n17866 & ~n17867;
  assign n17869 = ~n17849 & ~n17868;
  assign n17870 = n1442 & ~n16021;
  assign n17871 = pi341 & n17870;
  assign n17872 = ~n16014 & n16813;
  assign n17873 = n16014 & ~n16813;
  assign n17874 = ~n17872 & ~n17873;
  assign n17875 = ~n16031 & ~n17874;
  assign n17876 = n16014 & n16813;
  assign n17877 = ~n16014 & ~n16813;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = n16031 & ~n17878;
  assign n17880 = ~n17875 & ~n17879;
  assign n17881 = n16021 & ~n16819;
  assign n17882 = ~n17880 & ~n17881;
  assign n17883 = ~n17871 & ~n17882;
  assign n17884 = ~n17869 & n17883;
  assign n17885 = n17869 & ~n17883;
  assign n17886 = ~n17884 & ~n17885;
  assign n17887 = pi339 & n2464;
  assign n17888 = n16051 & n16675;
  assign n17889 = ~n16671 & ~n16701;
  assign n17890 = n16671 & n16701;
  assign n17891 = ~n17889 & ~n17890;
  assign n17892 = n6556 & ~n17891;
  assign n17893 = pi331 & n17892;
  assign n17894 = ~n16671 & n16701;
  assign n17895 = n16671 & ~n16701;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = ~n16642 & ~n17896;
  assign n17898 = ~n17893 & ~n17897;
  assign n17899 = ~n16641 & ~n17898;
  assign n17900 = n6556 & ~n17896;
  assign n17901 = pi331 & n17900;
  assign n17902 = ~n16642 & ~n17891;
  assign n17903 = ~n17901 & ~n17902;
  assign n17904 = ~n16717 & ~n17903;
  assign n17905 = ~n17899 & ~n17904;
  assign n17906 = ~n16051 & ~n16675;
  assign n17907 = n17905 & ~n17906;
  assign n17908 = ~n17888 & ~n17907;
  assign n17909 = n5257 & ~n16058;
  assign n17910 = pi335 & n17909;
  assign n17911 = n16051 & ~n16722;
  assign n17912 = ~n16051 & n16722;
  assign n17913 = ~n17911 & ~n17912;
  assign n17914 = ~n16074 & ~n17913;
  assign n17915 = n16051 & n16722;
  assign n17916 = ~n16051 & ~n16722;
  assign n17917 = ~n17915 & ~n17916;
  assign n17918 = n16074 & ~n17917;
  assign n17919 = ~n17914 & ~n17918;
  assign n17920 = n16058 & ~n16728;
  assign n17921 = ~n17919 & ~n17920;
  assign n17922 = ~n17910 & ~n17921;
  assign n17923 = ~n17908 & n17922;
  assign n17924 = n17908 & ~n17922;
  assign n17925 = ~n17923 & ~n17924;
  assign n17926 = pi333 & n5973;
  assign n17927 = ~n16078 & ~n16613;
  assign n17928 = n16078 & n16613;
  assign n17929 = n11366 & ~n17928;
  assign n17930 = pi328 & n17929;
  assign n17931 = ~n17927 & ~n17930;
  assign n17932 = n16091 & ~n16095;
  assign n17933 = ~n16091 & n16095;
  assign n17934 = ~n16078 & n16613;
  assign n17935 = n16078 & ~n16613;
  assign n17936 = ~n17934 & ~n17935;
  assign n17937 = n11366 & ~n17936;
  assign n17938 = pi328 & n17937;
  assign n17939 = ~n17927 & ~n17928;
  assign n17940 = ~n16619 & ~n17939;
  assign n17941 = ~n17938 & ~n17940;
  assign n17942 = ~n17933 & ~n17941;
  assign n17943 = ~n17932 & ~n17942;
  assign n17944 = n17931 & n17943;
  assign n17945 = ~n17931 & ~n17943;
  assign n17946 = ~n17944 & ~n17945;
  assign n17947 = pi329 & n11366;
  assign n17948 = ~n16099 & n16592;
  assign n17949 = n16099 & ~n16592;
  assign n17950 = ~n16599 & ~n17949;
  assign n17951 = ~n17948 & ~n17950;
  assign n17952 = ~n16099 & ~n16587;
  assign n17953 = n16099 & n16587;
  assign n17954 = ~n17952 & ~n17953;
  assign n17955 = n16119 & n16591;
  assign n17956 = ~n16574 & n16592;
  assign n17957 = n16574 & ~n16592;
  assign n17958 = ~n17956 & ~n17957;
  assign n17959 = ~n17955 & ~n17958;
  assign n17960 = ~n17954 & n17959;
  assign n17961 = ~n16099 & n16587;
  assign n17962 = n16099 & ~n16587;
  assign n17963 = ~n17961 & ~n17962;
  assign n17964 = n16574 & n16592;
  assign n17965 = ~n16574 & ~n16592;
  assign n17966 = ~n17964 & ~n17965;
  assign n17967 = ~n17955 & ~n17966;
  assign n17968 = ~n17963 & n17967;
  assign n17969 = ~n16119 & ~n16591;
  assign n17970 = ~n17968 & ~n17969;
  assign n17971 = ~n17960 & n17970;
  assign n17972 = n17951 & n17971;
  assign n17973 = ~n17951 & ~n17971;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~n16124 & ~n16543;
  assign n17976 = ~n16551 & ~n17975;
  assign n17977 = ~n16132 & n16554;
  assign n17978 = ~n16124 & ~n16552;
  assign n17979 = n16124 & ~n16551;
  assign n17980 = ~n16543 & n17979;
  assign n17981 = ~n17978 & ~n17980;
  assign n17982 = n16132 & ~n16554;
  assign n17983 = ~n17981 & ~n17982;
  assign n17984 = ~n17977 & ~n17983;
  assign n17985 = ~n17976 & n17984;
  assign n17986 = n17976 & ~n17984;
  assign n17987 = ~n17985 & ~n17986;
  assign n17988 = ~n15166 & ~n15621;
  assign n17989 = ~n15622 & ~n17988;
  assign n17990 = n16527 & n17989;
  assign n17991 = ~n16527 & ~n17989;
  assign n17992 = ~n17990 & ~n17991;
  assign n17993 = ~n15616 & ~n17992;
  assign n17994 = ~n16527 & n17989;
  assign n17995 = n16527 & ~n17989;
  assign n17996 = ~n17994 & ~n17995;
  assign n17997 = n15616 & ~n17996;
  assign n17998 = ~n17993 & ~n17997;
  assign n17999 = pi323 & ~n17998;
  assign n18000 = pi151 & pi258;
  assign n18001 = ~n16527 & n18000;
  assign n18002 = n16527 & ~n18000;
  assign n18003 = ~n18001 & ~n18002;
  assign n18004 = n16485 & n16490;
  assign n18005 = ~n16485 & ~n16490;
  assign n18006 = n16479 & ~n18005;
  assign n18007 = ~n18004 & ~n18006;
  assign n18008 = n16489 & n16505;
  assign n18009 = n16490 & ~n16522;
  assign n18010 = ~n16488 & ~n16490;
  assign n18011 = ~n18009 & ~n18010;
  assign n18012 = ~n16489 & ~n16505;
  assign n18013 = ~n18011 & ~n18012;
  assign n18014 = ~n18008 & ~n18013;
  assign n18015 = ~n18007 & ~n18014;
  assign n18016 = n18007 & n18014;
  assign n18017 = ~n18015 & ~n18016;
  assign n18018 = pi149 & pi260;
  assign n18019 = pi133 & pi276;
  assign n18020 = ~n16197 & ~n16204;
  assign n18021 = ~n15254 & n18020;
  assign n18022 = ~n16205 & ~n18021;
  assign n18023 = pi130 & pi279;
  assign n18024 = pi128 & pi281;
  assign n18025 = pi280 & ~n18024;
  assign n18026 = pi129 & n18025;
  assign n18027 = pi129 & pi280;
  assign n18028 = pi281 & ~n18027;
  assign n18029 = pi128 & n18028;
  assign n18030 = ~n18026 & ~n18029;
  assign n18031 = ~n16154 & ~n16157;
  assign n18032 = n16154 & n16157;
  assign n18033 = ~n16153 & ~n18032;
  assign n18034 = ~n18031 & ~n18033;
  assign n18035 = ~n18030 & ~n18034;
  assign n18036 = ~n16152 & ~n18031;
  assign n18037 = ~n15181 & n18036;
  assign n18038 = ~n18032 & ~n18037;
  assign n18039 = n18030 & ~n18038;
  assign n18040 = ~n18035 & ~n18039;
  assign n18041 = n18023 & ~n18040;
  assign n18042 = n18030 & ~n18034;
  assign n18043 = ~n18030 & ~n18038;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = ~n18023 & ~n18044;
  assign n18046 = ~n16153 & ~n16160;
  assign n18047 = ~n16152 & n16160;
  assign n18048 = ~n15181 & n18047;
  assign n18049 = ~n16161 & ~n18048;
  assign n18050 = ~n18046 & n18049;
  assign n18051 = ~n18046 & ~n18048;
  assign n18052 = pi278 & ~n18051;
  assign n18053 = pi130 & n18052;
  assign n18054 = ~n16177 & ~n18053;
  assign n18055 = ~n18050 & ~n18054;
  assign n18056 = ~n18045 & ~n18055;
  assign n18057 = ~n18041 & n18056;
  assign n18058 = ~n18041 & ~n18045;
  assign n18059 = n18055 & ~n18058;
  assign n18060 = ~n18057 & ~n18059;
  assign n18061 = pi278 & ~n18060;
  assign n18062 = pi131 & n18061;
  assign n18063 = pi131 & pi278;
  assign n18064 = ~n18057 & ~n18063;
  assign n18065 = ~n18059 & n18064;
  assign n18066 = ~n16181 & ~n16190;
  assign n18067 = ~n18065 & n18066;
  assign n18068 = ~n18062 & n18067;
  assign n18069 = ~n18062 & ~n18065;
  assign n18070 = ~n18066 & ~n18069;
  assign n18071 = ~n18068 & ~n18070;
  assign n18072 = pi277 & ~n18071;
  assign n18073 = pi132 & n18072;
  assign n18074 = pi132 & pi277;
  assign n18075 = ~n18068 & ~n18074;
  assign n18076 = ~n18070 & n18075;
  assign n18077 = ~n18073 & ~n18076;
  assign n18078 = ~n18022 & ~n18077;
  assign n18079 = n18022 & ~n18076;
  assign n18080 = ~n18073 & n18079;
  assign n18081 = ~n18078 & ~n18080;
  assign n18082 = ~n18019 & ~n18081;
  assign n18083 = n18022 & ~n18077;
  assign n18084 = ~n18022 & ~n18076;
  assign n18085 = ~n18073 & n18084;
  assign n18086 = ~n18083 & ~n18085;
  assign n18087 = pi276 & ~n18086;
  assign n18088 = pi133 & n18087;
  assign n18089 = ~n18082 & ~n18088;
  assign n18090 = n16192 & ~n16197;
  assign n18091 = ~n15254 & n18090;
  assign n18092 = ~n16192 & ~n16200;
  assign n18093 = ~n18091 & ~n18092;
  assign n18094 = ~n16145 & ~n18093;
  assign n18095 = ~n16192 & ~n16197;
  assign n18096 = ~n15254 & n18095;
  assign n18097 = n16192 & ~n16200;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = pi276 & ~n18098;
  assign n18100 = pi132 & n18099;
  assign n18101 = ~n18094 & ~n18100;
  assign n18102 = ~n15313 & n18101;
  assign n18103 = n16143 & n18102;
  assign n18104 = ~pi275 & ~n18101;
  assign n18105 = ~n16238 & ~n18104;
  assign n18106 = pi274 & n18105;
  assign n18107 = ~n16144 & ~n18101;
  assign n18108 = pi275 & ~n18107;
  assign n18109 = ~n18106 & ~n18108;
  assign n18110 = pi133 & ~n18109;
  assign n18111 = ~n18103 & ~n18110;
  assign n18112 = n18089 & n18111;
  assign n18113 = ~n18089 & ~n18111;
  assign n18114 = ~n18112 & ~n18113;
  assign n18115 = pi134 & pi275;
  assign n18116 = ~n15267 & ~n16144;
  assign n18117 = ~n16238 & ~n18116;
  assign n18118 = ~n16212 & ~n18117;
  assign n18119 = ~n16242 & ~n18118;
  assign n18120 = ~n16251 & ~n18119;
  assign n18121 = pi134 & pi274;
  assign n18122 = n16251 & n18119;
  assign n18123 = n18121 & ~n18122;
  assign n18124 = ~n18120 & ~n18123;
  assign n18125 = n18115 & ~n18124;
  assign n18126 = ~n18120 & ~n18121;
  assign n18127 = ~n18122 & ~n18126;
  assign n18128 = ~n18115 & ~n18127;
  assign n18129 = ~n18125 & ~n18128;
  assign n18130 = ~n18114 & ~n18129;
  assign n18131 = n18089 & ~n18111;
  assign n18132 = ~n18089 & n18111;
  assign n18133 = ~n18131 & ~n18132;
  assign n18134 = ~n18115 & ~n18124;
  assign n18135 = n18115 & ~n18127;
  assign n18136 = ~n18134 & ~n18135;
  assign n18137 = ~n18133 & ~n18136;
  assign n18138 = ~n18130 & ~n18137;
  assign n18139 = ~n16254 & ~n16255;
  assign n18140 = n16254 & n16255;
  assign n18141 = ~n16260 & ~n18140;
  assign n18142 = ~n18139 & ~n18141;
  assign n18143 = ~n18138 & n18142;
  assign n18144 = n18138 & ~n18142;
  assign n18145 = ~n18143 & ~n18144;
  assign n18146 = pi136 & pi273;
  assign n18147 = pi135 & pi274;
  assign n18148 = n18146 & n18147;
  assign n18149 = ~n18146 & ~n18147;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = ~n18145 & ~n18150;
  assign n18152 = n18138 & n18142;
  assign n18153 = ~n18138 & ~n18142;
  assign n18154 = ~n18152 & ~n18153;
  assign n18155 = pi273 & ~n18147;
  assign n18156 = pi136 & n18155;
  assign n18157 = pi274 & ~n18146;
  assign n18158 = pi135 & n18157;
  assign n18159 = ~n18156 & ~n18158;
  assign n18160 = ~n18154 & ~n18159;
  assign n18161 = ~n18151 & ~n18160;
  assign n18162 = ~n16287 & ~n16291;
  assign n18163 = ~n16292 & ~n18162;
  assign n18164 = n18161 & n18163;
  assign n18165 = ~n18161 & ~n18163;
  assign n18166 = ~n18164 & ~n18165;
  assign n18167 = pi137 & pi272;
  assign n18168 = n16271 & ~n16284;
  assign n18169 = ~n16280 & n18168;
  assign n18170 = ~n16271 & ~n16287;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = ~n16139 & ~n18171;
  assign n18173 = ~n16271 & ~n16284;
  assign n18174 = ~n16280 & n18173;
  assign n18175 = n16271 & ~n16287;
  assign n18176 = ~n18174 & ~n18175;
  assign n18177 = pi272 & ~n18176;
  assign n18178 = pi136 & n18177;
  assign n18179 = ~n18172 & ~n18178;
  assign n18180 = ~n16303 & ~n18179;
  assign n18181 = n16303 & n18179;
  assign n18182 = n16281 & ~n18181;
  assign n18183 = ~n18180 & ~n18182;
  assign n18184 = n18167 & ~n18183;
  assign n18185 = ~n16281 & ~n18180;
  assign n18186 = ~n18181 & ~n18185;
  assign n18187 = ~n18167 & ~n18186;
  assign n18188 = ~n18184 & ~n18187;
  assign n18189 = ~n18166 & ~n18188;
  assign n18190 = n18161 & ~n18163;
  assign n18191 = ~n18161 & n18163;
  assign n18192 = ~n18190 & ~n18191;
  assign n18193 = ~n18167 & ~n18183;
  assign n18194 = n18167 & ~n18186;
  assign n18195 = ~n18193 & ~n18194;
  assign n18196 = ~n18192 & ~n18195;
  assign n18197 = ~n18189 & ~n18196;
  assign n18198 = ~n16307 & ~n16318;
  assign n18199 = n16307 & n16318;
  assign n18200 = ~n16312 & ~n18199;
  assign n18201 = ~n18198 & ~n18200;
  assign n18202 = ~n18197 & n18201;
  assign n18203 = n18197 & ~n18201;
  assign n18204 = ~n18202 & ~n18203;
  assign n18205 = pi139 & pi270;
  assign n18206 = pi138 & pi271;
  assign n18207 = n18205 & n18206;
  assign n18208 = ~n18205 & ~n18206;
  assign n18209 = ~n18207 & ~n18208;
  assign n18210 = ~n18204 & ~n18209;
  assign n18211 = n18197 & n18201;
  assign n18212 = ~n18197 & ~n18201;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = pi270 & ~n18206;
  assign n18215 = pi139 & n18214;
  assign n18216 = pi271 & ~n18205;
  assign n18217 = pi138 & n18216;
  assign n18218 = ~n18215 & ~n18217;
  assign n18219 = ~n18213 & ~n18218;
  assign n18220 = ~n18210 & ~n18219;
  assign n18221 = ~n16336 & ~n16343;
  assign n18222 = ~n16331 & n18221;
  assign n18223 = ~n16344 & ~n18222;
  assign n18224 = n18220 & n18223;
  assign n18225 = ~n18220 & ~n18223;
  assign n18226 = ~n18224 & ~n18225;
  assign n18227 = pi140 & pi269;
  assign n18228 = ~n16323 & ~n16336;
  assign n18229 = ~n16331 & n18228;
  assign n18230 = n16323 & ~n16339;
  assign n18231 = ~n18229 & ~n18230;
  assign n18232 = ~n16138 & ~n18231;
  assign n18233 = n16323 & ~n16336;
  assign n18234 = ~n16331 & n18233;
  assign n18235 = ~n16323 & ~n16339;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = pi269 & ~n18236;
  assign n18238 = pi139 & n18237;
  assign n18239 = ~n18232 & ~n18238;
  assign n18240 = n16355 & n18239;
  assign n18241 = ~n16355 & ~n18239;
  assign n18242 = n16332 & ~n18241;
  assign n18243 = ~n18240 & ~n18242;
  assign n18244 = n18227 & ~n18243;
  assign n18245 = ~n16332 & ~n18240;
  assign n18246 = ~n18241 & ~n18245;
  assign n18247 = ~n18227 & ~n18246;
  assign n18248 = ~n18244 & ~n18247;
  assign n18249 = ~n18226 & ~n18248;
  assign n18250 = n18220 & ~n18223;
  assign n18251 = ~n18220 & n18223;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = ~n18227 & ~n18243;
  assign n18254 = n18227 & ~n18246;
  assign n18255 = ~n18253 & ~n18254;
  assign n18256 = ~n18252 & ~n18255;
  assign n18257 = ~n18249 & ~n18256;
  assign n18258 = ~n16359 & ~n16370;
  assign n18259 = n16359 & n16370;
  assign n18260 = ~n16364 & ~n18259;
  assign n18261 = ~n18258 & ~n18260;
  assign n18262 = ~n18257 & n18261;
  assign n18263 = n18257 & ~n18261;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = pi142 & pi267;
  assign n18266 = pi141 & pi268;
  assign n18267 = n18265 & n18266;
  assign n18268 = ~n18265 & ~n18266;
  assign n18269 = ~n18267 & ~n18268;
  assign n18270 = ~n18264 & ~n18269;
  assign n18271 = n18257 & n18261;
  assign n18272 = ~n18257 & ~n18261;
  assign n18273 = ~n18271 & ~n18272;
  assign n18274 = pi267 & ~n18266;
  assign n18275 = pi142 & n18274;
  assign n18276 = pi268 & ~n18265;
  assign n18277 = pi141 & n18276;
  assign n18278 = ~n18275 & ~n18277;
  assign n18279 = ~n18273 & ~n18278;
  assign n18280 = ~n18270 & ~n18279;
  assign n18281 = ~n16388 & ~n16395;
  assign n18282 = ~n16383 & n18281;
  assign n18283 = ~n16396 & ~n18282;
  assign n18284 = n18280 & ~n18283;
  assign n18285 = ~n18280 & n18283;
  assign n18286 = ~n18284 & ~n18285;
  assign n18287 = pi143 & pi266;
  assign n18288 = ~n16375 & ~n16388;
  assign n18289 = ~n16383 & n18288;
  assign n18290 = n16375 & ~n16391;
  assign n18291 = ~n18289 & ~n18290;
  assign n18292 = ~n16137 & ~n18291;
  assign n18293 = n16375 & ~n16388;
  assign n18294 = ~n16383 & n18293;
  assign n18295 = ~n16375 & ~n16391;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = pi266 & ~n18296;
  assign n18298 = pi142 & n18297;
  assign n18299 = ~n18292 & ~n18298;
  assign n18300 = n16407 & n18299;
  assign n18301 = ~n16407 & ~n18299;
  assign n18302 = n16384 & ~n18301;
  assign n18303 = ~n18300 & ~n18302;
  assign n18304 = n18287 & ~n18303;
  assign n18305 = ~n16384 & ~n18300;
  assign n18306 = ~n18301 & ~n18305;
  assign n18307 = ~n18287 & ~n18306;
  assign n18308 = ~n18304 & ~n18307;
  assign n18309 = ~n18286 & ~n18308;
  assign n18310 = n18280 & n18283;
  assign n18311 = ~n18280 & ~n18283;
  assign n18312 = ~n18310 & ~n18311;
  assign n18313 = ~n18287 & ~n18303;
  assign n18314 = n18287 & ~n18306;
  assign n18315 = ~n18313 & ~n18314;
  assign n18316 = ~n18312 & ~n18315;
  assign n18317 = ~n18309 & ~n18316;
  assign n18318 = n16411 & ~n16422;
  assign n18319 = ~n16411 & n16422;
  assign n18320 = ~n16413 & ~n18319;
  assign n18321 = ~n18318 & ~n18320;
  assign n18322 = ~n18317 & n18321;
  assign n18323 = n18317 & ~n18321;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = pi145 & pi264;
  assign n18326 = pi144 & pi265;
  assign n18327 = n18325 & n18326;
  assign n18328 = ~n18325 & ~n18326;
  assign n18329 = ~n18327 & ~n18328;
  assign n18330 = ~n18324 & ~n18329;
  assign n18331 = n18317 & n18321;
  assign n18332 = ~n18317 & ~n18321;
  assign n18333 = ~n18331 & ~n18332;
  assign n18334 = pi264 & ~n18326;
  assign n18335 = pi145 & n18334;
  assign n18336 = pi265 & ~n18325;
  assign n18337 = pi144 & n18336;
  assign n18338 = ~n18335 & ~n18337;
  assign n18339 = ~n18333 & ~n18338;
  assign n18340 = ~n18330 & ~n18339;
  assign n18341 = ~n16443 & ~n16447;
  assign n18342 = ~n16448 & ~n18341;
  assign n18343 = n18340 & ~n18342;
  assign n18344 = ~n18340 & n18342;
  assign n18345 = ~n18343 & ~n18344;
  assign n18346 = pi146 & pi263;
  assign n18347 = ~n16427 & ~n16440;
  assign n18348 = ~n16436 & n18347;
  assign n18349 = n16427 & ~n16443;
  assign n18350 = ~n18348 & ~n18349;
  assign n18351 = ~n16136 & ~n18350;
  assign n18352 = n16427 & ~n16440;
  assign n18353 = ~n16436 & n18352;
  assign n18354 = ~n16427 & ~n16443;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = pi263 & ~n18355;
  assign n18357 = pi145 & n18356;
  assign n18358 = ~n18351 & ~n18357;
  assign n18359 = n16459 & n18358;
  assign n18360 = ~n16459 & ~n18358;
  assign n18361 = n16437 & ~n18360;
  assign n18362 = ~n18359 & ~n18361;
  assign n18363 = n18346 & ~n18362;
  assign n18364 = ~n16437 & ~n18359;
  assign n18365 = ~n18360 & ~n18364;
  assign n18366 = ~n18346 & ~n18365;
  assign n18367 = ~n18363 & ~n18366;
  assign n18368 = ~n18345 & ~n18367;
  assign n18369 = n18340 & n18342;
  assign n18370 = ~n18340 & ~n18342;
  assign n18371 = ~n18369 & ~n18370;
  assign n18372 = ~n18346 & ~n18362;
  assign n18373 = n18346 & ~n18365;
  assign n18374 = ~n18372 & ~n18373;
  assign n18375 = ~n18371 & ~n18374;
  assign n18376 = ~n18368 & ~n18375;
  assign n18377 = n16463 & ~n16474;
  assign n18378 = ~n16463 & n16474;
  assign n18379 = ~n16465 & ~n18378;
  assign n18380 = ~n18377 & ~n18379;
  assign n18381 = ~n18376 & n18380;
  assign n18382 = n18376 & ~n18380;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = pi148 & pi261;
  assign n18385 = pi147 & pi262;
  assign n18386 = n18384 & n18385;
  assign n18387 = ~n18384 & ~n18385;
  assign n18388 = ~n18386 & ~n18387;
  assign n18389 = ~n18383 & ~n18388;
  assign n18390 = n18376 & n18380;
  assign n18391 = ~n18376 & ~n18380;
  assign n18392 = ~n18390 & ~n18391;
  assign n18393 = pi261 & ~n18385;
  assign n18394 = pi148 & n18393;
  assign n18395 = pi262 & ~n18384;
  assign n18396 = pi147 & n18395;
  assign n18397 = ~n18394 & ~n18396;
  assign n18398 = ~n18392 & ~n18397;
  assign n18399 = ~n18389 & ~n18398;
  assign n18400 = ~n18018 & n18399;
  assign n18401 = n18018 & ~n18399;
  assign n18402 = ~n18400 & ~n18401;
  assign n18403 = ~n16493 & n16505;
  assign n18404 = ~n16505 & ~n16513;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = ~n16522 & ~n18405;
  assign n18407 = n16505 & ~n16513;
  assign n18408 = ~n16493 & ~n16505;
  assign n18409 = ~n18407 & ~n18408;
  assign n18410 = ~n16488 & ~n18409;
  assign n18411 = ~n18406 & ~n18410;
  assign n18412 = n16506 & ~n18411;
  assign n18413 = pi150 & pi259;
  assign n18414 = n18412 & n18413;
  assign n18415 = ~n18412 & ~n18413;
  assign n18416 = ~n18414 & ~n18415;
  assign n18417 = ~n18402 & ~n18416;
  assign n18418 = n18018 & n18399;
  assign n18419 = ~n18018 & ~n18399;
  assign n18420 = ~n18418 & ~n18419;
  assign n18421 = ~n18412 & n18413;
  assign n18422 = n18412 & ~n18413;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = ~n18420 & ~n18423;
  assign n18425 = ~n18417 & ~n18424;
  assign n18426 = ~n18017 & ~n18425;
  assign n18427 = ~n18007 & n18014;
  assign n18428 = n18007 & ~n18014;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = ~n18416 & ~n18420;
  assign n18431 = ~n18402 & ~n18423;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = ~n18429 & ~n18432;
  assign n18434 = ~n18426 & ~n18433;
  assign n18435 = ~n15616 & ~n17990;
  assign n18436 = ~n17991 & ~n18435;
  assign n18437 = n18434 & ~n18436;
  assign n18438 = ~n18434 & n18436;
  assign n18439 = ~n18437 & ~n18438;
  assign n18440 = ~n18003 & ~n18439;
  assign n18441 = n18434 & n18436;
  assign n18442 = ~n18434 & ~n18436;
  assign n18443 = ~n18441 & ~n18442;
  assign n18444 = n16527 & n18000;
  assign n18445 = ~n16527 & ~n18000;
  assign n18446 = ~n18444 & ~n18445;
  assign n18447 = ~n18443 & ~n18446;
  assign n18448 = pi322 & ~n18447;
  assign n18449 = ~n18440 & n18448;
  assign n18450 = ~n17999 & ~n18449;
  assign n18451 = pi322 & ~n17998;
  assign n18452 = ~n18003 & ~n18443;
  assign n18453 = ~n18439 & ~n18446;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = n18451 & ~n18454;
  assign n18456 = pi323 & n18455;
  assign n18457 = ~n18450 & ~n18456;
  assign n18458 = pi325 & n13762;
  assign n18459 = ~n15166 & ~n15627;
  assign n18460 = n15166 & ~n15623;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = pi324 & n18461;
  assign n18463 = n18458 & n18462;
  assign n18464 = ~n18458 & ~n18462;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = ~n18457 & ~n18465;
  assign n18467 = ~n18458 & n18462;
  assign n18468 = n18458 & ~n18462;
  assign n18469 = ~n18467 & ~n18468;
  assign n18470 = ~n18456 & ~n18469;
  assign n18471 = ~n18450 & n18470;
  assign n18472 = ~n18466 & ~n18471;
  assign n18473 = ~n17987 & ~n18472;
  assign n18474 = ~n17976 & ~n17984;
  assign n18475 = n17976 & n17984;
  assign n18476 = ~n18474 & ~n18475;
  assign n18477 = ~n18457 & ~n18469;
  assign n18478 = ~n18456 & ~n18465;
  assign n18479 = ~n18450 & n18478;
  assign n18480 = ~n18477 & ~n18479;
  assign n18481 = ~n18476 & ~n18480;
  assign n18482 = ~n18473 & ~n18481;
  assign n18483 = n16553 & ~n16587;
  assign n18484 = ~n16554 & ~n17981;
  assign n18485 = n16124 & ~n16552;
  assign n18486 = ~n16124 & ~n16551;
  assign n18487 = ~n16543 & n18486;
  assign n18488 = ~n18485 & ~n18487;
  assign n18489 = n13762 & ~n18488;
  assign n18490 = pi324 & n18489;
  assign n18491 = ~n18484 & ~n18490;
  assign n18492 = n16132 & ~n18491;
  assign n18493 = ~n16132 & n18491;
  assign n18494 = ~n18492 & ~n18493;
  assign n18495 = ~n16553 & n16587;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = ~n18483 & ~n18496;
  assign n18498 = n18482 & n18497;
  assign n18499 = ~n18482 & ~n18497;
  assign n18500 = ~n18498 & ~n18499;
  assign n18501 = pi327 & n11711;
  assign n18502 = pi326 & n12917;
  assign n18503 = n18501 & n18502;
  assign n18504 = ~n18501 & ~n18502;
  assign n18505 = ~n18503 & ~n18504;
  assign n18506 = ~n18500 & ~n18505;
  assign n18507 = ~n18482 & n18497;
  assign n18508 = n18482 & ~n18497;
  assign n18509 = ~n18507 & ~n18508;
  assign n18510 = ~n18501 & n18502;
  assign n18511 = n18501 & ~n18502;
  assign n18512 = ~n18510 & ~n18511;
  assign n18513 = ~n18509 & ~n18512;
  assign n18514 = ~n18506 & ~n18513;
  assign n18515 = ~n17974 & ~n18514;
  assign n18516 = n17951 & ~n17971;
  assign n18517 = ~n17951 & n17971;
  assign n18518 = ~n18516 & ~n18517;
  assign n18519 = ~n18505 & ~n18509;
  assign n18520 = ~n18500 & ~n18512;
  assign n18521 = ~n18519 & ~n18520;
  assign n18522 = ~n18518 & ~n18521;
  assign n18523 = ~n18515 & ~n18522;
  assign n18524 = ~n17947 & n18523;
  assign n18525 = n17947 & ~n18523;
  assign n18526 = ~n18524 & ~n18525;
  assign n18527 = n11384 & ~n18526;
  assign n18528 = pi328 & n18527;
  assign n18529 = pi328 & n11384;
  assign n18530 = n17947 & n18523;
  assign n18531 = ~n17947 & ~n18523;
  assign n18532 = ~n18530 & ~n18531;
  assign n18533 = ~n18529 & ~n18532;
  assign n18534 = ~n18528 & ~n18533;
  assign n18535 = ~n17946 & ~n18534;
  assign n18536 = n17931 & ~n17943;
  assign n18537 = ~n17931 & n17943;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = n11384 & ~n18532;
  assign n18540 = pi328 & n18539;
  assign n18541 = ~n18526 & ~n18529;
  assign n18542 = ~n18540 & ~n18541;
  assign n18543 = ~n18538 & ~n18542;
  assign n18544 = ~n18535 & ~n18543;
  assign n18545 = ~n16638 & n16642;
  assign n18546 = n16638 & ~n16642;
  assign n18547 = n6556 & ~n16659;
  assign n18548 = ~n16660 & ~n18547;
  assign n18549 = n9205 & ~n18548;
  assign n18550 = pi330 & n18549;
  assign n18551 = ~n9205 & ~n18547;
  assign n18552 = pi330 & ~n18551;
  assign n18553 = ~n16660 & ~n18552;
  assign n18554 = ~n18550 & ~n18553;
  assign n18555 = n16634 & ~n18554;
  assign n18556 = ~n16634 & n18554;
  assign n18557 = ~n18555 & ~n18556;
  assign n18558 = ~n18546 & ~n18557;
  assign n18559 = ~n18545 & ~n18558;
  assign n18560 = n18544 & n18559;
  assign n18561 = ~n18544 & ~n18559;
  assign n18562 = ~n18560 & ~n18561;
  assign n18563 = pi331 & n9205;
  assign n18564 = n16634 & ~n18553;
  assign n18565 = ~n18550 & ~n18564;
  assign n18566 = n10561 & n18565;
  assign n18567 = pi330 & n18566;
  assign n18568 = pi330 & n10561;
  assign n18569 = ~n18565 & ~n18568;
  assign n18570 = ~n18567 & ~n18569;
  assign n18571 = ~n18563 & n18570;
  assign n18572 = n18563 & ~n18570;
  assign n18573 = ~n18571 & ~n18572;
  assign n18574 = pi332 & n6556;
  assign n18575 = n5973 & ~n16043;
  assign n18576 = pi331 & n18575;
  assign n18577 = ~n15085 & ~n16034;
  assign n18578 = ~n16679 & ~n18577;
  assign n18579 = ~n18576 & n18578;
  assign n18580 = ~n16685 & ~n18579;
  assign n18581 = n16680 & ~n18580;
  assign n18582 = ~n16674 & ~n18581;
  assign n18583 = ~n16717 & n18582;
  assign n18584 = ~n16680 & n18580;
  assign n18585 = ~n16708 & ~n18581;
  assign n18586 = ~n16641 & n18585;
  assign n18587 = ~n18584 & ~n18586;
  assign n18588 = ~n18583 & n18587;
  assign n18589 = n18574 & ~n18588;
  assign n18590 = ~n18574 & n18588;
  assign n18591 = ~n18589 & ~n18590;
  assign n18592 = ~n18573 & ~n18591;
  assign n18593 = n18563 & n18570;
  assign n18594 = ~n18563 & ~n18570;
  assign n18595 = ~n18593 & ~n18594;
  assign n18596 = ~n18574 & ~n18588;
  assign n18597 = n18574 & n18588;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = ~n18595 & ~n18598;
  assign n18600 = ~n18592 & ~n18599;
  assign n18601 = ~n18562 & ~n18600;
  assign n18602 = n18544 & ~n18559;
  assign n18603 = ~n18544 & n18559;
  assign n18604 = ~n18602 & ~n18603;
  assign n18605 = ~n18591 & ~n18595;
  assign n18606 = ~n18573 & ~n18598;
  assign n18607 = ~n18605 & ~n18606;
  assign n18608 = ~n18604 & ~n18607;
  assign n18609 = ~n18601 & ~n18608;
  assign n18610 = ~n17926 & n18609;
  assign n18611 = n17926 & ~n18609;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = pi335 & n5714;
  assign n18614 = pi334 & n5732;
  assign n18615 = n5257 & ~n16062;
  assign n18616 = ~n16063 & ~n18615;
  assign n18617 = n5714 & ~n18616;
  assign n18618 = pi334 & n18617;
  assign n18619 = ~n5714 & ~n18615;
  assign n18620 = pi334 & ~n18619;
  assign n18621 = ~n16063 & ~n18620;
  assign n18622 = ~n17917 & ~n18621;
  assign n18623 = ~n18618 & ~n18622;
  assign n18624 = ~n18614 & ~n18623;
  assign n18625 = n17913 & ~n18621;
  assign n18626 = n5732 & ~n18625;
  assign n18627 = pi334 & n18626;
  assign n18628 = ~n18618 & n18627;
  assign n18629 = ~n18624 & ~n18628;
  assign n18630 = n18613 & ~n18629;
  assign n18631 = ~n18613 & n18629;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = ~n18612 & ~n18632;
  assign n18634 = n17926 & n18609;
  assign n18635 = ~n17926 & ~n18609;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = ~n18613 & ~n18629;
  assign n18638 = n18613 & n18629;
  assign n18639 = ~n18637 & ~n18638;
  assign n18640 = ~n18636 & ~n18639;
  assign n18641 = ~n18633 & ~n18640;
  assign n18642 = ~n17925 & ~n18641;
  assign n18643 = ~n17908 & ~n17922;
  assign n18644 = n17908 & n17922;
  assign n18645 = ~n18643 & ~n18644;
  assign n18646 = ~n18632 & ~n18636;
  assign n18647 = ~n18612 & ~n18639;
  assign n18648 = ~n18646 & ~n18647;
  assign n18649 = ~n18645 & ~n18648;
  assign n18650 = ~n18642 & ~n18649;
  assign n18651 = ~n16747 & n16751;
  assign n18652 = ~n16743 & ~n16762;
  assign n18653 = n16743 & n16762;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = n16747 & ~n16751;
  assign n18656 = ~n18654 & ~n18655;
  assign n18657 = ~n18651 & ~n18656;
  assign n18658 = n18650 & n18657;
  assign n18659 = ~n18650 & ~n18657;
  assign n18660 = ~n18658 & ~n18659;
  assign n18661 = pi337 & n4596;
  assign n18662 = ~n16743 & ~n16757;
  assign n18663 = n16743 & n16757;
  assign n18664 = ~n4596 & ~n18663;
  assign n18665 = ~n18662 & ~n18664;
  assign n18666 = n5257 & ~n18665;
  assign n18667 = ~n5257 & ~n18662;
  assign n18668 = n4596 & n18667;
  assign n18669 = ~n18666 & ~n18668;
  assign n18670 = pi336 & ~n18669;
  assign n18671 = pi336 & n5257;
  assign n18672 = n16743 & ~n18671;
  assign n18673 = n16757 & n18672;
  assign n18674 = ~n18670 & ~n18673;
  assign n18675 = ~n18661 & n18674;
  assign n18676 = n18661 & ~n18674;
  assign n18677 = ~n18675 & ~n18676;
  assign n18678 = pi338 & n2887;
  assign n18679 = n2464 & ~n16006;
  assign n18680 = pi337 & n18679;
  assign n18681 = ~n15054 & ~n15997;
  assign n18682 = ~n16770 & ~n18681;
  assign n18683 = ~n18680 & n18682;
  assign n18684 = ~n16776 & ~n18683;
  assign n18685 = n16771 & ~n18684;
  assign n18686 = ~n16765 & ~n18685;
  assign n18687 = ~n16808 & n18686;
  assign n18688 = ~n16771 & n18684;
  assign n18689 = ~n16799 & ~n18685;
  assign n18690 = ~n16750 & n18689;
  assign n18691 = ~n18688 & ~n18690;
  assign n18692 = ~n18687 & n18691;
  assign n18693 = n18678 & ~n18692;
  assign n18694 = ~n18678 & n18692;
  assign n18695 = ~n18693 & ~n18694;
  assign n18696 = ~n18677 & ~n18695;
  assign n18697 = n18661 & n18674;
  assign n18698 = ~n18661 & ~n18674;
  assign n18699 = ~n18697 & ~n18698;
  assign n18700 = ~n18678 & ~n18692;
  assign n18701 = n18678 & n18692;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = ~n18699 & ~n18702;
  assign n18704 = ~n18696 & ~n18703;
  assign n18705 = ~n18660 & ~n18704;
  assign n18706 = n18650 & ~n18657;
  assign n18707 = ~n18650 & n18657;
  assign n18708 = ~n18706 & ~n18707;
  assign n18709 = ~n18695 & ~n18699;
  assign n18710 = ~n18677 & ~n18702;
  assign n18711 = ~n18709 & ~n18710;
  assign n18712 = ~n18708 & ~n18711;
  assign n18713 = ~n18705 & ~n18712;
  assign n18714 = ~n17887 & n18713;
  assign n18715 = n17887 & ~n18713;
  assign n18716 = ~n18714 & ~n18715;
  assign n18717 = pi341 & n1729;
  assign n18718 = pi340 & n2091;
  assign n18719 = n1729 & ~n16026;
  assign n18720 = pi340 & n18719;
  assign n18721 = ~n16025 & ~n16029;
  assign n18722 = ~n15889 & n18721;
  assign n18723 = ~n17878 & ~n18722;
  assign n18724 = ~n18720 & ~n18723;
  assign n18725 = ~n18718 & ~n18724;
  assign n18726 = n17874 & ~n18722;
  assign n18727 = ~n18720 & ~n18726;
  assign n18728 = n2091 & n18727;
  assign n18729 = pi340 & n18728;
  assign n18730 = ~n18725 & ~n18729;
  assign n18731 = n18717 & ~n18730;
  assign n18732 = ~n18717 & n18730;
  assign n18733 = ~n18731 & ~n18732;
  assign n18734 = ~n18716 & ~n18733;
  assign n18735 = n17887 & n18713;
  assign n18736 = ~n17887 & ~n18713;
  assign n18737 = ~n18735 & ~n18736;
  assign n18738 = ~n18717 & ~n18730;
  assign n18739 = n18717 & n18730;
  assign n18740 = ~n18738 & ~n18739;
  assign n18741 = ~n18737 & ~n18740;
  assign n18742 = ~n18734 & ~n18741;
  assign n18743 = ~n17886 & ~n18742;
  assign n18744 = ~n17869 & ~n17883;
  assign n18745 = n17869 & n17883;
  assign n18746 = ~n18744 & ~n18745;
  assign n18747 = ~n18733 & ~n18737;
  assign n18748 = ~n18716 & ~n18740;
  assign n18749 = ~n18747 & ~n18748;
  assign n18750 = ~n18746 & ~n18749;
  assign n18751 = ~n18743 & ~n18750;
  assign n18752 = ~n16842 & ~n16856;
  assign n18753 = ~n16843 & ~n18752;
  assign n18754 = n18751 & n18753;
  assign n18755 = ~n18751 & ~n18753;
  assign n18756 = ~n18754 & ~n18755;
  assign n18757 = n15989 & n16834;
  assign n18758 = ~n15989 & ~n16834;
  assign n18759 = ~n1256 & ~n18758;
  assign n18760 = ~n18757 & ~n18759;
  assign n18761 = n1442 & ~n18760;
  assign n18762 = pi342 & n18761;
  assign n18763 = ~n1442 & ~n18759;
  assign n18764 = pi342 & ~n18763;
  assign n18765 = ~n18757 & ~n18764;
  assign n18766 = ~n18762 & ~n18765;
  assign n18767 = ~n1256 & ~n18766;
  assign n18768 = pi343 & n18767;
  assign n18769 = pi343 & ~n1256;
  assign n18770 = ~n18765 & ~n18769;
  assign n18771 = ~n18762 & n18770;
  assign n18772 = ~n18768 & ~n18771;
  assign n18773 = ~n18756 & ~n18772;
  assign n18774 = n18751 & ~n18753;
  assign n18775 = ~n18751 & n18753;
  assign n18776 = ~n18774 & ~n18775;
  assign n18777 = ~n18766 & ~n18769;
  assign n18778 = n18766 & n18769;
  assign n18779 = ~n18777 & ~n18778;
  assign n18780 = ~n18776 & ~n18779;
  assign n18781 = ~n18773 & ~n18780;
  assign n18782 = n17848 & ~n18781;
  assign n18783 = ~n17848 & n18781;
  assign n18784 = ~n18782 & ~n18783;
  assign n18785 = ~n16862 & ~n17379;
  assign n18786 = n16862 & n17379;
  assign n18787 = ~pi280 & ~n18786;
  assign n18788 = ~n18785 & ~n18787;
  assign n18789 = ~pi281 & n18788;
  assign n18790 = pi281 & ~n18788;
  assign n18791 = ~n18789 & ~n18790;
  assign n18792 = n1156 & ~n18791;
  assign n18793 = pi345 & n18792;
  assign n18794 = pi345 & n1156;
  assign n18795 = ~pi281 & ~n18788;
  assign n18796 = pi281 & n18788;
  assign n18797 = ~n18795 & ~n18796;
  assign n18798 = ~n18794 & ~n18797;
  assign n18799 = ~n18793 & ~n18798;
  assign n18800 = ~n18784 & ~n18799;
  assign n18801 = n17848 & n18781;
  assign n18802 = ~n17848 & ~n18781;
  assign n18803 = ~n18801 & ~n18802;
  assign n18804 = n1156 & ~n18797;
  assign n18805 = pi345 & n18804;
  assign n18806 = ~n18791 & ~n18794;
  assign n18807 = ~n18805 & ~n18806;
  assign n18808 = ~n18803 & ~n18807;
  assign n18809 = ~n18800 & ~n18808;
  assign n18810 = ~n17839 & n18809;
  assign n18811 = n17839 & ~n18809;
  assign n18812 = ~n18810 & ~n18811;
  assign n18813 = pi298 & ~n18812;
  assign n18814 = pi128 & n18813;
  assign n18815 = pi128 & pi298;
  assign n18816 = n17839 & n18809;
  assign n18817 = ~n17839 & ~n18809;
  assign n18818 = ~n18816 & ~n18817;
  assign n18819 = ~n18815 & ~n18818;
  assign n18820 = ~n18814 & ~n18819;
  assign n18821 = ~n16866 & n17371;
  assign n18822 = n16866 & ~n17371;
  assign n18823 = ~n18785 & ~n18786;
  assign n18824 = pi280 & ~n18823;
  assign n18825 = n16862 & ~n17379;
  assign n18826 = ~n16862 & n17379;
  assign n18827 = ~n18825 & ~n18826;
  assign n18828 = ~pi280 & ~n18827;
  assign n18829 = ~n18824 & ~n18828;
  assign n18830 = ~n18822 & ~n18829;
  assign n18831 = ~n18821 & ~n18830;
  assign n18832 = n18820 & n18831;
  assign n18833 = ~n18820 & ~n18831;
  assign n18834 = ~n18832 & ~n18833;
  assign n18835 = ~n831 & ~n18834;
  assign n18836 = ~n17405 & ~n18835;
  assign n18837 = pi161 & ~n18836;
  assign n18838 = ~n17404 & ~n18837;
  assign po216 = ~pi160 & n18838;
  assign n18840 = ~pi088 & ~pi161;
  assign n18841 = ~pi282 & n831;
  assign n18842 = pi299 & n1515;
  assign n18843 = ~n17821 & ~n17835;
  assign n18844 = ~n17836 & ~n18843;
  assign n18845 = n18842 & ~n18844;
  assign n18846 = ~n17834 & ~n17836;
  assign n18847 = ~n17835 & ~n18846;
  assign n18848 = ~n18842 & ~n18847;
  assign n18849 = ~n18845 & ~n18848;
  assign n18850 = pi301 & n1533;
  assign n18851 = ~n17800 & ~n17804;
  assign n18852 = ~n17805 & ~n18851;
  assign n18853 = ~n18850 & ~n18852;
  assign n18854 = ~n17797 & ~n17805;
  assign n18855 = ~n17782 & n18854;
  assign n18856 = ~n17804 & ~n18855;
  assign n18857 = n18850 & ~n18856;
  assign n18858 = ~n18853 & ~n18857;
  assign n18859 = n17744 & ~n17748;
  assign n18860 = ~n17744 & n17748;
  assign n18861 = ~n18859 & ~n18860;
  assign n18862 = ~n17416 & ~n18861;
  assign n18863 = ~n17325 & ~n17329;
  assign n18864 = ~n17324 & ~n18863;
  assign n18865 = n17416 & n18861;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = ~n18862 & ~n18866;
  assign n18868 = pi305 & n3012;
  assign n18869 = ~n17730 & ~n17737;
  assign n18870 = ~n17738 & ~n18869;
  assign n18871 = ~n18868 & ~n18870;
  assign n18872 = ~n17733 & ~n17738;
  assign n18873 = ~n17737 & ~n18872;
  assign n18874 = n18868 & ~n18873;
  assign n18875 = ~n18871 & ~n18874;
  assign n18876 = ~n17430 & ~n17692;
  assign n18877 = ~n17253 & ~n17258;
  assign n18878 = ~n17254 & ~n18877;
  assign n18879 = n17430 & n17692;
  assign n18880 = ~n18878 & ~n18879;
  assign n18881 = ~n18876 & ~n18880;
  assign n18882 = pi309 & n5463;
  assign n18883 = ~n17671 & ~n17678;
  assign n18884 = ~n17679 & ~n18883;
  assign n18885 = ~n18882 & ~n18884;
  assign n18886 = ~n17674 & ~n17679;
  assign n18887 = ~n17678 & ~n18886;
  assign n18888 = n18882 & ~n18887;
  assign n18889 = ~n18885 & ~n18888;
  assign n18890 = ~n17604 & ~n17605;
  assign n18891 = n17604 & n17605;
  assign n18892 = ~n17610 & ~n18891;
  assign n18893 = ~n18890 & ~n18892;
  assign n18894 = pi313 & n9517;
  assign n18895 = ~n17583 & ~n17590;
  assign n18896 = ~n17591 & ~n18895;
  assign n18897 = ~n18894 & ~n18896;
  assign n18898 = ~n17586 & ~n17591;
  assign n18899 = ~n17590 & ~n18898;
  assign n18900 = n18894 & ~n18899;
  assign n18901 = ~n18897 & ~n18900;
  assign n18902 = ~n17550 & ~n17551;
  assign n18903 = n17550 & n17551;
  assign n18904 = ~n17117 & ~n18903;
  assign n18905 = ~n17111 & n18904;
  assign n18906 = ~n18902 & ~n18905;
  assign n18907 = ~n17506 & n17511;
  assign n18908 = ~n17505 & ~n17511;
  assign n18909 = ~n17502 & n18908;
  assign n18910 = ~n18907 & ~n18909;
  assign n18911 = ~n17532 & ~n18910;
  assign n18912 = pi317 & n14156;
  assign n18913 = ~pi152 & ~n16976;
  assign n18914 = pi151 & n18913;
  assign n18915 = ~pi151 & pi152;
  assign n18916 = pi150 & n18915;
  assign n18917 = ~n18914 & ~n18916;
  assign n18918 = pi149 & ~n18917;
  assign n18919 = pi151 & pi152;
  assign n18920 = ~pi150 & n18919;
  assign n18921 = ~pi152 & n16976;
  assign n18922 = ~pi151 & n18921;
  assign n18923 = ~n18920 & ~n18922;
  assign n18924 = ~pi149 & ~n18923;
  assign n18925 = pi151 & ~pi152;
  assign n18926 = pi152 & ~n16976;
  assign n18927 = ~pi151 & n18926;
  assign n18928 = ~n18925 & ~n18927;
  assign n18929 = pi150 & ~n18928;
  assign n18930 = ~pi151 & ~pi152;
  assign n18931 = pi152 & n16976;
  assign n18932 = pi151 & n18931;
  assign n18933 = ~n18930 & ~n18932;
  assign n18934 = ~pi150 & ~n18933;
  assign n18935 = ~n18929 & ~n18934;
  assign n18936 = ~n18924 & n18935;
  assign n18937 = ~n18918 & n18936;
  assign n18938 = n17455 & ~n17462;
  assign n18939 = ~pi320 & ~n18938;
  assign n18940 = ~n16985 & ~n17455;
  assign n18941 = pi320 & n18938;
  assign n18942 = ~n17465 & ~n18941;
  assign n18943 = ~n18940 & n18942;
  assign n18944 = ~n18939 & n18943;
  assign n18945 = n18937 & ~n18944;
  assign n18946 = ~n17462 & ~n18937;
  assign n18947 = ~pi320 & n17455;
  assign n18948 = n18946 & n18947;
  assign n18949 = ~n18945 & ~n18948;
  assign n18950 = pi321 & ~n18949;
  assign n18951 = n17462 & ~n18937;
  assign n18952 = ~n16985 & n18951;
  assign n18953 = ~pi321 & ~n17470;
  assign n18954 = ~n18952 & ~n18953;
  assign n18955 = n17455 & ~n18954;
  assign n18956 = pi321 & n18937;
  assign n18957 = ~n17462 & ~n18956;
  assign n18958 = ~n17455 & n18957;
  assign n18959 = n16985 & n18958;
  assign n18960 = ~n18955 & ~n18959;
  assign n18961 = pi320 & ~n18960;
  assign n18962 = ~n18950 & ~n18961;
  assign n18963 = pi319 & n16985;
  assign n18964 = n18962 & n18963;
  assign n18965 = ~n18962 & ~n18963;
  assign n18966 = ~n18964 & ~n18965;
  assign n18967 = ~n17008 & ~n17021;
  assign n18968 = ~n17007 & ~n18967;
  assign n18969 = ~n17478 & ~n18968;
  assign n18970 = ~n17477 & ~n18969;
  assign n18971 = n18966 & ~n18970;
  assign n18972 = ~n18966 & n18970;
  assign n18973 = ~n18971 & ~n18972;
  assign n18974 = pi318 & n14618;
  assign n18975 = ~n17484 & n17495;
  assign n18976 = n18974 & ~n18975;
  assign n18977 = ~n17487 & n18976;
  assign n18978 = ~n17487 & ~n18975;
  assign n18979 = ~n18974 & ~n18978;
  assign n18980 = ~n18977 & ~n18979;
  assign n18981 = ~n18973 & ~n18980;
  assign n18982 = n18966 & n18970;
  assign n18983 = ~n18966 & ~n18970;
  assign n18984 = ~n18982 & ~n18983;
  assign n18985 = ~n18974 & ~n18975;
  assign n18986 = ~n17487 & n18985;
  assign n18987 = n18974 & ~n18978;
  assign n18988 = ~n18986 & ~n18987;
  assign n18989 = ~n18984 & ~n18988;
  assign n18990 = ~n18981 & ~n18989;
  assign n18991 = ~n18912 & ~n18990;
  assign n18992 = n18912 & n18990;
  assign n18993 = ~n18991 & ~n18992;
  assign n18994 = pi316 & n11998;
  assign n18995 = ~n17505 & n17511;
  assign n18996 = ~n18994 & ~n18995;
  assign n18997 = ~n17502 & n18996;
  assign n18998 = ~n17502 & ~n18995;
  assign n18999 = n18994 & ~n18998;
  assign n19000 = ~n18997 & ~n18999;
  assign n19001 = ~n18993 & ~n19000;
  assign n19002 = ~n18912 & n18990;
  assign n19003 = n18912 & ~n18990;
  assign n19004 = ~n19002 & ~n19003;
  assign n19005 = n18994 & ~n18995;
  assign n19006 = ~n17502 & n19005;
  assign n19007 = ~n18994 & ~n18998;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = ~n19004 & ~n19008;
  assign n19010 = ~n19001 & ~n19009;
  assign n19011 = ~n10908 & ~n19010;
  assign n19012 = ~pi315 & ~n19010;
  assign n19013 = n10908 & n19010;
  assign n19014 = pi315 & n19013;
  assign n19015 = ~n19012 & ~n19014;
  assign n19016 = ~pi316 & ~n19015;
  assign n19017 = ~n19011 & ~n19016;
  assign n19018 = ~n18911 & ~n19017;
  assign n19019 = n10908 & n18910;
  assign n19020 = n17532 & n19010;
  assign n19021 = n19019 & n19020;
  assign n19022 = n10908 & n18911;
  assign n19023 = n17532 & ~n18910;
  assign n19024 = ~n17532 & n18910;
  assign n19025 = ~n19023 & ~n19024;
  assign n19026 = pi316 & ~n19025;
  assign n19027 = ~n19022 & ~n19026;
  assign n19028 = ~n19010 & ~n19027;
  assign n19029 = ~n19021 & ~n19028;
  assign n19030 = pi315 & ~n19029;
  assign n19031 = ~n17532 & n19010;
  assign n19032 = ~n10908 & ~n18910;
  assign n19033 = n19031 & n19032;
  assign n19034 = n17532 & ~n19010;
  assign n19035 = n18910 & n19034;
  assign n19036 = n17532 & n18910;
  assign n19037 = n10908 & ~n19036;
  assign n19038 = pi316 & n19037;
  assign n19039 = ~n18911 & ~n19038;
  assign n19040 = n19010 & ~n19039;
  assign n19041 = ~n19035 & ~n19040;
  assign n19042 = ~pi315 & ~n19041;
  assign n19043 = ~n19033 & ~n19042;
  assign n19044 = ~n19030 & n19043;
  assign n19045 = ~n19018 & n19044;
  assign n19046 = n17538 & ~n17541;
  assign n19047 = ~n17099 & n17104;
  assign n19048 = ~n17100 & ~n19047;
  assign n19049 = ~n17538 & n17541;
  assign n19050 = ~n19048 & ~n19049;
  assign n19051 = ~n19046 & ~n19050;
  assign n19052 = ~n19045 & n19051;
  assign n19053 = n19045 & ~n19051;
  assign n19054 = ~n19052 & ~n19053;
  assign n19055 = n9815 & ~n19054;
  assign n19056 = pi314 & n19055;
  assign n19057 = pi314 & n9815;
  assign n19058 = ~n19053 & ~n19057;
  assign n19059 = ~n19052 & n19058;
  assign n19060 = ~n19056 & ~n19059;
  assign n19061 = ~n18906 & ~n19060;
  assign n19062 = n18906 & ~n19059;
  assign n19063 = ~n19056 & n19062;
  assign n19064 = ~n19061 & ~n19063;
  assign n19065 = n18901 & ~n19064;
  assign n19066 = ~n18901 & n19064;
  assign n19067 = ~n19065 & ~n19066;
  assign n19068 = pi312 & n7874;
  assign n19069 = pi313 & ~n14735;
  assign n19070 = n17566 & ~n19069;
  assign n19071 = pi313 & ~n17566;
  assign n19072 = n14732 & n19071;
  assign n19073 = ~n19070 & ~n19072;
  assign n19074 = ~n17580 & ~n19073;
  assign n19075 = ~n7874 & n17566;
  assign n19076 = ~n17568 & ~n19075;
  assign n19077 = ~n17119 & ~n19076;
  assign n19078 = n17579 & n19077;
  assign n19079 = n14747 & ~n17566;
  assign n19080 = ~n7044 & ~n17119;
  assign n19081 = n7874 & ~n19080;
  assign n19082 = n17566 & n19081;
  assign n19083 = ~n19079 & ~n19082;
  assign n19084 = pi313 & ~n19083;
  assign n19085 = n17119 & n17590;
  assign n19086 = ~n19084 & ~n19085;
  assign n19087 = ~n17579 & ~n19086;
  assign n19088 = ~n7874 & ~n17566;
  assign n19089 = n7874 & n17566;
  assign n19090 = ~n19088 & ~n19089;
  assign n19091 = n7044 & ~n19090;
  assign n19092 = pi313 & n19091;
  assign n19093 = n17119 & n19092;
  assign n19094 = ~n19087 & ~n19093;
  assign n19095 = ~n19078 & n19094;
  assign n19096 = ~n19074 & n19095;
  assign n19097 = ~n17601 & ~n19096;
  assign n19098 = n17601 & n19096;
  assign n19099 = n17570 & ~n19098;
  assign n19100 = ~n19097 & ~n19099;
  assign n19101 = n19068 & ~n19100;
  assign n19102 = ~n17570 & ~n19097;
  assign n19103 = ~n19098 & ~n19102;
  assign n19104 = ~n19068 & ~n19103;
  assign n19105 = ~n19101 & ~n19104;
  assign n19106 = ~n19067 & ~n19105;
  assign n19107 = n18901 & n19064;
  assign n19108 = ~n18901 & ~n19064;
  assign n19109 = ~n19107 & ~n19108;
  assign n19110 = ~n19068 & ~n19100;
  assign n19111 = n19068 & ~n19103;
  assign n19112 = ~n19110 & ~n19111;
  assign n19113 = ~n19109 & ~n19112;
  assign n19114 = ~n19106 & ~n19113;
  assign n19115 = n18893 & ~n19114;
  assign n19116 = ~n18893 & n19114;
  assign n19117 = ~n19115 & ~n19116;
  assign n19118 = n7044 & ~n19117;
  assign n19119 = pi311 & n19118;
  assign n19120 = pi311 & n7044;
  assign n19121 = ~n18893 & ~n19114;
  assign n19122 = n18893 & n19114;
  assign n19123 = ~n19121 & ~n19122;
  assign n19124 = ~n19120 & ~n19123;
  assign n19125 = ~n19119 & ~n19124;
  assign n19126 = ~n5463 & ~n17621;
  assign n19127 = ~n17193 & ~n19126;
  assign n19128 = n4772 & n19127;
  assign n19129 = ~n17192 & ~n17621;
  assign n19130 = n5463 & ~n19129;
  assign n19131 = ~n19128 & ~n19130;
  assign n19132 = pi310 & ~n19131;
  assign n19133 = ~n17631 & ~n19132;
  assign n19134 = n19125 & ~n19133;
  assign n19135 = ~n19125 & n19133;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = n6777 & ~n19136;
  assign n19138 = pi310 & n19137;
  assign n19139 = pi310 & n6777;
  assign n19140 = ~n19125 & ~n19133;
  assign n19141 = n19125 & n19133;
  assign n19142 = ~n19140 & ~n19141;
  assign n19143 = ~n19139 & ~n19142;
  assign n19144 = ~n19138 & ~n19143;
  assign n19145 = n18889 & n19144;
  assign n19146 = ~n18889 & ~n19144;
  assign n19147 = ~n19145 & ~n19146;
  assign n19148 = pi308 & n4772;
  assign n19149 = pi309 & ~n9912;
  assign n19150 = n17653 & ~n19149;
  assign n19151 = pi309 & ~n17653;
  assign n19152 = n9909 & n19151;
  assign n19153 = ~n19150 & ~n19152;
  assign n19154 = ~n17668 & ~n19153;
  assign n19155 = ~n4772 & n17653;
  assign n19156 = ~n17679 & ~n19155;
  assign n19157 = n17202 & ~n19156;
  assign n19158 = n17667 & n19157;
  assign n19159 = n9924 & ~n17653;
  assign n19160 = ~n4086 & n17202;
  assign n19161 = n4772 & ~n19160;
  assign n19162 = n17653 & n19161;
  assign n19163 = ~n19159 & ~n19162;
  assign n19164 = pi309 & ~n19163;
  assign n19165 = ~n17202 & n17654;
  assign n19166 = ~n19164 & ~n19165;
  assign n19167 = ~n17667 & ~n19166;
  assign n19168 = ~n4772 & ~n17653;
  assign n19169 = n4772 & n17653;
  assign n19170 = ~n19168 & ~n19169;
  assign n19171 = n4086 & ~n19170;
  assign n19172 = pi309 & n19171;
  assign n19173 = ~n17202 & n19172;
  assign n19174 = ~n19167 & ~n19173;
  assign n19175 = ~n19158 & n19174;
  assign n19176 = ~n19154 & n19175;
  assign n19177 = n17689 & n19176;
  assign n19178 = ~n17689 & ~n19176;
  assign n19179 = n17657 & ~n19178;
  assign n19180 = ~n19177 & ~n19179;
  assign n19181 = n19148 & ~n19180;
  assign n19182 = ~n17657 & ~n19177;
  assign n19183 = ~n19178 & ~n19182;
  assign n19184 = ~n19148 & ~n19183;
  assign n19185 = ~n19181 & ~n19184;
  assign n19186 = ~n19147 & ~n19185;
  assign n19187 = n18889 & ~n19144;
  assign n19188 = ~n18889 & n19144;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~n19148 & ~n19180;
  assign n19191 = n19148 & ~n19183;
  assign n19192 = ~n19190 & ~n19191;
  assign n19193 = ~n19189 & ~n19192;
  assign n19194 = ~n19186 & ~n19193;
  assign n19195 = ~n18881 & ~n19194;
  assign n19196 = n18881 & n19194;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = n4086 & ~n19197;
  assign n19199 = pi307 & n19198;
  assign n19200 = pi307 & n4086;
  assign n19201 = n18881 & ~n19194;
  assign n19202 = ~n18881 & n19194;
  assign n19203 = ~n19201 & ~n19202;
  assign n19204 = ~n19200 & ~n19203;
  assign n19205 = ~n19199 & ~n19204;
  assign n19206 = n17696 & ~n17706;
  assign n19207 = ~n17696 & n17706;
  assign n19208 = ~n17697 & ~n19207;
  assign n19209 = ~n17268 & n19208;
  assign n19210 = ~n19206 & ~n19209;
  assign n19211 = ~n19205 & n19210;
  assign n19212 = n19205 & ~n19210;
  assign n19213 = ~n19211 & ~n19212;
  assign n19214 = n3552 & ~n19213;
  assign n19215 = pi306 & n19214;
  assign n19216 = pi306 & n3552;
  assign n19217 = n19205 & n19210;
  assign n19218 = ~n19205 & ~n19210;
  assign n19219 = ~n19217 & ~n19218;
  assign n19220 = ~n19216 & ~n19219;
  assign n19221 = ~n19215 & ~n19220;
  assign n19222 = n18875 & n19221;
  assign n19223 = ~n18875 & ~n19221;
  assign n19224 = ~n19222 & ~n19223;
  assign n19225 = pi304 & n2574;
  assign n19226 = pi305 & n17712;
  assign n19227 = n9627 & n19226;
  assign n19228 = pi305 & ~n9624;
  assign n19229 = ~n17712 & ~n19228;
  assign n19230 = ~n19227 & ~n19229;
  assign n19231 = ~n17727 & ~n19230;
  assign n19232 = ~n2574 & ~n17712;
  assign n19233 = ~n17738 & ~n19232;
  assign n19234 = ~n17273 & ~n19233;
  assign n19235 = n17726 & n19234;
  assign n19236 = n2574 & ~n17712;
  assign n19237 = ~n2574 & n17712;
  assign n19238 = ~n19236 & ~n19237;
  assign n19239 = n2183 & ~n19238;
  assign n19240 = pi305 & n19239;
  assign n19241 = n17273 & n19240;
  assign n19242 = ~n2183 & ~n17273;
  assign n19243 = n2574 & ~n19242;
  assign n19244 = ~n17712 & n19243;
  assign n19245 = n9636 & n17712;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = pi305 & ~n19246;
  assign n19248 = n17273 & n17713;
  assign n19249 = ~n19247 & ~n19248;
  assign n19250 = ~n17726 & ~n19249;
  assign n19251 = ~n19241 & ~n19250;
  assign n19252 = ~n19235 & n19251;
  assign n19253 = ~n19231 & n19252;
  assign n19254 = n17748 & n19253;
  assign n19255 = ~n17748 & ~n19253;
  assign n19256 = n17716 & ~n19255;
  assign n19257 = ~n19254 & ~n19256;
  assign n19258 = n19225 & ~n19257;
  assign n19259 = ~n17716 & ~n19254;
  assign n19260 = ~n19255 & ~n19259;
  assign n19261 = ~n19225 & ~n19260;
  assign n19262 = ~n19258 & ~n19261;
  assign n19263 = ~n19224 & ~n19262;
  assign n19264 = n18875 & ~n19221;
  assign n19265 = ~n18875 & n19221;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = ~n19225 & ~n19257;
  assign n19268 = n19225 & ~n19260;
  assign n19269 = ~n19267 & ~n19268;
  assign n19270 = ~n19266 & ~n19269;
  assign n19271 = ~n19263 & ~n19270;
  assign n19272 = ~n18867 & ~n19271;
  assign n19273 = n18867 & n19271;
  assign n19274 = ~n19272 & ~n19273;
  assign n19275 = n2183 & ~n19274;
  assign n19276 = pi303 & n19275;
  assign n19277 = pi303 & n2183;
  assign n19278 = n18867 & ~n19271;
  assign n19279 = ~n18867 & n19271;
  assign n19280 = ~n19278 & ~n19279;
  assign n19281 = ~n19277 & ~n19280;
  assign n19282 = ~n19276 & ~n19281;
  assign n19283 = ~n17754 & ~n17755;
  assign n19284 = n17754 & n17755;
  assign n19285 = ~n17342 & ~n19284;
  assign n19286 = ~n17336 & n19285;
  assign n19287 = ~n19283 & ~n19286;
  assign n19288 = ~n19282 & n19287;
  assign n19289 = n19282 & ~n19287;
  assign n19290 = ~n19288 & ~n19289;
  assign n19291 = n1840 & ~n19290;
  assign n19292 = pi302 & n19291;
  assign n19293 = pi302 & n1840;
  assign n19294 = n19282 & n19287;
  assign n19295 = ~n19282 & ~n19287;
  assign n19296 = ~n19294 & ~n19295;
  assign n19297 = ~n19293 & ~n19296;
  assign n19298 = ~n19292 & ~n19297;
  assign n19299 = n18858 & ~n19298;
  assign n19300 = ~n18858 & n19298;
  assign n19301 = ~n19299 & ~n19300;
  assign n19302 = pi300 & n1553;
  assign n19303 = n17770 & ~n17797;
  assign n19304 = ~n17782 & n19303;
  assign n19305 = ~n17770 & ~n17800;
  assign n19306 = ~n19304 & ~n19305;
  assign n19307 = ~n17406 & ~n19306;
  assign n19308 = ~n17770 & ~n17797;
  assign n19309 = ~n17782 & n19308;
  assign n19310 = n17770 & ~n17800;
  assign n19311 = ~n19309 & ~n19310;
  assign n19312 = n1553 & ~n19311;
  assign n19313 = pi301 & n19312;
  assign n19314 = ~n19307 & ~n19313;
  assign n19315 = ~n17818 & ~n19314;
  assign n19316 = n17818 & n19314;
  assign n19317 = n17783 & ~n19316;
  assign n19318 = ~n19315 & ~n19317;
  assign n19319 = n19302 & ~n19318;
  assign n19320 = ~n17783 & ~n19315;
  assign n19321 = ~n19316 & ~n19320;
  assign n19322 = ~n19302 & ~n19321;
  assign n19323 = ~n19319 & ~n19322;
  assign n19324 = ~n19301 & ~n19323;
  assign n19325 = n18858 & n19298;
  assign n19326 = ~n18858 & ~n19298;
  assign n19327 = ~n19325 & ~n19326;
  assign n19328 = ~n19302 & ~n19318;
  assign n19329 = n19302 & ~n19321;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = ~n19327 & ~n19330;
  assign n19332 = ~n19324 & ~n19331;
  assign n19333 = n18849 & ~n19332;
  assign n19334 = ~n18849 & n19332;
  assign n19335 = ~n19333 & ~n19334;
  assign n19336 = ~n17839 & n18815;
  assign n19337 = pi298 & ~n1568;
  assign n19338 = ~n19336 & ~n19337;
  assign n19339 = n19336 & n19337;
  assign n19340 = ~n19338 & ~n19339;
  assign n19341 = pi297 & ~n19340;
  assign n19342 = pi128 & n19341;
  assign n19343 = pi128 & pi297;
  assign n19344 = n19336 & ~n19337;
  assign n19345 = ~n19336 & n19337;
  assign n19346 = ~n19344 & ~n19345;
  assign n19347 = ~n19343 & ~n19346;
  assign n19348 = ~n19342 & ~n19347;
  assign n19349 = ~n19335 & ~n19348;
  assign n19350 = n18849 & n19332;
  assign n19351 = ~n18849 & ~n19332;
  assign n19352 = ~n19350 & ~n19351;
  assign n19353 = pi297 & ~n19346;
  assign n19354 = pi128 & n19353;
  assign n19355 = ~n19340 & ~n19343;
  assign n19356 = ~n19354 & ~n19355;
  assign n19357 = ~n19352 & ~n19356;
  assign n19358 = ~n19349 & ~n19357;
  assign n19359 = n1156 & ~n18784;
  assign n19360 = pi345 & n19359;
  assign n19361 = ~n18794 & ~n18803;
  assign n19362 = ~n19360 & ~n19361;
  assign n19363 = ~n18796 & ~n19362;
  assign n19364 = ~n18795 & ~n19363;
  assign n19365 = pi258 & ~n18803;
  assign n19366 = pi128 & n19365;
  assign n19367 = pi345 & n19366;
  assign n19368 = ~n17869 & n18713;
  assign n19369 = n17869 & ~n18713;
  assign n19370 = ~n19368 & ~n19369;
  assign n19371 = ~n17883 & n18717;
  assign n19372 = n17887 & ~n18730;
  assign n19373 = ~n17887 & n18730;
  assign n19374 = ~n19372 & ~n19373;
  assign n19375 = ~n19371 & ~n19374;
  assign n19376 = ~n19370 & n19375;
  assign n19377 = n17869 & n18713;
  assign n19378 = ~n17869 & ~n18713;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = ~n17887 & ~n18730;
  assign n19381 = n17887 & n18730;
  assign n19382 = ~n19380 & ~n19381;
  assign n19383 = ~n19371 & ~n19382;
  assign n19384 = ~n19379 & n19383;
  assign n19385 = n17883 & ~n18717;
  assign n19386 = ~n19384 & ~n19385;
  assign n19387 = ~n19376 & n19386;
  assign n19388 = ~n1256 & ~n18753;
  assign n19389 = pi343 & n19388;
  assign n19390 = n18753 & ~n18769;
  assign n19391 = ~n18751 & ~n18765;
  assign n19392 = ~n18762 & n19391;
  assign n19393 = n18751 & ~n18766;
  assign n19394 = ~n19392 & ~n19393;
  assign n19395 = ~n19390 & ~n19394;
  assign n19396 = ~n19389 & ~n19395;
  assign n19397 = n19387 & n19396;
  assign n19398 = ~n19387 & ~n19396;
  assign n19399 = ~n19397 & ~n19398;
  assign n19400 = pi341 & n2091;
  assign n19401 = n17908 & ~n18609;
  assign n19402 = ~n17908 & n18609;
  assign n19403 = ~n19401 & ~n19402;
  assign n19404 = ~n17922 & n18613;
  assign n19405 = n17926 & ~n18629;
  assign n19406 = ~n17926 & n18629;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = ~n19404 & ~n19407;
  assign n19409 = ~n19403 & n19408;
  assign n19410 = n17908 & n18609;
  assign n19411 = ~n17908 & ~n18609;
  assign n19412 = ~n19410 & ~n19411;
  assign n19413 = ~n17926 & ~n18629;
  assign n19414 = n17926 & n18629;
  assign n19415 = ~n19413 & ~n19414;
  assign n19416 = ~n19404 & ~n19415;
  assign n19417 = ~n19412 & n19416;
  assign n19418 = n17922 & ~n18613;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = ~n19409 & n19419;
  assign n19421 = ~n18657 & n18661;
  assign n19422 = ~n18650 & ~n18674;
  assign n19423 = n18650 & n18674;
  assign n19424 = ~n19422 & ~n19423;
  assign n19425 = n18657 & ~n18661;
  assign n19426 = ~n19424 & ~n19425;
  assign n19427 = ~n19421 & ~n19426;
  assign n19428 = n19420 & n19427;
  assign n19429 = ~n19420 & ~n19427;
  assign n19430 = ~n19428 & ~n19429;
  assign n19431 = n4596 & ~n18662;
  assign n19432 = pi336 & n19431;
  assign n19433 = ~n18663 & ~n19432;
  assign n19434 = ~n18650 & n19433;
  assign n19435 = n18650 & ~n19433;
  assign n19436 = ~n5257 & ~n19435;
  assign n19437 = ~n19434 & ~n19436;
  assign n19438 = n5714 & ~n19437;
  assign n19439 = ~n5714 & ~n19434;
  assign n19440 = n5257 & n19439;
  assign n19441 = ~n19438 & ~n19440;
  assign n19442 = pi336 & ~n19441;
  assign n19443 = pi336 & n5714;
  assign n19444 = n18650 & ~n19443;
  assign n19445 = ~n19433 & n19444;
  assign n19446 = ~n19442 & ~n19445;
  assign n19447 = ~n17943 & ~n17947;
  assign n19448 = n17943 & n17947;
  assign n19449 = ~n17931 & n18523;
  assign n19450 = n17931 & ~n18523;
  assign n19451 = ~n19449 & ~n19450;
  assign n19452 = n11384 & ~n19451;
  assign n19453 = pi328 & n19452;
  assign n19454 = ~n17931 & ~n18523;
  assign n19455 = n17931 & n18523;
  assign n19456 = ~n19454 & ~n19455;
  assign n19457 = ~n18529 & ~n19456;
  assign n19458 = ~n19453 & ~n19457;
  assign n19459 = ~n19448 & ~n19458;
  assign n19460 = ~n19447 & ~n19459;
  assign n19461 = ~n18559 & n18563;
  assign n19462 = ~n18544 & ~n18570;
  assign n19463 = n18544 & n18570;
  assign n19464 = ~n19462 & ~n19463;
  assign n19465 = n18559 & ~n18563;
  assign n19466 = ~n19464 & ~n19465;
  assign n19467 = ~n19461 & ~n19466;
  assign n19468 = n19460 & n19467;
  assign n19469 = ~n19460 & ~n19467;
  assign n19470 = ~n19468 & ~n19469;
  assign n19471 = ~n18544 & n18565;
  assign n19472 = n18544 & ~n18565;
  assign n19473 = ~n10561 & ~n19472;
  assign n19474 = ~n19471 & ~n19473;
  assign n19475 = n11366 & ~n19474;
  assign n19476 = ~n11366 & ~n19471;
  assign n19477 = n10561 & n19476;
  assign n19478 = ~n19475 & ~n19477;
  assign n19479 = pi330 & ~n19478;
  assign n19480 = pi330 & n11366;
  assign n19481 = n18544 & ~n19480;
  assign n19482 = ~n18565 & n19481;
  assign n19483 = ~n19479 & ~n19482;
  assign n19484 = ~n17951 & ~n18497;
  assign n19485 = n17951 & n18497;
  assign n19486 = ~n19484 & ~n19485;
  assign n19487 = n17971 & n18501;
  assign n19488 = ~n18482 & n18502;
  assign n19489 = n18482 & ~n18502;
  assign n19490 = ~n19488 & ~n19489;
  assign n19491 = ~n19487 & ~n19490;
  assign n19492 = ~n19486 & n19491;
  assign n19493 = ~n17951 & n18497;
  assign n19494 = n17951 & ~n18497;
  assign n19495 = ~n19493 & ~n19494;
  assign n19496 = n18482 & n18502;
  assign n19497 = ~n18482 & ~n18502;
  assign n19498 = ~n19496 & ~n19497;
  assign n19499 = ~n19487 & ~n19498;
  assign n19500 = ~n19495 & n19499;
  assign n19501 = ~n17971 & ~n18501;
  assign n19502 = ~n19500 & ~n19501;
  assign n19503 = ~n19492 & n19502;
  assign n19504 = n11384 & ~n19455;
  assign n19505 = pi328 & n19504;
  assign n19506 = ~n19454 & ~n19505;
  assign n19507 = n19503 & ~n19506;
  assign n19508 = ~n19503 & n19506;
  assign n19509 = ~n19507 & ~n19508;
  assign n19510 = pi327 & n12917;
  assign n19511 = n18458 & ~n18497;
  assign n19512 = ~n17976 & ~n18457;
  assign n19513 = n17976 & ~n18456;
  assign n19514 = ~n18450 & n19513;
  assign n19515 = ~n19512 & ~n19514;
  assign n19516 = ~n18462 & ~n19515;
  assign n19517 = n17976 & ~n18457;
  assign n19518 = ~n17976 & ~n18456;
  assign n19519 = ~n18450 & n19518;
  assign n19520 = ~n19517 & ~n19519;
  assign n19521 = n18461 & ~n19520;
  assign n19522 = pi324 & n19521;
  assign n19523 = ~n19516 & ~n19522;
  assign n19524 = n17984 & ~n19523;
  assign n19525 = ~n17984 & n19523;
  assign n19526 = ~n19524 & ~n19525;
  assign n19527 = ~n18458 & n18497;
  assign n19528 = ~n19526 & ~n19527;
  assign n19529 = ~n19511 & ~n19528;
  assign n19530 = ~n17951 & n18502;
  assign n19531 = n17951 & ~n18502;
  assign n19532 = ~n18509 & ~n19531;
  assign n19533 = ~n19530 & ~n19532;
  assign n19534 = n19529 & ~n19533;
  assign n19535 = ~n19529 & n19533;
  assign n19536 = ~n19534 & ~n19535;
  assign n19537 = ~n15616 & ~n17996;
  assign n19538 = n15616 & ~n17992;
  assign n19539 = ~n19537 & ~n19538;
  assign n19540 = pi324 & n19539;
  assign n19541 = ~n17976 & ~n18450;
  assign n19542 = ~n18456 & ~n19541;
  assign n19543 = ~n19540 & ~n19542;
  assign n19544 = n19540 & n19542;
  assign n19545 = ~n19543 & ~n19544;
  assign n19546 = ~n18000 & n18434;
  assign n19547 = n18000 & ~n18434;
  assign n19548 = ~n19546 & ~n19547;
  assign n19549 = n18436 & ~n19548;
  assign n19550 = ~n18436 & n19548;
  assign n19551 = ~n19549 & ~n19550;
  assign n19552 = ~n16527 & ~n19551;
  assign n19553 = ~n18436 & ~n19548;
  assign n19554 = n18436 & n19548;
  assign n19555 = ~n19553 & ~n19554;
  assign n19556 = n16527 & ~n19555;
  assign n19557 = ~n19552 & ~n19556;
  assign n19558 = pi323 & n19557;
  assign n19559 = ~n18014 & n18018;
  assign n19560 = n18014 & ~n18018;
  assign n19561 = pi262 & ~n18392;
  assign n19562 = pi147 & n19561;
  assign n19563 = ~n18383 & ~n18385;
  assign n19564 = ~n19562 & ~n19563;
  assign n19565 = pi261 & ~n19564;
  assign n19566 = pi148 & n19565;
  assign n19567 = ~n18384 & ~n19563;
  assign n19568 = ~n19562 & n19567;
  assign n19569 = ~n19566 & ~n19568;
  assign n19570 = ~n18007 & ~n19569;
  assign n19571 = n18007 & n19569;
  assign n19572 = ~n19570 & ~n19571;
  assign n19573 = ~n19560 & ~n19572;
  assign n19574 = ~n19559 & ~n19573;
  assign n19575 = ~n18402 & ~n18414;
  assign n19576 = ~n18017 & n19575;
  assign n19577 = ~n18414 & ~n18420;
  assign n19578 = ~n18429 & n19577;
  assign n19579 = ~n18415 & ~n19578;
  assign n19580 = ~n19576 & n19579;
  assign n19581 = n19574 & n19580;
  assign n19582 = ~n19574 & ~n19580;
  assign n19583 = ~n19581 & ~n19582;
  assign n19584 = pi149 & pi261;
  assign n19585 = pi145 & pi265;
  assign n19586 = pi142 & pi268;
  assign n19587 = pi139 & pi271;
  assign n19588 = pi136 & pi274;
  assign n19589 = pi133 & pi277;
  assign n19590 = ~n18041 & ~n18055;
  assign n19591 = n18024 & n18027;
  assign n19592 = ~n18024 & ~n18027;
  assign n19593 = ~n18038 & ~n19592;
  assign n19594 = ~n19591 & ~n19593;
  assign n19595 = pi128 & pi282;
  assign n19596 = pi281 & ~n19595;
  assign n19597 = pi129 & n19596;
  assign n19598 = pi129 & pi281;
  assign n19599 = pi282 & ~n19598;
  assign n19600 = pi128 & n19599;
  assign n19601 = ~n19597 & ~n19600;
  assign n19602 = ~n19594 & n19601;
  assign n19603 = n19594 & ~n19601;
  assign n19604 = ~n19602 & ~n19603;
  assign n19605 = pi280 & ~n19604;
  assign n19606 = pi130 & n19605;
  assign n19607 = pi130 & pi280;
  assign n19608 = ~n19603 & ~n19607;
  assign n19609 = ~n19602 & n19608;
  assign n19610 = ~n19606 & ~n19609;
  assign n19611 = ~n19590 & ~n19610;
  assign n19612 = ~n18045 & n19611;
  assign n19613 = ~n18045 & ~n19590;
  assign n19614 = ~n19609 & ~n19613;
  assign n19615 = ~n19606 & n19614;
  assign n19616 = ~n19612 & ~n19615;
  assign n19617 = pi279 & ~n19616;
  assign n19618 = pi131 & n19617;
  assign n19619 = pi131 & pi279;
  assign n19620 = ~n19615 & ~n19619;
  assign n19621 = ~n19612 & n19620;
  assign n19622 = ~n19618 & ~n19621;
  assign n19623 = ~n18065 & ~n18066;
  assign n19624 = ~n18062 & ~n19623;
  assign n19625 = ~n19622 & n19624;
  assign n19626 = n19622 & ~n19624;
  assign n19627 = ~n19625 & ~n19626;
  assign n19628 = pi132 & pi278;
  assign n19629 = n18022 & ~n18073;
  assign n19630 = n19628 & ~n19629;
  assign n19631 = ~n18076 & n19630;
  assign n19632 = ~n18076 & ~n19629;
  assign n19633 = ~n19628 & ~n19632;
  assign n19634 = ~n19631 & ~n19633;
  assign n19635 = ~n19627 & ~n19634;
  assign n19636 = ~n19622 & ~n19624;
  assign n19637 = n19622 & n19624;
  assign n19638 = ~n19636 & ~n19637;
  assign n19639 = ~n19628 & ~n19629;
  assign n19640 = ~n18076 & n19639;
  assign n19641 = n19628 & ~n19632;
  assign n19642 = ~n19640 & ~n19641;
  assign n19643 = ~n19638 & ~n19642;
  assign n19644 = ~n19635 & ~n19643;
  assign n19645 = ~n19589 & n19644;
  assign n19646 = n19589 & ~n19644;
  assign n19647 = ~n19645 & ~n19646;
  assign n19648 = pi276 & ~n18081;
  assign n19649 = pi133 & n19648;
  assign n19650 = pi134 & pi276;
  assign n19651 = ~n18019 & ~n18080;
  assign n19652 = ~n18078 & n19651;
  assign n19653 = ~n18111 & ~n19652;
  assign n19654 = ~n19650 & ~n19653;
  assign n19655 = ~n19649 & n19654;
  assign n19656 = ~n19649 & ~n19653;
  assign n19657 = n19650 & ~n19656;
  assign n19658 = ~n19655 & ~n19657;
  assign n19659 = ~n19647 & ~n19658;
  assign n19660 = ~n19589 & ~n19644;
  assign n19661 = n19589 & n19644;
  assign n19662 = ~n19660 & ~n19661;
  assign n19663 = n19650 & ~n19653;
  assign n19664 = ~n19649 & n19663;
  assign n19665 = ~n19650 & ~n19656;
  assign n19666 = ~n19664 & ~n19665;
  assign n19667 = ~n19662 & ~n19666;
  assign n19668 = ~n19659 & ~n19667;
  assign n19669 = n18115 & ~n18133;
  assign n19670 = ~n18115 & n18133;
  assign n19671 = ~n18124 & ~n19670;
  assign n19672 = ~n19669 & ~n19671;
  assign n19673 = n19668 & n19672;
  assign n19674 = ~n19668 & ~n19672;
  assign n19675 = ~n19673 & ~n19674;
  assign n19676 = pi135 & pi275;
  assign n19677 = n18147 & ~n18153;
  assign n19678 = ~n18152 & ~n19677;
  assign n19679 = n19676 & ~n19678;
  assign n19680 = ~n18147 & ~n18152;
  assign n19681 = ~n18153 & ~n19680;
  assign n19682 = ~n19676 & ~n19681;
  assign n19683 = ~n19679 & ~n19682;
  assign n19684 = ~n19675 & ~n19683;
  assign n19685 = n19668 & ~n19672;
  assign n19686 = ~n19668 & n19672;
  assign n19687 = ~n19685 & ~n19686;
  assign n19688 = ~n19676 & ~n19678;
  assign n19689 = n19676 & ~n19681;
  assign n19690 = ~n19688 & ~n19689;
  assign n19691 = ~n19687 & ~n19690;
  assign n19692 = ~n19684 & ~n19691;
  assign n19693 = ~n19588 & n19692;
  assign n19694 = n19588 & ~n19692;
  assign n19695 = ~n19693 & ~n19694;
  assign n19696 = pi274 & ~n18154;
  assign n19697 = pi135 & n19696;
  assign n19698 = ~n18145 & ~n18147;
  assign n19699 = ~n19697 & ~n19698;
  assign n19700 = pi273 & ~n19699;
  assign n19701 = pi136 & n19700;
  assign n19702 = pi137 & pi273;
  assign n19703 = ~n18146 & ~n19698;
  assign n19704 = ~n19697 & n19703;
  assign n19705 = ~n18163 & ~n19704;
  assign n19706 = ~n19702 & ~n19705;
  assign n19707 = ~n19701 & n19706;
  assign n19708 = ~n19701 & ~n19705;
  assign n19709 = n19702 & ~n19708;
  assign n19710 = ~n19707 & ~n19709;
  assign n19711 = ~n19695 & ~n19710;
  assign n19712 = ~n19588 & ~n19692;
  assign n19713 = n19588 & n19692;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = n19702 & ~n19705;
  assign n19716 = ~n19701 & n19715;
  assign n19717 = ~n19702 & ~n19708;
  assign n19718 = ~n19716 & ~n19717;
  assign n19719 = ~n19714 & ~n19718;
  assign n19720 = ~n19711 & ~n19719;
  assign n19721 = n18167 & ~n18192;
  assign n19722 = ~n18167 & n18192;
  assign n19723 = ~n18183 & ~n19722;
  assign n19724 = ~n19721 & ~n19723;
  assign n19725 = n19720 & ~n19724;
  assign n19726 = ~n19720 & n19724;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = pi138 & pi272;
  assign n19729 = n18206 & ~n18212;
  assign n19730 = ~n18211 & ~n19729;
  assign n19731 = n19728 & ~n19730;
  assign n19732 = ~n18206 & ~n18211;
  assign n19733 = ~n18212 & ~n19732;
  assign n19734 = ~n19728 & ~n19733;
  assign n19735 = ~n19731 & ~n19734;
  assign n19736 = ~n19727 & ~n19735;
  assign n19737 = n19720 & n19724;
  assign n19738 = ~n19720 & ~n19724;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = ~n19728 & ~n19730;
  assign n19741 = n19728 & ~n19733;
  assign n19742 = ~n19740 & ~n19741;
  assign n19743 = ~n19739 & ~n19742;
  assign n19744 = ~n19736 & ~n19743;
  assign n19745 = ~n19587 & ~n19744;
  assign n19746 = n19587 & n19744;
  assign n19747 = ~n19745 & ~n19746;
  assign n19748 = pi271 & ~n18213;
  assign n19749 = pi138 & n19748;
  assign n19750 = ~n18204 & ~n18206;
  assign n19751 = ~n18205 & ~n19750;
  assign n19752 = ~n19749 & n19751;
  assign n19753 = pi140 & pi270;
  assign n19754 = ~n19749 & ~n19750;
  assign n19755 = pi270 & ~n19754;
  assign n19756 = pi139 & n19755;
  assign n19757 = n18223 & ~n19756;
  assign n19758 = n19753 & ~n19757;
  assign n19759 = ~n19752 & n19758;
  assign n19760 = ~n19752 & ~n19757;
  assign n19761 = ~n19753 & ~n19760;
  assign n19762 = ~n19759 & ~n19761;
  assign n19763 = ~n19747 & ~n19762;
  assign n19764 = ~n19587 & n19744;
  assign n19765 = n19587 & ~n19744;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~n19753 & ~n19757;
  assign n19768 = ~n19752 & n19767;
  assign n19769 = n19753 & ~n19760;
  assign n19770 = ~n19768 & ~n19769;
  assign n19771 = ~n19766 & ~n19770;
  assign n19772 = ~n19763 & ~n19771;
  assign n19773 = ~n18226 & ~n18227;
  assign n19774 = n18226 & n18227;
  assign n19775 = ~n18246 & ~n19774;
  assign n19776 = ~n19773 & ~n19775;
  assign n19777 = n19772 & n19776;
  assign n19778 = ~n19772 & ~n19776;
  assign n19779 = ~n19777 & ~n19778;
  assign n19780 = pi141 & pi269;
  assign n19781 = n18266 & ~n18272;
  assign n19782 = ~n18271 & ~n19781;
  assign n19783 = n19780 & ~n19782;
  assign n19784 = ~n18266 & ~n18271;
  assign n19785 = ~n18272 & ~n19784;
  assign n19786 = ~n19780 & ~n19785;
  assign n19787 = ~n19783 & ~n19786;
  assign n19788 = ~n19779 & ~n19787;
  assign n19789 = n19772 & ~n19776;
  assign n19790 = ~n19772 & n19776;
  assign n19791 = ~n19789 & ~n19790;
  assign n19792 = ~n19780 & ~n19782;
  assign n19793 = n19780 & ~n19785;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = ~n19791 & ~n19794;
  assign n19796 = ~n19788 & ~n19795;
  assign n19797 = ~n19586 & ~n19796;
  assign n19798 = n19586 & n19796;
  assign n19799 = ~n19797 & ~n19798;
  assign n19800 = pi268 & ~n18273;
  assign n19801 = pi141 & n19800;
  assign n19802 = ~n18264 & ~n18266;
  assign n19803 = ~n18265 & ~n19802;
  assign n19804 = ~n19801 & n19803;
  assign n19805 = pi143 & pi267;
  assign n19806 = ~n19801 & ~n19802;
  assign n19807 = pi267 & ~n19806;
  assign n19808 = pi142 & n19807;
  assign n19809 = n18283 & ~n19808;
  assign n19810 = n19805 & ~n19809;
  assign n19811 = ~n19804 & n19810;
  assign n19812 = ~n19804 & ~n19809;
  assign n19813 = ~n19805 & ~n19812;
  assign n19814 = ~n19811 & ~n19813;
  assign n19815 = ~n19799 & ~n19814;
  assign n19816 = ~n19586 & n19796;
  assign n19817 = n19586 & ~n19796;
  assign n19818 = ~n19816 & ~n19817;
  assign n19819 = ~n19805 & ~n19809;
  assign n19820 = ~n19804 & n19819;
  assign n19821 = n19805 & ~n19812;
  assign n19822 = ~n19820 & ~n19821;
  assign n19823 = ~n19818 & ~n19822;
  assign n19824 = ~n19815 & ~n19823;
  assign n19825 = ~n18287 & ~n18312;
  assign n19826 = n18287 & n18312;
  assign n19827 = ~n18306 & ~n19826;
  assign n19828 = ~n19825 & ~n19827;
  assign n19829 = n19824 & ~n19828;
  assign n19830 = ~n19824 & n19828;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = pi144 & pi266;
  assign n19833 = n18326 & ~n18331;
  assign n19834 = ~n18332 & ~n19833;
  assign n19835 = n19832 & ~n19834;
  assign n19836 = ~n18326 & ~n18332;
  assign n19837 = ~n18331 & ~n19836;
  assign n19838 = ~n19832 & ~n19837;
  assign n19839 = ~n19835 & ~n19838;
  assign n19840 = ~n19831 & ~n19839;
  assign n19841 = n19824 & n19828;
  assign n19842 = ~n19824 & ~n19828;
  assign n19843 = ~n19841 & ~n19842;
  assign n19844 = ~n19832 & ~n19834;
  assign n19845 = n19832 & ~n19837;
  assign n19846 = ~n19844 & ~n19845;
  assign n19847 = ~n19843 & ~n19846;
  assign n19848 = ~n19840 & ~n19847;
  assign n19849 = ~n19585 & n19848;
  assign n19850 = n19585 & ~n19848;
  assign n19851 = ~n19849 & ~n19850;
  assign n19852 = pi265 & ~n18333;
  assign n19853 = pi144 & n19852;
  assign n19854 = ~n18324 & ~n18326;
  assign n19855 = ~n19853 & ~n19854;
  assign n19856 = pi264 & ~n19855;
  assign n19857 = pi145 & n19856;
  assign n19858 = pi146 & pi264;
  assign n19859 = ~n18325 & ~n19854;
  assign n19860 = ~n19853 & n19859;
  assign n19861 = ~n18342 & ~n19860;
  assign n19862 = ~n19858 & ~n19861;
  assign n19863 = ~n19857 & n19862;
  assign n19864 = ~n19857 & ~n19861;
  assign n19865 = n19858 & ~n19864;
  assign n19866 = ~n19863 & ~n19865;
  assign n19867 = ~n19851 & ~n19866;
  assign n19868 = ~n19585 & ~n19848;
  assign n19869 = n19585 & n19848;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = n19858 & ~n19861;
  assign n19872 = ~n19857 & n19871;
  assign n19873 = ~n19858 & ~n19864;
  assign n19874 = ~n19872 & ~n19873;
  assign n19875 = ~n19870 & ~n19874;
  assign n19876 = ~n19867 & ~n19875;
  assign n19877 = ~n18346 & ~n18371;
  assign n19878 = n18346 & n18371;
  assign n19879 = ~n18365 & ~n19878;
  assign n19880 = ~n19877 & ~n19879;
  assign n19881 = n19876 & ~n19880;
  assign n19882 = ~n19876 & n19880;
  assign n19883 = ~n19881 & ~n19882;
  assign n19884 = pi263 & ~n19883;
  assign n19885 = pi147 & n19884;
  assign n19886 = pi147 & pi263;
  assign n19887 = ~n19876 & ~n19880;
  assign n19888 = n19876 & n19880;
  assign n19889 = ~n19887 & ~n19888;
  assign n19890 = ~n19886 & ~n19889;
  assign n19891 = ~n19885 & ~n19890;
  assign n19892 = ~n18380 & n18385;
  assign n19893 = n18380 & ~n18385;
  assign n19894 = ~n18376 & ~n19893;
  assign n19895 = ~n19892 & ~n19894;
  assign n19896 = n19891 & ~n19895;
  assign n19897 = ~n19891 & n19895;
  assign n19898 = ~n19896 & ~n19897;
  assign n19899 = pi148 & pi262;
  assign n19900 = ~n18007 & ~n19568;
  assign n19901 = ~n19899 & ~n19900;
  assign n19902 = ~n19566 & n19901;
  assign n19903 = ~n19566 & ~n19900;
  assign n19904 = n19899 & ~n19903;
  assign n19905 = ~n19902 & ~n19904;
  assign n19906 = ~n19898 & ~n19905;
  assign n19907 = n19891 & n19895;
  assign n19908 = ~n19891 & ~n19895;
  assign n19909 = ~n19907 & ~n19908;
  assign n19910 = n19899 & ~n19900;
  assign n19911 = ~n19566 & n19910;
  assign n19912 = ~n19899 & ~n19903;
  assign n19913 = ~n19911 & ~n19912;
  assign n19914 = ~n19909 & ~n19913;
  assign n19915 = ~n19906 & ~n19914;
  assign n19916 = ~n19584 & n19915;
  assign n19917 = n19584 & ~n19915;
  assign n19918 = ~n19916 & ~n19917;
  assign n19919 = pi260 & ~n19918;
  assign n19920 = pi150 & n19919;
  assign n19921 = pi150 & pi260;
  assign n19922 = n19584 & n19915;
  assign n19923 = ~n19584 & ~n19915;
  assign n19924 = ~n19922 & ~n19923;
  assign n19925 = ~n19921 & ~n19924;
  assign n19926 = ~n19920 & ~n19925;
  assign n19927 = ~n19583 & ~n19926;
  assign n19928 = n19574 & ~n19580;
  assign n19929 = ~n19574 & n19580;
  assign n19930 = ~n19928 & ~n19929;
  assign n19931 = pi260 & ~n19924;
  assign n19932 = pi150 & n19931;
  assign n19933 = ~n19918 & ~n19921;
  assign n19934 = ~n19932 & ~n19933;
  assign n19935 = ~n19930 & ~n19934;
  assign n19936 = ~n19927 & ~n19935;
  assign n19937 = ~n16527 & ~n18436;
  assign n19938 = n16527 & n18436;
  assign n19939 = ~n19548 & ~n19938;
  assign n19940 = ~n19937 & ~n19939;
  assign n19941 = n19936 & n19940;
  assign n19942 = ~n19936 & ~n19940;
  assign n19943 = ~n19941 & ~n19942;
  assign n19944 = pi258 & n18434;
  assign n19945 = pi259 & ~n19944;
  assign n19946 = ~pi259 & n18434;
  assign n19947 = pi258 & n19946;
  assign n19948 = ~n19945 & ~n19947;
  assign n19949 = pi151 & ~n19948;
  assign n19950 = n19548 & ~n19949;
  assign n19951 = ~n19548 & n19949;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = pi258 & ~n19952;
  assign n19954 = pi152 & n19953;
  assign n19955 = pi152 & pi258;
  assign n19956 = ~n19548 & ~n19949;
  assign n19957 = n19548 & n19949;
  assign n19958 = ~n19956 & ~n19957;
  assign n19959 = ~n19955 & ~n19958;
  assign n19960 = ~n19954 & ~n19959;
  assign n19961 = ~n19943 & ~n19960;
  assign n19962 = n19936 & ~n19940;
  assign n19963 = ~n19936 & n19940;
  assign n19964 = ~n19962 & ~n19963;
  assign n19965 = pi258 & ~n19958;
  assign n19966 = pi152 & n19965;
  assign n19967 = ~n19952 & ~n19955;
  assign n19968 = ~n19966 & ~n19967;
  assign n19969 = ~n19964 & ~n19968;
  assign n19970 = ~n19961 & ~n19969;
  assign n19971 = pi322 & n19970;
  assign n19972 = ~n19558 & ~n19971;
  assign n19973 = n19557 & n19970;
  assign n19974 = n1445 & n19973;
  assign n19975 = ~n19972 & ~n19974;
  assign n19976 = ~n19545 & ~n19975;
  assign n19977 = ~n19540 & n19542;
  assign n19978 = n19540 & ~n19542;
  assign n19979 = ~n19977 & ~n19978;
  assign n19980 = ~n19558 & n19970;
  assign n19981 = pi322 & n19980;
  assign n19982 = n19557 & ~n19971;
  assign n19983 = pi323 & n19982;
  assign n19984 = ~n19981 & ~n19983;
  assign n19985 = ~n19979 & ~n19984;
  assign n19986 = ~n19976 & ~n19985;
  assign n19987 = ~n17984 & n18462;
  assign n19988 = n17984 & ~n18462;
  assign n19989 = ~n19515 & ~n19988;
  assign n19990 = ~n19987 & ~n19989;
  assign n19991 = n19986 & ~n19990;
  assign n19992 = ~n19986 & n19990;
  assign n19993 = ~n19991 & ~n19992;
  assign n19994 = pi326 & n13762;
  assign n19995 = pi325 & n18461;
  assign n19996 = n19994 & n19995;
  assign n19997 = ~n19994 & ~n19995;
  assign n19998 = ~n19996 & ~n19997;
  assign n19999 = ~n19993 & ~n19998;
  assign n20000 = ~n19986 & ~n19990;
  assign n20001 = n19986 & n19990;
  assign n20002 = ~n20000 & ~n20001;
  assign n20003 = ~n19994 & n19995;
  assign n20004 = n19994 & ~n19995;
  assign n20005 = ~n20003 & ~n20004;
  assign n20006 = ~n20002 & ~n20005;
  assign n20007 = ~n19999 & ~n20006;
  assign n20008 = ~n19536 & ~n20007;
  assign n20009 = n19529 & n19533;
  assign n20010 = ~n19529 & ~n19533;
  assign n20011 = ~n20009 & ~n20010;
  assign n20012 = ~n19998 & ~n20002;
  assign n20013 = ~n19993 & ~n20005;
  assign n20014 = ~n20012 & ~n20013;
  assign n20015 = ~n20011 & ~n20014;
  assign n20016 = ~n20008 & ~n20015;
  assign n20017 = ~n19510 & n20016;
  assign n20018 = n19510 & ~n20016;
  assign n20019 = ~n20017 & ~n20018;
  assign n20020 = pi329 & n11384;
  assign n20021 = pi328 & n11711;
  assign n20022 = n20020 & n20021;
  assign n20023 = ~n20020 & ~n20021;
  assign n20024 = ~n20022 & ~n20023;
  assign n20025 = ~n20019 & ~n20024;
  assign n20026 = n19510 & n20016;
  assign n20027 = ~n19510 & ~n20016;
  assign n20028 = ~n20026 & ~n20027;
  assign n20029 = ~n20020 & n20021;
  assign n20030 = n20020 & ~n20021;
  assign n20031 = ~n20029 & ~n20030;
  assign n20032 = ~n20028 & ~n20031;
  assign n20033 = ~n20025 & ~n20032;
  assign n20034 = ~n19509 & ~n20033;
  assign n20035 = n19503 & n19506;
  assign n20036 = ~n19503 & ~n19506;
  assign n20037 = ~n20035 & ~n20036;
  assign n20038 = ~n20024 & ~n20028;
  assign n20039 = ~n20019 & ~n20031;
  assign n20040 = ~n20038 & ~n20039;
  assign n20041 = ~n20037 & ~n20040;
  assign n20042 = ~n20034 & ~n20041;
  assign n20043 = n19483 & n20042;
  assign n20044 = ~n19483 & ~n20042;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = n10561 & ~n20045;
  assign n20047 = pi331 & n20046;
  assign n20048 = pi331 & n10561;
  assign n20049 = ~n19483 & n20042;
  assign n20050 = n19483 & ~n20042;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = ~n20048 & ~n20051;
  assign n20053 = ~n20047 & ~n20052;
  assign n20054 = ~n19470 & ~n20053;
  assign n20055 = n19460 & ~n19467;
  assign n20056 = ~n19460 & n19467;
  assign n20057 = ~n20055 & ~n20056;
  assign n20058 = n10561 & ~n20051;
  assign n20059 = pi331 & n20058;
  assign n20060 = ~n20045 & ~n20048;
  assign n20061 = ~n20059 & ~n20060;
  assign n20062 = ~n20057 & ~n20061;
  assign n20063 = ~n20054 & ~n20062;
  assign n20064 = ~n17908 & n17926;
  assign n20065 = n17908 & ~n17926;
  assign n20066 = n18609 & ~n20065;
  assign n20067 = ~n20064 & ~n20066;
  assign n20068 = n20063 & n20067;
  assign n20069 = ~n20063 & ~n20067;
  assign n20070 = ~n20068 & ~n20069;
  assign n20071 = pi333 & n6556;
  assign n20072 = ~n18573 & ~n18597;
  assign n20073 = ~n18604 & n20072;
  assign n20074 = ~n18595 & ~n18597;
  assign n20075 = ~n18562 & n20074;
  assign n20076 = ~n18596 & ~n20075;
  assign n20077 = ~n20073 & n20076;
  assign n20078 = pi332 & n9205;
  assign n20079 = n20077 & ~n20078;
  assign n20080 = n9205 & ~n20077;
  assign n20081 = pi332 & n20080;
  assign n20082 = ~n20079 & ~n20081;
  assign n20083 = ~n20071 & n20082;
  assign n20084 = n20071 & ~n20082;
  assign n20085 = ~n20083 & ~n20084;
  assign n20086 = pi335 & n5732;
  assign n20087 = pi334 & n5973;
  assign n20088 = ~n18618 & ~n18625;
  assign n20089 = ~n18614 & n20088;
  assign n20090 = ~n20087 & ~n20089;
  assign n20091 = n17926 & n20090;
  assign n20092 = n18614 & ~n20088;
  assign n20093 = n20087 & ~n20092;
  assign n20094 = ~n17926 & n20093;
  assign n20095 = ~n20091 & ~n20094;
  assign n20096 = ~n19403 & ~n20095;
  assign n20097 = n17926 & n20093;
  assign n20098 = ~n17926 & n20090;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~n19412 & ~n20099;
  assign n20101 = ~n20087 & ~n20088;
  assign n20102 = n18614 & n20101;
  assign n20103 = n20087 & n20088;
  assign n20104 = ~n18614 & n20103;
  assign n20105 = ~n20102 & ~n20104;
  assign n20106 = ~n20100 & n20105;
  assign n20107 = ~n20096 & n20106;
  assign n20108 = n20086 & ~n20107;
  assign n20109 = ~n20086 & n20107;
  assign n20110 = ~n20108 & ~n20109;
  assign n20111 = ~n20085 & ~n20110;
  assign n20112 = n20071 & n20082;
  assign n20113 = ~n20071 & ~n20082;
  assign n20114 = ~n20112 & ~n20113;
  assign n20115 = ~n20086 & ~n20107;
  assign n20116 = n20086 & n20107;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = ~n20114 & ~n20117;
  assign n20119 = ~n20111 & ~n20118;
  assign n20120 = ~n20070 & ~n20119;
  assign n20121 = n20063 & ~n20067;
  assign n20122 = ~n20063 & n20067;
  assign n20123 = ~n20121 & ~n20122;
  assign n20124 = ~n20110 & ~n20114;
  assign n20125 = ~n20085 & ~n20117;
  assign n20126 = ~n20124 & ~n20125;
  assign n20127 = ~n20123 & ~n20126;
  assign n20128 = ~n20120 & ~n20127;
  assign n20129 = n19446 & n20128;
  assign n20130 = ~n19446 & ~n20128;
  assign n20131 = ~n20129 & ~n20130;
  assign n20132 = n5257 & ~n20131;
  assign n20133 = pi337 & n20132;
  assign n20134 = pi337 & n5257;
  assign n20135 = ~n19446 & n20128;
  assign n20136 = n19446 & ~n20128;
  assign n20137 = ~n20135 & ~n20136;
  assign n20138 = ~n20134 & ~n20137;
  assign n20139 = ~n20133 & ~n20138;
  assign n20140 = ~n19430 & ~n20139;
  assign n20141 = n19420 & ~n19427;
  assign n20142 = ~n19420 & n19427;
  assign n20143 = ~n20141 & ~n20142;
  assign n20144 = n5257 & ~n20137;
  assign n20145 = pi337 & n20144;
  assign n20146 = ~n20131 & ~n20134;
  assign n20147 = ~n20145 & ~n20146;
  assign n20148 = ~n20143 & ~n20147;
  assign n20149 = ~n20140 & ~n20148;
  assign n20150 = ~n17869 & n17887;
  assign n20151 = n17869 & ~n17887;
  assign n20152 = n18713 & ~n20151;
  assign n20153 = ~n20150 & ~n20152;
  assign n20154 = n20149 & n20153;
  assign n20155 = ~n20149 & ~n20153;
  assign n20156 = ~n20154 & ~n20155;
  assign n20157 = pi339 & n2887;
  assign n20158 = ~n18677 & ~n18701;
  assign n20159 = ~n18708 & n20158;
  assign n20160 = ~n18699 & ~n18701;
  assign n20161 = ~n18660 & n20160;
  assign n20162 = ~n18700 & ~n20161;
  assign n20163 = ~n20159 & n20162;
  assign n20164 = pi338 & n4596;
  assign n20165 = n20163 & ~n20164;
  assign n20166 = n4596 & ~n20163;
  assign n20167 = pi338 & n20166;
  assign n20168 = ~n20165 & ~n20167;
  assign n20169 = ~n20157 & n20168;
  assign n20170 = n20157 & ~n20168;
  assign n20171 = ~n20169 & ~n20170;
  assign n20172 = pi340 & n2464;
  assign n20173 = n2091 & ~n18727;
  assign n20174 = pi340 & n20173;
  assign n20175 = n17887 & ~n19370;
  assign n20176 = ~n17887 & ~n19379;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = ~n18718 & n18727;
  assign n20179 = ~n20177 & ~n20178;
  assign n20180 = ~n20174 & ~n20179;
  assign n20181 = n20172 & n20180;
  assign n20182 = ~n20172 & ~n20180;
  assign n20183 = ~n20181 & ~n20182;
  assign n20184 = ~n20171 & ~n20183;
  assign n20185 = n20157 & n20168;
  assign n20186 = ~n20157 & ~n20168;
  assign n20187 = ~n20185 & ~n20186;
  assign n20188 = ~n20172 & n20180;
  assign n20189 = n20172 & ~n20180;
  assign n20190 = ~n20188 & ~n20189;
  assign n20191 = ~n20187 & ~n20190;
  assign n20192 = ~n20184 & ~n20191;
  assign n20193 = ~n20156 & ~n20192;
  assign n20194 = n20149 & ~n20153;
  assign n20195 = ~n20149 & n20153;
  assign n20196 = ~n20194 & ~n20195;
  assign n20197 = ~n20183 & ~n20187;
  assign n20198 = ~n20171 & ~n20190;
  assign n20199 = ~n20197 & ~n20198;
  assign n20200 = ~n20196 & ~n20199;
  assign n20201 = ~n20193 & ~n20200;
  assign n20202 = ~n19400 & n20201;
  assign n20203 = n19400 & ~n20201;
  assign n20204 = ~n20202 & ~n20203;
  assign n20205 = pi343 & n1442;
  assign n20206 = pi342 & n1729;
  assign n20207 = n18751 & ~n18765;
  assign n20208 = ~n18762 & ~n20207;
  assign n20209 = ~n20206 & ~n20208;
  assign n20210 = n1729 & ~n20207;
  assign n20211 = pi342 & n20210;
  assign n20212 = ~n18762 & n20211;
  assign n20213 = ~n20209 & ~n20212;
  assign n20214 = n20205 & ~n20213;
  assign n20215 = ~n20205 & n20213;
  assign n20216 = ~n20214 & ~n20215;
  assign n20217 = ~n20204 & ~n20216;
  assign n20218 = n19400 & n20201;
  assign n20219 = ~n19400 & ~n20201;
  assign n20220 = ~n20218 & ~n20219;
  assign n20221 = ~n20205 & ~n20213;
  assign n20222 = n20205 & n20213;
  assign n20223 = ~n20221 & ~n20222;
  assign n20224 = ~n20220 & ~n20223;
  assign n20225 = ~n20217 & ~n20224;
  assign n20226 = ~n19399 & ~n20225;
  assign n20227 = n19387 & ~n19396;
  assign n20228 = ~n19387 & n19396;
  assign n20229 = ~n20227 & ~n20228;
  assign n20230 = ~n20216 & ~n20220;
  assign n20231 = ~n20204 & ~n20223;
  assign n20232 = ~n20230 & ~n20231;
  assign n20233 = ~n20229 & ~n20232;
  assign n20234 = ~n20226 & ~n20233;
  assign n20235 = n19367 & n20234;
  assign n20236 = ~n19367 & ~n20234;
  assign n20237 = ~n20235 & ~n20236;
  assign n20238 = n17844 & n18781;
  assign n20239 = ~n17844 & ~n18781;
  assign n20240 = ~n1154 & ~n20239;
  assign n20241 = ~n20238 & ~n20240;
  assign n20242 = ~n1256 & ~n20241;
  assign n20243 = pi344 & n20242;
  assign n20244 = ~n1154 & n18781;
  assign n20245 = n1256 & ~n20244;
  assign n20246 = pi344 & ~n20245;
  assign n20247 = n1154 & ~n18781;
  assign n20248 = n17844 & ~n20247;
  assign n20249 = ~n20246 & ~n20248;
  assign n20250 = ~n20243 & ~n20249;
  assign n20251 = ~n1154 & ~n20250;
  assign n20252 = pi345 & n20251;
  assign n20253 = pi345 & ~n1154;
  assign n20254 = ~n20249 & ~n20253;
  assign n20255 = ~n20243 & n20254;
  assign n20256 = ~n20252 & ~n20255;
  assign n20257 = ~n20237 & ~n20256;
  assign n20258 = n19367 & ~n20234;
  assign n20259 = ~n19367 & n20234;
  assign n20260 = ~n20258 & ~n20259;
  assign n20261 = ~n20250 & ~n20253;
  assign n20262 = n20250 & n20253;
  assign n20263 = ~n20261 & ~n20262;
  assign n20264 = ~n20260 & ~n20263;
  assign n20265 = ~n20257 & ~n20264;
  assign n20266 = pi346 & n1156;
  assign n20267 = ~n20265 & ~n20266;
  assign n20268 = pi346 & n20265;
  assign n20269 = n1156 & n20268;
  assign n20270 = ~n20267 & ~n20269;
  assign n20271 = pi282 & ~n20270;
  assign n20272 = ~pi282 & n20270;
  assign n20273 = ~n20271 & ~n20272;
  assign n20274 = ~n19364 & ~n20273;
  assign n20275 = n19364 & n20273;
  assign n20276 = ~n20274 & ~n20275;
  assign n20277 = ~n19358 & ~n20276;
  assign n20278 = ~n19364 & n20273;
  assign n20279 = n19364 & ~n20273;
  assign n20280 = ~n20278 & ~n20279;
  assign n20281 = n19358 & ~n20280;
  assign n20282 = ~n20277 & ~n20281;
  assign n20283 = ~n18809 & ~n18831;
  assign n20284 = n18809 & n18831;
  assign n20285 = n17839 & ~n18815;
  assign n20286 = ~n19336 & ~n20285;
  assign n20287 = ~n20284 & ~n20286;
  assign n20288 = ~n20283 & ~n20287;
  assign n20289 = n20282 & n20288;
  assign n20290 = ~n20282 & ~n20288;
  assign n20291 = ~n20289 & ~n20290;
  assign n20292 = ~n831 & ~n20291;
  assign n20293 = ~n18841 & ~n20292;
  assign n20294 = pi161 & ~n20293;
  assign n20295 = ~n18840 & ~n20294;
  assign po217 = ~pi160 & n20295;
  assign n20297 = pi283 & n831;
  assign n20298 = ~n19340 & ~n19352;
  assign n20299 = ~n19335 & ~n19346;
  assign n20300 = ~n20298 & ~n20299;
  assign n20301 = pi297 & ~n20300;
  assign n20302 = pi128 & n20301;
  assign n20303 = ~pi128 & pi297;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = pi129 & ~n20304;
  assign n20306 = pi297 & ~n20302;
  assign n20307 = n1567 & n20306;
  assign n20308 = ~n20305 & ~n20307;
  assign n20309 = pi301 & n1840;
  assign n20310 = pi305 & n3552;
  assign n20311 = pi309 & n6777;
  assign n20312 = pi313 & n9815;
  assign n20313 = ~n18973 & n18974;
  assign n20314 = n18973 & ~n18974;
  assign n20315 = ~n18975 & ~n20314;
  assign n20316 = ~n17487 & n20315;
  assign n20317 = ~n20313 & ~n20316;
  assign n20318 = pi152 & ~pi153;
  assign n20319 = pi150 & n20318;
  assign n20320 = pi153 & ~n16976;
  assign n20321 = n18925 & n20320;
  assign n20322 = ~n20319 & ~n20321;
  assign n20323 = pi149 & ~n20322;
  assign n20324 = pi153 & n16976;
  assign n20325 = n18915 & n20324;
  assign n20326 = ~pi152 & ~pi153;
  assign n20327 = ~pi150 & n20326;
  assign n20328 = ~n20325 & ~n20327;
  assign n20329 = ~pi149 & ~n20328;
  assign n20330 = ~pi152 & pi153;
  assign n20331 = pi151 & n20330;
  assign n20332 = ~pi153 & ~n16976;
  assign n20333 = pi152 & n20332;
  assign n20334 = ~n20331 & ~n20333;
  assign n20335 = pi150 & ~n20334;
  assign n20336 = pi152 & pi153;
  assign n20337 = ~pi151 & n20336;
  assign n20338 = ~pi153 & n16976;
  assign n20339 = ~pi152 & n20338;
  assign n20340 = ~n20337 & ~n20339;
  assign n20341 = ~pi150 & ~n20340;
  assign n20342 = ~n18919 & ~n18930;
  assign n20343 = ~pi153 & ~n20342;
  assign n20344 = ~n20341 & ~n20343;
  assign n20345 = ~n20335 & n20344;
  assign n20346 = ~n20329 & n20345;
  assign n20347 = ~n20323 & n20346;
  assign n20348 = pi321 & n20347;
  assign n20349 = ~n17462 & n18937;
  assign n20350 = ~n17455 & ~n20349;
  assign n20351 = n16985 & ~n20350;
  assign n20352 = n17455 & ~n18951;
  assign n20353 = ~n20351 & ~n20352;
  assign n20354 = pi321 & ~n20353;
  assign n20355 = n16985 & n18938;
  assign n20356 = ~n20354 & ~n20355;
  assign n20357 = pi320 & ~n20356;
  assign n20358 = n17456 & n20349;
  assign n20359 = ~n20357 & ~n20358;
  assign n20360 = pi320 & n18937;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = n18937 & n20359;
  assign n20363 = pi320 & n20362;
  assign n20364 = ~n20361 & ~n20363;
  assign n20365 = ~n20348 & ~n20364;
  assign n20366 = n20359 & ~n20360;
  assign n20367 = n18937 & ~n20359;
  assign n20368 = pi320 & n20367;
  assign n20369 = ~n20366 & ~n20368;
  assign n20370 = n20347 & ~n20369;
  assign n20371 = pi321 & n20370;
  assign n20372 = ~n20365 & ~n20371;
  assign n20373 = pi319 & n17455;
  assign n20374 = ~n20372 & ~n20373;
  assign n20375 = n17455 & n20372;
  assign n20376 = pi319 & n20375;
  assign n20377 = ~n20374 & ~n20376;
  assign n20378 = n18962 & ~n18963;
  assign n20379 = ~n18962 & n18963;
  assign n20380 = ~n17442 & ~n17478;
  assign n20381 = ~n20379 & ~n20380;
  assign n20382 = ~n17477 & n20381;
  assign n20383 = ~n20378 & ~n20382;
  assign n20384 = n20377 & n20383;
  assign n20385 = ~n20377 & ~n20383;
  assign n20386 = ~n20384 & ~n20385;
  assign n20387 = n16985 & ~n20386;
  assign n20388 = pi318 & n20387;
  assign n20389 = pi318 & n16985;
  assign n20390 = ~n20385 & ~n20389;
  assign n20391 = ~n20384 & n20390;
  assign n20392 = ~n20388 & ~n20391;
  assign n20393 = ~n20317 & ~n20392;
  assign n20394 = n20317 & n20392;
  assign n20395 = ~n20393 & ~n20394;
  assign n20396 = n14618 & ~n20395;
  assign n20397 = pi317 & n20396;
  assign n20398 = pi317 & n14618;
  assign n20399 = ~n20394 & ~n20398;
  assign n20400 = ~n20393 & n20399;
  assign n20401 = ~n20397 & ~n20400;
  assign n20402 = ~n18998 & ~n19002;
  assign n20403 = ~n19003 & ~n20402;
  assign n20404 = pi316 & n14156;
  assign n20405 = ~n20403 & ~n20404;
  assign n20406 = n14156 & n20403;
  assign n20407 = pi316 & n20406;
  assign n20408 = ~n20405 & ~n20407;
  assign n20409 = ~n20401 & ~n20408;
  assign n20410 = n20403 & ~n20404;
  assign n20411 = n14156 & ~n20403;
  assign n20412 = pi316 & n20411;
  assign n20413 = ~n20410 & ~n20412;
  assign n20414 = ~n20400 & ~n20413;
  assign n20415 = ~n20397 & n20414;
  assign n20416 = ~n20409 & ~n20415;
  assign n20417 = ~n18990 & ~n18995;
  assign n20418 = ~n17502 & n20417;
  assign n20419 = n18990 & ~n18998;
  assign n20420 = ~n20418 & ~n20419;
  assign n20421 = ~n18912 & ~n20420;
  assign n20422 = n18990 & ~n18995;
  assign n20423 = ~n17502 & n20422;
  assign n20424 = ~n18990 & ~n18998;
  assign n20425 = ~n20423 & ~n20424;
  assign n20426 = n14156 & ~n20425;
  assign n20427 = pi317 & n20426;
  assign n20428 = ~n20421 & ~n20427;
  assign n20429 = ~n17532 & ~n20428;
  assign n20430 = ~n18910 & n20429;
  assign n20431 = ~n11998 & n20428;
  assign n20432 = ~n19036 & ~n20431;
  assign n20433 = n10908 & n20432;
  assign n20434 = ~n18911 & n20428;
  assign n20435 = n11998 & ~n20434;
  assign n20436 = ~n20433 & ~n20435;
  assign n20437 = pi316 & ~n20436;
  assign n20438 = ~n20430 & ~n20437;
  assign n20439 = n20416 & n20438;
  assign n20440 = ~n20416 & ~n20438;
  assign n20441 = ~n20439 & ~n20440;
  assign n20442 = n11998 & ~n20441;
  assign n20443 = pi315 & n20442;
  assign n20444 = pi315 & n11998;
  assign n20445 = ~n20416 & n20438;
  assign n20446 = n20416 & ~n20438;
  assign n20447 = ~n20445 & ~n20446;
  assign n20448 = ~n20444 & ~n20447;
  assign n20449 = ~n20443 & ~n20448;
  assign n20450 = pi315 & n10908;
  assign n20451 = ~n19051 & n20450;
  assign n20452 = ~n17512 & ~n18911;
  assign n20453 = ~n19036 & ~n20452;
  assign n20454 = ~n19010 & ~n20453;
  assign n20455 = ~n19040 & ~n20454;
  assign n20456 = n19051 & ~n20450;
  assign n20457 = ~n20455 & ~n20456;
  assign n20458 = ~n20451 & ~n20457;
  assign n20459 = n20449 & n20458;
  assign n20460 = ~n20449 & ~n20458;
  assign n20461 = ~n20459 & ~n20460;
  assign n20462 = pi314 & n10908;
  assign n20463 = ~n19062 & ~n20462;
  assign n20464 = ~n19056 & n20463;
  assign n20465 = ~n19056 & ~n19062;
  assign n20466 = n20462 & ~n20465;
  assign n20467 = ~n20464 & ~n20466;
  assign n20468 = ~n20461 & ~n20467;
  assign n20469 = n20449 & ~n20458;
  assign n20470 = ~n20449 & n20458;
  assign n20471 = ~n20469 & ~n20470;
  assign n20472 = ~n19062 & n20462;
  assign n20473 = ~n19056 & n20472;
  assign n20474 = ~n20462 & ~n20465;
  assign n20475 = ~n20473 & ~n20474;
  assign n20476 = ~n20471 & ~n20475;
  assign n20477 = ~n20468 & ~n20476;
  assign n20478 = ~n20312 & n20477;
  assign n20479 = n20312 & ~n20477;
  assign n20480 = ~n20478 & ~n20479;
  assign n20481 = pi312 & n9517;
  assign n20482 = n17119 & ~n17590;
  assign n20483 = n7044 & ~n19088;
  assign n20484 = pi313 & n20483;
  assign n20485 = ~n20482 & ~n20484;
  assign n20486 = ~n17579 & ~n20485;
  assign n20487 = n17119 & n20483;
  assign n20488 = ~n19089 & ~n20487;
  assign n20489 = pi313 & ~n20488;
  assign n20490 = ~n20486 & ~n20489;
  assign n20491 = n19064 & ~n20490;
  assign n20492 = ~n19064 & n20490;
  assign n20493 = n18894 & ~n20492;
  assign n20494 = ~n20491 & ~n20493;
  assign n20495 = n20481 & ~n20494;
  assign n20496 = ~n18894 & ~n20491;
  assign n20497 = ~n20492 & ~n20496;
  assign n20498 = ~n20481 & ~n20497;
  assign n20499 = ~n20495 & ~n20498;
  assign n20500 = ~n20480 & ~n20499;
  assign n20501 = ~n20312 & ~n20477;
  assign n20502 = n20312 & n20477;
  assign n20503 = ~n20501 & ~n20502;
  assign n20504 = ~n20481 & ~n20494;
  assign n20505 = n20481 & ~n20497;
  assign n20506 = ~n20504 & ~n20505;
  assign n20507 = ~n20503 & ~n20506;
  assign n20508 = ~n20500 & ~n20507;
  assign n20509 = n19068 & ~n19109;
  assign n20510 = ~n19068 & n19109;
  assign n20511 = ~n19100 & ~n20510;
  assign n20512 = ~n20509 & ~n20511;
  assign n20513 = n20508 & n20512;
  assign n20514 = ~n20508 & ~n20512;
  assign n20515 = ~n20513 & ~n20514;
  assign n20516 = pi311 & n7874;
  assign n20517 = n19120 & ~n19121;
  assign n20518 = ~n19122 & ~n20517;
  assign n20519 = n20516 & ~n20518;
  assign n20520 = ~n19120 & ~n19122;
  assign n20521 = ~n19121 & ~n20520;
  assign n20522 = ~n20516 & ~n20521;
  assign n20523 = ~n20519 & ~n20522;
  assign n20524 = ~n20515 & ~n20523;
  assign n20525 = n20508 & ~n20512;
  assign n20526 = ~n20508 & n20512;
  assign n20527 = ~n20525 & ~n20526;
  assign n20528 = ~n20516 & ~n20518;
  assign n20529 = n20516 & ~n20521;
  assign n20530 = ~n20528 & ~n20529;
  assign n20531 = ~n20527 & ~n20530;
  assign n20532 = ~n20524 & ~n20531;
  assign n20533 = ~pi310 & n20532;
  assign n20534 = ~n7044 & n20532;
  assign n20535 = n7044 & ~n20532;
  assign n20536 = pi310 & n20535;
  assign n20537 = ~n20534 & ~n20536;
  assign n20538 = ~n6777 & ~n20537;
  assign n20539 = ~n20533 & ~n20538;
  assign n20540 = ~n19134 & ~n20539;
  assign n20541 = ~n19133 & n20532;
  assign n20542 = n19125 & n20541;
  assign n20543 = n19133 & ~n20532;
  assign n20544 = ~n19125 & n20543;
  assign n20545 = ~n20542 & ~n20544;
  assign n20546 = pi310 & ~n20545;
  assign n20547 = ~n19142 & n20532;
  assign n20548 = n6777 & n20547;
  assign n20549 = ~n20546 & ~n20548;
  assign n20550 = n7044 & ~n20549;
  assign n20551 = ~n19133 & ~n20532;
  assign n20552 = ~pi310 & n19125;
  assign n20553 = n20551 & n20552;
  assign n20554 = n19133 & n20532;
  assign n20555 = ~n19125 & n20554;
  assign n20556 = n6777 & ~n19135;
  assign n20557 = pi310 & n20556;
  assign n20558 = ~n19134 & ~n20557;
  assign n20559 = ~n20532 & ~n20558;
  assign n20560 = ~n20555 & ~n20559;
  assign n20561 = ~n7044 & ~n20560;
  assign n20562 = ~n20553 & ~n20561;
  assign n20563 = ~n20550 & n20562;
  assign n20564 = ~n20540 & n20563;
  assign n20565 = ~n20311 & ~n20564;
  assign n20566 = n20311 & n20564;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = pi308 & n5463;
  assign n20569 = n4086 & ~n19155;
  assign n20570 = pi309 & n20569;
  assign n20571 = ~n17202 & ~n17678;
  assign n20572 = ~n20570 & ~n20571;
  assign n20573 = ~n17667 & ~n20572;
  assign n20574 = n4772 & ~n17653;
  assign n20575 = ~n17202 & n20569;
  assign n20576 = ~n20574 & ~n20575;
  assign n20577 = pi309 & ~n20576;
  assign n20578 = ~n20573 & ~n20577;
  assign n20579 = ~n19144 & ~n20578;
  assign n20580 = n19144 & n20578;
  assign n20581 = n18882 & ~n20580;
  assign n20582 = ~n20579 & ~n20581;
  assign n20583 = n20568 & ~n20582;
  assign n20584 = ~n18882 & ~n20579;
  assign n20585 = ~n20580 & ~n20584;
  assign n20586 = ~n20568 & ~n20585;
  assign n20587 = ~n20583 & ~n20586;
  assign n20588 = ~n20567 & ~n20587;
  assign n20589 = ~n20311 & n20564;
  assign n20590 = n20311 & ~n20564;
  assign n20591 = ~n20589 & ~n20590;
  assign n20592 = ~n20568 & ~n20582;
  assign n20593 = n20568 & ~n20585;
  assign n20594 = ~n20592 & ~n20593;
  assign n20595 = ~n20591 & ~n20594;
  assign n20596 = ~n20588 & ~n20595;
  assign n20597 = ~n19147 & ~n19148;
  assign n20598 = n19147 & n19148;
  assign n20599 = ~n19183 & ~n20598;
  assign n20600 = ~n20597 & ~n20599;
  assign n20601 = n20596 & n20600;
  assign n20602 = ~n20596 & ~n20600;
  assign n20603 = ~n20601 & ~n20602;
  assign n20604 = pi307 & n4772;
  assign n20605 = ~n19195 & n19200;
  assign n20606 = ~n19196 & ~n20605;
  assign n20607 = n20604 & ~n20606;
  assign n20608 = ~n19196 & ~n19200;
  assign n20609 = ~n19195 & ~n20608;
  assign n20610 = ~n20604 & ~n20609;
  assign n20611 = ~n20607 & ~n20610;
  assign n20612 = ~n20603 & ~n20611;
  assign n20613 = n20596 & ~n20600;
  assign n20614 = ~n20596 & n20600;
  assign n20615 = ~n20613 & ~n20614;
  assign n20616 = ~n20604 & ~n20606;
  assign n20617 = n20604 & ~n20609;
  assign n20618 = ~n20616 & ~n20617;
  assign n20619 = ~n20615 & ~n20618;
  assign n20620 = ~n20612 & ~n20619;
  assign n20621 = ~pi306 & n20620;
  assign n20622 = ~n4086 & n20620;
  assign n20623 = n4086 & ~n20620;
  assign n20624 = pi306 & n20623;
  assign n20625 = ~n20622 & ~n20624;
  assign n20626 = ~n3552 & ~n20625;
  assign n20627 = ~n20621 & ~n20626;
  assign n20628 = ~n19218 & ~n20627;
  assign n20629 = ~n19210 & n20620;
  assign n20630 = ~n19205 & n20629;
  assign n20631 = n19210 & ~n20620;
  assign n20632 = n19205 & n20631;
  assign n20633 = ~n20630 & ~n20632;
  assign n20634 = pi306 & ~n20633;
  assign n20635 = ~n19213 & n20620;
  assign n20636 = n3552 & n20635;
  assign n20637 = ~n20634 & ~n20636;
  assign n20638 = n4086 & ~n20637;
  assign n20639 = ~pi306 & ~n19205;
  assign n20640 = ~n19210 & ~n20620;
  assign n20641 = n20639 & n20640;
  assign n20642 = n19210 & n20620;
  assign n20643 = n19205 & n20642;
  assign n20644 = n3552 & ~n19217;
  assign n20645 = pi306 & n20644;
  assign n20646 = ~n19218 & ~n20645;
  assign n20647 = ~n20620 & ~n20646;
  assign n20648 = ~n20643 & ~n20647;
  assign n20649 = ~n4086 & ~n20648;
  assign n20650 = ~n20641 & ~n20649;
  assign n20651 = ~n20638 & n20650;
  assign n20652 = ~n20628 & n20651;
  assign n20653 = ~n20310 & n20652;
  assign n20654 = n20310 & ~n20652;
  assign n20655 = ~n20653 & ~n20654;
  assign n20656 = pi304 & n3012;
  assign n20657 = n17273 & ~n17737;
  assign n20658 = n2183 & ~n19232;
  assign n20659 = pi305 & n20658;
  assign n20660 = ~n20657 & ~n20659;
  assign n20661 = ~n17726 & ~n20660;
  assign n20662 = n2574 & n17712;
  assign n20663 = n17273 & n20658;
  assign n20664 = ~n20662 & ~n20663;
  assign n20665 = pi305 & ~n20664;
  assign n20666 = ~n20661 & ~n20665;
  assign n20667 = n19221 & ~n20666;
  assign n20668 = ~n19221 & n20666;
  assign n20669 = n18868 & ~n20668;
  assign n20670 = ~n20667 & ~n20669;
  assign n20671 = n20656 & ~n20670;
  assign n20672 = ~n18868 & ~n20667;
  assign n20673 = ~n20668 & ~n20672;
  assign n20674 = ~n20656 & ~n20673;
  assign n20675 = ~n20671 & ~n20674;
  assign n20676 = ~n20655 & ~n20675;
  assign n20677 = ~n20310 & ~n20652;
  assign n20678 = n20310 & n20652;
  assign n20679 = ~n20677 & ~n20678;
  assign n20680 = ~n20656 & ~n20670;
  assign n20681 = n20656 & ~n20673;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20679 & ~n20682;
  assign n20684 = ~n20676 & ~n20683;
  assign n20685 = ~n19225 & ~n19266;
  assign n20686 = n19225 & n19266;
  assign n20687 = ~n19260 & ~n20686;
  assign n20688 = ~n20685 & ~n20687;
  assign n20689 = n20684 & ~n20688;
  assign n20690 = ~n20684 & n20688;
  assign n20691 = ~n20689 & ~n20690;
  assign n20692 = pi303 & n2574;
  assign n20693 = n19277 & ~n19279;
  assign n20694 = ~n19278 & ~n20693;
  assign n20695 = n20692 & ~n20694;
  assign n20696 = ~n19277 & ~n19278;
  assign n20697 = ~n19279 & ~n20696;
  assign n20698 = ~n20692 & ~n20697;
  assign n20699 = ~n20695 & ~n20698;
  assign n20700 = ~n20691 & ~n20699;
  assign n20701 = n20684 & n20688;
  assign n20702 = ~n20684 & ~n20688;
  assign n20703 = ~n20701 & ~n20702;
  assign n20704 = ~n20692 & ~n20694;
  assign n20705 = n20692 & ~n20697;
  assign n20706 = ~n20704 & ~n20705;
  assign n20707 = ~n20703 & ~n20706;
  assign n20708 = ~n20700 & ~n20707;
  assign n20709 = ~pi302 & ~n20708;
  assign n20710 = ~n2183 & ~n20708;
  assign n20711 = n2183 & n20708;
  assign n20712 = pi302 & n20711;
  assign n20713 = ~n20710 & ~n20712;
  assign n20714 = ~n1840 & ~n20713;
  assign n20715 = ~n20709 & ~n20714;
  assign n20716 = ~n19294 & ~n20715;
  assign n20717 = ~n19290 & ~n20708;
  assign n20718 = n1840 & n20717;
  assign n20719 = ~n19287 & n20708;
  assign n20720 = ~n19282 & n20719;
  assign n20721 = n19287 & ~n20708;
  assign n20722 = n19282 & n20721;
  assign n20723 = ~n20720 & ~n20722;
  assign n20724 = pi302 & ~n20723;
  assign n20725 = ~n20718 & ~n20724;
  assign n20726 = n2183 & ~n20725;
  assign n20727 = ~n19287 & ~n20708;
  assign n20728 = ~n19282 & n20727;
  assign n20729 = n1840 & ~n19295;
  assign n20730 = pi302 & n20729;
  assign n20731 = ~n19294 & ~n20730;
  assign n20732 = n20708 & ~n20731;
  assign n20733 = ~n20728 & ~n20732;
  assign n20734 = ~n2183 & ~n20733;
  assign n20735 = n19287 & n20708;
  assign n20736 = ~pi302 & n19282;
  assign n20737 = n20735 & n20736;
  assign n20738 = ~n20734 & ~n20737;
  assign n20739 = ~n20726 & n20738;
  assign n20740 = ~n20716 & n20739;
  assign n20741 = ~n20309 & n20740;
  assign n20742 = n20309 & ~n20740;
  assign n20743 = ~n20741 & ~n20742;
  assign n20744 = pi300 & n1533;
  assign n20745 = ~n18852 & n19298;
  assign n20746 = n18852 & ~n19298;
  assign n20747 = n18850 & ~n20746;
  assign n20748 = ~n20745 & ~n20747;
  assign n20749 = n20744 & ~n20748;
  assign n20750 = ~n18850 & ~n20745;
  assign n20751 = ~n20746 & ~n20750;
  assign n20752 = ~n20744 & ~n20751;
  assign n20753 = ~n20749 & ~n20752;
  assign n20754 = ~n20743 & ~n20753;
  assign n20755 = ~n20309 & ~n20740;
  assign n20756 = n20309 & n20740;
  assign n20757 = ~n20755 & ~n20756;
  assign n20758 = ~n20744 & ~n20748;
  assign n20759 = n20744 & ~n20751;
  assign n20760 = ~n20758 & ~n20759;
  assign n20761 = ~n20757 & ~n20760;
  assign n20762 = ~n20754 & ~n20761;
  assign n20763 = n19302 & ~n19327;
  assign n20764 = ~n19302 & n19327;
  assign n20765 = ~n19318 & ~n20764;
  assign n20766 = ~n20763 & ~n20765;
  assign n20767 = ~n20762 & ~n20766;
  assign n20768 = n20762 & n20766;
  assign n20769 = ~n20767 & ~n20768;
  assign n20770 = ~n17839 & n19337;
  assign n20771 = n18815 & n20770;
  assign n20772 = ~n19338 & ~n19352;
  assign n20773 = ~n20771 & ~n20772;
  assign n20774 = n20769 & ~n20773;
  assign n20775 = ~n20769 & n20773;
  assign n20776 = ~n20774 & ~n20775;
  assign n20777 = ~n1515 & ~n19332;
  assign n20778 = n1515 & n19332;
  assign n20779 = n18847 & ~n20778;
  assign n20780 = ~n20777 & ~n20779;
  assign n20781 = n1553 & ~n20780;
  assign n20782 = n18847 & ~n19332;
  assign n20783 = ~n1553 & ~n20782;
  assign n20784 = n1515 & n20783;
  assign n20785 = ~n20781 & ~n20784;
  assign n20786 = pi299 & ~n20785;
  assign n20787 = pi299 & n1553;
  assign n20788 = n19332 & ~n20787;
  assign n20789 = ~n18847 & n20788;
  assign n20790 = ~n20786 & ~n20789;
  assign n20791 = pi298 & n1515;
  assign n20792 = n20790 & ~n20791;
  assign n20793 = n1515 & ~n20790;
  assign n20794 = pi298 & n20793;
  assign n20795 = ~n20792 & ~n20794;
  assign n20796 = ~n20776 & ~n20795;
  assign n20797 = ~n20769 & ~n20773;
  assign n20798 = n20769 & n20773;
  assign n20799 = ~n20797 & ~n20798;
  assign n20800 = ~n20790 & ~n20791;
  assign n20801 = n1515 & n20790;
  assign n20802 = pi298 & n20801;
  assign n20803 = ~n20800 & ~n20802;
  assign n20804 = ~n20799 & ~n20803;
  assign n20805 = ~n20796 & ~n20804;
  assign n20806 = n20308 & n20805;
  assign n20807 = ~n20308 & ~n20805;
  assign n20808 = ~n20806 & ~n20807;
  assign n20809 = pi296 & ~n20808;
  assign n20810 = pi128 & n20809;
  assign n20811 = pi128 & pi296;
  assign n20812 = ~n20807 & ~n20811;
  assign n20813 = ~n20806 & n20812;
  assign n20814 = ~n20810 & ~n20813;
  assign n20815 = ~n19364 & ~n20270;
  assign n20816 = n19364 & n20270;
  assign n20817 = ~pi282 & ~n20816;
  assign n20818 = ~n20815 & ~n20817;
  assign n20819 = n1154 & ~n20265;
  assign n20820 = n1156 & n20819;
  assign n20821 = n1156 & ~n20265;
  assign n20822 = ~n1154 & ~n20821;
  assign n20823 = ~n20820 & ~n20822;
  assign n20824 = pi346 & ~n20823;
  assign n20825 = n19387 & n19400;
  assign n20826 = ~n19387 & ~n19400;
  assign n20827 = n20201 & ~n20826;
  assign n20828 = ~n20825 & ~n20827;
  assign n20829 = ~n19387 & n20201;
  assign n20830 = n19387 & ~n20201;
  assign n20831 = ~n20829 & ~n20830;
  assign n20832 = n19400 & ~n20213;
  assign n20833 = ~n19400 & n20213;
  assign n20834 = ~n20832 & ~n20833;
  assign n20835 = n19396 & ~n20205;
  assign n20836 = ~n20834 & ~n20835;
  assign n20837 = ~n20831 & n20836;
  assign n20838 = ~n19396 & n20205;
  assign n20839 = ~n19387 & ~n20201;
  assign n20840 = n19387 & n20201;
  assign n20841 = ~n20839 & ~n20840;
  assign n20842 = ~n19400 & ~n20213;
  assign n20843 = n19400 & n20213;
  assign n20844 = ~n20842 & ~n20843;
  assign n20845 = ~n20835 & ~n20844;
  assign n20846 = ~n20841 & n20845;
  assign n20847 = ~n20838 & ~n20846;
  assign n20848 = ~n20837 & n20847;
  assign n20849 = ~n20828 & n20848;
  assign n20850 = n20828 & ~n20848;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = pi341 & n2464;
  assign n20853 = n19420 & n20086;
  assign n20854 = ~n20082 & ~n20107;
  assign n20855 = n20082 & n20107;
  assign n20856 = ~n20854 & ~n20855;
  assign n20857 = n6556 & ~n20856;
  assign n20858 = pi333 & n20857;
  assign n20859 = ~n20082 & n20107;
  assign n20860 = n20082 & ~n20107;
  assign n20861 = ~n20859 & ~n20860;
  assign n20862 = ~n20071 & ~n20861;
  assign n20863 = ~n20858 & ~n20862;
  assign n20864 = ~n20070 & ~n20863;
  assign n20865 = n6556 & ~n20861;
  assign n20866 = pi333 & n20865;
  assign n20867 = ~n20071 & ~n20856;
  assign n20868 = ~n20866 & ~n20867;
  assign n20869 = ~n20123 & ~n20868;
  assign n20870 = ~n20864 & ~n20869;
  assign n20871 = ~n19420 & ~n20086;
  assign n20872 = n20870 & ~n20871;
  assign n20873 = ~n20853 & ~n20872;
  assign n20874 = ~n19420 & n20128;
  assign n20875 = n19420 & ~n20128;
  assign n20876 = ~n20874 & ~n20875;
  assign n20877 = ~n19446 & ~n20876;
  assign n20878 = n19420 & n20128;
  assign n20879 = ~n19420 & ~n20128;
  assign n20880 = ~n20878 & ~n20879;
  assign n20881 = n19446 & ~n20880;
  assign n20882 = ~n20877 & ~n20881;
  assign n20883 = n19427 & ~n20134;
  assign n20884 = ~n20882 & ~n20883;
  assign n20885 = n5257 & ~n19427;
  assign n20886 = pi337 & n20885;
  assign n20887 = ~n20884 & ~n20886;
  assign n20888 = ~n20873 & n20887;
  assign n20889 = n20873 & ~n20887;
  assign n20890 = ~n20888 & ~n20889;
  assign n20891 = pi335 & n5973;
  assign n20892 = n19503 & ~n20016;
  assign n20893 = ~n19503 & n20016;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = ~n19510 & ~n20021;
  assign n20896 = n19510 & n20021;
  assign n20897 = ~n20895 & ~n20896;
  assign n20898 = ~n20894 & ~n20897;
  assign n20899 = ~n19503 & ~n20016;
  assign n20900 = n19503 & n20016;
  assign n20901 = ~n20899 & ~n20900;
  assign n20902 = n11711 & ~n19510;
  assign n20903 = pi328 & n20902;
  assign n20904 = n12917 & ~n20021;
  assign n20905 = pi327 & n20904;
  assign n20906 = ~n20903 & ~n20905;
  assign n20907 = ~n20901 & ~n20906;
  assign n20908 = ~n20898 & ~n20907;
  assign n20909 = ~n19506 & n20908;
  assign n20910 = n19506 & ~n20908;
  assign n20911 = ~n20909 & ~n20910;
  assign n20912 = ~n19460 & ~n20020;
  assign n20913 = ~n20911 & ~n20912;
  assign n20914 = n19460 & n20020;
  assign n20915 = ~n20913 & ~n20914;
  assign n20916 = n19460 & ~n20042;
  assign n20917 = ~n19460 & n20042;
  assign n20918 = ~n20916 & ~n20917;
  assign n20919 = ~n19483 & ~n20918;
  assign n20920 = n19460 & n20042;
  assign n20921 = ~n19460 & ~n20042;
  assign n20922 = ~n20920 & ~n20921;
  assign n20923 = n19483 & ~n20922;
  assign n20924 = ~n20919 & ~n20923;
  assign n20925 = n19467 & ~n20048;
  assign n20926 = ~n20924 & ~n20925;
  assign n20927 = n10561 & ~n19467;
  assign n20928 = pi331 & n20927;
  assign n20929 = ~n20926 & ~n20928;
  assign n20930 = ~n20915 & n20929;
  assign n20931 = n20915 & ~n20929;
  assign n20932 = ~n20930 & ~n20931;
  assign n20933 = pi329 & n11711;
  assign n20934 = n19503 & n19510;
  assign n20935 = ~n19503 & ~n19510;
  assign n20936 = n20016 & ~n20935;
  assign n20937 = ~n20934 & ~n20936;
  assign n20938 = ~n19506 & n20021;
  assign n20939 = n19510 & ~n20901;
  assign n20940 = ~n19510 & ~n20894;
  assign n20941 = ~n20939 & ~n20940;
  assign n20942 = n19506 & ~n20021;
  assign n20943 = ~n20941 & ~n20942;
  assign n20944 = ~n20938 & ~n20943;
  assign n20945 = ~n20937 & ~n20944;
  assign n20946 = n20937 & n20944;
  assign n20947 = ~n20945 & ~n20946;
  assign n20948 = n19540 & ~n19990;
  assign n20949 = ~n19542 & ~n19971;
  assign n20950 = n19542 & n19970;
  assign n20951 = pi322 & n20950;
  assign n20952 = ~n20949 & ~n20951;
  assign n20953 = ~n19558 & ~n20952;
  assign n20954 = n19542 & ~n19971;
  assign n20955 = ~n19542 & n19970;
  assign n20956 = pi322 & n20955;
  assign n20957 = ~n20954 & ~n20956;
  assign n20958 = n19557 & ~n20957;
  assign n20959 = pi323 & n20958;
  assign n20960 = ~n20953 & ~n20959;
  assign n20961 = ~n19540 & n19990;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = ~n20948 & ~n20962;
  assign n20964 = ~n19529 & n19995;
  assign n20965 = n19529 & ~n19995;
  assign n20966 = ~n19993 & ~n20965;
  assign n20967 = ~n20964 & ~n20966;
  assign n20968 = ~n20963 & n20967;
  assign n20969 = n20963 & ~n20967;
  assign n20970 = ~n20968 & ~n20969;
  assign n20971 = pi324 & n19557;
  assign n20972 = pi323 & n19970;
  assign n20973 = ~n19542 & n19557;
  assign n20974 = pi323 & n20973;
  assign n20975 = n19542 & ~n19558;
  assign n20976 = n19970 & ~n20975;
  assign n20977 = pi322 & n20976;
  assign n20978 = ~n20974 & ~n20977;
  assign n20979 = n19936 & n19944;
  assign n20980 = ~n19936 & ~n19944;
  assign n20981 = pi259 & ~n20980;
  assign n20982 = ~n20979 & ~n20981;
  assign n20983 = ~pi260 & ~n20982;
  assign n20984 = ~pi259 & ~n19936;
  assign n20985 = pi259 & n19936;
  assign n20986 = ~n19944 & ~n20985;
  assign n20987 = ~n20984 & ~n20986;
  assign n20988 = pi260 & ~n20987;
  assign n20989 = ~n20983 & ~n20988;
  assign n20990 = pi151 & ~n20989;
  assign n20991 = pi131 & pi280;
  assign n20992 = ~n19594 & n19595;
  assign n20993 = pi129 & pi282;
  assign n20994 = pi283 & ~n20993;
  assign n20995 = pi128 & n20994;
  assign n20996 = pi128 & pi283;
  assign n20997 = pi282 & ~n20996;
  assign n20998 = pi129 & n20997;
  assign n20999 = ~n20995 & ~n20998;
  assign n21000 = ~pi281 & ~n20999;
  assign n21001 = ~pi130 & ~n20999;
  assign n21002 = pi281 & n20999;
  assign n21003 = pi130 & n21002;
  assign n21004 = ~n21001 & ~n21003;
  assign n21005 = ~pi129 & ~n21004;
  assign n21006 = ~n21000 & ~n21005;
  assign n21007 = ~n20992 & ~n21006;
  assign n21008 = n19594 & n19595;
  assign n21009 = ~n19594 & ~n19595;
  assign n21010 = ~n21008 & ~n21009;
  assign n21011 = pi129 & ~n21010;
  assign n21012 = pi281 & n20992;
  assign n21013 = ~n21011 & ~n21012;
  assign n21014 = ~n20999 & ~n21013;
  assign n21015 = pi281 & n19594;
  assign n21016 = ~n19595 & n20999;
  assign n21017 = n21015 & n21016;
  assign n21018 = ~n21014 & ~n21017;
  assign n21019 = pi130 & ~n21018;
  assign n21020 = ~n19595 & ~n20999;
  assign n21021 = n19594 & n21020;
  assign n21022 = n19594 & ~n19595;
  assign n21023 = pi281 & ~n21022;
  assign n21024 = pi129 & n21023;
  assign n21025 = ~n20992 & ~n21024;
  assign n21026 = n20999 & ~n21025;
  assign n21027 = ~n21021 & ~n21026;
  assign n21028 = ~pi130 & ~n21027;
  assign n21029 = n19595 & n20999;
  assign n21030 = ~pi281 & ~n19594;
  assign n21031 = n21029 & n21030;
  assign n21032 = ~n21028 & ~n21031;
  assign n21033 = ~n21019 & n21032;
  assign n21034 = ~n21007 & n21033;
  assign n21035 = ~n19606 & ~n19613;
  assign n21036 = ~n19609 & ~n21035;
  assign n21037 = ~n21034 & ~n21036;
  assign n21038 = n21034 & ~n21035;
  assign n21039 = ~n19609 & n21038;
  assign n21040 = ~n21037 & ~n21039;
  assign n21041 = n20991 & ~n21040;
  assign n21042 = n21034 & ~n21036;
  assign n21043 = ~n21034 & ~n21035;
  assign n21044 = ~n19609 & n21043;
  assign n21045 = ~n21042 & ~n21044;
  assign n21046 = ~n20991 & ~n21045;
  assign n21047 = ~n19621 & ~n19624;
  assign n21048 = ~n19618 & ~n21047;
  assign n21049 = ~n21046 & n21048;
  assign n21050 = ~n21041 & n21049;
  assign n21051 = ~n21041 & ~n21046;
  assign n21052 = ~n21048 & ~n21051;
  assign n21053 = ~n21050 & ~n21052;
  assign n21054 = pi279 & ~n21053;
  assign n21055 = pi132 & n21054;
  assign n21056 = pi132 & pi279;
  assign n21057 = ~n21050 & ~n21056;
  assign n21058 = ~n21052 & n21057;
  assign n21059 = ~n21055 & ~n21058;
  assign n21060 = n19628 & ~n19638;
  assign n21061 = ~n19628 & n19638;
  assign n21062 = ~n19629 & ~n21061;
  assign n21063 = ~n18076 & n21062;
  assign n21064 = ~n21060 & ~n21063;
  assign n21065 = pi133 & pi278;
  assign n21066 = ~n21064 & ~n21065;
  assign n21067 = pi278 & n21064;
  assign n21068 = pi133 & n21067;
  assign n21069 = ~n21066 & ~n21068;
  assign n21070 = ~n21059 & ~n21069;
  assign n21071 = n21064 & ~n21065;
  assign n21072 = pi278 & ~n21064;
  assign n21073 = pi133 & n21072;
  assign n21074 = ~n21071 & ~n21073;
  assign n21075 = ~n21058 & ~n21074;
  assign n21076 = ~n21055 & n21075;
  assign n21077 = ~n21070 & ~n21076;
  assign n21078 = ~n19656 & ~n19660;
  assign n21079 = ~n19661 & ~n21078;
  assign n21080 = n21077 & n21079;
  assign n21081 = ~n21077 & ~n21079;
  assign n21082 = ~n21080 & ~n21081;
  assign n21083 = pi134 & pi277;
  assign n21084 = n19644 & ~n19653;
  assign n21085 = ~n19649 & n21084;
  assign n21086 = ~n19644 & ~n19656;
  assign n21087 = ~n21085 & ~n21086;
  assign n21088 = ~n19589 & ~n21087;
  assign n21089 = ~n19644 & ~n19653;
  assign n21090 = ~n19649 & n21089;
  assign n21091 = n19644 & ~n19656;
  assign n21092 = ~n21090 & ~n21091;
  assign n21093 = pi277 & ~n21092;
  assign n21094 = pi133 & n21093;
  assign n21095 = ~n21088 & ~n21094;
  assign n21096 = ~n19672 & ~n21095;
  assign n21097 = n19672 & n21095;
  assign n21098 = n19650 & ~n21097;
  assign n21099 = ~n21096 & ~n21098;
  assign n21100 = n21083 & ~n21099;
  assign n21101 = ~n19650 & ~n21096;
  assign n21102 = ~n21097 & ~n21101;
  assign n21103 = ~n21083 & ~n21102;
  assign n21104 = ~n21100 & ~n21103;
  assign n21105 = ~n21082 & ~n21104;
  assign n21106 = n21077 & ~n21079;
  assign n21107 = ~n21077 & n21079;
  assign n21108 = ~n21106 & ~n21107;
  assign n21109 = ~n21083 & ~n21099;
  assign n21110 = n21083 & ~n21102;
  assign n21111 = ~n21109 & ~n21110;
  assign n21112 = ~n21108 & ~n21111;
  assign n21113 = ~n21105 & ~n21112;
  assign n21114 = ~n19675 & ~n19676;
  assign n21115 = n19675 & n19676;
  assign n21116 = ~n19681 & ~n21115;
  assign n21117 = ~n21114 & ~n21116;
  assign n21118 = ~n21113 & n21117;
  assign n21119 = n21113 & ~n21117;
  assign n21120 = ~n21118 & ~n21119;
  assign n21121 = pi136 & pi275;
  assign n21122 = pi135 & pi276;
  assign n21123 = n21121 & n21122;
  assign n21124 = ~n21121 & ~n21122;
  assign n21125 = ~n21123 & ~n21124;
  assign n21126 = ~n21120 & ~n21125;
  assign n21127 = n21113 & n21117;
  assign n21128 = ~n21113 & ~n21117;
  assign n21129 = ~n21127 & ~n21128;
  assign n21130 = pi275 & ~n21122;
  assign n21131 = pi136 & n21130;
  assign n21132 = pi276 & ~n21121;
  assign n21133 = pi135 & n21132;
  assign n21134 = ~n21131 & ~n21133;
  assign n21135 = ~n21129 & ~n21134;
  assign n21136 = ~n21126 & ~n21135;
  assign n21137 = ~n19708 & ~n19712;
  assign n21138 = ~n19713 & ~n21137;
  assign n21139 = n21136 & n21138;
  assign n21140 = ~n21136 & ~n21138;
  assign n21141 = ~n21139 & ~n21140;
  assign n21142 = pi137 & pi274;
  assign n21143 = n19692 & ~n19705;
  assign n21144 = ~n19701 & n21143;
  assign n21145 = ~n19692 & ~n19708;
  assign n21146 = ~n21144 & ~n21145;
  assign n21147 = ~n19588 & ~n21146;
  assign n21148 = ~n19692 & ~n19705;
  assign n21149 = ~n19701 & n21148;
  assign n21150 = n19692 & ~n19708;
  assign n21151 = ~n21149 & ~n21150;
  assign n21152 = pi274 & ~n21151;
  assign n21153 = pi136 & n21152;
  assign n21154 = ~n21147 & ~n21153;
  assign n21155 = ~n19724 & ~n21154;
  assign n21156 = n19724 & n21154;
  assign n21157 = n19702 & ~n21156;
  assign n21158 = ~n21155 & ~n21157;
  assign n21159 = n21142 & ~n21158;
  assign n21160 = ~n19702 & ~n21155;
  assign n21161 = ~n21156 & ~n21160;
  assign n21162 = ~n21142 & ~n21161;
  assign n21163 = ~n21159 & ~n21162;
  assign n21164 = ~n21141 & ~n21163;
  assign n21165 = n21136 & ~n21138;
  assign n21166 = ~n21136 & n21138;
  assign n21167 = ~n21165 & ~n21166;
  assign n21168 = ~n21142 & ~n21158;
  assign n21169 = n21142 & ~n21161;
  assign n21170 = ~n21168 & ~n21169;
  assign n21171 = ~n21167 & ~n21170;
  assign n21172 = ~n21164 & ~n21171;
  assign n21173 = ~n19728 & ~n19739;
  assign n21174 = n19728 & n19739;
  assign n21175 = ~n19733 & ~n21174;
  assign n21176 = ~n21173 & ~n21175;
  assign n21177 = ~n21172 & n21176;
  assign n21178 = n21172 & ~n21176;
  assign n21179 = ~n21177 & ~n21178;
  assign n21180 = pi139 & pi272;
  assign n21181 = pi138 & pi273;
  assign n21182 = n21180 & n21181;
  assign n21183 = ~n21180 & ~n21181;
  assign n21184 = ~n21182 & ~n21183;
  assign n21185 = ~n21179 & ~n21184;
  assign n21186 = n21172 & n21176;
  assign n21187 = ~n21172 & ~n21176;
  assign n21188 = ~n21186 & ~n21187;
  assign n21189 = pi272 & ~n21181;
  assign n21190 = pi139 & n21189;
  assign n21191 = pi273 & ~n21180;
  assign n21192 = pi138 & n21191;
  assign n21193 = ~n21190 & ~n21192;
  assign n21194 = ~n21188 & ~n21193;
  assign n21195 = ~n21185 & ~n21194;
  assign n21196 = ~n19757 & ~n19764;
  assign n21197 = ~n19752 & n21196;
  assign n21198 = ~n19765 & ~n21197;
  assign n21199 = n21195 & n21198;
  assign n21200 = ~n21195 & ~n21198;
  assign n21201 = ~n21199 & ~n21200;
  assign n21202 = pi140 & pi271;
  assign n21203 = ~n19744 & ~n19757;
  assign n21204 = ~n19752 & n21203;
  assign n21205 = n19744 & ~n19760;
  assign n21206 = ~n21204 & ~n21205;
  assign n21207 = ~n19587 & ~n21206;
  assign n21208 = n19744 & ~n19757;
  assign n21209 = ~n19752 & n21208;
  assign n21210 = ~n19744 & ~n19760;
  assign n21211 = ~n21209 & ~n21210;
  assign n21212 = pi271 & ~n21211;
  assign n21213 = pi139 & n21212;
  assign n21214 = ~n21207 & ~n21213;
  assign n21215 = n19776 & n21214;
  assign n21216 = ~n19776 & ~n21214;
  assign n21217 = n19753 & ~n21216;
  assign n21218 = ~n21215 & ~n21217;
  assign n21219 = n21202 & ~n21218;
  assign n21220 = ~n19753 & ~n21215;
  assign n21221 = ~n21216 & ~n21220;
  assign n21222 = ~n21202 & ~n21221;
  assign n21223 = ~n21219 & ~n21222;
  assign n21224 = ~n21201 & ~n21223;
  assign n21225 = n21195 & ~n21198;
  assign n21226 = ~n21195 & n21198;
  assign n21227 = ~n21225 & ~n21226;
  assign n21228 = ~n21202 & ~n21218;
  assign n21229 = n21202 & ~n21221;
  assign n21230 = ~n21228 & ~n21229;
  assign n21231 = ~n21227 & ~n21230;
  assign n21232 = ~n21224 & ~n21231;
  assign n21233 = ~n19780 & ~n19791;
  assign n21234 = n19780 & n19791;
  assign n21235 = ~n19785 & ~n21234;
  assign n21236 = ~n21233 & ~n21235;
  assign n21237 = ~n21232 & n21236;
  assign n21238 = n21232 & ~n21236;
  assign n21239 = ~n21237 & ~n21238;
  assign n21240 = pi142 & pi269;
  assign n21241 = pi141 & pi270;
  assign n21242 = n21240 & n21241;
  assign n21243 = ~n21240 & ~n21241;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = ~n21239 & ~n21244;
  assign n21246 = n21232 & n21236;
  assign n21247 = ~n21232 & ~n21236;
  assign n21248 = ~n21246 & ~n21247;
  assign n21249 = pi269 & ~n21241;
  assign n21250 = pi142 & n21249;
  assign n21251 = pi270 & ~n21240;
  assign n21252 = pi141 & n21251;
  assign n21253 = ~n21250 & ~n21252;
  assign n21254 = ~n21248 & ~n21253;
  assign n21255 = ~n21245 & ~n21254;
  assign n21256 = ~n19809 & ~n19816;
  assign n21257 = ~n19804 & n21256;
  assign n21258 = ~n19817 & ~n21257;
  assign n21259 = n21255 & ~n21258;
  assign n21260 = ~n21255 & n21258;
  assign n21261 = ~n21259 & ~n21260;
  assign n21262 = pi143 & pi268;
  assign n21263 = ~n19796 & ~n19809;
  assign n21264 = ~n19804 & n21263;
  assign n21265 = n19796 & ~n19812;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = ~n19586 & ~n21266;
  assign n21268 = n19796 & ~n19809;
  assign n21269 = ~n19804 & n21268;
  assign n21270 = ~n19796 & ~n19812;
  assign n21271 = ~n21269 & ~n21270;
  assign n21272 = pi268 & ~n21271;
  assign n21273 = pi142 & n21272;
  assign n21274 = ~n21267 & ~n21273;
  assign n21275 = n19828 & n21274;
  assign n21276 = ~n19828 & ~n21274;
  assign n21277 = n19805 & ~n21276;
  assign n21278 = ~n21275 & ~n21277;
  assign n21279 = n21262 & ~n21278;
  assign n21280 = ~n19805 & ~n21275;
  assign n21281 = ~n21276 & ~n21280;
  assign n21282 = ~n21262 & ~n21281;
  assign n21283 = ~n21279 & ~n21282;
  assign n21284 = ~n21261 & ~n21283;
  assign n21285 = n21255 & n21258;
  assign n21286 = ~n21255 & ~n21258;
  assign n21287 = ~n21285 & ~n21286;
  assign n21288 = ~n21262 & ~n21278;
  assign n21289 = n21262 & ~n21281;
  assign n21290 = ~n21288 & ~n21289;
  assign n21291 = ~n21287 & ~n21290;
  assign n21292 = ~n21284 & ~n21291;
  assign n21293 = n19832 & ~n19843;
  assign n21294 = ~n19832 & n19843;
  assign n21295 = ~n19834 & ~n21294;
  assign n21296 = ~n21293 & ~n21295;
  assign n21297 = ~n21292 & n21296;
  assign n21298 = n21292 & ~n21296;
  assign n21299 = ~n21297 & ~n21298;
  assign n21300 = pi145 & pi266;
  assign n21301 = pi144 & pi267;
  assign n21302 = n21300 & n21301;
  assign n21303 = ~n21300 & ~n21301;
  assign n21304 = ~n21302 & ~n21303;
  assign n21305 = ~n21299 & ~n21304;
  assign n21306 = n21292 & n21296;
  assign n21307 = ~n21292 & ~n21296;
  assign n21308 = ~n21306 & ~n21307;
  assign n21309 = pi266 & ~n21301;
  assign n21310 = pi145 & n21309;
  assign n21311 = pi267 & ~n21300;
  assign n21312 = pi144 & n21311;
  assign n21313 = ~n21310 & ~n21312;
  assign n21314 = ~n21308 & ~n21313;
  assign n21315 = ~n21305 & ~n21314;
  assign n21316 = ~n19864 & ~n19868;
  assign n21317 = ~n19869 & ~n21316;
  assign n21318 = n21315 & ~n21317;
  assign n21319 = ~n21315 & n21317;
  assign n21320 = ~n21318 & ~n21319;
  assign n21321 = pi146 & pi265;
  assign n21322 = ~n19848 & ~n19861;
  assign n21323 = ~n19857 & n21322;
  assign n21324 = n19848 & ~n19864;
  assign n21325 = ~n21323 & ~n21324;
  assign n21326 = ~n19585 & ~n21325;
  assign n21327 = n19848 & ~n19861;
  assign n21328 = ~n19857 & n21327;
  assign n21329 = ~n19848 & ~n19864;
  assign n21330 = ~n21328 & ~n21329;
  assign n21331 = pi265 & ~n21330;
  assign n21332 = pi145 & n21331;
  assign n21333 = ~n21326 & ~n21332;
  assign n21334 = n19880 & n21333;
  assign n21335 = ~n19880 & ~n21333;
  assign n21336 = n19858 & ~n21335;
  assign n21337 = ~n21334 & ~n21336;
  assign n21338 = n21321 & ~n21337;
  assign n21339 = ~n19858 & ~n21334;
  assign n21340 = ~n21335 & ~n21339;
  assign n21341 = ~n21321 & ~n21340;
  assign n21342 = ~n21338 & ~n21341;
  assign n21343 = ~n21320 & ~n21342;
  assign n21344 = n21315 & n21317;
  assign n21345 = ~n21315 & ~n21317;
  assign n21346 = ~n21344 & ~n21345;
  assign n21347 = ~n21321 & ~n21337;
  assign n21348 = n21321 & ~n21340;
  assign n21349 = ~n21347 & ~n21348;
  assign n21350 = ~n21346 & ~n21349;
  assign n21351 = ~n21343 & ~n21350;
  assign n21352 = n19886 & ~n19889;
  assign n21353 = n18385 & ~n18390;
  assign n21354 = ~n18391 & ~n21353;
  assign n21355 = ~n19886 & n19889;
  assign n21356 = ~n21354 & ~n21355;
  assign n21357 = ~n21352 & ~n21356;
  assign n21358 = ~n21351 & n21357;
  assign n21359 = n21351 & ~n21357;
  assign n21360 = ~n21358 & ~n21359;
  assign n21361 = pi148 & pi263;
  assign n21362 = pi147 & pi264;
  assign n21363 = n21361 & n21362;
  assign n21364 = ~n21361 & ~n21362;
  assign n21365 = ~n21363 & ~n21364;
  assign n21366 = ~n21360 & ~n21365;
  assign n21367 = n21351 & n21357;
  assign n21368 = ~n21351 & ~n21357;
  assign n21369 = ~n21367 & ~n21368;
  assign n21370 = pi263 & ~n21362;
  assign n21371 = pi148 & n21370;
  assign n21372 = pi264 & ~n21361;
  assign n21373 = pi147 & n21372;
  assign n21374 = ~n21371 & ~n21373;
  assign n21375 = ~n21369 & ~n21374;
  assign n21376 = ~n21366 & ~n21375;
  assign n21377 = ~n19899 & ~n19909;
  assign n21378 = n19899 & n19909;
  assign n21379 = ~n19900 & ~n21378;
  assign n21380 = ~n19566 & n21379;
  assign n21381 = ~n21377 & ~n21380;
  assign n21382 = n21376 & ~n21381;
  assign n21383 = ~n21376 & n21381;
  assign n21384 = ~n21382 & ~n21383;
  assign n21385 = pi149 & pi262;
  assign n21386 = ~n19574 & ~n19915;
  assign n21387 = n19574 & n19915;
  assign n21388 = n19584 & ~n21387;
  assign n21389 = ~n21386 & ~n21388;
  assign n21390 = n21385 & ~n21389;
  assign n21391 = ~n19584 & ~n21386;
  assign n21392 = ~n21387 & ~n21391;
  assign n21393 = ~n21385 & ~n21392;
  assign n21394 = ~n21390 & ~n21393;
  assign n21395 = ~n21384 & ~n21394;
  assign n21396 = n21376 & n21381;
  assign n21397 = ~n21376 & ~n21381;
  assign n21398 = ~n21396 & ~n21397;
  assign n21399 = ~n21385 & ~n21389;
  assign n21400 = n21385 & ~n21392;
  assign n21401 = ~n21399 & ~n21400;
  assign n21402 = ~n21398 & ~n21401;
  assign n21403 = ~n21395 & ~n21402;
  assign n21404 = pi260 & n19580;
  assign n21405 = pi150 & n21404;
  assign n21406 = ~n19580 & ~n19921;
  assign n21407 = ~n19574 & n19915;
  assign n21408 = n19574 & ~n19915;
  assign n21409 = ~n21407 & ~n21408;
  assign n21410 = ~n19584 & ~n21409;
  assign n21411 = ~n21386 & ~n21387;
  assign n21412 = n19584 & ~n21411;
  assign n21413 = ~n21410 & ~n21412;
  assign n21414 = ~n21406 & ~n21413;
  assign n21415 = ~n21405 & ~n21414;
  assign n21416 = n21403 & n21415;
  assign n21417 = ~n21403 & ~n21415;
  assign n21418 = ~n21416 & ~n21417;
  assign n21419 = pi261 & ~n21418;
  assign n21420 = pi150 & n21419;
  assign n21421 = pi150 & pi261;
  assign n21422 = ~n21403 & n21415;
  assign n21423 = n21403 & ~n21415;
  assign n21424 = ~n21422 & ~n21423;
  assign n21425 = ~n21421 & ~n21424;
  assign n21426 = ~n21420 & ~n21425;
  assign n21427 = ~n20990 & n21426;
  assign n21428 = n20990 & ~n21426;
  assign n21429 = ~n21427 & ~n21428;
  assign n21430 = pi153 & pi258;
  assign n21431 = pi152 & pi259;
  assign n21432 = ~n21430 & ~n21431;
  assign n21433 = n21430 & n21431;
  assign n21434 = ~n21432 & ~n21433;
  assign n21435 = n19936 & ~n19949;
  assign n21436 = ~n19936 & n19949;
  assign n21437 = ~n21435 & ~n21436;
  assign n21438 = pi258 & ~n21437;
  assign n21439 = pi152 & n21438;
  assign n21440 = n19936 & n19949;
  assign n21441 = ~n19936 & ~n19949;
  assign n21442 = ~n21440 & ~n21441;
  assign n21443 = pi258 & ~n21442;
  assign n21444 = pi152 & n21443;
  assign n21445 = ~n19955 & ~n21437;
  assign n21446 = ~n21444 & ~n21445;
  assign n21447 = n21439 & ~n21446;
  assign n21448 = ~n21439 & n21446;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = ~n21434 & ~n21449;
  assign n21451 = n21430 & ~n21431;
  assign n21452 = ~n21430 & n21431;
  assign n21453 = ~n21451 & ~n21452;
  assign n21454 = ~n21439 & ~n21446;
  assign n21455 = n21439 & n21446;
  assign n21456 = ~n21454 & ~n21455;
  assign n21457 = ~n21453 & ~n21456;
  assign n21458 = ~n21450 & ~n21457;
  assign n21459 = ~n21429 & ~n21458;
  assign n21460 = ~n20990 & ~n21426;
  assign n21461 = n20990 & n21426;
  assign n21462 = ~n21460 & ~n21461;
  assign n21463 = ~n21449 & ~n21453;
  assign n21464 = ~n21434 & ~n21456;
  assign n21465 = ~n21463 & ~n21464;
  assign n21466 = ~n21462 & ~n21465;
  assign n21467 = ~n21459 & ~n21466;
  assign n21468 = ~n19940 & ~n21446;
  assign n21469 = n19940 & n21446;
  assign n21470 = ~n19548 & ~n21469;
  assign n21471 = ~n21468 & ~n21470;
  assign n21472 = n21467 & ~n21471;
  assign n21473 = ~n21467 & n21471;
  assign n21474 = ~n21472 & ~n21473;
  assign n21475 = n20978 & ~n21474;
  assign n21476 = pi322 & n21475;
  assign n21477 = ~n21467 & ~n21471;
  assign n21478 = n21467 & n21471;
  assign n21479 = ~n21477 & ~n21478;
  assign n21480 = pi322 & n21479;
  assign n21481 = ~n20978 & ~n21480;
  assign n21482 = ~n21476 & ~n21481;
  assign n21483 = ~n20972 & ~n21482;
  assign n21484 = ~n20978 & ~n21474;
  assign n21485 = pi322 & n21484;
  assign n21486 = n20978 & ~n21480;
  assign n21487 = ~n21485 & ~n21486;
  assign n21488 = n19970 & ~n21487;
  assign n21489 = pi323 & n21488;
  assign n21490 = ~n21483 & ~n21489;
  assign n21491 = ~n20971 & n21490;
  assign n21492 = n20971 & ~n21490;
  assign n21493 = ~n21491 & ~n21492;
  assign n21494 = pi326 & n18461;
  assign n21495 = pi325 & n19539;
  assign n21496 = n21494 & n21495;
  assign n21497 = ~n21494 & ~n21495;
  assign n21498 = ~n21496 & ~n21497;
  assign n21499 = ~n21493 & ~n21498;
  assign n21500 = n20971 & n21490;
  assign n21501 = ~n20971 & ~n21490;
  assign n21502 = ~n21500 & ~n21501;
  assign n21503 = ~n21494 & n21495;
  assign n21504 = n21494 & ~n21495;
  assign n21505 = ~n21503 & ~n21504;
  assign n21506 = ~n21502 & ~n21505;
  assign n21507 = ~n21499 & ~n21506;
  assign n21508 = ~n20970 & ~n21507;
  assign n21509 = ~n20963 & ~n20967;
  assign n21510 = n20963 & n20967;
  assign n21511 = ~n21509 & ~n21510;
  assign n21512 = ~n21498 & ~n21502;
  assign n21513 = ~n21493 & ~n21505;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = ~n21511 & ~n21514;
  assign n21516 = ~n21508 & ~n21515;
  assign n21517 = ~n19529 & n19990;
  assign n21518 = n19529 & ~n19990;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = ~n19986 & n19995;
  assign n21521 = n19986 & ~n19995;
  assign n21522 = ~n21520 & ~n21521;
  assign n21523 = n19533 & ~n19994;
  assign n21524 = ~n21522 & ~n21523;
  assign n21525 = ~n21519 & n21524;
  assign n21526 = ~n19533 & n19994;
  assign n21527 = ~n19529 & ~n19990;
  assign n21528 = n19529 & n19990;
  assign n21529 = ~n21527 & ~n21528;
  assign n21530 = n19986 & n19995;
  assign n21531 = ~n19986 & ~n19995;
  assign n21532 = ~n21530 & ~n21531;
  assign n21533 = ~n21523 & ~n21532;
  assign n21534 = ~n21529 & n21533;
  assign n21535 = ~n21526 & ~n21534;
  assign n21536 = ~n21525 & n21535;
  assign n21537 = n21516 & n21536;
  assign n21538 = ~n21516 & ~n21536;
  assign n21539 = ~n21537 & ~n21538;
  assign n21540 = pi328 & n12917;
  assign n21541 = pi327 & n13762;
  assign n21542 = n21540 & n21541;
  assign n21543 = ~n21540 & ~n21541;
  assign n21544 = ~n21542 & ~n21543;
  assign n21545 = ~n21539 & ~n21544;
  assign n21546 = ~n21516 & n21536;
  assign n21547 = n21516 & ~n21536;
  assign n21548 = ~n21546 & ~n21547;
  assign n21549 = ~n21540 & n21541;
  assign n21550 = n21540 & ~n21541;
  assign n21551 = ~n21549 & ~n21550;
  assign n21552 = ~n21548 & ~n21551;
  assign n21553 = ~n21545 & ~n21552;
  assign n21554 = ~n20947 & ~n21553;
  assign n21555 = ~n20937 & n20944;
  assign n21556 = n20937 & ~n20944;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 = ~n21544 & ~n21548;
  assign n21559 = ~n21539 & ~n21551;
  assign n21560 = ~n21558 & ~n21559;
  assign n21561 = ~n21557 & ~n21560;
  assign n21562 = ~n21554 & ~n21561;
  assign n21563 = ~n20933 & n21562;
  assign n21564 = n20933 & ~n21562;
  assign n21565 = ~n21563 & ~n21564;
  assign n21566 = pi331 & n11366;
  assign n21567 = pi330 & n11384;
  assign n21568 = n10561 & ~n19471;
  assign n21569 = ~n19472 & ~n21568;
  assign n21570 = n11366 & ~n21569;
  assign n21571 = pi330 & n21570;
  assign n21572 = ~n11366 & ~n21568;
  assign n21573 = pi330 & ~n21572;
  assign n21574 = ~n19472 & ~n21573;
  assign n21575 = ~n20922 & ~n21574;
  assign n21576 = ~n21571 & ~n21575;
  assign n21577 = ~n21567 & ~n21576;
  assign n21578 = n20918 & ~n21574;
  assign n21579 = n11384 & ~n21578;
  assign n21580 = pi330 & n21579;
  assign n21581 = ~n21571 & n21580;
  assign n21582 = ~n21577 & ~n21581;
  assign n21583 = n21566 & ~n21582;
  assign n21584 = ~n21566 & n21582;
  assign n21585 = ~n21583 & ~n21584;
  assign n21586 = ~n21565 & ~n21585;
  assign n21587 = n20933 & n21562;
  assign n21588 = ~n20933 & ~n21562;
  assign n21589 = ~n21587 & ~n21588;
  assign n21590 = ~n21566 & ~n21582;
  assign n21591 = n21566 & n21582;
  assign n21592 = ~n21590 & ~n21591;
  assign n21593 = ~n21589 & ~n21592;
  assign n21594 = ~n21586 & ~n21593;
  assign n21595 = ~n20932 & ~n21594;
  assign n21596 = ~n20915 & ~n20929;
  assign n21597 = n20915 & n20929;
  assign n21598 = ~n21596 & ~n21597;
  assign n21599 = ~n21585 & ~n21589;
  assign n21600 = ~n21565 & ~n21592;
  assign n21601 = ~n21599 & ~n21600;
  assign n21602 = ~n21598 & ~n21601;
  assign n21603 = ~n21595 & ~n21602;
  assign n21604 = ~n20067 & n20071;
  assign n21605 = ~n20063 & ~n20082;
  assign n21606 = n20063 & n20082;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = n20067 & ~n20071;
  assign n21609 = ~n21607 & ~n21608;
  assign n21610 = ~n21604 & ~n21609;
  assign n21611 = n21603 & n21610;
  assign n21612 = ~n21603 & ~n21610;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 = pi333 & n9205;
  assign n21615 = ~n20063 & ~n20077;
  assign n21616 = n20063 & n20077;
  assign n21617 = ~n9205 & ~n21616;
  assign n21618 = ~n21615 & ~n21617;
  assign n21619 = n10561 & ~n21618;
  assign n21620 = ~n10561 & ~n21615;
  assign n21621 = n9205 & n21620;
  assign n21622 = ~n21619 & ~n21621;
  assign n21623 = pi332 & ~n21622;
  assign n21624 = pi332 & n10561;
  assign n21625 = n20063 & ~n21624;
  assign n21626 = n20077 & n21625;
  assign n21627 = ~n21623 & ~n21626;
  assign n21628 = ~n21614 & n21627;
  assign n21629 = n21614 & ~n21627;
  assign n21630 = ~n21628 & ~n21629;
  assign n21631 = pi334 & n6556;
  assign n21632 = n17926 & ~n19403;
  assign n21633 = ~n17926 & ~n19412;
  assign n21634 = ~n21632 & ~n21633;
  assign n21635 = ~n20089 & ~n21634;
  assign n21636 = ~n20092 & ~n21635;
  assign n21637 = n20087 & ~n21636;
  assign n21638 = ~n20085 & ~n21637;
  assign n21639 = ~n20123 & n21638;
  assign n21640 = ~n20087 & n21636;
  assign n21641 = ~n20114 & ~n21637;
  assign n21642 = ~n20070 & n21641;
  assign n21643 = ~n21640 & ~n21642;
  assign n21644 = ~n21639 & n21643;
  assign n21645 = n21631 & ~n21644;
  assign n21646 = ~n21631 & n21644;
  assign n21647 = ~n21645 & ~n21646;
  assign n21648 = ~n21630 & ~n21647;
  assign n21649 = n21614 & n21627;
  assign n21650 = ~n21614 & ~n21627;
  assign n21651 = ~n21649 & ~n21650;
  assign n21652 = ~n21631 & ~n21644;
  assign n21653 = n21631 & n21644;
  assign n21654 = ~n21652 & ~n21653;
  assign n21655 = ~n21651 & ~n21654;
  assign n21656 = ~n21648 & ~n21655;
  assign n21657 = ~n21613 & ~n21656;
  assign n21658 = n21603 & ~n21610;
  assign n21659 = ~n21603 & n21610;
  assign n21660 = ~n21658 & ~n21659;
  assign n21661 = ~n21647 & ~n21651;
  assign n21662 = ~n21630 & ~n21654;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = ~n21660 & ~n21663;
  assign n21665 = ~n21657 & ~n21664;
  assign n21666 = ~n20891 & n21665;
  assign n21667 = n20891 & ~n21665;
  assign n21668 = ~n21666 & ~n21667;
  assign n21669 = pi337 & n5714;
  assign n21670 = n5257 & ~n19434;
  assign n21671 = pi336 & n21670;
  assign n21672 = ~n19435 & ~n21671;
  assign n21673 = ~pi336 & ~n21672;
  assign n21674 = ~n19443 & n21672;
  assign n21675 = ~n5732 & ~n21674;
  assign n21676 = ~n21673 & ~n21675;
  assign n21677 = ~n20880 & ~n21676;
  assign n21678 = ~n5732 & ~n21672;
  assign n21679 = n5714 & n21678;
  assign n21680 = ~n5714 & n21672;
  assign n21681 = n5714 & ~n21672;
  assign n21682 = ~n20876 & ~n21681;
  assign n21683 = ~n21680 & ~n21682;
  assign n21684 = n5732 & ~n21683;
  assign n21685 = ~n21679 & ~n21684;
  assign n21686 = pi336 & ~n21685;
  assign n21687 = ~n21677 & ~n21686;
  assign n21688 = n21669 & ~n21687;
  assign n21689 = ~n21669 & n21687;
  assign n21690 = ~n21688 & ~n21689;
  assign n21691 = ~n21668 & ~n21690;
  assign n21692 = n20891 & n21665;
  assign n21693 = ~n20891 & ~n21665;
  assign n21694 = ~n21692 & ~n21693;
  assign n21695 = ~n21669 & ~n21687;
  assign n21696 = n21669 & n21687;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = ~n21694 & ~n21697;
  assign n21699 = ~n21691 & ~n21698;
  assign n21700 = ~n20890 & ~n21699;
  assign n21701 = ~n20873 & ~n20887;
  assign n21702 = n20873 & n20887;
  assign n21703 = ~n21701 & ~n21702;
  assign n21704 = ~n21690 & ~n21694;
  assign n21705 = ~n21668 & ~n21697;
  assign n21706 = ~n21704 & ~n21705;
  assign n21707 = ~n21703 & ~n21706;
  assign n21708 = ~n21700 & ~n21707;
  assign n21709 = ~n20153 & n20157;
  assign n21710 = ~n20149 & ~n20168;
  assign n21711 = n20149 & n20168;
  assign n21712 = ~n21710 & ~n21711;
  assign n21713 = n20153 & ~n20157;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = ~n21709 & ~n21714;
  assign n21716 = n21708 & n21715;
  assign n21717 = ~n21708 & ~n21715;
  assign n21718 = ~n21716 & ~n21717;
  assign n21719 = pi339 & n4596;
  assign n21720 = ~n20149 & ~n20163;
  assign n21721 = n20149 & n20163;
  assign n21722 = ~n4596 & ~n21721;
  assign n21723 = ~n21720 & ~n21722;
  assign n21724 = n5257 & ~n21723;
  assign n21725 = ~n5257 & ~n21720;
  assign n21726 = n4596 & n21725;
  assign n21727 = ~n21724 & ~n21726;
  assign n21728 = pi338 & ~n21727;
  assign n21729 = pi338 & n5257;
  assign n21730 = n20149 & ~n21729;
  assign n21731 = n20163 & n21730;
  assign n21732 = ~n21728 & ~n21731;
  assign n21733 = ~n21719 & n21732;
  assign n21734 = n21719 & ~n21732;
  assign n21735 = ~n21733 & ~n21734;
  assign n21736 = pi340 & n2887;
  assign n21737 = ~n20171 & ~n20189;
  assign n21738 = ~n20196 & n21737;
  assign n21739 = ~n20187 & ~n20189;
  assign n21740 = ~n20156 & n21739;
  assign n21741 = ~n20188 & ~n21740;
  assign n21742 = ~n21738 & n21741;
  assign n21743 = n21736 & ~n21742;
  assign n21744 = ~n21736 & n21742;
  assign n21745 = ~n21743 & ~n21744;
  assign n21746 = ~n21735 & ~n21745;
  assign n21747 = n21719 & n21732;
  assign n21748 = ~n21719 & ~n21732;
  assign n21749 = ~n21747 & ~n21748;
  assign n21750 = ~n21736 & ~n21742;
  assign n21751 = n21736 & n21742;
  assign n21752 = ~n21750 & ~n21751;
  assign n21753 = ~n21749 & ~n21752;
  assign n21754 = ~n21746 & ~n21753;
  assign n21755 = ~n21718 & ~n21754;
  assign n21756 = n21708 & ~n21715;
  assign n21757 = ~n21708 & n21715;
  assign n21758 = ~n21756 & ~n21757;
  assign n21759 = ~n21745 & ~n21749;
  assign n21760 = ~n21735 & ~n21752;
  assign n21761 = ~n21759 & ~n21760;
  assign n21762 = ~n21758 & ~n21761;
  assign n21763 = ~n21755 & ~n21762;
  assign n21764 = ~n20852 & n21763;
  assign n21765 = n20852 & ~n21763;
  assign n21766 = ~n21764 & ~n21765;
  assign n21767 = pi343 & n1729;
  assign n21768 = pi342 & n2091;
  assign n21769 = ~n20206 & n20208;
  assign n21770 = ~n21768 & ~n21769;
  assign n21771 = n19400 & n21770;
  assign n21772 = n20206 & ~n20208;
  assign n21773 = n21768 & ~n21772;
  assign n21774 = ~n19400 & n21773;
  assign n21775 = ~n21771 & ~n21774;
  assign n21776 = ~n20841 & ~n21775;
  assign n21777 = n19400 & n21773;
  assign n21778 = ~n19400 & n21770;
  assign n21779 = ~n21777 & ~n21778;
  assign n21780 = ~n20831 & ~n21779;
  assign n21781 = ~n20208 & ~n21768;
  assign n21782 = n20206 & n21781;
  assign n21783 = n20208 & n21768;
  assign n21784 = ~n20206 & n21783;
  assign n21785 = ~n21782 & ~n21784;
  assign n21786 = ~n21780 & n21785;
  assign n21787 = ~n21776 & n21786;
  assign n21788 = n21767 & ~n21787;
  assign n21789 = ~n21767 & n21787;
  assign n21790 = ~n21788 & ~n21789;
  assign n21791 = ~n21766 & ~n21790;
  assign n21792 = n20852 & n21763;
  assign n21793 = ~n20852 & ~n21763;
  assign n21794 = ~n21792 & ~n21793;
  assign n21795 = ~n21767 & ~n21787;
  assign n21796 = n21767 & n21787;
  assign n21797 = ~n21795 & ~n21796;
  assign n21798 = ~n21794 & ~n21797;
  assign n21799 = ~n21791 & ~n21798;
  assign n21800 = ~n20851 & ~n21799;
  assign n21801 = ~n20828 & ~n20848;
  assign n21802 = n20828 & n20848;
  assign n21803 = ~n21801 & ~n21802;
  assign n21804 = ~n21790 & ~n21794;
  assign n21805 = ~n21766 & ~n21797;
  assign n21806 = ~n21804 & ~n21805;
  assign n21807 = ~n21803 & ~n21806;
  assign n21808 = ~n21800 & ~n21807;
  assign n21809 = ~n1154 & n19367;
  assign n21810 = pi345 & n21809;
  assign n21811 = ~n19367 & ~n20253;
  assign n21812 = ~n20234 & ~n20249;
  assign n21813 = ~n20243 & n21812;
  assign n21814 = n20234 & ~n20250;
  assign n21815 = ~n21813 & ~n21814;
  assign n21816 = ~n21811 & ~n21815;
  assign n21817 = ~n21810 & ~n21816;
  assign n21818 = n21808 & ~n21817;
  assign n21819 = ~n21808 & n21817;
  assign n21820 = ~n21818 & ~n21819;
  assign n21821 = n20234 & ~n20249;
  assign n21822 = ~n20243 & ~n21821;
  assign n21823 = n1442 & ~n21822;
  assign n21824 = pi344 & n21823;
  assign n21825 = pi344 & n1442;
  assign n21826 = ~n21821 & ~n21825;
  assign n21827 = ~n20243 & n21826;
  assign n21828 = ~n21824 & ~n21827;
  assign n21829 = ~n1256 & ~n21828;
  assign n21830 = pi345 & n21829;
  assign n21831 = pi345 & ~n1256;
  assign n21832 = ~n21827 & ~n21831;
  assign n21833 = ~n21824 & n21832;
  assign n21834 = ~n21830 & ~n21833;
  assign n21835 = ~n21820 & ~n21834;
  assign n21836 = n21808 & n21817;
  assign n21837 = ~n21808 & ~n21817;
  assign n21838 = ~n21836 & ~n21837;
  assign n21839 = ~n21828 & ~n21831;
  assign n21840 = n21828 & n21831;
  assign n21841 = ~n21839 & ~n21840;
  assign n21842 = ~n21838 & ~n21841;
  assign n21843 = ~n21835 & ~n21842;
  assign n21844 = n20824 & ~n21843;
  assign n21845 = ~n20824 & n21843;
  assign n21846 = ~n21844 & ~n21845;
  assign n21847 = pi258 & ~n21846;
  assign n21848 = pi128 & n21847;
  assign n21849 = pi347 & n21848;
  assign n21850 = n20824 & n21843;
  assign n21851 = ~n20824 & ~n21843;
  assign n21852 = ~n21850 & ~n21851;
  assign n21853 = pi347 & n1156;
  assign n21854 = ~n21852 & ~n21853;
  assign n21855 = ~n21849 & ~n21854;
  assign n21856 = pi283 & ~n21855;
  assign n21857 = ~pi283 & n21855;
  assign n21858 = ~n21856 & ~n21857;
  assign n21859 = ~n20818 & n21858;
  assign n21860 = n20818 & ~n21858;
  assign n21861 = ~n21859 & ~n21860;
  assign n21862 = ~n20814 & ~n21861;
  assign n21863 = n20818 & n21858;
  assign n21864 = ~n20818 & ~n21858;
  assign n21865 = ~n21863 & ~n21864;
  assign n21866 = ~n20813 & ~n21865;
  assign n21867 = ~n20810 & n21866;
  assign n21868 = ~n21862 & ~n21867;
  assign n21869 = n19358 & ~n20288;
  assign n21870 = ~n19358 & n20288;
  assign n21871 = ~n20276 & ~n21870;
  assign n21872 = ~n21869 & ~n21871;
  assign n21873 = n21868 & ~n21872;
  assign n21874 = ~n21868 & n21872;
  assign n21875 = ~n21873 & ~n21874;
  assign n21876 = ~n831 & ~n21875;
  assign n21877 = ~n20297 & ~n21876;
  assign n21878 = pi161 & ~n21877;
  assign n21879 = pi089 & ~pi161;
  assign n21880 = ~n21878 & ~n21879;
  assign po218 = ~pi160 & ~n21880;
  assign n21882 = pi090 & ~pi161;
  assign n21883 = ~n1154 & ~n21843;
  assign n21884 = n1154 & n21843;
  assign n21885 = ~n20265 & ~n21884;
  assign n21886 = n1156 & n21885;
  assign n21887 = ~n21883 & ~n21886;
  assign n21888 = n1256 & ~n21887;
  assign n21889 = ~n20821 & ~n21883;
  assign n21890 = ~n21884 & ~n21889;
  assign n21891 = ~n1256 & ~n21890;
  assign n21892 = ~n21888 & ~n21891;
  assign n21893 = pi346 & ~n21892;
  assign n21894 = ~n20828 & ~n21763;
  assign n21895 = n20828 & n21763;
  assign n21896 = ~n21894 & ~n21895;
  assign n21897 = n20852 & ~n21787;
  assign n21898 = ~n20852 & n21787;
  assign n21899 = ~n21897 & ~n21898;
  assign n21900 = n20848 & ~n21767;
  assign n21901 = ~n21899 & ~n21900;
  assign n21902 = ~n21896 & n21901;
  assign n21903 = ~n20848 & n21767;
  assign n21904 = ~n20828 & n21763;
  assign n21905 = n20828 & ~n21763;
  assign n21906 = ~n21904 & ~n21905;
  assign n21907 = ~n20852 & ~n21787;
  assign n21908 = n20852 & n21787;
  assign n21909 = ~n21907 & ~n21908;
  assign n21910 = ~n21900 & ~n21909;
  assign n21911 = ~n21906 & n21910;
  assign n21912 = ~n21903 & ~n21911;
  assign n21913 = ~n21902 & n21912;
  assign n21914 = ~n1256 & ~n21817;
  assign n21915 = pi345 & n21914;
  assign n21916 = ~n21808 & ~n21827;
  assign n21917 = ~n21824 & n21916;
  assign n21918 = n21808 & ~n21828;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = n21817 & ~n21831;
  assign n21921 = ~n21919 & ~n21920;
  assign n21922 = ~n21915 & ~n21921;
  assign n21923 = n21913 & ~n21922;
  assign n21924 = ~n21913 & n21922;
  assign n21925 = ~n21923 & ~n21924;
  assign n21926 = pi343 & n2091;
  assign n21927 = n20873 & n21665;
  assign n21928 = ~n20873 & ~n21665;
  assign n21929 = ~n21927 & ~n21928;
  assign n21930 = n20891 & ~n21687;
  assign n21931 = ~n20891 & n21687;
  assign n21932 = ~n21930 & ~n21931;
  assign n21933 = n20887 & ~n21669;
  assign n21934 = ~n21932 & ~n21933;
  assign n21935 = ~n21929 & n21934;
  assign n21936 = ~n20887 & n21669;
  assign n21937 = ~n20873 & n21665;
  assign n21938 = n20873 & ~n21665;
  assign n21939 = ~n21937 & ~n21938;
  assign n21940 = ~n20891 & ~n21687;
  assign n21941 = n20891 & n21687;
  assign n21942 = ~n21940 & ~n21941;
  assign n21943 = ~n21933 & ~n21942;
  assign n21944 = ~n21939 & n21943;
  assign n21945 = ~n21936 & ~n21944;
  assign n21946 = ~n21935 & n21945;
  assign n21947 = ~n21715 & n21719;
  assign n21948 = n21715 & ~n21719;
  assign n21949 = n4596 & ~n21720;
  assign n21950 = ~n21721 & ~n21949;
  assign n21951 = n5257 & ~n21950;
  assign n21952 = pi338 & n21951;
  assign n21953 = ~n5257 & ~n21949;
  assign n21954 = pi338 & ~n21953;
  assign n21955 = ~n21721 & ~n21954;
  assign n21956 = ~n21952 & ~n21955;
  assign n21957 = n21708 & ~n21956;
  assign n21958 = ~n21708 & n21956;
  assign n21959 = ~n21957 & ~n21958;
  assign n21960 = ~n21948 & ~n21959;
  assign n21961 = ~n21947 & ~n21960;
  assign n21962 = n21946 & ~n21961;
  assign n21963 = ~n21946 & n21961;
  assign n21964 = ~n21962 & ~n21963;
  assign n21965 = pi337 & n5732;
  assign n21966 = n20915 & n21562;
  assign n21967 = ~n20915 & ~n21562;
  assign n21968 = ~n21966 & ~n21967;
  assign n21969 = n20933 & ~n21582;
  assign n21970 = ~n20933 & n21582;
  assign n21971 = ~n21969 & ~n21970;
  assign n21972 = n20929 & ~n21566;
  assign n21973 = ~n21971 & ~n21972;
  assign n21974 = ~n21968 & n21973;
  assign n21975 = ~n20929 & n21566;
  assign n21976 = n20915 & ~n21562;
  assign n21977 = ~n20915 & n21562;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~n20933 & ~n21582;
  assign n21980 = n20933 & n21582;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = ~n21972 & ~n21981;
  assign n21983 = ~n21978 & n21982;
  assign n21984 = ~n21975 & ~n21983;
  assign n21985 = ~n21974 & n21984;
  assign n21986 = ~n21610 & n21614;
  assign n21987 = n21610 & ~n21614;
  assign n21988 = n9205 & ~n21615;
  assign n21989 = ~n21616 & ~n21988;
  assign n21990 = n10561 & ~n21989;
  assign n21991 = pi332 & n21990;
  assign n21992 = ~n10561 & ~n21988;
  assign n21993 = pi332 & ~n21992;
  assign n21994 = ~n21616 & ~n21993;
  assign n21995 = ~n21991 & ~n21994;
  assign n21996 = n21603 & ~n21995;
  assign n21997 = ~n21603 & n21995;
  assign n21998 = ~n21996 & ~n21997;
  assign n21999 = ~n21987 & ~n21998;
  assign n22000 = ~n21986 & ~n21999;
  assign n22001 = n21985 & ~n22000;
  assign n22002 = ~n21985 & n22000;
  assign n22003 = ~n22001 & ~n22002;
  assign n22004 = pi331 & n11384;
  assign n22005 = n20937 & ~n21536;
  assign n22006 = ~n20937 & n21536;
  assign n22007 = ~n22005 & ~n22006;
  assign n22008 = ~n21516 & n21541;
  assign n22009 = n21516 & ~n21541;
  assign n22010 = ~n22008 & ~n22009;
  assign n22011 = n20944 & ~n21540;
  assign n22012 = ~n22010 & ~n22011;
  assign n22013 = ~n22007 & n22012;
  assign n22014 = ~n20944 & n21540;
  assign n22015 = n20937 & n21536;
  assign n22016 = ~n20937 & ~n21536;
  assign n22017 = ~n22015 & ~n22016;
  assign n22018 = n21516 & n21541;
  assign n22019 = ~n21516 & ~n21541;
  assign n22020 = ~n22018 & ~n22019;
  assign n22021 = ~n22011 & ~n22020;
  assign n22022 = ~n22017 & n22021;
  assign n22023 = ~n22014 & ~n22022;
  assign n22024 = ~n22013 & n22023;
  assign n22025 = ~n20915 & n20933;
  assign n22026 = n20915 & ~n20933;
  assign n22027 = n21562 & ~n22026;
  assign n22028 = ~n22025 & ~n22027;
  assign n22029 = n22024 & ~n22028;
  assign n22030 = ~n22024 & n22028;
  assign n22031 = ~n22029 & ~n22030;
  assign n22032 = pi328 & n13762;
  assign n22033 = n21494 & ~n21536;
  assign n22034 = n19539 & ~n21493;
  assign n22035 = pi325 & n22034;
  assign n22036 = ~n21495 & ~n21502;
  assign n22037 = ~n22035 & ~n22036;
  assign n22038 = ~n21511 & ~n22037;
  assign n22039 = n19539 & ~n21502;
  assign n22040 = pi325 & n22039;
  assign n22041 = ~n21493 & ~n21495;
  assign n22042 = ~n22040 & ~n22041;
  assign n22043 = ~n20970 & ~n22042;
  assign n22044 = ~n22038 & ~n22043;
  assign n22045 = ~n21494 & n21536;
  assign n22046 = ~n22044 & ~n22045;
  assign n22047 = ~n22033 & ~n22046;
  assign n22048 = n20937 & ~n21541;
  assign n22049 = ~n21548 & ~n22048;
  assign n22050 = ~n20937 & n21541;
  assign n22051 = ~n22049 & ~n22050;
  assign n22052 = n22047 & ~n22051;
  assign n22053 = ~n22047 & n22051;
  assign n22054 = ~n22052 & ~n22053;
  assign n22055 = n19970 & ~n20978;
  assign n22056 = pi323 & n22055;
  assign n22057 = ~n20972 & n20978;
  assign n22058 = n21479 & ~n22057;
  assign n22059 = pi322 & n22058;
  assign n22060 = ~n22056 & ~n22059;
  assign n22061 = ~n20963 & n20971;
  assign n22062 = n20963 & ~n20971;
  assign n22063 = ~n21490 & ~n22062;
  assign n22064 = ~n22061 & ~n22063;
  assign n22065 = ~n22060 & n22064;
  assign n22066 = n22060 & ~n22064;
  assign n22067 = ~n22065 & ~n22066;
  assign n22068 = pi151 & pi261;
  assign n22069 = pi148 & pi264;
  assign n22070 = pi145 & pi267;
  assign n22071 = pi142 & pi270;
  assign n22072 = pi139 & pi273;
  assign n22073 = pi136 & pi276;
  assign n22074 = ~n21059 & n21064;
  assign n22075 = ~n21058 & ~n21064;
  assign n22076 = ~n21055 & n22075;
  assign n22077 = ~n22074 & ~n22076;
  assign n22078 = ~n21079 & n22077;
  assign n22079 = pi133 & pi279;
  assign n22080 = pi283 & ~n19594;
  assign n22081 = pi282 & n22080;
  assign n22082 = ~pi283 & n19594;
  assign n22083 = pi282 & ~n22082;
  assign n22084 = ~pi282 & ~n22080;
  assign n22085 = pi281 & ~n22084;
  assign n22086 = ~n22083 & ~n22085;
  assign n22087 = pi129 & ~n22086;
  assign n22088 = ~n22081 & ~n22087;
  assign n22089 = pi128 & ~n22088;
  assign n22090 = pi282 & ~n19594;
  assign n22091 = n19598 & n22090;
  assign n22092 = ~n22089 & ~n22091;
  assign n22093 = pi128 & pi284;
  assign n22094 = pi283 & ~n22093;
  assign n22095 = pi129 & n22094;
  assign n22096 = pi129 & pi283;
  assign n22097 = pi284 & ~n22096;
  assign n22098 = pi128 & n22097;
  assign n22099 = ~n22095 & ~n22098;
  assign n22100 = n22092 & n22099;
  assign n22101 = ~n22092 & ~n22099;
  assign n22102 = ~n22100 & ~n22101;
  assign n22103 = pi282 & ~n22102;
  assign n22104 = pi130 & n22103;
  assign n22105 = pi130 & pi282;
  assign n22106 = ~n22092 & n22099;
  assign n22107 = n22092 & ~n22099;
  assign n22108 = ~n22106 & ~n22107;
  assign n22109 = ~n22105 & ~n22108;
  assign n22110 = ~n22104 & ~n22109;
  assign n22111 = pi130 & pi281;
  assign n22112 = ~n20999 & ~n21025;
  assign n22113 = ~n19598 & ~n20992;
  assign n22114 = ~n21022 & ~n22113;
  assign n22115 = n20999 & ~n22114;
  assign n22116 = ~n22112 & ~n22115;
  assign n22117 = n22111 & n22116;
  assign n22118 = ~n22111 & ~n22116;
  assign n22119 = ~n21035 & ~n22118;
  assign n22120 = ~n19609 & n22119;
  assign n22121 = ~n22117 & ~n22120;
  assign n22122 = ~n22110 & n22121;
  assign n22123 = n22110 & ~n22121;
  assign n22124 = ~n22122 & ~n22123;
  assign n22125 = pi281 & ~n22124;
  assign n22126 = pi131 & n22125;
  assign n22127 = pi131 & pi281;
  assign n22128 = ~n22123 & ~n22127;
  assign n22129 = ~n22122 & n22128;
  assign n22130 = ~n22126 & ~n22129;
  assign n22131 = ~n21046 & ~n21048;
  assign n22132 = ~n21041 & ~n22131;
  assign n22133 = pi280 & ~n22132;
  assign n22134 = pi132 & n22133;
  assign n22135 = pi132 & pi280;
  assign n22136 = ~n22131 & ~n22135;
  assign n22137 = ~n21041 & n22136;
  assign n22138 = ~n22134 & ~n22137;
  assign n22139 = ~n22130 & ~n22138;
  assign n22140 = n22132 & n22135;
  assign n22141 = ~n22132 & ~n22135;
  assign n22142 = ~n22140 & ~n22141;
  assign n22143 = ~n22129 & ~n22142;
  assign n22144 = ~n22126 & n22143;
  assign n22145 = ~n22139 & ~n22144;
  assign n22146 = ~n21055 & n21064;
  assign n22147 = ~n22145 & ~n22146;
  assign n22148 = ~n21058 & n22147;
  assign n22149 = ~n21058 & ~n22146;
  assign n22150 = n22145 & ~n22149;
  assign n22151 = ~n22148 & ~n22150;
  assign n22152 = ~n22079 & ~n22151;
  assign n22153 = n22145 & ~n22146;
  assign n22154 = ~n21058 & n22153;
  assign n22155 = ~n22145 & ~n22149;
  assign n22156 = ~n22154 & ~n22155;
  assign n22157 = pi279 & ~n22156;
  assign n22158 = pi133 & n22157;
  assign n22159 = ~n22152 & ~n22158;
  assign n22160 = ~pi278 & ~n22159;
  assign n22161 = ~pi134 & ~n22159;
  assign n22162 = pi278 & n22159;
  assign n22163 = pi134 & n22162;
  assign n22164 = ~n22161 & ~n22163;
  assign n22165 = ~pi133 & ~n22164;
  assign n22166 = ~n22160 & ~n22165;
  assign n22167 = ~n22078 & ~n22166;
  assign n22168 = n21079 & n22159;
  assign n22169 = pi278 & ~n22077;
  assign n22170 = n22168 & n22169;
  assign n22171 = n21079 & n22077;
  assign n22172 = ~n21079 & ~n22077;
  assign n22173 = ~n22171 & ~n22172;
  assign n22174 = pi133 & ~n22173;
  assign n22175 = pi278 & n22078;
  assign n22176 = ~n22174 & ~n22175;
  assign n22177 = ~n22159 & ~n22176;
  assign n22178 = ~n22170 & ~n22177;
  assign n22179 = pi134 & ~n22178;
  assign n22180 = ~pi278 & n22077;
  assign n22181 = ~n21079 & n22159;
  assign n22182 = n22180 & n22181;
  assign n22183 = n21079 & ~n22159;
  assign n22184 = ~n22077 & n22183;
  assign n22185 = n21079 & ~n22077;
  assign n22186 = pi278 & ~n22185;
  assign n22187 = pi133 & n22186;
  assign n22188 = ~n22078 & ~n22187;
  assign n22189 = n22159 & ~n22188;
  assign n22190 = ~n22184 & ~n22189;
  assign n22191 = ~pi134 & ~n22190;
  assign n22192 = ~n22182 & ~n22191;
  assign n22193 = ~n22179 & n22192;
  assign n22194 = ~n22167 & n22193;
  assign n22195 = n21083 & ~n21108;
  assign n22196 = ~n21083 & n21108;
  assign n22197 = ~n21099 & ~n22196;
  assign n22198 = ~n22195 & ~n22197;
  assign n22199 = n22194 & n22198;
  assign n22200 = ~n22194 & ~n22198;
  assign n22201 = ~n22199 & ~n22200;
  assign n22202 = pi135 & pi277;
  assign n22203 = n21122 & ~n21128;
  assign n22204 = ~n21127 & ~n22203;
  assign n22205 = n22202 & ~n22204;
  assign n22206 = ~n21122 & ~n21127;
  assign n22207 = ~n21128 & ~n22206;
  assign n22208 = ~n22202 & ~n22207;
  assign n22209 = ~n22205 & ~n22208;
  assign n22210 = ~n22201 & ~n22209;
  assign n22211 = n22194 & ~n22198;
  assign n22212 = ~n22194 & n22198;
  assign n22213 = ~n22211 & ~n22212;
  assign n22214 = ~n22202 & ~n22204;
  assign n22215 = n22202 & ~n22207;
  assign n22216 = ~n22214 & ~n22215;
  assign n22217 = ~n22213 & ~n22216;
  assign n22218 = ~n22210 & ~n22217;
  assign n22219 = ~n22073 & n22218;
  assign n22220 = n22073 & ~n22218;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = pi276 & ~n21129;
  assign n22223 = pi135 & n22222;
  assign n22224 = ~n21120 & ~n21122;
  assign n22225 = ~n22223 & ~n22224;
  assign n22226 = pi275 & ~n22225;
  assign n22227 = pi136 & n22226;
  assign n22228 = pi137 & pi275;
  assign n22229 = ~n21121 & ~n22224;
  assign n22230 = ~n22223 & n22229;
  assign n22231 = ~n21138 & ~n22230;
  assign n22232 = ~n22228 & ~n22231;
  assign n22233 = ~n22227 & n22232;
  assign n22234 = ~n22227 & ~n22231;
  assign n22235 = n22228 & ~n22234;
  assign n22236 = ~n22233 & ~n22235;
  assign n22237 = ~n22221 & ~n22236;
  assign n22238 = ~n22073 & ~n22218;
  assign n22239 = n22073 & n22218;
  assign n22240 = ~n22238 & ~n22239;
  assign n22241 = n22228 & ~n22231;
  assign n22242 = ~n22227 & n22241;
  assign n22243 = ~n22228 & ~n22234;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = ~n22240 & ~n22244;
  assign n22246 = ~n22237 & ~n22245;
  assign n22247 = n21142 & ~n21167;
  assign n22248 = ~n21142 & n21167;
  assign n22249 = ~n21158 & ~n22248;
  assign n22250 = ~n22247 & ~n22249;
  assign n22251 = n22246 & ~n22250;
  assign n22252 = ~n22246 & n22250;
  assign n22253 = ~n22251 & ~n22252;
  assign n22254 = pi138 & pi274;
  assign n22255 = n21181 & ~n21187;
  assign n22256 = ~n21186 & ~n22255;
  assign n22257 = n22254 & ~n22256;
  assign n22258 = ~n21181 & ~n21186;
  assign n22259 = ~n21187 & ~n22258;
  assign n22260 = ~n22254 & ~n22259;
  assign n22261 = ~n22257 & ~n22260;
  assign n22262 = ~n22253 & ~n22261;
  assign n22263 = n22246 & n22250;
  assign n22264 = ~n22246 & ~n22250;
  assign n22265 = ~n22263 & ~n22264;
  assign n22266 = ~n22254 & ~n22256;
  assign n22267 = n22254 & ~n22259;
  assign n22268 = ~n22266 & ~n22267;
  assign n22269 = ~n22265 & ~n22268;
  assign n22270 = ~n22262 & ~n22269;
  assign n22271 = ~n22072 & ~n22270;
  assign n22272 = n22072 & n22270;
  assign n22273 = ~n22271 & ~n22272;
  assign n22274 = pi273 & ~n21188;
  assign n22275 = pi138 & n22274;
  assign n22276 = ~n21179 & ~n21181;
  assign n22277 = ~n21180 & ~n22276;
  assign n22278 = ~n22275 & n22277;
  assign n22279 = pi140 & pi272;
  assign n22280 = ~n22275 & ~n22276;
  assign n22281 = pi272 & ~n22280;
  assign n22282 = pi139 & n22281;
  assign n22283 = n21198 & ~n22282;
  assign n22284 = n22279 & ~n22283;
  assign n22285 = ~n22278 & n22284;
  assign n22286 = ~n22278 & ~n22283;
  assign n22287 = ~n22279 & ~n22286;
  assign n22288 = ~n22285 & ~n22287;
  assign n22289 = ~n22273 & ~n22288;
  assign n22290 = ~n22072 & n22270;
  assign n22291 = n22072 & ~n22270;
  assign n22292 = ~n22290 & ~n22291;
  assign n22293 = ~n22279 & ~n22283;
  assign n22294 = ~n22278 & n22293;
  assign n22295 = n22279 & ~n22286;
  assign n22296 = ~n22294 & ~n22295;
  assign n22297 = ~n22292 & ~n22296;
  assign n22298 = ~n22289 & ~n22297;
  assign n22299 = ~n21201 & ~n21202;
  assign n22300 = n21201 & n21202;
  assign n22301 = ~n21221 & ~n22300;
  assign n22302 = ~n22299 & ~n22301;
  assign n22303 = n22298 & n22302;
  assign n22304 = ~n22298 & ~n22302;
  assign n22305 = ~n22303 & ~n22304;
  assign n22306 = pi141 & pi271;
  assign n22307 = n21241 & ~n21247;
  assign n22308 = ~n21246 & ~n22307;
  assign n22309 = n22306 & ~n22308;
  assign n22310 = ~n21241 & ~n21246;
  assign n22311 = ~n21247 & ~n22310;
  assign n22312 = ~n22306 & ~n22311;
  assign n22313 = ~n22309 & ~n22312;
  assign n22314 = ~n22305 & ~n22313;
  assign n22315 = n22298 & ~n22302;
  assign n22316 = ~n22298 & n22302;
  assign n22317 = ~n22315 & ~n22316;
  assign n22318 = ~n22306 & ~n22308;
  assign n22319 = n22306 & ~n22311;
  assign n22320 = ~n22318 & ~n22319;
  assign n22321 = ~n22317 & ~n22320;
  assign n22322 = ~n22314 & ~n22321;
  assign n22323 = ~n22071 & ~n22322;
  assign n22324 = n22071 & n22322;
  assign n22325 = ~n22323 & ~n22324;
  assign n22326 = pi270 & ~n21248;
  assign n22327 = pi141 & n22326;
  assign n22328 = ~n21239 & ~n21241;
  assign n22329 = ~n21240 & ~n22328;
  assign n22330 = ~n22327 & n22329;
  assign n22331 = pi143 & pi269;
  assign n22332 = ~n22327 & ~n22328;
  assign n22333 = pi269 & ~n22332;
  assign n22334 = pi142 & n22333;
  assign n22335 = n21258 & ~n22334;
  assign n22336 = n22331 & ~n22335;
  assign n22337 = ~n22330 & n22336;
  assign n22338 = ~n22330 & ~n22335;
  assign n22339 = ~n22331 & ~n22338;
  assign n22340 = ~n22337 & ~n22339;
  assign n22341 = ~n22325 & ~n22340;
  assign n22342 = ~n22071 & n22322;
  assign n22343 = n22071 & ~n22322;
  assign n22344 = ~n22342 & ~n22343;
  assign n22345 = ~n22331 & ~n22335;
  assign n22346 = ~n22330 & n22345;
  assign n22347 = n22331 & ~n22338;
  assign n22348 = ~n22346 & ~n22347;
  assign n22349 = ~n22344 & ~n22348;
  assign n22350 = ~n22341 & ~n22349;
  assign n22351 = ~n21262 & ~n21287;
  assign n22352 = n21262 & n21287;
  assign n22353 = ~n21281 & ~n22352;
  assign n22354 = ~n22351 & ~n22353;
  assign n22355 = n22350 & ~n22354;
  assign n22356 = ~n22350 & n22354;
  assign n22357 = ~n22355 & ~n22356;
  assign n22358 = pi144 & pi268;
  assign n22359 = n21301 & ~n21306;
  assign n22360 = ~n21307 & ~n22359;
  assign n22361 = n22358 & ~n22360;
  assign n22362 = ~n21301 & ~n21307;
  assign n22363 = ~n21306 & ~n22362;
  assign n22364 = ~n22358 & ~n22363;
  assign n22365 = ~n22361 & ~n22364;
  assign n22366 = ~n22357 & ~n22365;
  assign n22367 = n22350 & n22354;
  assign n22368 = ~n22350 & ~n22354;
  assign n22369 = ~n22367 & ~n22368;
  assign n22370 = ~n22358 & ~n22360;
  assign n22371 = n22358 & ~n22363;
  assign n22372 = ~n22370 & ~n22371;
  assign n22373 = ~n22369 & ~n22372;
  assign n22374 = ~n22366 & ~n22373;
  assign n22375 = ~n22070 & n22374;
  assign n22376 = n22070 & ~n22374;
  assign n22377 = ~n22375 & ~n22376;
  assign n22378 = pi267 & ~n21308;
  assign n22379 = pi144 & n22378;
  assign n22380 = ~n21299 & ~n21301;
  assign n22381 = ~n22379 & ~n22380;
  assign n22382 = pi266 & ~n22381;
  assign n22383 = pi145 & n22382;
  assign n22384 = pi146 & pi266;
  assign n22385 = ~n21300 & ~n22380;
  assign n22386 = ~n22379 & n22385;
  assign n22387 = ~n21317 & ~n22386;
  assign n22388 = ~n22384 & ~n22387;
  assign n22389 = ~n22383 & n22388;
  assign n22390 = ~n22383 & ~n22387;
  assign n22391 = n22384 & ~n22390;
  assign n22392 = ~n22389 & ~n22391;
  assign n22393 = ~n22377 & ~n22392;
  assign n22394 = ~n22070 & ~n22374;
  assign n22395 = n22070 & n22374;
  assign n22396 = ~n22394 & ~n22395;
  assign n22397 = n22384 & ~n22387;
  assign n22398 = ~n22383 & n22397;
  assign n22399 = ~n22384 & ~n22390;
  assign n22400 = ~n22398 & ~n22399;
  assign n22401 = ~n22396 & ~n22400;
  assign n22402 = ~n22393 & ~n22401;
  assign n22403 = ~n21321 & ~n21346;
  assign n22404 = n21321 & n21346;
  assign n22405 = ~n21340 & ~n22404;
  assign n22406 = ~n22403 & ~n22405;
  assign n22407 = n22402 & ~n22406;
  assign n22408 = ~n22402 & n22406;
  assign n22409 = ~n22407 & ~n22408;
  assign n22410 = pi147 & pi265;
  assign n22411 = n21362 & ~n21367;
  assign n22412 = ~n21368 & ~n22411;
  assign n22413 = n22410 & ~n22412;
  assign n22414 = ~n21362 & ~n21368;
  assign n22415 = ~n21367 & ~n22414;
  assign n22416 = ~n22410 & ~n22415;
  assign n22417 = ~n22413 & ~n22416;
  assign n22418 = ~n22409 & ~n22417;
  assign n22419 = n22402 & n22406;
  assign n22420 = ~n22402 & ~n22406;
  assign n22421 = ~n22419 & ~n22420;
  assign n22422 = ~n22410 & ~n22412;
  assign n22423 = n22410 & ~n22415;
  assign n22424 = ~n22422 & ~n22423;
  assign n22425 = ~n22421 & ~n22424;
  assign n22426 = ~n22418 & ~n22425;
  assign n22427 = ~n22069 & n22426;
  assign n22428 = n22069 & ~n22426;
  assign n22429 = ~n22427 & ~n22428;
  assign n22430 = pi264 & ~n21369;
  assign n22431 = pi147 & n22430;
  assign n22432 = ~n21360 & ~n21362;
  assign n22433 = ~n22431 & ~n22432;
  assign n22434 = pi263 & ~n22433;
  assign n22435 = pi148 & n22434;
  assign n22436 = pi149 & pi263;
  assign n22437 = ~n21361 & ~n22432;
  assign n22438 = ~n22431 & n22437;
  assign n22439 = n21381 & ~n22438;
  assign n22440 = ~n22436 & ~n22439;
  assign n22441 = ~n22435 & n22440;
  assign n22442 = ~n22435 & ~n22439;
  assign n22443 = n22436 & ~n22442;
  assign n22444 = ~n22441 & ~n22443;
  assign n22445 = ~n22429 & ~n22444;
  assign n22446 = ~n22069 & ~n22426;
  assign n22447 = n22069 & n22426;
  assign n22448 = ~n22446 & ~n22447;
  assign n22449 = n22436 & ~n22439;
  assign n22450 = ~n22435 & n22449;
  assign n22451 = ~n22436 & ~n22442;
  assign n22452 = ~n22450 & ~n22451;
  assign n22453 = ~n22448 & ~n22452;
  assign n22454 = ~n22445 & ~n22453;
  assign n22455 = n21385 & ~n21398;
  assign n22456 = ~n21385 & n21398;
  assign n22457 = ~n21389 & ~n22456;
  assign n22458 = ~n22455 & ~n22457;
  assign n22459 = n22454 & n22458;
  assign n22460 = ~n22454 & ~n22458;
  assign n22461 = ~n22459 & ~n22460;
  assign n22462 = pi150 & pi262;
  assign n22463 = n21421 & ~n21422;
  assign n22464 = ~n21423 & ~n22463;
  assign n22465 = n22462 & ~n22464;
  assign n22466 = ~n21421 & ~n21423;
  assign n22467 = ~n21422 & ~n22466;
  assign n22468 = ~n22462 & ~n22467;
  assign n22469 = ~n22465 & ~n22468;
  assign n22470 = ~n22461 & ~n22469;
  assign n22471 = n22454 & ~n22458;
  assign n22472 = ~n22454 & n22458;
  assign n22473 = ~n22471 & ~n22472;
  assign n22474 = ~n22462 & ~n22464;
  assign n22475 = n22462 & ~n22467;
  assign n22476 = ~n22474 & ~n22475;
  assign n22477 = ~n22473 & ~n22476;
  assign n22478 = ~n22470 & ~n22477;
  assign n22479 = ~n22068 & n22478;
  assign n22480 = n22068 & ~n22478;
  assign n22481 = ~n22479 & ~n22480;
  assign n22482 = pi152 & pi260;
  assign n22483 = pi151 & ~n20982;
  assign n22484 = n21426 & n22483;
  assign n22485 = pi151 & pi260;
  assign n22486 = ~n21426 & ~n22483;
  assign n22487 = n22485 & ~n22486;
  assign n22488 = ~n22484 & ~n22487;
  assign n22489 = n22482 & ~n22488;
  assign n22490 = ~n22484 & ~n22485;
  assign n22491 = ~n22486 & ~n22490;
  assign n22492 = ~n22482 & ~n22491;
  assign n22493 = ~n22489 & ~n22492;
  assign n22494 = ~n22481 & ~n22493;
  assign n22495 = ~n22068 & ~n22478;
  assign n22496 = n22068 & n22478;
  assign n22497 = ~n22495 & ~n22496;
  assign n22498 = ~n22482 & ~n22488;
  assign n22499 = n22482 & ~n22491;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = ~n22497 & ~n22500;
  assign n22502 = ~n22494 & ~n22501;
  assign n22503 = n21431 & n21439;
  assign n22504 = ~n21431 & ~n21439;
  assign n22505 = ~n21429 & ~n22504;
  assign n22506 = ~n22503 & ~n22505;
  assign n22507 = n22502 & ~n22506;
  assign n22508 = ~n22502 & n22506;
  assign n22509 = ~n22507 & ~n22508;
  assign n22510 = ~n22503 & ~n22504;
  assign n22511 = ~n21429 & ~n22510;
  assign n22512 = n21431 & ~n21439;
  assign n22513 = ~n21431 & n21439;
  assign n22514 = ~n22512 & ~n22513;
  assign n22515 = ~n21462 & ~n22514;
  assign n22516 = ~n22511 & ~n22515;
  assign n22517 = pi258 & ~n22516;
  assign n22518 = pi153 & n22517;
  assign n22519 = pi154 & pi258;
  assign n22520 = n22518 & ~n22519;
  assign n22521 = ~n22518 & n22519;
  assign n22522 = pi153 & n22521;
  assign n22523 = ~n22520 & ~n22522;
  assign n22524 = pi259 & ~n22523;
  assign n22525 = ~n22518 & ~n22519;
  assign n22526 = n22518 & n22519;
  assign n22527 = ~n22525 & ~n22526;
  assign n22528 = ~pi259 & ~n22527;
  assign n22529 = ~pi153 & n22525;
  assign n22530 = ~n22528 & ~n22529;
  assign n22531 = ~n22524 & n22530;
  assign n22532 = ~n22509 & ~n22531;
  assign n22533 = n22502 & n22506;
  assign n22534 = ~n22502 & ~n22506;
  assign n22535 = ~n22533 & ~n22534;
  assign n22536 = pi153 & n22525;
  assign n22537 = ~n22526 & ~n22536;
  assign n22538 = pi259 & ~n22537;
  assign n22539 = ~n22520 & ~n22521;
  assign n22540 = ~pi259 & ~n22539;
  assign n22541 = ~pi153 & n22521;
  assign n22542 = ~n22540 & ~n22541;
  assign n22543 = ~n22538 & n22542;
  assign n22544 = ~n22535 & ~n22543;
  assign n22545 = ~n22532 & ~n22544;
  assign n22546 = n21471 & ~n22545;
  assign n22547 = pi258 & ~n22510;
  assign n22548 = pi153 & n22547;
  assign n22549 = ~n21430 & ~n22514;
  assign n22550 = ~n22548 & ~n22549;
  assign n22551 = ~n21462 & ~n22550;
  assign n22552 = pi258 & ~n22514;
  assign n22553 = pi153 & n22552;
  assign n22554 = ~n21430 & ~n22510;
  assign n22555 = ~n22553 & ~n22554;
  assign n22556 = ~n21429 & ~n22555;
  assign n22557 = ~n22551 & ~n22556;
  assign n22558 = ~n21471 & n22545;
  assign n22559 = n22557 & n22558;
  assign n22560 = ~n22546 & ~n22559;
  assign n22561 = ~n21446 & ~n22560;
  assign n22562 = ~n21471 & ~n22545;
  assign n22563 = n21471 & n22545;
  assign n22564 = ~n22557 & n22563;
  assign n22565 = ~n22562 & ~n22564;
  assign n22566 = n21446 & ~n22565;
  assign n22567 = ~n21471 & ~n22557;
  assign n22568 = n21471 & n22557;
  assign n22569 = ~n22567 & ~n22568;
  assign n22570 = ~n22545 & ~n22569;
  assign n22571 = ~n22566 & ~n22570;
  assign n22572 = ~n22561 & n22571;
  assign n22573 = pi322 & ~n22572;
  assign n22574 = ~n21471 & n22557;
  assign n22575 = n21471 & ~n22557;
  assign n22576 = ~n22574 & ~n22575;
  assign n22577 = n21446 & ~n22576;
  assign n22578 = ~n21446 & ~n22569;
  assign n22579 = ~n22577 & ~n22578;
  assign n22580 = pi323 & ~n22579;
  assign n22581 = ~n22573 & ~n22580;
  assign n22582 = n21446 & n22574;
  assign n22583 = ~n22578 & ~n22582;
  assign n22584 = ~n22545 & ~n22583;
  assign n22585 = n21446 & ~n22557;
  assign n22586 = n22563 & n22585;
  assign n22587 = ~n22584 & ~n22586;
  assign n22588 = pi323 & ~n22587;
  assign n22589 = pi322 & n22588;
  assign n22590 = ~n22581 & ~n22589;
  assign n22591 = pi325 & n19557;
  assign n22592 = pi324 & n19970;
  assign n22593 = n22591 & n22592;
  assign n22594 = ~n22591 & ~n22592;
  assign n22595 = ~n22593 & ~n22594;
  assign n22596 = ~n22590 & ~n22595;
  assign n22597 = ~n22591 & n22592;
  assign n22598 = n22591 & ~n22592;
  assign n22599 = ~n22597 & ~n22598;
  assign n22600 = ~n22589 & ~n22599;
  assign n22601 = ~n22581 & n22600;
  assign n22602 = ~n22596 & ~n22601;
  assign n22603 = ~n22067 & ~n22602;
  assign n22604 = ~n22060 & ~n22064;
  assign n22605 = n22060 & n22064;
  assign n22606 = ~n22604 & ~n22605;
  assign n22607 = ~n22590 & ~n22599;
  assign n22608 = ~n22589 & ~n22595;
  assign n22609 = ~n22581 & n22608;
  assign n22610 = ~n22607 & ~n22609;
  assign n22611 = ~n22606 & ~n22610;
  assign n22612 = ~n22603 & ~n22611;
  assign n22613 = ~n20967 & n21495;
  assign n22614 = ~n20963 & ~n21490;
  assign n22615 = n20963 & n21490;
  assign n22616 = ~n22614 & ~n22615;
  assign n22617 = n20971 & ~n22616;
  assign n22618 = n20963 & ~n21490;
  assign n22619 = ~n20963 & n21490;
  assign n22620 = ~n22618 & ~n22619;
  assign n22621 = ~n20971 & ~n22620;
  assign n22622 = ~n22617 & ~n22621;
  assign n22623 = n20967 & ~n21495;
  assign n22624 = ~n22622 & ~n22623;
  assign n22625 = ~n22613 & ~n22624;
  assign n22626 = n22612 & n22625;
  assign n22627 = ~n22612 & ~n22625;
  assign n22628 = ~n22626 & ~n22627;
  assign n22629 = pi327 & n18461;
  assign n22630 = pi326 & n19539;
  assign n22631 = n22629 & n22630;
  assign n22632 = ~n22629 & ~n22630;
  assign n22633 = ~n22631 & ~n22632;
  assign n22634 = ~n22628 & ~n22633;
  assign n22635 = ~n22612 & n22625;
  assign n22636 = n22612 & ~n22625;
  assign n22637 = ~n22635 & ~n22636;
  assign n22638 = ~n22629 & n22630;
  assign n22639 = n22629 & ~n22630;
  assign n22640 = ~n22638 & ~n22639;
  assign n22641 = ~n22637 & ~n22640;
  assign n22642 = ~n22634 & ~n22641;
  assign n22643 = ~n22054 & ~n22642;
  assign n22644 = n22047 & n22051;
  assign n22645 = ~n22047 & ~n22051;
  assign n22646 = ~n22644 & ~n22645;
  assign n22647 = ~n22633 & ~n22637;
  assign n22648 = ~n22628 & ~n22640;
  assign n22649 = ~n22647 & ~n22648;
  assign n22650 = ~n22646 & ~n22649;
  assign n22651 = ~n22643 & ~n22650;
  assign n22652 = ~n22032 & n22651;
  assign n22653 = n22032 & ~n22651;
  assign n22654 = ~n22652 & ~n22653;
  assign n22655 = pi330 & n11711;
  assign n22656 = ~n21571 & ~n21578;
  assign n22657 = ~n21567 & n22656;
  assign n22658 = ~n22655 & ~n22657;
  assign n22659 = n20933 & n22658;
  assign n22660 = n21567 & ~n22656;
  assign n22661 = n22655 & ~n22660;
  assign n22662 = ~n20933 & n22661;
  assign n22663 = ~n22659 & ~n22662;
  assign n22664 = ~n21978 & ~n22663;
  assign n22665 = n20933 & n22661;
  assign n22666 = ~n20933 & n22658;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = ~n21968 & ~n22667;
  assign n22669 = ~n22655 & ~n22656;
  assign n22670 = n21567 & n22669;
  assign n22671 = n22655 & n22656;
  assign n22672 = ~n21567 & n22671;
  assign n22673 = ~n22670 & ~n22672;
  assign n22674 = ~n22668 & n22673;
  assign n22675 = ~n22664 & n22674;
  assign n22676 = pi329 & n12917;
  assign n22677 = ~n22675 & n22676;
  assign n22678 = n22675 & ~n22676;
  assign n22679 = ~n22677 & ~n22678;
  assign n22680 = ~n22654 & ~n22679;
  assign n22681 = n22032 & n22651;
  assign n22682 = ~n22032 & ~n22651;
  assign n22683 = ~n22681 & ~n22682;
  assign n22684 = n22675 & n22676;
  assign n22685 = ~n22675 & ~n22676;
  assign n22686 = ~n22684 & ~n22685;
  assign n22687 = ~n22683 & ~n22686;
  assign n22688 = ~n22680 & ~n22687;
  assign n22689 = ~n22031 & ~n22688;
  assign n22690 = n22024 & n22028;
  assign n22691 = ~n22024 & ~n22028;
  assign n22692 = ~n22690 & ~n22691;
  assign n22693 = ~n22679 & ~n22683;
  assign n22694 = ~n22654 & ~n22686;
  assign n22695 = ~n22693 & ~n22694;
  assign n22696 = ~n22692 & ~n22695;
  assign n22697 = ~n22689 & ~n22696;
  assign n22698 = ~n22004 & n22697;
  assign n22699 = n22004 & ~n22697;
  assign n22700 = ~n22698 & ~n22699;
  assign n22701 = pi333 & n10561;
  assign n22702 = pi332 & n11366;
  assign n22703 = n21603 & ~n21994;
  assign n22704 = ~n21991 & ~n22703;
  assign n22705 = ~n22702 & ~n22704;
  assign n22706 = n11366 & ~n22703;
  assign n22707 = pi332 & n22706;
  assign n22708 = ~n21991 & n22707;
  assign n22709 = ~n22705 & ~n22708;
  assign n22710 = n22701 & ~n22709;
  assign n22711 = ~n22701 & n22709;
  assign n22712 = ~n22710 & ~n22711;
  assign n22713 = ~n22700 & ~n22712;
  assign n22714 = n22004 & n22697;
  assign n22715 = ~n22004 & ~n22697;
  assign n22716 = ~n22714 & ~n22715;
  assign n22717 = ~n22701 & ~n22709;
  assign n22718 = n22701 & n22709;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = ~n22716 & ~n22719;
  assign n22721 = ~n22713 & ~n22720;
  assign n22722 = ~n22003 & ~n22721;
  assign n22723 = n21985 & n22000;
  assign n22724 = ~n21985 & ~n22000;
  assign n22725 = ~n22723 & ~n22724;
  assign n22726 = ~n22712 & ~n22716;
  assign n22727 = ~n22700 & ~n22719;
  assign n22728 = ~n22726 & ~n22727;
  assign n22729 = ~n22725 & ~n22728;
  assign n22730 = ~n22722 & ~n22729;
  assign n22731 = ~n20873 & n20891;
  assign n22732 = n20873 & ~n20891;
  assign n22733 = n21665 & ~n22732;
  assign n22734 = ~n22731 & ~n22733;
  assign n22735 = n22730 & n22734;
  assign n22736 = ~n22730 & ~n22734;
  assign n22737 = ~n22735 & ~n22736;
  assign n22738 = pi335 & n6556;
  assign n22739 = ~n21630 & ~n21653;
  assign n22740 = ~n21660 & n22739;
  assign n22741 = ~n21651 & ~n21653;
  assign n22742 = ~n21613 & n22741;
  assign n22743 = ~n21652 & ~n22742;
  assign n22744 = ~n22740 & n22743;
  assign n22745 = pi334 & n9205;
  assign n22746 = n22744 & ~n22745;
  assign n22747 = n9205 & ~n22744;
  assign n22748 = pi334 & n22747;
  assign n22749 = ~n22746 & ~n22748;
  assign n22750 = ~n22738 & n22749;
  assign n22751 = n22738 & ~n22749;
  assign n22752 = ~n22750 & ~n22751;
  assign n22753 = pi336 & n5973;
  assign n22754 = pi336 & n21681;
  assign n22755 = ~n20880 & ~n21674;
  assign n22756 = ~n22754 & ~n22755;
  assign n22757 = n5732 & ~n22756;
  assign n22758 = pi336 & n22757;
  assign n22759 = n20891 & ~n21939;
  assign n22760 = ~n20891 & ~n21929;
  assign n22761 = ~n22759 & ~n22760;
  assign n22762 = pi336 & n5732;
  assign n22763 = n22756 & ~n22762;
  assign n22764 = ~n22761 & ~n22763;
  assign n22765 = ~n22758 & ~n22764;
  assign n22766 = n22753 & n22765;
  assign n22767 = ~n22753 & ~n22765;
  assign n22768 = ~n22766 & ~n22767;
  assign n22769 = ~n22752 & ~n22768;
  assign n22770 = n22738 & n22749;
  assign n22771 = ~n22738 & ~n22749;
  assign n22772 = ~n22770 & ~n22771;
  assign n22773 = ~n22753 & n22765;
  assign n22774 = n22753 & ~n22765;
  assign n22775 = ~n22773 & ~n22774;
  assign n22776 = ~n22772 & ~n22775;
  assign n22777 = ~n22769 & ~n22776;
  assign n22778 = ~n22737 & ~n22777;
  assign n22779 = n22730 & ~n22734;
  assign n22780 = ~n22730 & n22734;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = ~n22768 & ~n22772;
  assign n22783 = ~n22752 & ~n22775;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = ~n22781 & ~n22784;
  assign n22786 = ~n22778 & ~n22785;
  assign n22787 = ~n21965 & n22786;
  assign n22788 = n21965 & ~n22786;
  assign n22789 = ~n22787 & ~n22788;
  assign n22790 = pi339 & n5257;
  assign n22791 = pi338 & n5714;
  assign n22792 = n21708 & ~n21955;
  assign n22793 = ~n21952 & ~n22792;
  assign n22794 = ~n22791 & ~n22793;
  assign n22795 = n5714 & ~n22792;
  assign n22796 = pi338 & n22795;
  assign n22797 = ~n21952 & n22796;
  assign n22798 = ~n22794 & ~n22797;
  assign n22799 = n22790 & ~n22798;
  assign n22800 = ~n22790 & n22798;
  assign n22801 = ~n22799 & ~n22800;
  assign n22802 = ~n22789 & ~n22801;
  assign n22803 = n21965 & n22786;
  assign n22804 = ~n21965 & ~n22786;
  assign n22805 = ~n22803 & ~n22804;
  assign n22806 = ~n22790 & ~n22798;
  assign n22807 = n22790 & n22798;
  assign n22808 = ~n22806 & ~n22807;
  assign n22809 = ~n22805 & ~n22808;
  assign n22810 = ~n22802 & ~n22809;
  assign n22811 = ~n21964 & ~n22810;
  assign n22812 = n21946 & n21961;
  assign n22813 = ~n21946 & ~n21961;
  assign n22814 = ~n22812 & ~n22813;
  assign n22815 = ~n22801 & ~n22805;
  assign n22816 = ~n22789 & ~n22808;
  assign n22817 = ~n22815 & ~n22816;
  assign n22818 = ~n22814 & ~n22817;
  assign n22819 = ~n22811 & ~n22818;
  assign n22820 = ~n20828 & n20852;
  assign n22821 = n20828 & ~n20852;
  assign n22822 = n21763 & ~n22821;
  assign n22823 = ~n22820 & ~n22822;
  assign n22824 = n22819 & n22823;
  assign n22825 = ~n22819 & ~n22823;
  assign n22826 = ~n22824 & ~n22825;
  assign n22827 = pi341 & n2887;
  assign n22828 = ~n21735 & ~n21751;
  assign n22829 = ~n21758 & n22828;
  assign n22830 = ~n21749 & ~n21751;
  assign n22831 = ~n21718 & n22830;
  assign n22832 = ~n21750 & ~n22831;
  assign n22833 = ~n22829 & n22832;
  assign n22834 = pi340 & n4596;
  assign n22835 = n22833 & ~n22834;
  assign n22836 = n4596 & ~n22833;
  assign n22837 = pi340 & n22836;
  assign n22838 = ~n22835 & ~n22837;
  assign n22839 = ~n22827 & n22838;
  assign n22840 = n22827 & ~n22838;
  assign n22841 = ~n22839 & ~n22840;
  assign n22842 = pi342 & n2464;
  assign n22843 = n20852 & ~n21906;
  assign n22844 = ~n20852 & ~n21896;
  assign n22845 = ~n22843 & ~n22844;
  assign n22846 = n19400 & ~n20841;
  assign n22847 = ~n19400 & ~n20831;
  assign n22848 = ~n22846 & ~n22847;
  assign n22849 = ~n21769 & ~n22848;
  assign n22850 = ~n21772 & ~n22849;
  assign n22851 = ~n21768 & n22850;
  assign n22852 = ~n22845 & ~n22851;
  assign n22853 = n21768 & ~n22850;
  assign n22854 = ~n22852 & ~n22853;
  assign n22855 = n22842 & n22854;
  assign n22856 = ~n22842 & ~n22854;
  assign n22857 = ~n22855 & ~n22856;
  assign n22858 = ~n22841 & ~n22857;
  assign n22859 = n22827 & n22838;
  assign n22860 = ~n22827 & ~n22838;
  assign n22861 = ~n22859 & ~n22860;
  assign n22862 = ~n22842 & n22854;
  assign n22863 = n22842 & ~n22854;
  assign n22864 = ~n22862 & ~n22863;
  assign n22865 = ~n22861 & ~n22864;
  assign n22866 = ~n22858 & ~n22865;
  assign n22867 = ~n22826 & ~n22866;
  assign n22868 = n22819 & ~n22823;
  assign n22869 = ~n22819 & n22823;
  assign n22870 = ~n22868 & ~n22869;
  assign n22871 = ~n22857 & ~n22861;
  assign n22872 = ~n22841 & ~n22864;
  assign n22873 = ~n22871 & ~n22872;
  assign n22874 = ~n22870 & ~n22873;
  assign n22875 = ~n22867 & ~n22874;
  assign n22876 = ~n21926 & n22875;
  assign n22877 = n21926 & ~n22875;
  assign n22878 = ~n22876 & ~n22877;
  assign n22879 = pi345 & n1442;
  assign n22880 = n21808 & ~n21827;
  assign n22881 = ~n21824 & ~n22880;
  assign n22882 = n1729 & n22881;
  assign n22883 = pi344 & n22882;
  assign n22884 = pi344 & n1729;
  assign n22885 = ~n22881 & ~n22884;
  assign n22886 = ~n22883 & ~n22885;
  assign n22887 = n22879 & ~n22886;
  assign n22888 = ~n22879 & n22886;
  assign n22889 = ~n22887 & ~n22888;
  assign n22890 = ~n22878 & ~n22889;
  assign n22891 = n21926 & n22875;
  assign n22892 = ~n21926 & ~n22875;
  assign n22893 = ~n22891 & ~n22892;
  assign n22894 = ~n22879 & ~n22886;
  assign n22895 = n22879 & n22886;
  assign n22896 = ~n22894 & ~n22895;
  assign n22897 = ~n22893 & ~n22896;
  assign n22898 = ~n22890 & ~n22897;
  assign n22899 = ~n21925 & ~n22898;
  assign n22900 = n21913 & n21922;
  assign n22901 = ~n21913 & ~n21922;
  assign n22902 = ~n22900 & ~n22901;
  assign n22903 = ~n22889 & ~n22893;
  assign n22904 = ~n22878 & ~n22896;
  assign n22905 = ~n22903 & ~n22904;
  assign n22906 = ~n22902 & ~n22905;
  assign n22907 = ~n22899 & ~n22906;
  assign n22908 = ~n21893 & n22907;
  assign n22909 = n21893 & ~n22907;
  assign n22910 = ~n22908 & ~n22909;
  assign n22911 = pi258 & ~n21852;
  assign n22912 = pi128 & n22911;
  assign n22913 = pi347 & n22912;
  assign n22914 = pi347 & ~n1154;
  assign n22915 = ~n22913 & ~n22914;
  assign n22916 = n22913 & n22914;
  assign n22917 = ~n22915 & ~n22916;
  assign n22918 = n1156 & ~n22917;
  assign n22919 = pi348 & n22918;
  assign n22920 = pi348 & n1156;
  assign n22921 = n22913 & ~n22914;
  assign n22922 = ~n22913 & n22914;
  assign n22923 = ~n22921 & ~n22922;
  assign n22924 = ~n22920 & ~n22923;
  assign n22925 = ~n22919 & ~n22924;
  assign n22926 = ~n22910 & ~n22925;
  assign n22927 = ~n21893 & ~n22907;
  assign n22928 = n21893 & n22907;
  assign n22929 = ~n22927 & ~n22928;
  assign n22930 = n1156 & ~n22923;
  assign n22931 = pi348 & n22930;
  assign n22932 = ~n22917 & ~n22920;
  assign n22933 = ~n22931 & ~n22932;
  assign n22934 = ~n22929 & ~n22933;
  assign n22935 = ~n22926 & ~n22934;
  assign n22936 = ~n20814 & ~n21872;
  assign n22937 = ~n21861 & ~n22936;
  assign n22938 = ~n20813 & n21872;
  assign n22939 = ~n20810 & n22938;
  assign n22940 = ~n22937 & ~n22939;
  assign n22941 = n22935 & ~n22940;
  assign n22942 = ~n22935 & n22940;
  assign n22943 = ~n22941 & ~n22942;
  assign n22944 = pi130 & pi297;
  assign n22945 = ~pi129 & ~n22944;
  assign n22946 = pi297 & ~n12284;
  assign n22947 = ~n1514 & n22946;
  assign n22948 = n20805 & ~n22947;
  assign n22949 = ~n22945 & ~n22948;
  assign n22950 = n20302 & ~n22949;
  assign n22951 = ~pi130 & n20805;
  assign n22952 = ~pi129 & n22951;
  assign n22953 = pi130 & ~n20805;
  assign n22954 = pi129 & n22953;
  assign n22955 = ~n22952 & ~n22954;
  assign n22956 = pi128 & ~n22955;
  assign n22957 = ~n20302 & n20805;
  assign n22958 = pi130 & n22957;
  assign n22959 = ~pi130 & ~n20805;
  assign n22960 = pi129 & n22959;
  assign n22961 = ~n22958 & ~n22960;
  assign n22962 = ~pi128 & ~n22961;
  assign n22963 = pi129 & n20805;
  assign n22964 = ~pi129 & ~n20805;
  assign n22965 = ~n22963 & ~n22964;
  assign n22966 = ~n20302 & ~n22965;
  assign n22967 = pi130 & n22966;
  assign n22968 = ~n22962 & ~n22967;
  assign n22969 = ~n22956 & n22968;
  assign n22970 = pi297 & ~n22969;
  assign n22971 = ~n22950 & ~n22970;
  assign n22972 = n20769 & n20790;
  assign n22973 = ~n20769 & ~n20790;
  assign n22974 = ~n22972 & ~n22973;
  assign n22975 = n20773 & ~n20791;
  assign n22976 = ~n22974 & ~n22975;
  assign n22977 = n1515 & ~n20773;
  assign n22978 = pi298 & n22977;
  assign n22979 = ~n22976 & ~n22978;
  assign n22980 = ~n20769 & ~n20787;
  assign n22981 = ~n18847 & n19332;
  assign n22982 = ~n18842 & ~n22981;
  assign n22983 = ~n20782 & ~n22982;
  assign n22984 = n20769 & n20787;
  assign n22985 = ~n22983 & ~n22984;
  assign n22986 = ~n22980 & ~n22985;
  assign n22987 = pi301 & n2183;
  assign n22988 = ~n20748 & ~n20755;
  assign n22989 = ~n20756 & ~n22988;
  assign n22990 = ~n22987 & ~n22989;
  assign n22991 = ~n20751 & ~n20756;
  assign n22992 = ~n20755 & ~n22991;
  assign n22993 = n22987 & ~n22992;
  assign n22994 = ~n22990 & ~n22993;
  assign n22995 = n19282 & n20735;
  assign n22996 = ~n19295 & ~n20710;
  assign n22997 = n1840 & n22996;
  assign n22998 = ~n19294 & ~n20708;
  assign n22999 = n2183 & ~n22998;
  assign n23000 = ~n22997 & ~n22999;
  assign n23001 = pi302 & ~n23000;
  assign n23002 = ~n22995 & ~n23001;
  assign n23003 = ~n20691 & ~n20692;
  assign n23004 = n20691 & n20692;
  assign n23005 = ~n20697 & ~n23004;
  assign n23006 = ~n23003 & ~n23005;
  assign n23007 = pi305 & n4086;
  assign n23008 = ~n20670 & ~n20677;
  assign n23009 = ~n20678 & ~n23008;
  assign n23010 = ~n23007 & ~n23009;
  assign n23011 = ~n20673 & ~n20678;
  assign n23012 = ~n20677 & ~n23011;
  assign n23013 = n23007 & ~n23012;
  assign n23014 = ~n23010 & ~n23013;
  assign n23015 = ~n20604 & ~n20615;
  assign n23016 = n20604 & n20615;
  assign n23017 = ~n20609 & ~n23016;
  assign n23018 = ~n23015 & ~n23017;
  assign n23019 = pi309 & n7044;
  assign n23020 = ~n20582 & ~n20589;
  assign n23021 = ~n20590 & ~n23020;
  assign n23022 = ~n23019 & ~n23021;
  assign n23023 = ~n20585 & ~n20590;
  assign n23024 = ~n20589 & ~n23023;
  assign n23025 = n23019 & ~n23024;
  assign n23026 = ~n23022 & ~n23025;
  assign n23027 = ~n20515 & ~n20516;
  assign n23028 = n20515 & n20516;
  assign n23029 = ~n20521 & ~n23028;
  assign n23030 = ~n23027 & ~n23029;
  assign n23031 = pi313 & n10908;
  assign n23032 = ~n20494 & ~n20501;
  assign n23033 = ~n20502 & ~n23032;
  assign n23034 = ~n23031 & ~n23033;
  assign n23035 = ~n20497 & ~n20502;
  assign n23036 = ~n20501 & ~n23035;
  assign n23037 = n23031 & ~n23036;
  assign n23038 = ~n23034 & ~n23037;
  assign n23039 = ~n20461 & ~n20462;
  assign n23040 = n20461 & n20462;
  assign n23041 = ~n19062 & ~n23040;
  assign n23042 = ~n19056 & n23041;
  assign n23043 = ~n23039 & ~n23042;
  assign n23044 = ~n20401 & ~n20403;
  assign n23045 = ~n20400 & n20403;
  assign n23046 = ~n20397 & n23045;
  assign n23047 = ~n23044 & ~n23046;
  assign n23048 = ~n20438 & ~n23047;
  assign n23049 = ~n20372 & n20383;
  assign n23050 = pi150 & pi152;
  assign n23051 = pi151 & n20320;
  assign n23052 = ~n23050 & ~n23051;
  assign n23053 = pi149 & ~n23052;
  assign n23054 = pi151 & pi153;
  assign n23055 = ~n18926 & ~n23054;
  assign n23056 = pi150 & ~n23055;
  assign n23057 = ~pi151 & ~pi153;
  assign n23058 = pi152 & ~n23057;
  assign n23059 = ~n23056 & ~n23058;
  assign n23060 = ~n23053 & n23059;
  assign n23061 = pi154 & n23060;
  assign n23062 = ~pi154 & ~n23060;
  assign n23063 = ~n23061 & ~n23062;
  assign n23064 = pi153 & ~n23063;
  assign n23065 = pi154 & ~n23060;
  assign n23066 = ~pi154 & n23060;
  assign n23067 = ~n23065 & ~n23066;
  assign n23068 = ~pi153 & ~n23067;
  assign n23069 = ~n23064 & ~n23068;
  assign n23070 = n20347 & ~n20359;
  assign n23071 = ~pi320 & ~n23070;
  assign n23072 = ~n18937 & ~n20347;
  assign n23073 = pi320 & n23070;
  assign n23074 = ~n20362 & ~n23073;
  assign n23075 = ~n23072 & n23074;
  assign n23076 = ~n23071 & n23075;
  assign n23077 = n23069 & ~n23076;
  assign n23078 = ~n20359 & ~n23069;
  assign n23079 = ~pi320 & n20347;
  assign n23080 = n23078 & n23079;
  assign n23081 = ~n23077 & ~n23080;
  assign n23082 = pi321 & ~n23081;
  assign n23083 = n20359 & ~n23069;
  assign n23084 = ~n18937 & n23083;
  assign n23085 = ~pi321 & ~n20367;
  assign n23086 = ~n23084 & ~n23085;
  assign n23087 = n20347 & ~n23086;
  assign n23088 = pi321 & n23069;
  assign n23089 = ~n20359 & ~n23088;
  assign n23090 = ~n20347 & n23089;
  assign n23091 = n18937 & n23090;
  assign n23092 = ~n23087 & ~n23091;
  assign n23093 = pi320 & ~n23092;
  assign n23094 = ~n23082 & ~n23093;
  assign n23095 = ~pi319 & ~n23094;
  assign n23096 = ~n18937 & ~n23094;
  assign n23097 = n18937 & n23094;
  assign n23098 = pi319 & n23097;
  assign n23099 = ~n23096 & ~n23098;
  assign n23100 = ~n17455 & ~n23099;
  assign n23101 = ~n23095 & ~n23100;
  assign n23102 = ~n23049 & ~n23101;
  assign n23103 = ~n20383 & n23094;
  assign n23104 = n20372 & n23103;
  assign n23105 = n20383 & ~n23094;
  assign n23106 = ~n20372 & n23105;
  assign n23107 = ~n23104 & ~n23106;
  assign n23108 = pi319 & ~n23107;
  assign n23109 = ~n20372 & ~n20383;
  assign n23110 = n20372 & n20383;
  assign n23111 = ~n23109 & ~n23110;
  assign n23112 = ~n23094 & ~n23111;
  assign n23113 = n17455 & n23112;
  assign n23114 = ~n23108 & ~n23113;
  assign n23115 = n18937 & ~n23114;
  assign n23116 = ~n20383 & ~n23094;
  assign n23117 = n20372 & n23116;
  assign n23118 = n20372 & ~n20383;
  assign n23119 = n17455 & ~n23118;
  assign n23120 = pi319 & n23119;
  assign n23121 = ~n23049 & ~n23120;
  assign n23122 = n23094 & ~n23121;
  assign n23123 = ~n23117 & ~n23122;
  assign n23124 = ~n18937 & ~n23123;
  assign n23125 = ~pi319 & ~n20372;
  assign n23126 = n20383 & n23094;
  assign n23127 = n23125 & n23126;
  assign n23128 = ~n23124 & ~n23127;
  assign n23129 = ~n23115 & n23128;
  assign n23130 = ~n23102 & n23129;
  assign n23131 = pi318 & n17455;
  assign n23132 = ~n23130 & ~n23131;
  assign n23133 = n17455 & n23130;
  assign n23134 = pi318 & n23133;
  assign n23135 = ~n23132 & ~n23134;
  assign n23136 = n20317 & ~n20388;
  assign n23137 = ~n20391 & ~n23136;
  assign n23138 = n23135 & n23137;
  assign n23139 = ~n23135 & ~n23137;
  assign n23140 = ~n23138 & ~n23139;
  assign n23141 = pi317 & n16985;
  assign n23142 = ~n20400 & ~n20403;
  assign n23143 = ~n23141 & ~n23142;
  assign n23144 = ~n20397 & n23143;
  assign n23145 = ~n20397 & ~n23142;
  assign n23146 = n23141 & ~n23145;
  assign n23147 = ~n23144 & ~n23146;
  assign n23148 = ~n23140 & ~n23147;
  assign n23149 = n23135 & ~n23137;
  assign n23150 = ~n23135 & n23137;
  assign n23151 = ~n23149 & ~n23150;
  assign n23152 = n23141 & ~n23142;
  assign n23153 = ~n20397 & n23152;
  assign n23154 = ~n23141 & ~n23145;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = ~n23151 & ~n23155;
  assign n23157 = ~n23148 & ~n23156;
  assign n23158 = ~pi316 & ~n23157;
  assign n23159 = ~n14618 & ~n23157;
  assign n23160 = n14618 & n23157;
  assign n23161 = pi316 & n23160;
  assign n23162 = ~n23159 & ~n23161;
  assign n23163 = ~n14156 & ~n23162;
  assign n23164 = ~n23158 & ~n23163;
  assign n23165 = ~n23048 & ~n23164;
  assign n23166 = n20438 & n23157;
  assign n23167 = n23047 & n23166;
  assign n23168 = ~n20438 & ~n23157;
  assign n23169 = ~n23047 & n23168;
  assign n23170 = ~n23167 & ~n23169;
  assign n23171 = pi316 & ~n23170;
  assign n23172 = n20438 & ~n23047;
  assign n23173 = ~n20438 & n23047;
  assign n23174 = ~n23172 & ~n23173;
  assign n23175 = ~n23157 & ~n23174;
  assign n23176 = n14156 & n23175;
  assign n23177 = ~n23171 & ~n23176;
  assign n23178 = n14618 & ~n23177;
  assign n23179 = n20438 & ~n23157;
  assign n23180 = n23047 & n23179;
  assign n23181 = n20438 & n23047;
  assign n23182 = n14156 & ~n23181;
  assign n23183 = pi316 & n23182;
  assign n23184 = ~n23048 & ~n23183;
  assign n23185 = n23157 & ~n23184;
  assign n23186 = ~n23180 & ~n23185;
  assign n23187 = ~n14618 & ~n23186;
  assign n23188 = ~pi316 & ~n23047;
  assign n23189 = ~n20438 & n23157;
  assign n23190 = n23188 & n23189;
  assign n23191 = ~n23187 & ~n23190;
  assign n23192 = ~n23178 & n23191;
  assign n23193 = ~n23165 & n23192;
  assign n23194 = n20444 & ~n20447;
  assign n23195 = ~n19051 & ~n20455;
  assign n23196 = n19051 & n20455;
  assign n23197 = n20450 & ~n23196;
  assign n23198 = ~n23195 & ~n23197;
  assign n23199 = ~n20444 & n20447;
  assign n23200 = ~n23198 & ~n23199;
  assign n23201 = ~n23194 & ~n23200;
  assign n23202 = n23193 & n23201;
  assign n23203 = ~n23193 & ~n23201;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = n14156 & ~n23204;
  assign n23206 = pi315 & n23205;
  assign n23207 = pi315 & n14156;
  assign n23208 = ~n23193 & n23201;
  assign n23209 = n23193 & ~n23201;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~n23207 & ~n23210;
  assign n23212 = ~n23206 & ~n23211;
  assign n23213 = n11998 & ~n23212;
  assign n23214 = pi314 & n23213;
  assign n23215 = pi314 & n11998;
  assign n23216 = ~n23211 & ~n23215;
  assign n23217 = ~n23206 & n23216;
  assign n23218 = ~n23214 & ~n23217;
  assign n23219 = ~n23043 & ~n23218;
  assign n23220 = n23043 & ~n23217;
  assign n23221 = ~n23214 & n23220;
  assign n23222 = ~n23219 & ~n23221;
  assign n23223 = n23038 & ~n23222;
  assign n23224 = ~n23038 & n23222;
  assign n23225 = ~n23223 & ~n23224;
  assign n23226 = pi312 & n9815;
  assign n23227 = ~n9517 & ~n9815;
  assign n23228 = pi313 & ~n23227;
  assign n23229 = n20477 & ~n23228;
  assign n23230 = ~n9517 & n9815;
  assign n23231 = pi313 & ~n20477;
  assign n23232 = n23230 & n23231;
  assign n23233 = ~n23229 & ~n23232;
  assign n23234 = ~n20491 & ~n23233;
  assign n23235 = ~n9815 & n20477;
  assign n23236 = ~n20479 & ~n23235;
  assign n23237 = ~n19064 & ~n23236;
  assign n23238 = n20490 & n23237;
  assign n23239 = n9517 & ~n9815;
  assign n23240 = ~n20477 & n23239;
  assign n23241 = ~n9517 & ~n19064;
  assign n23242 = n9815 & ~n23241;
  assign n23243 = n20477 & n23242;
  assign n23244 = ~n23240 & ~n23243;
  assign n23245 = pi313 & ~n23244;
  assign n23246 = n19064 & n20501;
  assign n23247 = ~n23245 & ~n23246;
  assign n23248 = ~n20490 & ~n23247;
  assign n23249 = ~n9815 & ~n20477;
  assign n23250 = n9815 & n20477;
  assign n23251 = ~n23249 & ~n23250;
  assign n23252 = n9517 & ~n23251;
  assign n23253 = pi313 & n23252;
  assign n23254 = n19064 & n23253;
  assign n23255 = ~n23248 & ~n23254;
  assign n23256 = ~n23238 & n23255;
  assign n23257 = ~n23234 & n23256;
  assign n23258 = ~n20512 & ~n23257;
  assign n23259 = n20512 & n23257;
  assign n23260 = n20481 & ~n23259;
  assign n23261 = ~n23258 & ~n23260;
  assign n23262 = n23226 & ~n23261;
  assign n23263 = ~n20481 & ~n23258;
  assign n23264 = ~n23259 & ~n23263;
  assign n23265 = ~n23226 & ~n23264;
  assign n23266 = ~n23262 & ~n23265;
  assign n23267 = ~n23225 & ~n23266;
  assign n23268 = n23038 & n23222;
  assign n23269 = ~n23038 & ~n23222;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = ~n23226 & ~n23261;
  assign n23272 = n23226 & ~n23264;
  assign n23273 = ~n23271 & ~n23272;
  assign n23274 = ~n23270 & ~n23273;
  assign n23275 = ~n23267 & ~n23274;
  assign n23276 = n23030 & ~n23275;
  assign n23277 = ~n23030 & n23275;
  assign n23278 = ~n23276 & ~n23277;
  assign n23279 = n9517 & ~n23278;
  assign n23280 = pi311 & n23279;
  assign n23281 = pi311 & n9517;
  assign n23282 = ~n23030 & ~n23275;
  assign n23283 = n23030 & n23275;
  assign n23284 = ~n23282 & ~n23283;
  assign n23285 = ~n23281 & ~n23284;
  assign n23286 = ~n23280 & ~n23285;
  assign n23287 = ~n7044 & ~n20532;
  assign n23288 = ~n19135 & ~n23287;
  assign n23289 = n6777 & n23288;
  assign n23290 = ~n19134 & ~n20532;
  assign n23291 = n7044 & ~n23290;
  assign n23292 = ~n23289 & ~n23291;
  assign n23293 = pi310 & ~n23292;
  assign n23294 = ~n20542 & ~n23293;
  assign n23295 = n23286 & ~n23294;
  assign n23296 = ~n23286 & n23294;
  assign n23297 = ~n23295 & ~n23296;
  assign n23298 = n7874 & ~n23297;
  assign n23299 = pi310 & n23298;
  assign n23300 = pi310 & n7874;
  assign n23301 = ~n23286 & ~n23294;
  assign n23302 = n23286 & n23294;
  assign n23303 = ~n23301 & ~n23302;
  assign n23304 = ~n23300 & ~n23303;
  assign n23305 = ~n23299 & ~n23304;
  assign n23306 = n23026 & n23305;
  assign n23307 = ~n23026 & ~n23305;
  assign n23308 = ~n23306 & ~n23307;
  assign n23309 = pi308 & n6777;
  assign n23310 = pi309 & ~n17124;
  assign n23311 = n20564 & ~n23310;
  assign n23312 = pi309 & ~n20564;
  assign n23313 = n17127 & n23312;
  assign n23314 = ~n23311 & ~n23313;
  assign n23315 = ~n20579 & ~n23314;
  assign n23316 = ~n6777 & n20564;
  assign n23317 = ~n20590 & ~n23316;
  assign n23318 = n19144 & ~n23317;
  assign n23319 = n20578 & n23318;
  assign n23320 = n17136 & ~n20564;
  assign n23321 = ~n5463 & n19144;
  assign n23322 = n6777 & ~n23321;
  assign n23323 = n20564 & n23322;
  assign n23324 = ~n23320 & ~n23323;
  assign n23325 = pi309 & ~n23324;
  assign n23326 = ~n19144 & n20565;
  assign n23327 = ~n23325 & ~n23326;
  assign n23328 = ~n20578 & ~n23327;
  assign n23329 = ~n6777 & ~n20564;
  assign n23330 = n6777 & n20564;
  assign n23331 = ~n23329 & ~n23330;
  assign n23332 = n5463 & ~n23331;
  assign n23333 = pi309 & n23332;
  assign n23334 = ~n19144 & n23333;
  assign n23335 = ~n23328 & ~n23334;
  assign n23336 = ~n23319 & n23335;
  assign n23337 = ~n23315 & n23336;
  assign n23338 = n20600 & n23337;
  assign n23339 = ~n20600 & ~n23337;
  assign n23340 = n20568 & ~n23339;
  assign n23341 = ~n23338 & ~n23340;
  assign n23342 = n23309 & ~n23341;
  assign n23343 = ~n20568 & ~n23338;
  assign n23344 = ~n23339 & ~n23343;
  assign n23345 = ~n23309 & ~n23344;
  assign n23346 = ~n23342 & ~n23345;
  assign n23347 = ~n23308 & ~n23346;
  assign n23348 = n23026 & ~n23305;
  assign n23349 = ~n23026 & n23305;
  assign n23350 = ~n23348 & ~n23349;
  assign n23351 = ~n23309 & ~n23341;
  assign n23352 = n23309 & ~n23344;
  assign n23353 = ~n23351 & ~n23352;
  assign n23354 = ~n23350 & ~n23353;
  assign n23355 = ~n23347 & ~n23354;
  assign n23356 = ~n23018 & ~n23355;
  assign n23357 = n23018 & n23355;
  assign n23358 = ~n23356 & ~n23357;
  assign n23359 = n5463 & ~n23358;
  assign n23360 = pi307 & n23359;
  assign n23361 = pi307 & n5463;
  assign n23362 = n23018 & ~n23355;
  assign n23363 = ~n23018 & n23355;
  assign n23364 = ~n23362 & ~n23363;
  assign n23365 = ~n23361 & ~n23364;
  assign n23366 = ~n23360 & ~n23365;
  assign n23367 = ~n19205 & n20640;
  assign n23368 = ~n19217 & ~n20622;
  assign n23369 = n3552 & n23368;
  assign n23370 = ~n19218 & n20620;
  assign n23371 = n4086 & ~n23370;
  assign n23372 = ~n23369 & ~n23371;
  assign n23373 = pi306 & ~n23372;
  assign n23374 = ~n23367 & ~n23373;
  assign n23375 = ~n23366 & n23374;
  assign n23376 = n23366 & ~n23374;
  assign n23377 = ~n23375 & ~n23376;
  assign n23378 = n4772 & ~n23377;
  assign n23379 = pi306 & n23378;
  assign n23380 = pi306 & n4772;
  assign n23381 = n23366 & n23374;
  assign n23382 = ~n23366 & ~n23374;
  assign n23383 = ~n23381 & ~n23382;
  assign n23384 = ~n23380 & ~n23383;
  assign n23385 = ~n23379 & ~n23384;
  assign n23386 = n23014 & n23385;
  assign n23387 = ~n23014 & ~n23385;
  assign n23388 = ~n23386 & ~n23387;
  assign n23389 = pi304 & n3552;
  assign n23390 = pi305 & n20652;
  assign n23391 = n11045 & n23390;
  assign n23392 = pi305 & ~n11042;
  assign n23393 = ~n20652 & ~n23392;
  assign n23394 = ~n23391 & ~n23393;
  assign n23395 = ~n20667 & ~n23394;
  assign n23396 = ~n3552 & ~n20652;
  assign n23397 = ~n20678 & ~n23396;
  assign n23398 = ~n19221 & ~n23397;
  assign n23399 = n20666 & n23398;
  assign n23400 = n3552 & ~n20652;
  assign n23401 = ~n3552 & n20652;
  assign n23402 = ~n23400 & ~n23401;
  assign n23403 = n3012 & ~n23402;
  assign n23404 = pi305 & n23403;
  assign n23405 = n19221 & n23404;
  assign n23406 = ~n3012 & ~n19221;
  assign n23407 = n3552 & ~n23406;
  assign n23408 = ~n20652 & n23407;
  assign n23409 = n11054 & n20652;
  assign n23410 = ~n23408 & ~n23409;
  assign n23411 = pi305 & ~n23410;
  assign n23412 = n19221 & n20653;
  assign n23413 = ~n23411 & ~n23412;
  assign n23414 = ~n20666 & ~n23413;
  assign n23415 = ~n23405 & ~n23414;
  assign n23416 = ~n23399 & n23415;
  assign n23417 = ~n23395 & n23416;
  assign n23418 = n20688 & n23417;
  assign n23419 = ~n20688 & ~n23417;
  assign n23420 = n20656 & ~n23419;
  assign n23421 = ~n23418 & ~n23420;
  assign n23422 = n23389 & ~n23421;
  assign n23423 = ~n20656 & ~n23418;
  assign n23424 = ~n23419 & ~n23423;
  assign n23425 = ~n23389 & ~n23424;
  assign n23426 = ~n23422 & ~n23425;
  assign n23427 = ~n23388 & ~n23426;
  assign n23428 = n23014 & ~n23385;
  assign n23429 = ~n23014 & n23385;
  assign n23430 = ~n23428 & ~n23429;
  assign n23431 = ~n23389 & ~n23421;
  assign n23432 = n23389 & ~n23424;
  assign n23433 = ~n23431 & ~n23432;
  assign n23434 = ~n23430 & ~n23433;
  assign n23435 = ~n23427 & ~n23434;
  assign n23436 = ~n23006 & n23435;
  assign n23437 = n23006 & ~n23435;
  assign n23438 = ~n23436 & ~n23437;
  assign n23439 = n3012 & ~n23438;
  assign n23440 = pi303 & n23439;
  assign n23441 = pi303 & n3012;
  assign n23442 = n23006 & n23435;
  assign n23443 = ~n23006 & ~n23435;
  assign n23444 = ~n23442 & ~n23443;
  assign n23445 = ~n23441 & ~n23444;
  assign n23446 = ~n23440 & ~n23445;
  assign n23447 = n2574 & ~n23446;
  assign n23448 = pi302 & n23447;
  assign n23449 = pi302 & n2574;
  assign n23450 = ~n23445 & ~n23449;
  assign n23451 = ~n23440 & n23450;
  assign n23452 = ~n23448 & ~n23451;
  assign n23453 = n23002 & ~n23452;
  assign n23454 = ~n23002 & ~n23451;
  assign n23455 = ~n23448 & n23454;
  assign n23456 = ~n23453 & ~n23455;
  assign n23457 = n22994 & ~n23456;
  assign n23458 = ~n22994 & n23456;
  assign n23459 = ~n23457 & ~n23458;
  assign n23460 = pi300 & n1840;
  assign n23461 = pi301 & ~n6883;
  assign n23462 = n20740 & ~n23461;
  assign n23463 = pi301 & ~n20740;
  assign n23464 = n6886 & n23463;
  assign n23465 = ~n23462 & ~n23464;
  assign n23466 = ~n20745 & ~n23465;
  assign n23467 = ~n1840 & n20740;
  assign n23468 = ~n20742 & ~n23467;
  assign n23469 = ~n19298 & ~n23468;
  assign n23470 = n18852 & n23469;
  assign n23471 = n6897 & ~n20740;
  assign n23472 = ~n1533 & ~n19298;
  assign n23473 = n1840 & ~n23472;
  assign n23474 = n20740 & n23473;
  assign n23475 = ~n23471 & ~n23474;
  assign n23476 = pi301 & ~n23475;
  assign n23477 = n19298 & n20755;
  assign n23478 = ~n23476 & ~n23477;
  assign n23479 = ~n18852 & ~n23478;
  assign n23480 = ~n1840 & ~n20740;
  assign n23481 = n1840 & n20740;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = n1533 & ~n23482;
  assign n23484 = pi301 & n23483;
  assign n23485 = n19298 & n23484;
  assign n23486 = ~n23479 & ~n23485;
  assign n23487 = ~n23470 & n23486;
  assign n23488 = ~n23466 & n23487;
  assign n23489 = ~n20766 & ~n23488;
  assign n23490 = n20766 & n23488;
  assign n23491 = n20744 & ~n23490;
  assign n23492 = ~n23489 & ~n23491;
  assign n23493 = n23460 & ~n23492;
  assign n23494 = ~n20744 & ~n23489;
  assign n23495 = ~n23490 & ~n23494;
  assign n23496 = ~n23460 & ~n23495;
  assign n23497 = ~n23493 & ~n23496;
  assign n23498 = ~n23459 & ~n23497;
  assign n23499 = n22994 & n23456;
  assign n23500 = ~n22994 & ~n23456;
  assign n23501 = ~n23499 & ~n23500;
  assign n23502 = ~n23460 & ~n23492;
  assign n23503 = n23460 & ~n23495;
  assign n23504 = ~n23502 & ~n23503;
  assign n23505 = ~n23501 & ~n23504;
  assign n23506 = ~n23498 & ~n23505;
  assign n23507 = n22986 & n23506;
  assign n23508 = ~n22986 & ~n23506;
  assign n23509 = ~n23507 & ~n23508;
  assign n23510 = n1533 & ~n23509;
  assign n23511 = pi299 & n23510;
  assign n23512 = pi299 & n1533;
  assign n23513 = ~n22986 & n23506;
  assign n23514 = n22986 & ~n23506;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = ~n23512 & ~n23515;
  assign n23517 = ~n23511 & ~n23516;
  assign n23518 = n1553 & ~n23517;
  assign n23519 = pi298 & n23518;
  assign n23520 = pi298 & n1553;
  assign n23521 = ~n23516 & ~n23520;
  assign n23522 = ~n23511 & n23521;
  assign n23523 = ~n23519 & ~n23522;
  assign n23524 = ~n22979 & ~n23523;
  assign n23525 = n22979 & ~n23522;
  assign n23526 = ~n23519 & n23525;
  assign n23527 = ~n23524 & ~n23526;
  assign n23528 = n22971 & n23527;
  assign n23529 = ~n22971 & ~n23527;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = pi296 & ~n1568;
  assign n23532 = ~n20810 & ~n23531;
  assign n23533 = n20810 & n23531;
  assign n23534 = ~n23532 & ~n23533;
  assign n23535 = pi295 & ~n23534;
  assign n23536 = pi128 & n23535;
  assign n23537 = pi128 & pi295;
  assign n23538 = n20810 & ~n23531;
  assign n23539 = ~n20810 & n23531;
  assign n23540 = ~n23538 & ~n23539;
  assign n23541 = ~n23537 & ~n23540;
  assign n23542 = ~n23536 & ~n23541;
  assign n23543 = ~n23530 & ~n23542;
  assign n23544 = n22971 & ~n23527;
  assign n23545 = ~n22971 & n23527;
  assign n23546 = ~n23544 & ~n23545;
  assign n23547 = pi295 & ~n23540;
  assign n23548 = pi128 & n23547;
  assign n23549 = ~n23534 & ~n23537;
  assign n23550 = ~n23548 & ~n23549;
  assign n23551 = ~n23546 & ~n23550;
  assign n23552 = ~n23543 & ~n23551;
  assign n23553 = ~n20818 & ~n21855;
  assign n23554 = n20818 & n21855;
  assign n23555 = ~pi283 & ~n23554;
  assign n23556 = ~n23553 & ~n23555;
  assign n23557 = n23552 & n23556;
  assign n23558 = ~n23552 & ~n23556;
  assign n23559 = ~n23557 & ~n23558;
  assign n23560 = pi284 & ~n23559;
  assign n23561 = ~n23552 & n23556;
  assign n23562 = n23552 & ~n23556;
  assign n23563 = ~n23561 & ~n23562;
  assign n23564 = ~pi284 & ~n23563;
  assign n23565 = ~n23560 & ~n23564;
  assign n23566 = ~n22943 & ~n23565;
  assign n23567 = n22935 & n22940;
  assign n23568 = ~n22935 & ~n22940;
  assign n23569 = ~n23567 & ~n23568;
  assign n23570 = pi284 & ~n23563;
  assign n23571 = ~pi284 & ~n23559;
  assign n23572 = ~n23570 & ~n23571;
  assign n23573 = ~n23569 & ~n23572;
  assign n23574 = ~n23566 & ~n23573;
  assign n23575 = ~n831 & ~n23574;
  assign n23576 = ~pi284 & n831;
  assign n23577 = ~n23575 & ~n23576;
  assign n23578 = pi161 & n23577;
  assign n23579 = ~n21882 & ~n23578;
  assign po219 = ~pi160 & ~n23579;
  assign n23581 = ~pi091 & ~pi161;
  assign n23582 = ~pi285 & n831;
  assign n23583 = pi297 & n1553;
  assign n23584 = ~n1533 & ~n23506;
  assign n23585 = n1533 & n23506;
  assign n23586 = ~n22986 & ~n23585;
  assign n23587 = ~n23584 & ~n23586;
  assign n23588 = n1840 & ~n23587;
  assign n23589 = ~n1840 & ~n23508;
  assign n23590 = n1533 & n23589;
  assign n23591 = ~n23588 & ~n23590;
  assign n23592 = pi299 & ~n23591;
  assign n23593 = pi299 & n1840;
  assign n23594 = n23506 & ~n23593;
  assign n23595 = n22986 & n23594;
  assign n23596 = ~n23592 & ~n23595;
  assign n23597 = pi301 & n2574;
  assign n23598 = ~n3012 & n23435;
  assign n23599 = n3012 & ~n23435;
  assign n23600 = ~n23006 & ~n23599;
  assign n23601 = ~n23598 & ~n23600;
  assign n23602 = n3552 & ~n23601;
  assign n23603 = ~n3552 & ~n23436;
  assign n23604 = n3012 & n23603;
  assign n23605 = ~n23602 & ~n23604;
  assign n23606 = pi303 & ~n23605;
  assign n23607 = pi303 & n3552;
  assign n23608 = ~n23435 & ~n23607;
  assign n23609 = n23006 & n23608;
  assign n23610 = ~n23606 & ~n23609;
  assign n23611 = pi305 & n4772;
  assign n23612 = pi309 & n7874;
  assign n23613 = pi313 & n11998;
  assign n23614 = ~pi155 & n23060;
  assign n23615 = pi155 & ~n23060;
  assign n23616 = ~pi154 & n23615;
  assign n23617 = ~n23614 & ~n23616;
  assign n23618 = pi153 & ~n23617;
  assign n23619 = ~pi155 & ~n23060;
  assign n23620 = pi155 & n23060;
  assign n23621 = pi154 & n23620;
  assign n23622 = ~n23619 & ~n23621;
  assign n23623 = ~pi153 & ~n23622;
  assign n23624 = ~pi155 & ~n23067;
  assign n23625 = ~n23623 & ~n23624;
  assign n23626 = ~n23618 & n23625;
  assign n23627 = ~n20348 & n20359;
  assign n23628 = n18937 & ~n23627;
  assign n23629 = pi320 & n23628;
  assign n23630 = pi321 & n23070;
  assign n23631 = ~n23629 & ~n23630;
  assign n23632 = n23069 & ~n23631;
  assign n23633 = ~pi320 & ~n23632;
  assign n23634 = ~n20347 & ~n23069;
  assign n23635 = n20347 & n23631;
  assign n23636 = pi320 & n23632;
  assign n23637 = ~n23635 & ~n23636;
  assign n23638 = ~n23634 & n23637;
  assign n23639 = ~n23633 & n23638;
  assign n23640 = n23626 & ~n23639;
  assign n23641 = ~n23626 & ~n23631;
  assign n23642 = ~pi320 & n23069;
  assign n23643 = n23641 & n23642;
  assign n23644 = ~n23640 & ~n23643;
  assign n23645 = pi321 & ~n23644;
  assign n23646 = ~n23626 & n23631;
  assign n23647 = ~n20347 & n23646;
  assign n23648 = n20347 & ~n23631;
  assign n23649 = ~pi321 & ~n23648;
  assign n23650 = ~n23647 & ~n23649;
  assign n23651 = n23069 & ~n23650;
  assign n23652 = pi321 & n23626;
  assign n23653 = ~n23631 & ~n23652;
  assign n23654 = ~n23069 & n23653;
  assign n23655 = n20347 & n23654;
  assign n23656 = ~n23651 & ~n23655;
  assign n23657 = pi320 & ~n23656;
  assign n23658 = ~n23645 & ~n23657;
  assign n23659 = pi319 & n20347;
  assign n23660 = ~n23658 & ~n23659;
  assign n23661 = n20347 & n23658;
  assign n23662 = pi319 & n23661;
  assign n23663 = ~n23660 & ~n23662;
  assign n23664 = ~n18937 & n23094;
  assign n23665 = ~n23118 & ~n23664;
  assign n23666 = n17455 & n23665;
  assign n23667 = ~n23049 & n23094;
  assign n23668 = n18937 & ~n23667;
  assign n23669 = ~n23666 & ~n23668;
  assign n23670 = pi319 & ~n23669;
  assign n23671 = ~n23106 & ~n23670;
  assign n23672 = ~n23663 & ~n23671;
  assign n23673 = n23663 & n23671;
  assign n23674 = ~n23672 & ~n23673;
  assign n23675 = n18937 & ~n23674;
  assign n23676 = pi318 & n23675;
  assign n23677 = pi318 & n18937;
  assign n23678 = n23663 & ~n23671;
  assign n23679 = ~n23663 & n23671;
  assign n23680 = ~n23678 & ~n23679;
  assign n23681 = ~n23677 & ~n23680;
  assign n23682 = ~n23676 & ~n23681;
  assign n23683 = n17455 & ~n23130;
  assign n23684 = pi318 & n23683;
  assign n23685 = n23130 & ~n23131;
  assign n23686 = ~n23136 & ~n23685;
  assign n23687 = ~n20391 & n23686;
  assign n23688 = ~n23684 & ~n23687;
  assign n23689 = ~n23682 & n23688;
  assign n23690 = n23682 & ~n23688;
  assign n23691 = ~n23689 & ~n23690;
  assign n23692 = n17455 & ~n23691;
  assign n23693 = pi317 & n23692;
  assign n23694 = pi317 & n17455;
  assign n23695 = ~n23690 & ~n23694;
  assign n23696 = ~n23689 & n23695;
  assign n23697 = ~n23693 & ~n23696;
  assign n23698 = ~n23141 & ~n23151;
  assign n23699 = n23141 & n23151;
  assign n23700 = ~n23142 & ~n23699;
  assign n23701 = ~n20397 & n23700;
  assign n23702 = ~n23698 & ~n23701;
  assign n23703 = pi316 & n16985;
  assign n23704 = n23702 & ~n23703;
  assign n23705 = n16985 & ~n23702;
  assign n23706 = pi316 & n23705;
  assign n23707 = ~n23704 & ~n23706;
  assign n23708 = ~n23697 & ~n23707;
  assign n23709 = ~n23702 & ~n23703;
  assign n23710 = n16985 & n23702;
  assign n23711 = pi316 & n23710;
  assign n23712 = ~n23709 & ~n23711;
  assign n23713 = ~n23696 & ~n23712;
  assign n23714 = ~n23693 & n23713;
  assign n23715 = ~n23708 & ~n23714;
  assign n23716 = ~n14618 & n23157;
  assign n23717 = ~n23181 & ~n23716;
  assign n23718 = n14156 & n23717;
  assign n23719 = ~n23048 & n23157;
  assign n23720 = n14618 & ~n23719;
  assign n23721 = ~n23718 & ~n23720;
  assign n23722 = pi316 & ~n23721;
  assign n23723 = ~n23169 & ~n23722;
  assign n23724 = n23715 & n23723;
  assign n23725 = ~n23715 & ~n23723;
  assign n23726 = ~n23724 & ~n23725;
  assign n23727 = n14618 & ~n23726;
  assign n23728 = pi315 & n23727;
  assign n23729 = pi315 & n14618;
  assign n23730 = ~n23715 & n23723;
  assign n23731 = n23715 & ~n23723;
  assign n23732 = ~n23730 & ~n23731;
  assign n23733 = ~n23729 & ~n23732;
  assign n23734 = ~n23728 & ~n23733;
  assign n23735 = ~n23201 & n23207;
  assign n23736 = n23201 & ~n23207;
  assign n23737 = ~n23193 & ~n23736;
  assign n23738 = ~n23735 & ~n23737;
  assign n23739 = n23734 & n23738;
  assign n23740 = ~n23734 & ~n23738;
  assign n23741 = ~n23739 & ~n23740;
  assign n23742 = pi314 & n14156;
  assign n23743 = ~n23220 & ~n23742;
  assign n23744 = ~n23214 & n23743;
  assign n23745 = ~n23214 & ~n23220;
  assign n23746 = n23742 & ~n23745;
  assign n23747 = ~n23744 & ~n23746;
  assign n23748 = ~n23741 & ~n23747;
  assign n23749 = n23734 & ~n23738;
  assign n23750 = ~n23734 & n23738;
  assign n23751 = ~n23749 & ~n23750;
  assign n23752 = ~n23220 & n23742;
  assign n23753 = ~n23214 & n23752;
  assign n23754 = ~n23742 & ~n23745;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = ~n23751 & ~n23755;
  assign n23757 = ~n23748 & ~n23756;
  assign n23758 = ~n23613 & n23757;
  assign n23759 = n23613 & ~n23757;
  assign n23760 = ~n23758 & ~n23759;
  assign n23761 = pi312 & n10908;
  assign n23762 = n19064 & ~n20501;
  assign n23763 = n9517 & ~n23249;
  assign n23764 = pi313 & n23763;
  assign n23765 = ~n23762 & ~n23764;
  assign n23766 = ~n20490 & ~n23765;
  assign n23767 = n19064 & n23763;
  assign n23768 = ~n23250 & ~n23767;
  assign n23769 = pi313 & ~n23768;
  assign n23770 = ~n23766 & ~n23769;
  assign n23771 = n23222 & ~n23770;
  assign n23772 = ~n23222 & n23770;
  assign n23773 = n23031 & ~n23772;
  assign n23774 = ~n23771 & ~n23773;
  assign n23775 = n23761 & ~n23774;
  assign n23776 = ~n23031 & ~n23771;
  assign n23777 = ~n23772 & ~n23776;
  assign n23778 = ~n23761 & ~n23777;
  assign n23779 = ~n23775 & ~n23778;
  assign n23780 = ~n23760 & ~n23779;
  assign n23781 = ~n23613 & ~n23757;
  assign n23782 = n23613 & n23757;
  assign n23783 = ~n23781 & ~n23782;
  assign n23784 = ~n23761 & ~n23774;
  assign n23785 = n23761 & ~n23777;
  assign n23786 = ~n23784 & ~n23785;
  assign n23787 = ~n23783 & ~n23786;
  assign n23788 = ~n23780 & ~n23787;
  assign n23789 = n23226 & ~n23270;
  assign n23790 = ~n23226 & n23270;
  assign n23791 = ~n23261 & ~n23790;
  assign n23792 = ~n23789 & ~n23791;
  assign n23793 = n23788 & n23792;
  assign n23794 = ~n23788 & ~n23792;
  assign n23795 = ~n23793 & ~n23794;
  assign n23796 = pi311 & n9815;
  assign n23797 = n23281 & ~n23282;
  assign n23798 = ~n23283 & ~n23797;
  assign n23799 = n23796 & ~n23798;
  assign n23800 = ~n23281 & ~n23283;
  assign n23801 = ~n23282 & ~n23800;
  assign n23802 = ~n23796 & ~n23801;
  assign n23803 = ~n23799 & ~n23802;
  assign n23804 = ~n23795 & ~n23803;
  assign n23805 = n23788 & ~n23792;
  assign n23806 = ~n23788 & n23792;
  assign n23807 = ~n23805 & ~n23806;
  assign n23808 = ~n23796 & ~n23798;
  assign n23809 = n23796 & ~n23801;
  assign n23810 = ~n23808 & ~n23809;
  assign n23811 = ~n23807 & ~n23810;
  assign n23812 = ~n23804 & ~n23811;
  assign n23813 = ~pi310 & n23812;
  assign n23814 = ~n9517 & n23812;
  assign n23815 = n9517 & ~n23812;
  assign n23816 = pi310 & n23815;
  assign n23817 = ~n23814 & ~n23816;
  assign n23818 = ~n7874 & ~n23817;
  assign n23819 = ~n23813 & ~n23818;
  assign n23820 = ~n23295 & ~n23819;
  assign n23821 = ~n23294 & n23812;
  assign n23822 = n23286 & n23821;
  assign n23823 = n23294 & ~n23812;
  assign n23824 = ~n23286 & n23823;
  assign n23825 = ~n23822 & ~n23824;
  assign n23826 = pi310 & ~n23825;
  assign n23827 = ~n23303 & n23812;
  assign n23828 = n7874 & n23827;
  assign n23829 = ~n23826 & ~n23828;
  assign n23830 = n9517 & ~n23829;
  assign n23831 = ~n23294 & ~n23812;
  assign n23832 = ~pi310 & n23286;
  assign n23833 = n23831 & n23832;
  assign n23834 = n23294 & n23812;
  assign n23835 = ~n23286 & n23834;
  assign n23836 = n7874 & ~n23296;
  assign n23837 = pi310 & n23836;
  assign n23838 = ~n23295 & ~n23837;
  assign n23839 = ~n23812 & ~n23838;
  assign n23840 = ~n23835 & ~n23839;
  assign n23841 = ~n9517 & ~n23840;
  assign n23842 = ~n23833 & ~n23841;
  assign n23843 = ~n23830 & n23842;
  assign n23844 = ~n23820 & n23843;
  assign n23845 = ~n23612 & ~n23844;
  assign n23846 = n23612 & n23844;
  assign n23847 = ~n23845 & ~n23846;
  assign n23848 = pi308 & n7044;
  assign n23849 = n5463 & ~n23316;
  assign n23850 = pi309 & n23849;
  assign n23851 = ~n19144 & ~n20589;
  assign n23852 = ~n23850 & ~n23851;
  assign n23853 = ~n20578 & ~n23852;
  assign n23854 = n6777 & ~n20564;
  assign n23855 = ~n19144 & n23849;
  assign n23856 = ~n23854 & ~n23855;
  assign n23857 = pi309 & ~n23856;
  assign n23858 = ~n23853 & ~n23857;
  assign n23859 = ~n23305 & ~n23858;
  assign n23860 = n23305 & n23858;
  assign n23861 = n23019 & ~n23860;
  assign n23862 = ~n23859 & ~n23861;
  assign n23863 = n23848 & ~n23862;
  assign n23864 = ~n23019 & ~n23859;
  assign n23865 = ~n23860 & ~n23864;
  assign n23866 = ~n23848 & ~n23865;
  assign n23867 = ~n23863 & ~n23866;
  assign n23868 = ~n23847 & ~n23867;
  assign n23869 = ~n23612 & n23844;
  assign n23870 = n23612 & ~n23844;
  assign n23871 = ~n23869 & ~n23870;
  assign n23872 = ~n23848 & ~n23862;
  assign n23873 = n23848 & ~n23865;
  assign n23874 = ~n23872 & ~n23873;
  assign n23875 = ~n23871 & ~n23874;
  assign n23876 = ~n23868 & ~n23875;
  assign n23877 = ~n23308 & ~n23309;
  assign n23878 = n23308 & n23309;
  assign n23879 = ~n23344 & ~n23878;
  assign n23880 = ~n23877 & ~n23879;
  assign n23881 = n23876 & n23880;
  assign n23882 = ~n23876 & ~n23880;
  assign n23883 = ~n23881 & ~n23882;
  assign n23884 = pi307 & n6777;
  assign n23885 = ~n23356 & n23361;
  assign n23886 = ~n23357 & ~n23885;
  assign n23887 = n23884 & ~n23886;
  assign n23888 = ~n23357 & ~n23361;
  assign n23889 = ~n23356 & ~n23888;
  assign n23890 = ~n23884 & ~n23889;
  assign n23891 = ~n23887 & ~n23890;
  assign n23892 = ~n23883 & ~n23891;
  assign n23893 = n23876 & ~n23880;
  assign n23894 = ~n23876 & n23880;
  assign n23895 = ~n23893 & ~n23894;
  assign n23896 = ~n23884 & ~n23886;
  assign n23897 = n23884 & ~n23889;
  assign n23898 = ~n23896 & ~n23897;
  assign n23899 = ~n23895 & ~n23898;
  assign n23900 = ~n23892 & ~n23899;
  assign n23901 = ~pi306 & n23900;
  assign n23902 = ~n5463 & n23900;
  assign n23903 = n5463 & ~n23900;
  assign n23904 = pi306 & n23903;
  assign n23905 = ~n23902 & ~n23904;
  assign n23906 = ~n4772 & ~n23905;
  assign n23907 = ~n23901 & ~n23906;
  assign n23908 = ~n23382 & ~n23907;
  assign n23909 = ~n23374 & n23900;
  assign n23910 = ~n23366 & n23909;
  assign n23911 = n23374 & ~n23900;
  assign n23912 = n23366 & n23911;
  assign n23913 = ~n23910 & ~n23912;
  assign n23914 = pi306 & ~n23913;
  assign n23915 = ~n23377 & n23900;
  assign n23916 = n4772 & n23915;
  assign n23917 = ~n23914 & ~n23916;
  assign n23918 = n5463 & ~n23917;
  assign n23919 = ~pi306 & ~n23366;
  assign n23920 = ~n23374 & ~n23900;
  assign n23921 = n23919 & n23920;
  assign n23922 = n23374 & n23900;
  assign n23923 = n23366 & n23922;
  assign n23924 = n4772 & ~n23381;
  assign n23925 = pi306 & n23924;
  assign n23926 = ~n23382 & ~n23925;
  assign n23927 = ~n23900 & ~n23926;
  assign n23928 = ~n23923 & ~n23927;
  assign n23929 = ~n5463 & ~n23928;
  assign n23930 = ~n23921 & ~n23929;
  assign n23931 = ~n23918 & n23930;
  assign n23932 = ~n23908 & n23931;
  assign n23933 = ~n23611 & n23932;
  assign n23934 = n23611 & ~n23932;
  assign n23935 = ~n23933 & ~n23934;
  assign n23936 = pi304 & n4086;
  assign n23937 = n19221 & ~n20677;
  assign n23938 = n3012 & ~n23396;
  assign n23939 = pi305 & n23938;
  assign n23940 = ~n23937 & ~n23939;
  assign n23941 = ~n20666 & ~n23940;
  assign n23942 = n3552 & n20652;
  assign n23943 = n19221 & n23938;
  assign n23944 = ~n23942 & ~n23943;
  assign n23945 = pi305 & ~n23944;
  assign n23946 = ~n23941 & ~n23945;
  assign n23947 = n23385 & ~n23946;
  assign n23948 = ~n23385 & n23946;
  assign n23949 = n23007 & ~n23948;
  assign n23950 = ~n23947 & ~n23949;
  assign n23951 = n23936 & ~n23950;
  assign n23952 = ~n23007 & ~n23947;
  assign n23953 = ~n23948 & ~n23952;
  assign n23954 = ~n23936 & ~n23953;
  assign n23955 = ~n23951 & ~n23954;
  assign n23956 = ~n23935 & ~n23955;
  assign n23957 = ~n23611 & ~n23932;
  assign n23958 = n23611 & n23932;
  assign n23959 = ~n23957 & ~n23958;
  assign n23960 = ~n23936 & ~n23950;
  assign n23961 = n23936 & ~n23953;
  assign n23962 = ~n23960 & ~n23961;
  assign n23963 = ~n23959 & ~n23962;
  assign n23964 = ~n23956 & ~n23963;
  assign n23965 = ~n23389 & ~n23430;
  assign n23966 = n23389 & n23430;
  assign n23967 = ~n23424 & ~n23966;
  assign n23968 = ~n23965 & ~n23967;
  assign n23969 = ~n23964 & ~n23968;
  assign n23970 = n23964 & n23968;
  assign n23971 = ~n23969 & ~n23970;
  assign n23972 = n23610 & n23971;
  assign n23973 = ~n23610 & ~n23971;
  assign n23974 = ~n23972 & ~n23973;
  assign n23975 = pi302 & n3012;
  assign n23976 = ~n23454 & ~n23975;
  assign n23977 = ~n23448 & n23976;
  assign n23978 = ~n23448 & ~n23454;
  assign n23979 = n23975 & ~n23978;
  assign n23980 = ~n23977 & ~n23979;
  assign n23981 = ~n23974 & ~n23980;
  assign n23982 = n23610 & ~n23971;
  assign n23983 = ~n23610 & n23971;
  assign n23984 = ~n23982 & ~n23983;
  assign n23985 = ~n23454 & n23975;
  assign n23986 = ~n23448 & n23985;
  assign n23987 = ~n23975 & ~n23978;
  assign n23988 = ~n23986 & ~n23987;
  assign n23989 = ~n23984 & ~n23988;
  assign n23990 = ~n23981 & ~n23989;
  assign n23991 = ~n23597 & n23990;
  assign n23992 = n23597 & ~n23990;
  assign n23993 = ~n23991 & ~n23992;
  assign n23994 = pi300 & n2183;
  assign n23995 = n19298 & ~n20755;
  assign n23996 = n1533 & ~n23480;
  assign n23997 = pi301 & n23996;
  assign n23998 = ~n23995 & ~n23997;
  assign n23999 = ~n18852 & ~n23998;
  assign n24000 = n19298 & n23996;
  assign n24001 = ~n23481 & ~n24000;
  assign n24002 = pi301 & ~n24001;
  assign n24003 = ~n23999 & ~n24002;
  assign n24004 = n23456 & ~n24003;
  assign n24005 = ~n23456 & n24003;
  assign n24006 = n22987 & ~n24005;
  assign n24007 = ~n24004 & ~n24006;
  assign n24008 = n23994 & ~n24007;
  assign n24009 = ~n22987 & ~n24004;
  assign n24010 = ~n24005 & ~n24009;
  assign n24011 = ~n23994 & ~n24010;
  assign n24012 = ~n24008 & ~n24011;
  assign n24013 = ~n23993 & ~n24012;
  assign n24014 = ~n23597 & ~n23990;
  assign n24015 = n23597 & n23990;
  assign n24016 = ~n24014 & ~n24015;
  assign n24017 = ~n23994 & ~n24007;
  assign n24018 = n23994 & ~n24010;
  assign n24019 = ~n24017 & ~n24018;
  assign n24020 = ~n24016 & ~n24019;
  assign n24021 = ~n24013 & ~n24020;
  assign n24022 = n23460 & ~n23501;
  assign n24023 = ~n23460 & n23501;
  assign n24024 = ~n23492 & ~n24023;
  assign n24025 = ~n24022 & ~n24024;
  assign n24026 = ~n24021 & ~n24025;
  assign n24027 = n24021 & n24025;
  assign n24028 = ~n24026 & ~n24027;
  assign n24029 = n23596 & n24028;
  assign n24030 = ~n23596 & ~n24028;
  assign n24031 = ~n24029 & ~n24030;
  assign n24032 = pi298 & n1533;
  assign n24033 = ~n22979 & ~n23522;
  assign n24034 = ~n24032 & ~n24033;
  assign n24035 = ~n23519 & n24034;
  assign n24036 = ~n23519 & ~n24033;
  assign n24037 = n24032 & ~n24036;
  assign n24038 = ~n24035 & ~n24037;
  assign n24039 = ~n24031 & ~n24038;
  assign n24040 = n23596 & ~n24028;
  assign n24041 = ~n23596 & n24028;
  assign n24042 = ~n24040 & ~n24041;
  assign n24043 = n24032 & ~n24033;
  assign n24044 = ~n23519 & n24043;
  assign n24045 = ~n24032 & ~n24036;
  assign n24046 = ~n24044 & ~n24045;
  assign n24047 = ~n24042 & ~n24046;
  assign n24048 = ~n24039 & ~n24047;
  assign n24049 = ~n23583 & ~n24048;
  assign n24050 = n23583 & n24048;
  assign n24051 = ~n24049 & ~n24050;
  assign n24052 = n1335 & n22951;
  assign n24053 = ~pi129 & n20302;
  assign n24054 = pi129 & ~n20302;
  assign n24055 = n20805 & ~n24054;
  assign n24056 = pi128 & n24055;
  assign n24057 = ~n24053 & ~n24056;
  assign n24058 = pi130 & ~n24057;
  assign n24059 = ~n24052 & ~n24058;
  assign n24060 = pi297 & ~n24059;
  assign n24061 = pi296 & n1515;
  assign n24062 = n20302 & n20805;
  assign n24063 = ~pi130 & ~n24062;
  assign n24064 = pi128 & n24063;
  assign n24065 = pi297 & ~n11201;
  assign n24066 = ~n20805 & ~n24065;
  assign n24067 = ~n24064 & ~n24066;
  assign n24068 = pi129 & ~n24067;
  assign n24069 = pi128 & n20805;
  assign n24070 = ~pi130 & ~n24069;
  assign n24071 = ~pi129 & n24070;
  assign n24072 = pi297 & ~n24071;
  assign n24073 = ~n20302 & ~n24072;
  assign n24074 = ~n24068 & ~n24073;
  assign n24075 = ~n23527 & n24074;
  assign n24076 = ~n24061 & ~n24075;
  assign n24077 = ~n24060 & n24076;
  assign n24078 = ~n24060 & ~n24075;
  assign n24079 = n24061 & ~n24078;
  assign n24080 = ~n24077 & ~n24079;
  assign n24081 = ~n24051 & ~n24080;
  assign n24082 = ~n23583 & n24048;
  assign n24083 = n23583 & ~n24048;
  assign n24084 = ~n24082 & ~n24083;
  assign n24085 = n24061 & ~n24075;
  assign n24086 = ~n24060 & n24085;
  assign n24087 = ~n24061 & ~n24078;
  assign n24088 = ~n24086 & ~n24087;
  assign n24089 = ~n24084 & ~n24088;
  assign n24090 = ~n24081 & ~n24089;
  assign n24091 = ~n24060 & n24074;
  assign n24092 = ~n23527 & ~n24091;
  assign n24093 = n23527 & n24091;
  assign n24094 = ~n24092 & ~n24093;
  assign n24095 = ~n23532 & ~n24094;
  assign n24096 = ~n23533 & ~n24095;
  assign n24097 = ~n24090 & ~n24096;
  assign n24098 = n24090 & n24096;
  assign n24099 = ~n24097 & ~n24098;
  assign n24100 = ~n23534 & ~n23546;
  assign n24101 = ~n23530 & ~n23540;
  assign n24102 = ~n24100 & ~n24101;
  assign n24103 = pi295 & ~n24102;
  assign n24104 = pi128 & n24103;
  assign n24105 = pi129 & n24104;
  assign n24106 = pi295 & ~n1568;
  assign n24107 = ~n24104 & n24106;
  assign n24108 = ~n24105 & ~n24107;
  assign n24109 = ~n24099 & ~n24108;
  assign n24110 = n24090 & ~n24096;
  assign n24111 = ~n24090 & n24096;
  assign n24112 = ~n24110 & ~n24111;
  assign n24113 = ~pi129 & n24104;
  assign n24114 = ~n24104 & ~n24106;
  assign n24115 = ~n24113 & ~n24114;
  assign n24116 = ~n24112 & ~n24115;
  assign n24117 = ~n24109 & ~n24116;
  assign n24118 = ~n22917 & ~n22929;
  assign n24119 = ~n22910 & ~n22923;
  assign n24120 = ~n24118 & ~n24119;
  assign n24121 = n1156 & ~n24120;
  assign n24122 = pi348 & n24121;
  assign n24123 = n1154 & n24122;
  assign n24124 = ~n1154 & ~n24122;
  assign n24125 = pi348 & n24124;
  assign n24126 = ~n24123 & ~n24125;
  assign n24127 = n21913 & n22875;
  assign n24128 = ~n21913 & ~n22875;
  assign n24129 = ~n24127 & ~n24128;
  assign n24130 = ~n21922 & n22879;
  assign n24131 = n21926 & ~n22886;
  assign n24132 = ~n21926 & n22886;
  assign n24133 = ~n24131 & ~n24132;
  assign n24134 = ~n24130 & ~n24133;
  assign n24135 = ~n24129 & n24134;
  assign n24136 = ~n21913 & n22875;
  assign n24137 = n21913 & ~n22875;
  assign n24138 = ~n24136 & ~n24137;
  assign n24139 = ~n21926 & ~n22886;
  assign n24140 = n21926 & n22886;
  assign n24141 = ~n24139 & ~n24140;
  assign n24142 = ~n24130 & ~n24141;
  assign n24143 = ~n24138 & n24142;
  assign n24144 = n21922 & ~n22879;
  assign n24145 = ~n24143 & ~n24144;
  assign n24146 = ~n24135 & n24145;
  assign n24147 = ~n1256 & ~n21887;
  assign n24148 = pi346 & n24147;
  assign n24149 = n1256 & ~n21883;
  assign n24150 = ~n21886 & n24149;
  assign n24151 = pi346 & ~n24150;
  assign n24152 = ~n24148 & n24151;
  assign n24153 = ~n22907 & ~n24152;
  assign n24154 = n22907 & n24152;
  assign n24155 = ~n24153 & ~n24154;
  assign n24156 = ~n22915 & ~n24155;
  assign n24157 = ~n22916 & ~n24156;
  assign n24158 = n24146 & n24157;
  assign n24159 = ~n24146 & ~n24157;
  assign n24160 = ~n24158 & ~n24159;
  assign n24161 = pi345 & n1729;
  assign n24162 = ~n21946 & ~n22786;
  assign n24163 = n21946 & n22786;
  assign n24164 = ~n24162 & ~n24163;
  assign n24165 = ~n21961 & n22790;
  assign n24166 = n21965 & ~n22798;
  assign n24167 = ~n21965 & n22798;
  assign n24168 = ~n24166 & ~n24167;
  assign n24169 = ~n24165 & ~n24168;
  assign n24170 = ~n24164 & n24169;
  assign n24171 = ~n21946 & n22786;
  assign n24172 = n21946 & ~n22786;
  assign n24173 = ~n24171 & ~n24172;
  assign n24174 = ~n21965 & ~n22798;
  assign n24175 = n21965 & n22798;
  assign n24176 = ~n24174 & ~n24175;
  assign n24177 = ~n24165 & ~n24176;
  assign n24178 = ~n24173 & n24177;
  assign n24179 = n21961 & ~n22790;
  assign n24180 = ~n24178 & ~n24179;
  assign n24181 = ~n24170 & n24180;
  assign n24182 = ~n22819 & n22838;
  assign n24183 = n22819 & ~n22838;
  assign n24184 = ~n24182 & ~n24183;
  assign n24185 = n22823 & ~n22827;
  assign n24186 = ~n24184 & ~n24185;
  assign n24187 = ~n22823 & n22827;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = n24181 & n24188;
  assign n24190 = ~n24181 & ~n24188;
  assign n24191 = ~n24189 & ~n24190;
  assign n24192 = n22819 & ~n22833;
  assign n24193 = ~n22819 & n22833;
  assign n24194 = ~n4596 & ~n24193;
  assign n24195 = ~n24192 & ~n24194;
  assign n24196 = n5257 & ~n24195;
  assign n24197 = ~n5257 & ~n24192;
  assign n24198 = n4596 & n24197;
  assign n24199 = ~n24196 & ~n24198;
  assign n24200 = pi340 & ~n24199;
  assign n24201 = pi340 & n5257;
  assign n24202 = ~n22819 & ~n24201;
  assign n24203 = n22833 & n24202;
  assign n24204 = ~n24200 & ~n24203;
  assign n24205 = ~n21985 & ~n22697;
  assign n24206 = n21985 & n22697;
  assign n24207 = ~n24205 & ~n24206;
  assign n24208 = ~n22000 & n22701;
  assign n24209 = n22004 & ~n22709;
  assign n24210 = ~n22004 & n22709;
  assign n24211 = ~n24209 & ~n24210;
  assign n24212 = ~n24208 & ~n24211;
  assign n24213 = ~n24207 & n24212;
  assign n24214 = ~n21985 & n22697;
  assign n24215 = n21985 & ~n22697;
  assign n24216 = ~n24214 & ~n24215;
  assign n24217 = ~n22004 & ~n22709;
  assign n24218 = n22004 & n22709;
  assign n24219 = ~n24217 & ~n24218;
  assign n24220 = ~n24208 & ~n24219;
  assign n24221 = ~n24216 & n24220;
  assign n24222 = n22000 & ~n22701;
  assign n24223 = ~n24221 & ~n24222;
  assign n24224 = ~n24213 & n24223;
  assign n24225 = ~n22730 & n22749;
  assign n24226 = n22730 & ~n22749;
  assign n24227 = ~n24225 & ~n24226;
  assign n24228 = n22734 & ~n22738;
  assign n24229 = ~n24227 & ~n24228;
  assign n24230 = ~n22734 & n22738;
  assign n24231 = ~n24229 & ~n24230;
  assign n24232 = n24224 & n24231;
  assign n24233 = ~n24224 & ~n24231;
  assign n24234 = ~n24232 & ~n24233;
  assign n24235 = n22730 & ~n22744;
  assign n24236 = ~n22730 & n22744;
  assign n24237 = ~n9205 & ~n24236;
  assign n24238 = ~n24235 & ~n24237;
  assign n24239 = n10561 & ~n24238;
  assign n24240 = ~n10561 & ~n24235;
  assign n24241 = n9205 & n24240;
  assign n24242 = ~n24239 & ~n24241;
  assign n24243 = pi334 & ~n24242;
  assign n24244 = pi334 & n10561;
  assign n24245 = ~n22730 & ~n24244;
  assign n24246 = n22744 & n24245;
  assign n24247 = ~n24243 & ~n24246;
  assign n24248 = ~n22024 & n22032;
  assign n24249 = n22024 & ~n22032;
  assign n24250 = ~n22651 & ~n24249;
  assign n24251 = ~n24248 & ~n24250;
  assign n24252 = ~n22028 & n22676;
  assign n24253 = ~n22024 & ~n22651;
  assign n24254 = n22024 & n22651;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = n22032 & ~n24255;
  assign n24257 = n22024 & ~n22651;
  assign n24258 = ~n22024 & n22651;
  assign n24259 = ~n24257 & ~n24258;
  assign n24260 = ~n22032 & ~n24259;
  assign n24261 = ~n24256 & ~n24260;
  assign n24262 = n22028 & ~n22676;
  assign n24263 = ~n24261 & ~n24262;
  assign n24264 = ~n24252 & ~n24263;
  assign n24265 = n24251 & ~n24264;
  assign n24266 = ~n24251 & n24264;
  assign n24267 = ~n24265 & ~n24266;
  assign n24268 = pi329 & n13762;
  assign n24269 = ~n22047 & n22630;
  assign n24270 = n22047 & ~n22630;
  assign n24271 = ~n22637 & ~n24270;
  assign n24272 = ~n24269 & ~n24271;
  assign n24273 = ~n22047 & ~n22625;
  assign n24274 = n22047 & n22625;
  assign n24275 = ~n24273 & ~n24274;
  assign n24276 = ~n22051 & n22629;
  assign n24277 = ~n22612 & n22630;
  assign n24278 = n22612 & ~n22630;
  assign n24279 = ~n24277 & ~n24278;
  assign n24280 = ~n24276 & ~n24279;
  assign n24281 = ~n24275 & n24280;
  assign n24282 = ~n22047 & n22625;
  assign n24283 = n22047 & ~n22625;
  assign n24284 = ~n24282 & ~n24283;
  assign n24285 = n22612 & n22630;
  assign n24286 = ~n22612 & ~n22630;
  assign n24287 = ~n24285 & ~n24286;
  assign n24288 = ~n24276 & ~n24287;
  assign n24289 = ~n24284 & n24288;
  assign n24290 = n22051 & ~n22629;
  assign n24291 = ~n24289 & ~n24290;
  assign n24292 = ~n24281 & n24291;
  assign n24293 = n24272 & n24292;
  assign n24294 = ~n24272 & ~n24292;
  assign n24295 = ~n24293 & ~n24294;
  assign n24296 = ~n22060 & ~n22581;
  assign n24297 = ~n22589 & ~n24296;
  assign n24298 = ~n22064 & n22592;
  assign n24299 = ~n22060 & ~n22590;
  assign n24300 = n22060 & ~n22589;
  assign n24301 = ~n22581 & n24300;
  assign n24302 = ~n24299 & ~n24301;
  assign n24303 = n22064 & ~n22592;
  assign n24304 = ~n24302 & ~n24303;
  assign n24305 = ~n24298 & ~n24304;
  assign n24306 = ~n24297 & n24305;
  assign n24307 = n24297 & ~n24305;
  assign n24308 = ~n24306 & ~n24307;
  assign n24309 = ~n21446 & ~n22568;
  assign n24310 = ~n22567 & ~n24309;
  assign n24311 = pi133 & pi280;
  assign n24312 = ~n22130 & ~n22132;
  assign n24313 = ~n21041 & ~n22126;
  assign n24314 = ~n22129 & ~n22131;
  assign n24315 = n24313 & n24314;
  assign n24316 = ~n22135 & ~n24315;
  assign n24317 = ~n24312 & n24316;
  assign n24318 = ~n24312 & ~n24315;
  assign n24319 = pi280 & ~n24318;
  assign n24320 = pi132 & n24319;
  assign n24321 = ~n22149 & ~n24320;
  assign n24322 = ~n24317 & ~n24321;
  assign n24323 = pi132 & pi281;
  assign n24324 = n22102 & ~n22121;
  assign n24325 = ~n22092 & n22093;
  assign n24326 = pi129 & pi284;
  assign n24327 = pi285 & ~n24326;
  assign n24328 = pi128 & n24327;
  assign n24329 = pi128 & pi285;
  assign n24330 = pi284 & ~n24329;
  assign n24331 = pi129 & n24330;
  assign n24332 = ~n24328 & ~n24331;
  assign n24333 = ~pi283 & ~n24332;
  assign n24334 = ~pi130 & ~n24332;
  assign n24335 = pi283 & n24332;
  assign n24336 = pi130 & n24335;
  assign n24337 = ~n24334 & ~n24336;
  assign n24338 = ~pi129 & ~n24337;
  assign n24339 = ~n24333 & ~n24338;
  assign n24340 = ~n24325 & ~n24339;
  assign n24341 = n22092 & n22093;
  assign n24342 = ~n22092 & ~n22093;
  assign n24343 = ~n24341 & ~n24342;
  assign n24344 = pi129 & ~n24343;
  assign n24345 = pi283 & n24325;
  assign n24346 = ~n24344 & ~n24345;
  assign n24347 = ~n24332 & ~n24346;
  assign n24348 = pi283 & n22092;
  assign n24349 = ~n22093 & n24332;
  assign n24350 = n24348 & n24349;
  assign n24351 = ~n24347 & ~n24350;
  assign n24352 = pi130 & ~n24351;
  assign n24353 = ~n22093 & ~n24332;
  assign n24354 = n22092 & n24353;
  assign n24355 = n22092 & ~n22093;
  assign n24356 = pi283 & ~n24355;
  assign n24357 = pi129 & n24356;
  assign n24358 = ~n24325 & ~n24357;
  assign n24359 = n24332 & ~n24358;
  assign n24360 = ~n24354 & ~n24359;
  assign n24361 = ~pi130 & ~n24360;
  assign n24362 = n22093 & n24332;
  assign n24363 = ~pi283 & ~n22092;
  assign n24364 = n24362 & n24363;
  assign n24365 = ~n24361 & ~n24364;
  assign n24366 = ~n24352 & n24365;
  assign n24367 = ~n24340 & n24366;
  assign n24368 = ~pi282 & ~n24367;
  assign n24369 = ~pi131 & ~n24367;
  assign n24370 = pi282 & n24367;
  assign n24371 = pi131 & n24370;
  assign n24372 = ~n24369 & ~n24371;
  assign n24373 = ~pi130 & ~n24372;
  assign n24374 = ~n24368 & ~n24373;
  assign n24375 = ~n24324 & ~n24374;
  assign n24376 = pi282 & n24324;
  assign n24377 = ~n22102 & ~n22121;
  assign n24378 = n22102 & n22121;
  assign n24379 = ~n24377 & ~n24378;
  assign n24380 = pi130 & ~n24379;
  assign n24381 = ~n24376 & ~n24380;
  assign n24382 = ~n24367 & ~n24381;
  assign n24383 = n22121 & n24367;
  assign n24384 = n22103 & n24383;
  assign n24385 = ~n24382 & ~n24384;
  assign n24386 = pi131 & ~n24385;
  assign n24387 = ~n22102 & n22121;
  assign n24388 = pi282 & ~n24387;
  assign n24389 = pi130 & n24388;
  assign n24390 = ~n24324 & ~n24389;
  assign n24391 = n24367 & ~n24390;
  assign n24392 = n22121 & ~n24367;
  assign n24393 = ~n22102 & n24392;
  assign n24394 = ~n24391 & ~n24393;
  assign n24395 = ~pi131 & ~n24394;
  assign n24396 = ~pi282 & n22102;
  assign n24397 = ~n22121 & n24367;
  assign n24398 = n24396 & n24397;
  assign n24399 = ~n24395 & ~n24398;
  assign n24400 = ~n24386 & n24399;
  assign n24401 = ~n24375 & n24400;
  assign n24402 = ~n22129 & ~n22132;
  assign n24403 = ~n22126 & ~n24402;
  assign n24404 = n24401 & ~n24403;
  assign n24405 = ~n24401 & ~n24402;
  assign n24406 = ~n22126 & n24405;
  assign n24407 = ~n24404 & ~n24406;
  assign n24408 = n24323 & ~n24407;
  assign n24409 = n24401 & ~n24402;
  assign n24410 = ~n22126 & n24409;
  assign n24411 = ~n24401 & ~n24403;
  assign n24412 = ~n24410 & ~n24411;
  assign n24413 = ~n24323 & ~n24412;
  assign n24414 = ~n24408 & ~n24413;
  assign n24415 = n24322 & ~n24414;
  assign n24416 = ~n24322 & ~n24413;
  assign n24417 = ~n24408 & n24416;
  assign n24418 = ~n24415 & ~n24417;
  assign n24419 = ~n24311 & ~n24418;
  assign n24420 = ~n24322 & ~n24414;
  assign n24421 = n24322 & ~n24413;
  assign n24422 = ~n24408 & n24421;
  assign n24423 = ~n24420 & ~n24422;
  assign n24424 = pi280 & ~n24423;
  assign n24425 = pi133 & n24424;
  assign n24426 = ~n24419 & ~n24425;
  assign n24427 = ~n24317 & ~n24320;
  assign n24428 = ~n22149 & ~n24427;
  assign n24429 = ~n22146 & ~n24317;
  assign n24430 = ~n24320 & n24429;
  assign n24431 = ~n21058 & n24430;
  assign n24432 = ~n24428 & ~n24431;
  assign n24433 = ~n21079 & n24432;
  assign n24434 = n22077 & n24433;
  assign n24435 = ~pi279 & ~n24432;
  assign n24436 = ~n22185 & ~n24435;
  assign n24437 = pi278 & n24436;
  assign n24438 = ~n22078 & ~n24432;
  assign n24439 = pi279 & ~n24438;
  assign n24440 = ~n24437 & ~n24439;
  assign n24441 = pi133 & ~n24440;
  assign n24442 = ~n24434 & ~n24441;
  assign n24443 = n24426 & n24442;
  assign n24444 = ~n24426 & ~n24442;
  assign n24445 = ~n24443 & ~n24444;
  assign n24446 = ~n22159 & ~n22188;
  assign n24447 = ~pi133 & ~n22078;
  assign n24448 = ~n22185 & ~n24447;
  assign n24449 = n22159 & ~n24448;
  assign n24450 = ~n24446 & ~n24449;
  assign n24451 = ~pi134 & ~n24450;
  assign n24452 = ~n21079 & ~n22159;
  assign n24453 = n22077 & n24452;
  assign n24454 = ~n22078 & n22159;
  assign n24455 = ~n24453 & ~n24454;
  assign n24456 = ~pi278 & ~n24455;
  assign n24457 = ~n24451 & ~n24456;
  assign n24458 = pi134 & pi279;
  assign n24459 = pi133 & ~n22185;
  assign n24460 = ~n22078 & ~n24459;
  assign n24461 = n22159 & ~n24460;
  assign n24462 = ~n22159 & ~n24448;
  assign n24463 = ~n24461 & ~n24462;
  assign n24464 = pi278 & ~n24463;
  assign n24465 = pi134 & n24464;
  assign n24466 = n22198 & ~n24465;
  assign n24467 = n24458 & ~n24466;
  assign n24468 = n24457 & n24467;
  assign n24469 = n24457 & ~n24466;
  assign n24470 = ~n24458 & ~n24469;
  assign n24471 = ~n24468 & ~n24470;
  assign n24472 = ~n24445 & ~n24471;
  assign n24473 = n24426 & ~n24442;
  assign n24474 = ~n24426 & n24442;
  assign n24475 = ~n24473 & ~n24474;
  assign n24476 = ~n24458 & ~n24466;
  assign n24477 = n24457 & n24476;
  assign n24478 = n24458 & ~n24469;
  assign n24479 = ~n24477 & ~n24478;
  assign n24480 = ~n24475 & ~n24479;
  assign n24481 = ~n24472 & ~n24480;
  assign n24482 = ~n22201 & ~n22202;
  assign n24483 = n22201 & n22202;
  assign n24484 = ~n22207 & ~n24483;
  assign n24485 = ~n24482 & ~n24484;
  assign n24486 = n24481 & ~n24485;
  assign n24487 = ~n24481 & n24485;
  assign n24488 = ~n24486 & ~n24487;
  assign n24489 = pi136 & pi277;
  assign n24490 = pi135 & pi278;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = n24489 & n24490;
  assign n24493 = ~n24491 & ~n24492;
  assign n24494 = ~n24488 & ~n24493;
  assign n24495 = ~n24481 & ~n24485;
  assign n24496 = n24481 & n24485;
  assign n24497 = ~n24495 & ~n24496;
  assign n24498 = pi277 & ~n24490;
  assign n24499 = pi136 & n24498;
  assign n24500 = pi278 & ~n24489;
  assign n24501 = pi135 & n24500;
  assign n24502 = ~n24499 & ~n24501;
  assign n24503 = ~n24497 & ~n24502;
  assign n24504 = ~n24494 & ~n24503;
  assign n24505 = ~n22234 & ~n22238;
  assign n24506 = ~n22239 & ~n24505;
  assign n24507 = n24504 & n24506;
  assign n24508 = ~n24504 & ~n24506;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = pi137 & pi276;
  assign n24511 = n22218 & ~n22231;
  assign n24512 = ~n22227 & n24511;
  assign n24513 = ~n22218 & ~n22234;
  assign n24514 = ~n24512 & ~n24513;
  assign n24515 = ~n22073 & ~n24514;
  assign n24516 = ~n22218 & ~n22231;
  assign n24517 = ~n22227 & n24516;
  assign n24518 = n22218 & ~n22234;
  assign n24519 = ~n24517 & ~n24518;
  assign n24520 = pi276 & ~n24519;
  assign n24521 = pi136 & n24520;
  assign n24522 = ~n24515 & ~n24521;
  assign n24523 = ~n22250 & ~n24522;
  assign n24524 = n22250 & n24522;
  assign n24525 = n22228 & ~n24524;
  assign n24526 = ~n24523 & ~n24525;
  assign n24527 = n24510 & ~n24526;
  assign n24528 = ~n22228 & ~n24523;
  assign n24529 = ~n24524 & ~n24528;
  assign n24530 = ~n24510 & ~n24529;
  assign n24531 = ~n24527 & ~n24530;
  assign n24532 = ~n24509 & ~n24531;
  assign n24533 = n24504 & ~n24506;
  assign n24534 = ~n24504 & n24506;
  assign n24535 = ~n24533 & ~n24534;
  assign n24536 = ~n24510 & ~n24526;
  assign n24537 = n24510 & ~n24529;
  assign n24538 = ~n24536 & ~n24537;
  assign n24539 = ~n24535 & ~n24538;
  assign n24540 = ~n24532 & ~n24539;
  assign n24541 = ~n22254 & ~n22265;
  assign n24542 = n22254 & n22265;
  assign n24543 = ~n22259 & ~n24542;
  assign n24544 = ~n24541 & ~n24543;
  assign n24545 = ~n24540 & n24544;
  assign n24546 = n24540 & ~n24544;
  assign n24547 = ~n24545 & ~n24546;
  assign n24548 = pi139 & pi274;
  assign n24549 = pi138 & pi275;
  assign n24550 = n24548 & n24549;
  assign n24551 = ~n24548 & ~n24549;
  assign n24552 = ~n24550 & ~n24551;
  assign n24553 = ~n24547 & ~n24552;
  assign n24554 = n24540 & n24544;
  assign n24555 = ~n24540 & ~n24544;
  assign n24556 = ~n24554 & ~n24555;
  assign n24557 = pi274 & ~n24549;
  assign n24558 = pi139 & n24557;
  assign n24559 = pi275 & ~n24548;
  assign n24560 = pi138 & n24559;
  assign n24561 = ~n24558 & ~n24560;
  assign n24562 = ~n24556 & ~n24561;
  assign n24563 = ~n24553 & ~n24562;
  assign n24564 = ~n22283 & ~n22290;
  assign n24565 = ~n22278 & n24564;
  assign n24566 = ~n22291 & ~n24565;
  assign n24567 = n24563 & n24566;
  assign n24568 = ~n24563 & ~n24566;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = pi140 & pi273;
  assign n24571 = ~n22270 & ~n22283;
  assign n24572 = ~n22278 & n24571;
  assign n24573 = n22270 & ~n22286;
  assign n24574 = ~n24572 & ~n24573;
  assign n24575 = ~n22072 & ~n24574;
  assign n24576 = n22270 & ~n22283;
  assign n24577 = ~n22278 & n24576;
  assign n24578 = ~n22270 & ~n22286;
  assign n24579 = ~n24577 & ~n24578;
  assign n24580 = pi273 & ~n24579;
  assign n24581 = pi139 & n24580;
  assign n24582 = ~n24575 & ~n24581;
  assign n24583 = n22302 & n24582;
  assign n24584 = ~n22302 & ~n24582;
  assign n24585 = n22279 & ~n24584;
  assign n24586 = ~n24583 & ~n24585;
  assign n24587 = n24570 & ~n24586;
  assign n24588 = ~n22279 & ~n24583;
  assign n24589 = ~n24584 & ~n24588;
  assign n24590 = ~n24570 & ~n24589;
  assign n24591 = ~n24587 & ~n24590;
  assign n24592 = ~n24569 & ~n24591;
  assign n24593 = n24563 & ~n24566;
  assign n24594 = ~n24563 & n24566;
  assign n24595 = ~n24593 & ~n24594;
  assign n24596 = ~n24570 & ~n24586;
  assign n24597 = n24570 & ~n24589;
  assign n24598 = ~n24596 & ~n24597;
  assign n24599 = ~n24595 & ~n24598;
  assign n24600 = ~n24592 & ~n24599;
  assign n24601 = ~n22306 & ~n22317;
  assign n24602 = n22306 & n22317;
  assign n24603 = ~n22311 & ~n24602;
  assign n24604 = ~n24601 & ~n24603;
  assign n24605 = ~n24600 & n24604;
  assign n24606 = n24600 & ~n24604;
  assign n24607 = ~n24605 & ~n24606;
  assign n24608 = pi142 & pi271;
  assign n24609 = pi141 & pi272;
  assign n24610 = n24608 & n24609;
  assign n24611 = ~n24608 & ~n24609;
  assign n24612 = ~n24610 & ~n24611;
  assign n24613 = ~n24607 & ~n24612;
  assign n24614 = n24600 & n24604;
  assign n24615 = ~n24600 & ~n24604;
  assign n24616 = ~n24614 & ~n24615;
  assign n24617 = pi271 & ~n24609;
  assign n24618 = pi142 & n24617;
  assign n24619 = pi272 & ~n24608;
  assign n24620 = pi141 & n24619;
  assign n24621 = ~n24618 & ~n24620;
  assign n24622 = ~n24616 & ~n24621;
  assign n24623 = ~n24613 & ~n24622;
  assign n24624 = ~n22335 & ~n22342;
  assign n24625 = ~n22330 & n24624;
  assign n24626 = ~n22343 & ~n24625;
  assign n24627 = n24623 & ~n24626;
  assign n24628 = ~n24623 & n24626;
  assign n24629 = ~n24627 & ~n24628;
  assign n24630 = pi143 & pi270;
  assign n24631 = ~n22322 & ~n22335;
  assign n24632 = ~n22330 & n24631;
  assign n24633 = n22322 & ~n22338;
  assign n24634 = ~n24632 & ~n24633;
  assign n24635 = ~n22071 & ~n24634;
  assign n24636 = n22322 & ~n22335;
  assign n24637 = ~n22330 & n24636;
  assign n24638 = ~n22322 & ~n22338;
  assign n24639 = ~n24637 & ~n24638;
  assign n24640 = pi270 & ~n24639;
  assign n24641 = pi142 & n24640;
  assign n24642 = ~n24635 & ~n24641;
  assign n24643 = n22354 & n24642;
  assign n24644 = ~n22354 & ~n24642;
  assign n24645 = n22331 & ~n24644;
  assign n24646 = ~n24643 & ~n24645;
  assign n24647 = n24630 & ~n24646;
  assign n24648 = ~n22331 & ~n24643;
  assign n24649 = ~n24644 & ~n24648;
  assign n24650 = ~n24630 & ~n24649;
  assign n24651 = ~n24647 & ~n24650;
  assign n24652 = ~n24629 & ~n24651;
  assign n24653 = n24623 & n24626;
  assign n24654 = ~n24623 & ~n24626;
  assign n24655 = ~n24653 & ~n24654;
  assign n24656 = ~n24630 & ~n24646;
  assign n24657 = n24630 & ~n24649;
  assign n24658 = ~n24656 & ~n24657;
  assign n24659 = ~n24655 & ~n24658;
  assign n24660 = ~n24652 & ~n24659;
  assign n24661 = n22358 & ~n22369;
  assign n24662 = ~n22358 & n22369;
  assign n24663 = ~n22360 & ~n24662;
  assign n24664 = ~n24661 & ~n24663;
  assign n24665 = ~n24660 & n24664;
  assign n24666 = n24660 & ~n24664;
  assign n24667 = ~n24665 & ~n24666;
  assign n24668 = pi145 & pi268;
  assign n24669 = pi144 & pi269;
  assign n24670 = n24668 & n24669;
  assign n24671 = ~n24668 & ~n24669;
  assign n24672 = ~n24670 & ~n24671;
  assign n24673 = ~n24667 & ~n24672;
  assign n24674 = n24660 & n24664;
  assign n24675 = ~n24660 & ~n24664;
  assign n24676 = ~n24674 & ~n24675;
  assign n24677 = pi268 & ~n24669;
  assign n24678 = pi145 & n24677;
  assign n24679 = pi269 & ~n24668;
  assign n24680 = pi144 & n24679;
  assign n24681 = ~n24678 & ~n24680;
  assign n24682 = ~n24676 & ~n24681;
  assign n24683 = ~n24673 & ~n24682;
  assign n24684 = ~n22390 & ~n22394;
  assign n24685 = ~n22395 & ~n24684;
  assign n24686 = n24683 & ~n24685;
  assign n24687 = ~n24683 & n24685;
  assign n24688 = ~n24686 & ~n24687;
  assign n24689 = pi146 & pi267;
  assign n24690 = ~n22374 & ~n22387;
  assign n24691 = ~n22383 & n24690;
  assign n24692 = n22374 & ~n22390;
  assign n24693 = ~n24691 & ~n24692;
  assign n24694 = ~n22070 & ~n24693;
  assign n24695 = n22374 & ~n22387;
  assign n24696 = ~n22383 & n24695;
  assign n24697 = ~n22374 & ~n22390;
  assign n24698 = ~n24696 & ~n24697;
  assign n24699 = pi267 & ~n24698;
  assign n24700 = pi145 & n24699;
  assign n24701 = ~n24694 & ~n24700;
  assign n24702 = n22406 & n24701;
  assign n24703 = ~n22406 & ~n24701;
  assign n24704 = n22384 & ~n24703;
  assign n24705 = ~n24702 & ~n24704;
  assign n24706 = n24689 & ~n24705;
  assign n24707 = ~n22384 & ~n24702;
  assign n24708 = ~n24703 & ~n24707;
  assign n24709 = ~n24689 & ~n24708;
  assign n24710 = ~n24706 & ~n24709;
  assign n24711 = ~n24688 & ~n24710;
  assign n24712 = n24683 & n24685;
  assign n24713 = ~n24683 & ~n24685;
  assign n24714 = ~n24712 & ~n24713;
  assign n24715 = ~n24689 & ~n24705;
  assign n24716 = n24689 & ~n24708;
  assign n24717 = ~n24715 & ~n24716;
  assign n24718 = ~n24714 & ~n24717;
  assign n24719 = ~n24711 & ~n24718;
  assign n24720 = n22410 & ~n22421;
  assign n24721 = ~n22410 & n22421;
  assign n24722 = ~n22412 & ~n24721;
  assign n24723 = ~n24720 & ~n24722;
  assign n24724 = ~n24719 & n24723;
  assign n24725 = n24719 & ~n24723;
  assign n24726 = ~n24724 & ~n24725;
  assign n24727 = pi148 & pi265;
  assign n24728 = pi147 & pi266;
  assign n24729 = n24727 & n24728;
  assign n24730 = ~n24727 & ~n24728;
  assign n24731 = ~n24729 & ~n24730;
  assign n24732 = ~n24726 & ~n24731;
  assign n24733 = n24719 & n24723;
  assign n24734 = ~n24719 & ~n24723;
  assign n24735 = ~n24733 & ~n24734;
  assign n24736 = pi265 & ~n24728;
  assign n24737 = pi148 & n24736;
  assign n24738 = pi266 & ~n24727;
  assign n24739 = pi147 & n24738;
  assign n24740 = ~n24737 & ~n24739;
  assign n24741 = ~n24735 & ~n24740;
  assign n24742 = ~n24732 & ~n24741;
  assign n24743 = ~n22442 & ~n22446;
  assign n24744 = ~n22447 & ~n24743;
  assign n24745 = n24742 & n24744;
  assign n24746 = ~n24742 & ~n24744;
  assign n24747 = ~n24745 & ~n24746;
  assign n24748 = pi149 & pi264;
  assign n24749 = n22426 & ~n22439;
  assign n24750 = ~n22435 & n24749;
  assign n24751 = ~n22426 & ~n22442;
  assign n24752 = ~n24750 & ~n24751;
  assign n24753 = ~n22069 & ~n24752;
  assign n24754 = ~n22426 & ~n22439;
  assign n24755 = ~n22435 & n24754;
  assign n24756 = n22426 & ~n22442;
  assign n24757 = ~n24755 & ~n24756;
  assign n24758 = pi264 & ~n24757;
  assign n24759 = pi148 & n24758;
  assign n24760 = ~n24753 & ~n24759;
  assign n24761 = ~n22458 & ~n24760;
  assign n24762 = n22458 & n24760;
  assign n24763 = n22436 & ~n24762;
  assign n24764 = ~n24761 & ~n24763;
  assign n24765 = n24748 & ~n24764;
  assign n24766 = ~n22436 & ~n24761;
  assign n24767 = ~n24762 & ~n24766;
  assign n24768 = ~n24748 & ~n24767;
  assign n24769 = ~n24765 & ~n24768;
  assign n24770 = ~n24747 & ~n24769;
  assign n24771 = n24742 & ~n24744;
  assign n24772 = ~n24742 & n24744;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = ~n24748 & ~n24764;
  assign n24775 = n24748 & ~n24767;
  assign n24776 = ~n24774 & ~n24775;
  assign n24777 = ~n24773 & ~n24776;
  assign n24778 = ~n24770 & ~n24777;
  assign n24779 = ~n22461 & ~n22462;
  assign n24780 = n22461 & n22462;
  assign n24781 = ~n22467 & ~n24780;
  assign n24782 = ~n24779 & ~n24781;
  assign n24783 = ~n24778 & n24782;
  assign n24784 = n24778 & ~n24782;
  assign n24785 = ~n24783 & ~n24784;
  assign n24786 = pi151 & pi262;
  assign n24787 = pi150 & pi263;
  assign n24788 = n24786 & n24787;
  assign n24789 = ~n24786 & ~n24787;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = ~n24785 & ~n24790;
  assign n24792 = n24778 & n24782;
  assign n24793 = ~n24778 & ~n24782;
  assign n24794 = ~n24792 & ~n24793;
  assign n24795 = pi262 & ~n24787;
  assign n24796 = pi151 & n24795;
  assign n24797 = pi263 & ~n24786;
  assign n24798 = pi150 & n24797;
  assign n24799 = ~n24796 & ~n24798;
  assign n24800 = ~n24794 & ~n24799;
  assign n24801 = ~n24791 & ~n24800;
  assign n24802 = ~pi261 & ~n22478;
  assign n24803 = pi260 & ~n24802;
  assign n24804 = pi151 & n24803;
  assign n24805 = n21426 & ~n22495;
  assign n24806 = ~n24804 & ~n24805;
  assign n24807 = n22483 & ~n24806;
  assign n24808 = pi261 & n22478;
  assign n24809 = n21426 & n24803;
  assign n24810 = ~n24808 & ~n24809;
  assign n24811 = pi151 & ~n24810;
  assign n24812 = ~n24807 & ~n24811;
  assign n24813 = n24801 & n24812;
  assign n24814 = ~n24801 & ~n24812;
  assign n24815 = ~n24813 & ~n24814;
  assign n24816 = pi152 & pi261;
  assign n24817 = pi151 & ~n1377;
  assign n24818 = n22478 & ~n24817;
  assign n24819 = ~pi260 & pi261;
  assign n24820 = pi151 & ~n22478;
  assign n24821 = n24819 & n24820;
  assign n24822 = ~n24818 & ~n24821;
  assign n24823 = ~n22484 & ~n24822;
  assign n24824 = ~pi261 & n22478;
  assign n24825 = ~n22480 & ~n24824;
  assign n24826 = ~n21426 & ~n24825;
  assign n24827 = ~n22483 & n24826;
  assign n24828 = pi260 & ~pi261;
  assign n24829 = ~n22478 & n24828;
  assign n24830 = ~pi260 & ~n21426;
  assign n24831 = pi261 & ~n24830;
  assign n24832 = n22478 & n24831;
  assign n24833 = ~n24829 & ~n24832;
  assign n24834 = pi151 & ~n24833;
  assign n24835 = n21426 & n22495;
  assign n24836 = ~n24834 & ~n24835;
  assign n24837 = n22483 & ~n24836;
  assign n24838 = ~n24802 & ~n24808;
  assign n24839 = pi260 & ~n24838;
  assign n24840 = pi151 & n24839;
  assign n24841 = n21426 & n24840;
  assign n24842 = ~n24837 & ~n24841;
  assign n24843 = ~n24827 & n24842;
  assign n24844 = ~n24823 & n24843;
  assign n24845 = ~n22506 & ~n24844;
  assign n24846 = n22506 & n24844;
  assign n24847 = n22482 & ~n24846;
  assign n24848 = ~n24845 & ~n24847;
  assign n24849 = n24816 & ~n24848;
  assign n24850 = ~n22482 & ~n24845;
  assign n24851 = ~n24846 & ~n24850;
  assign n24852 = ~n24816 & ~n24851;
  assign n24853 = ~n24849 & ~n24852;
  assign n24854 = ~n24815 & ~n24853;
  assign n24855 = n24801 & ~n24812;
  assign n24856 = ~n24801 & n24812;
  assign n24857 = ~n24855 & ~n24856;
  assign n24858 = ~n24816 & ~n24848;
  assign n24859 = n24816 & ~n24851;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = ~n24857 & ~n24860;
  assign n24862 = ~n24854 & ~n24861;
  assign n24863 = pi259 & n22518;
  assign n24864 = pi153 & pi259;
  assign n24865 = ~n22518 & ~n24864;
  assign n24866 = ~n22509 & ~n24865;
  assign n24867 = ~n24863 & ~n24866;
  assign n24868 = n24862 & n24867;
  assign n24869 = ~n24862 & ~n24867;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = pi154 & pi259;
  assign n24872 = pi153 & pi260;
  assign n24873 = ~n24871 & ~n24872;
  assign n24874 = n24871 & n24872;
  assign n24875 = ~n24873 & ~n24874;
  assign n24876 = ~pi259 & n22518;
  assign n24877 = pi259 & ~n22518;
  assign n24878 = pi153 & n24877;
  assign n24879 = ~n24876 & ~n24878;
  assign n24880 = ~n22535 & ~n24879;
  assign n24881 = ~n24863 & ~n24865;
  assign n24882 = ~n22509 & ~n24881;
  assign n24883 = ~n24880 & ~n24882;
  assign n24884 = n22519 & ~n24883;
  assign n24885 = pi155 & pi258;
  assign n24886 = n24884 & n24885;
  assign n24887 = ~n24884 & ~n24885;
  assign n24888 = ~n24886 & ~n24887;
  assign n24889 = ~n24875 & ~n24888;
  assign n24890 = n24871 & ~n24872;
  assign n24891 = ~n24871 & n24872;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n24884 & n24885;
  assign n24894 = n24884 & ~n24885;
  assign n24895 = ~n24893 & ~n24894;
  assign n24896 = ~n24892 & ~n24895;
  assign n24897 = ~n24889 & ~n24896;
  assign n24898 = ~n24870 & ~n24897;
  assign n24899 = n24862 & ~n24867;
  assign n24900 = ~n24862 & n24867;
  assign n24901 = ~n24899 & ~n24900;
  assign n24902 = ~n24888 & ~n24892;
  assign n24903 = ~n24875 & ~n24895;
  assign n24904 = ~n24902 & ~n24903;
  assign n24905 = ~n24901 & ~n24904;
  assign n24906 = ~n24898 & ~n24905;
  assign n24907 = n24310 & ~n24906;
  assign n24908 = ~n24310 & n24906;
  assign n24909 = n22545 & n24908;
  assign n24910 = ~n24907 & ~n24909;
  assign n24911 = ~n22557 & ~n24910;
  assign n24912 = ~n24310 & ~n24906;
  assign n24913 = n24310 & n24906;
  assign n24914 = ~n22545 & n24913;
  assign n24915 = ~n24912 & ~n24914;
  assign n24916 = n22557 & ~n24915;
  assign n24917 = ~n22545 & ~n24310;
  assign n24918 = n22545 & n24310;
  assign n24919 = ~n24917 & ~n24918;
  assign n24920 = ~n24906 & ~n24919;
  assign n24921 = ~n24916 & ~n24920;
  assign n24922 = ~n24911 & n24921;
  assign n24923 = pi322 & ~n24922;
  assign n24924 = n22545 & ~n24310;
  assign n24925 = ~n22545 & n24310;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = n22557 & ~n24926;
  assign n24928 = ~n22557 & ~n24919;
  assign n24929 = ~n24927 & ~n24928;
  assign n24930 = pi323 & ~n24929;
  assign n24931 = ~n24923 & ~n24930;
  assign n24932 = n22557 & n24924;
  assign n24933 = ~n24928 & ~n24932;
  assign n24934 = ~n24906 & ~n24933;
  assign n24935 = ~n22545 & n22557;
  assign n24936 = n24913 & n24935;
  assign n24937 = ~n24934 & ~n24936;
  assign n24938 = pi323 & ~n24937;
  assign n24939 = pi322 & n24938;
  assign n24940 = ~n24931 & ~n24939;
  assign n24941 = pi325 & n19970;
  assign n24942 = pi324 & n21479;
  assign n24943 = n24941 & n24942;
  assign n24944 = ~n24941 & ~n24942;
  assign n24945 = ~n24943 & ~n24944;
  assign n24946 = ~n24940 & ~n24945;
  assign n24947 = ~n24941 & n24942;
  assign n24948 = n24941 & ~n24942;
  assign n24949 = ~n24947 & ~n24948;
  assign n24950 = ~n24939 & ~n24949;
  assign n24951 = ~n24931 & n24950;
  assign n24952 = ~n24946 & ~n24951;
  assign n24953 = ~n24308 & ~n24952;
  assign n24954 = ~n24297 & ~n24305;
  assign n24955 = n24297 & n24305;
  assign n24956 = ~n24954 & ~n24955;
  assign n24957 = ~n24940 & ~n24949;
  assign n24958 = ~n24939 & ~n24945;
  assign n24959 = ~n24931 & n24958;
  assign n24960 = ~n24957 & ~n24959;
  assign n24961 = ~n24956 & ~n24960;
  assign n24962 = ~n24953 & ~n24961;
  assign n24963 = n22591 & ~n22625;
  assign n24964 = ~n22589 & ~n22592;
  assign n24965 = ~n22581 & n24964;
  assign n24966 = n19970 & ~n22590;
  assign n24967 = pi324 & n24966;
  assign n24968 = ~n24965 & ~n24967;
  assign n24969 = ~n22606 & ~n24968;
  assign n24970 = ~n22590 & ~n22592;
  assign n24971 = n22590 & n22592;
  assign n24972 = ~n24970 & ~n24971;
  assign n24973 = ~n22067 & ~n24972;
  assign n24974 = ~n24969 & ~n24973;
  assign n24975 = ~n22591 & n22625;
  assign n24976 = ~n24974 & ~n24975;
  assign n24977 = ~n24963 & ~n24976;
  assign n24978 = n24962 & n24977;
  assign n24979 = ~n24962 & ~n24977;
  assign n24980 = ~n24978 & ~n24979;
  assign n24981 = pi327 & n19539;
  assign n24982 = pi326 & n19557;
  assign n24983 = n24981 & n24982;
  assign n24984 = ~n24981 & ~n24982;
  assign n24985 = ~n24983 & ~n24984;
  assign n24986 = ~n24980 & ~n24985;
  assign n24987 = ~n24962 & n24977;
  assign n24988 = n24962 & ~n24977;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 = ~n24981 & n24982;
  assign n24991 = n24981 & ~n24982;
  assign n24992 = ~n24990 & ~n24991;
  assign n24993 = ~n24989 & ~n24992;
  assign n24994 = ~n24986 & ~n24993;
  assign n24995 = ~n24295 & ~n24994;
  assign n24996 = n24272 & ~n24292;
  assign n24997 = ~n24272 & n24292;
  assign n24998 = ~n24996 & ~n24997;
  assign n24999 = ~n24985 & ~n24989;
  assign n25000 = ~n24980 & ~n24992;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = ~n24998 & ~n25001;
  assign n25003 = ~n24995 & ~n25002;
  assign n25004 = ~n24268 & n25003;
  assign n25005 = n24268 & ~n25003;
  assign n25006 = ~n25004 & ~n25005;
  assign n25007 = n18461 & ~n25006;
  assign n25008 = pi328 & n25007;
  assign n25009 = pi328 & n18461;
  assign n25010 = n24268 & n25003;
  assign n25011 = ~n24268 & ~n25003;
  assign n25012 = ~n25010 & ~n25011;
  assign n25013 = ~n25009 & ~n25012;
  assign n25014 = ~n25008 & ~n25013;
  assign n25015 = ~n24267 & ~n25014;
  assign n25016 = n24251 & n24264;
  assign n25017 = ~n24251 & ~n24264;
  assign n25018 = ~n25016 & ~n25017;
  assign n25019 = n18461 & ~n25012;
  assign n25020 = pi328 & n25019;
  assign n25021 = ~n25006 & ~n25009;
  assign n25022 = ~n25020 & ~n25021;
  assign n25023 = ~n25018 & ~n25022;
  assign n25024 = ~n25015 & ~n25023;
  assign n25025 = ~n21985 & n22004;
  assign n25026 = n21985 & ~n22004;
  assign n25027 = ~n22697 & ~n25026;
  assign n25028 = ~n25025 & ~n25027;
  assign n25029 = n25024 & n25028;
  assign n25030 = ~n25024 & ~n25028;
  assign n25031 = ~n25029 & ~n25030;
  assign n25032 = pi331 & n11711;
  assign n25033 = n20933 & ~n21978;
  assign n25034 = ~n20933 & ~n21968;
  assign n25035 = ~n25033 & ~n25034;
  assign n25036 = ~n22657 & ~n25035;
  assign n25037 = ~n22660 & ~n25036;
  assign n25038 = n12917 & ~n22654;
  assign n25039 = pi329 & n25038;
  assign n25040 = ~n22676 & ~n22683;
  assign n25041 = ~n25039 & ~n25040;
  assign n25042 = ~n22031 & ~n25041;
  assign n25043 = n12917 & ~n22683;
  assign n25044 = pi329 & n25043;
  assign n25045 = ~n22654 & ~n22676;
  assign n25046 = ~n25044 & ~n25045;
  assign n25047 = ~n22692 & ~n25046;
  assign n25048 = ~n25042 & ~n25047;
  assign n25049 = n25037 & ~n25048;
  assign n25050 = ~n25037 & n25048;
  assign n25051 = ~n11711 & ~n25050;
  assign n25052 = ~n25049 & ~n25051;
  assign n25053 = n12917 & ~n25052;
  assign n25054 = ~n12917 & ~n25049;
  assign n25055 = n11711 & n25054;
  assign n25056 = ~n25053 & ~n25055;
  assign n25057 = pi330 & ~n25056;
  assign n25058 = pi330 & n12917;
  assign n25059 = n25048 & ~n25058;
  assign n25060 = ~n25037 & n25059;
  assign n25061 = ~n25057 & ~n25060;
  assign n25062 = ~n25032 & n25061;
  assign n25063 = n25032 & ~n25061;
  assign n25064 = ~n25062 & ~n25063;
  assign n25065 = pi333 & n11366;
  assign n25066 = pi332 & n11384;
  assign n25067 = ~n22702 & n22704;
  assign n25068 = ~n25066 & ~n25067;
  assign n25069 = n22004 & n25068;
  assign n25070 = n22702 & ~n22704;
  assign n25071 = n25066 & ~n25070;
  assign n25072 = ~n22004 & n25071;
  assign n25073 = ~n25069 & ~n25072;
  assign n25074 = ~n24207 & ~n25073;
  assign n25075 = n22004 & n25071;
  assign n25076 = ~n22004 & n25068;
  assign n25077 = ~n25075 & ~n25076;
  assign n25078 = ~n24216 & ~n25077;
  assign n25079 = ~n22704 & ~n25066;
  assign n25080 = n22702 & n25079;
  assign n25081 = n22704 & n25066;
  assign n25082 = ~n22702 & n25081;
  assign n25083 = ~n25080 & ~n25082;
  assign n25084 = ~n25078 & n25083;
  assign n25085 = ~n25074 & n25084;
  assign n25086 = n25065 & ~n25085;
  assign n25087 = ~n25065 & n25085;
  assign n25088 = ~n25086 & ~n25087;
  assign n25089 = ~n25064 & ~n25088;
  assign n25090 = n25032 & n25061;
  assign n25091 = ~n25032 & ~n25061;
  assign n25092 = ~n25090 & ~n25091;
  assign n25093 = ~n25065 & ~n25085;
  assign n25094 = n25065 & n25085;
  assign n25095 = ~n25093 & ~n25094;
  assign n25096 = ~n25092 & ~n25095;
  assign n25097 = ~n25089 & ~n25096;
  assign n25098 = ~n25031 & ~n25097;
  assign n25099 = n25024 & ~n25028;
  assign n25100 = ~n25024 & n25028;
  assign n25101 = ~n25099 & ~n25100;
  assign n25102 = ~n25088 & ~n25092;
  assign n25103 = ~n25064 & ~n25095;
  assign n25104 = ~n25102 & ~n25103;
  assign n25105 = ~n25101 & ~n25104;
  assign n25106 = ~n25098 & ~n25105;
  assign n25107 = n24247 & n25106;
  assign n25108 = ~n24247 & ~n25106;
  assign n25109 = ~n25107 & ~n25108;
  assign n25110 = n9205 & ~n25109;
  assign n25111 = pi335 & n25110;
  assign n25112 = pi335 & n9205;
  assign n25113 = ~n24247 & n25106;
  assign n25114 = n24247 & ~n25106;
  assign n25115 = ~n25113 & ~n25114;
  assign n25116 = ~n25112 & ~n25115;
  assign n25117 = ~n25111 & ~n25116;
  assign n25118 = ~n24234 & ~n25117;
  assign n25119 = n24224 & ~n24231;
  assign n25120 = ~n24224 & n24231;
  assign n25121 = ~n25119 & ~n25120;
  assign n25122 = n9205 & ~n25115;
  assign n25123 = pi335 & n25122;
  assign n25124 = ~n25109 & ~n25112;
  assign n25125 = ~n25123 & ~n25124;
  assign n25126 = ~n25121 & ~n25125;
  assign n25127 = ~n25118 & ~n25126;
  assign n25128 = ~n21946 & n21965;
  assign n25129 = n21946 & ~n21965;
  assign n25130 = ~n22786 & ~n25129;
  assign n25131 = ~n25128 & ~n25130;
  assign n25132 = n25127 & n25131;
  assign n25133 = ~n25127 & ~n25131;
  assign n25134 = ~n25132 & ~n25133;
  assign n25135 = pi337 & n5973;
  assign n25136 = ~n22752 & ~n22774;
  assign n25137 = ~n22737 & n25136;
  assign n25138 = ~n22772 & ~n22774;
  assign n25139 = ~n22781 & n25138;
  assign n25140 = ~n22773 & ~n25139;
  assign n25141 = ~n25137 & n25140;
  assign n25142 = pi336 & n6556;
  assign n25143 = n25141 & ~n25142;
  assign n25144 = n6556 & ~n25141;
  assign n25145 = pi336 & n25144;
  assign n25146 = ~n25143 & ~n25145;
  assign n25147 = ~n25135 & n25146;
  assign n25148 = n25135 & ~n25146;
  assign n25149 = ~n25147 & ~n25148;
  assign n25150 = pi339 & n5714;
  assign n25151 = pi338 & n5732;
  assign n25152 = ~n22791 & n22793;
  assign n25153 = ~n25151 & ~n25152;
  assign n25154 = n21965 & n25153;
  assign n25155 = n22791 & ~n22793;
  assign n25156 = n25151 & ~n25155;
  assign n25157 = ~n21965 & n25156;
  assign n25158 = ~n25154 & ~n25157;
  assign n25159 = ~n24164 & ~n25158;
  assign n25160 = n21965 & n25156;
  assign n25161 = ~n21965 & n25153;
  assign n25162 = ~n25160 & ~n25161;
  assign n25163 = ~n24173 & ~n25162;
  assign n25164 = ~n22793 & ~n25151;
  assign n25165 = n22791 & n25164;
  assign n25166 = n22793 & n25151;
  assign n25167 = ~n22791 & n25166;
  assign n25168 = ~n25165 & ~n25167;
  assign n25169 = ~n25163 & n25168;
  assign n25170 = ~n25159 & n25169;
  assign n25171 = n25150 & ~n25170;
  assign n25172 = ~n25150 & n25170;
  assign n25173 = ~n25171 & ~n25172;
  assign n25174 = ~n25149 & ~n25173;
  assign n25175 = n25135 & n25146;
  assign n25176 = ~n25135 & ~n25146;
  assign n25177 = ~n25175 & ~n25176;
  assign n25178 = ~n25150 & ~n25170;
  assign n25179 = n25150 & n25170;
  assign n25180 = ~n25178 & ~n25179;
  assign n25181 = ~n25177 & ~n25180;
  assign n25182 = ~n25174 & ~n25181;
  assign n25183 = ~n25134 & ~n25182;
  assign n25184 = n25127 & ~n25131;
  assign n25185 = ~n25127 & n25131;
  assign n25186 = ~n25184 & ~n25185;
  assign n25187 = ~n25173 & ~n25177;
  assign n25188 = ~n25149 & ~n25180;
  assign n25189 = ~n25187 & ~n25188;
  assign n25190 = ~n25186 & ~n25189;
  assign n25191 = ~n25183 & ~n25190;
  assign n25192 = n24204 & n25191;
  assign n25193 = ~n24204 & ~n25191;
  assign n25194 = ~n25192 & ~n25193;
  assign n25195 = n4596 & ~n25194;
  assign n25196 = pi341 & n25195;
  assign n25197 = pi341 & n4596;
  assign n25198 = ~n24204 & n25191;
  assign n25199 = n24204 & ~n25191;
  assign n25200 = ~n25198 & ~n25199;
  assign n25201 = ~n25197 & ~n25200;
  assign n25202 = ~n25196 & ~n25201;
  assign n25203 = ~n24191 & ~n25202;
  assign n25204 = n24181 & ~n24188;
  assign n25205 = ~n24181 & n24188;
  assign n25206 = ~n25204 & ~n25205;
  assign n25207 = n4596 & ~n25200;
  assign n25208 = pi341 & n25207;
  assign n25209 = ~n25194 & ~n25197;
  assign n25210 = ~n25208 & ~n25209;
  assign n25211 = ~n25206 & ~n25210;
  assign n25212 = ~n25203 & ~n25211;
  assign n25213 = ~n21913 & n21926;
  assign n25214 = n21913 & ~n21926;
  assign n25215 = ~n22875 & ~n25214;
  assign n25216 = ~n25213 & ~n25215;
  assign n25217 = n25212 & n25216;
  assign n25218 = ~n25212 & ~n25216;
  assign n25219 = ~n25217 & ~n25218;
  assign n25220 = pi343 & n2464;
  assign n25221 = ~n22841 & ~n22863;
  assign n25222 = ~n22826 & n25221;
  assign n25223 = ~n22861 & ~n22863;
  assign n25224 = ~n22870 & n25223;
  assign n25225 = ~n22862 & ~n25224;
  assign n25226 = ~n25222 & n25225;
  assign n25227 = pi342 & n2887;
  assign n25228 = n25226 & ~n25227;
  assign n25229 = n2887 & ~n25226;
  assign n25230 = pi342 & n25229;
  assign n25231 = ~n25228 & ~n25230;
  assign n25232 = ~n25220 & n25231;
  assign n25233 = n25220 & ~n25231;
  assign n25234 = ~n25232 & ~n25233;
  assign n25235 = pi344 & n2091;
  assign n25236 = n1729 & ~n22881;
  assign n25237 = pi344 & n25236;
  assign n25238 = n21926 & ~n24129;
  assign n25239 = ~n21926 & ~n24138;
  assign n25240 = ~n25238 & ~n25239;
  assign n25241 = n22881 & ~n22884;
  assign n25242 = ~n25240 & ~n25241;
  assign n25243 = ~n25237 & ~n25242;
  assign n25244 = n25235 & n25243;
  assign n25245 = ~n25235 & ~n25243;
  assign n25246 = ~n25244 & ~n25245;
  assign n25247 = ~n25234 & ~n25246;
  assign n25248 = n25220 & n25231;
  assign n25249 = ~n25220 & ~n25231;
  assign n25250 = ~n25248 & ~n25249;
  assign n25251 = ~n25235 & n25243;
  assign n25252 = n25235 & ~n25243;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = ~n25250 & ~n25253;
  assign n25255 = ~n25247 & ~n25254;
  assign n25256 = ~n25219 & ~n25255;
  assign n25257 = n25212 & ~n25216;
  assign n25258 = ~n25212 & n25216;
  assign n25259 = ~n25257 & ~n25258;
  assign n25260 = ~n25246 & ~n25250;
  assign n25261 = ~n25234 & ~n25253;
  assign n25262 = ~n25260 & ~n25261;
  assign n25263 = ~n25259 & ~n25262;
  assign n25264 = ~n25256 & ~n25263;
  assign n25265 = ~n24161 & n25264;
  assign n25266 = n24161 & ~n25264;
  assign n25267 = ~n25265 & ~n25266;
  assign n25268 = pi347 & ~n1256;
  assign n25269 = ~n22907 & n24151;
  assign n25270 = ~n24148 & ~n25269;
  assign n25271 = n1442 & n25270;
  assign n25272 = pi346 & n25271;
  assign n25273 = pi346 & n1442;
  assign n25274 = ~n25270 & ~n25273;
  assign n25275 = ~n25272 & ~n25274;
  assign n25276 = n25268 & ~n25275;
  assign n25277 = ~n25268 & n25275;
  assign n25278 = ~n25276 & ~n25277;
  assign n25279 = ~n25267 & ~n25278;
  assign n25280 = n24161 & n25264;
  assign n25281 = ~n24161 & ~n25264;
  assign n25282 = ~n25280 & ~n25281;
  assign n25283 = ~n25268 & ~n25275;
  assign n25284 = n25268 & n25275;
  assign n25285 = ~n25283 & ~n25284;
  assign n25286 = ~n25282 & ~n25285;
  assign n25287 = ~n25279 & ~n25286;
  assign n25288 = ~n24160 & ~n25287;
  assign n25289 = n24146 & ~n24157;
  assign n25290 = ~n24146 & n24157;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = ~n25278 & ~n25282;
  assign n25293 = ~n25267 & ~n25285;
  assign n25294 = ~n25292 & ~n25293;
  assign n25295 = ~n25291 & ~n25294;
  assign n25296 = ~n25288 & ~n25295;
  assign n25297 = n24126 & ~n25296;
  assign n25298 = ~n24126 & n25296;
  assign n25299 = ~n25297 & ~n25298;
  assign n25300 = ~n22935 & ~n23556;
  assign n25301 = n22935 & n23556;
  assign n25302 = ~pi284 & ~n25301;
  assign n25303 = ~n25300 & ~n25302;
  assign n25304 = ~pi285 & n25303;
  assign n25305 = pi285 & ~n25303;
  assign n25306 = ~n25304 & ~n25305;
  assign n25307 = n1156 & ~n25306;
  assign n25308 = pi349 & n25307;
  assign n25309 = pi349 & n1156;
  assign n25310 = ~pi285 & ~n25303;
  assign n25311 = pi285 & n25303;
  assign n25312 = ~n25310 & ~n25311;
  assign n25313 = ~n25309 & ~n25312;
  assign n25314 = ~n25308 & ~n25313;
  assign n25315 = ~n25299 & ~n25314;
  assign n25316 = n24126 & n25296;
  assign n25317 = ~n24126 & ~n25296;
  assign n25318 = ~n25316 & ~n25317;
  assign n25319 = n1156 & ~n25312;
  assign n25320 = pi349 & n25319;
  assign n25321 = ~n25306 & ~n25309;
  assign n25322 = ~n25320 & ~n25321;
  assign n25323 = ~n25318 & ~n25322;
  assign n25324 = ~n25315 & ~n25323;
  assign n25325 = ~n24117 & n25324;
  assign n25326 = n24117 & ~n25324;
  assign n25327 = ~n25325 & ~n25326;
  assign n25328 = pi294 & ~n25327;
  assign n25329 = pi128 & n25328;
  assign n25330 = pi128 & pi294;
  assign n25331 = n24117 & n25324;
  assign n25332 = ~n24117 & ~n25324;
  assign n25333 = ~n25331 & ~n25332;
  assign n25334 = ~n25330 & ~n25333;
  assign n25335 = ~n25329 & ~n25334;
  assign n25336 = n22940 & n23552;
  assign n25337 = ~n22940 & ~n23552;
  assign n25338 = ~n25300 & ~n25301;
  assign n25339 = pi284 & ~n25338;
  assign n25340 = n22935 & ~n23556;
  assign n25341 = ~n22935 & n23556;
  assign n25342 = ~n25340 & ~n25341;
  assign n25343 = ~pi284 & ~n25342;
  assign n25344 = ~n25339 & ~n25343;
  assign n25345 = ~n25337 & ~n25344;
  assign n25346 = ~n25336 & ~n25345;
  assign n25347 = n25335 & n25346;
  assign n25348 = ~n25335 & ~n25346;
  assign n25349 = ~n25347 & ~n25348;
  assign n25350 = ~n831 & ~n25349;
  assign n25351 = ~n23582 & ~n25350;
  assign n25352 = pi161 & ~n25351;
  assign n25353 = ~n23581 & ~n25352;
  assign po220 = ~pi160 & n25353;
  assign n25355 = ~pi092 & ~pi161;
  assign n25356 = ~pi286 & n831;
  assign n25357 = pi295 & n1515;
  assign n25358 = ~n24099 & ~n24113;
  assign n25359 = ~n24114 & ~n25358;
  assign n25360 = n25357 & ~n25359;
  assign n25361 = ~n24112 & ~n24114;
  assign n25362 = ~n24113 & ~n25361;
  assign n25363 = ~n25357 & ~n25362;
  assign n25364 = ~n25360 & ~n25363;
  assign n25365 = pi297 & n1533;
  assign n25366 = ~n24078 & ~n24082;
  assign n25367 = ~n24083 & ~n25366;
  assign n25368 = ~n25365 & ~n25367;
  assign n25369 = ~n24075 & ~n24083;
  assign n25370 = ~n24060 & n25369;
  assign n25371 = ~n24082 & ~n25370;
  assign n25372 = n25365 & ~n25371;
  assign n25373 = ~n25368 & ~n25372;
  assign n25374 = ~n23593 & ~n24028;
  assign n25375 = ~n23507 & ~n23512;
  assign n25376 = ~n23508 & ~n25375;
  assign n25377 = n23593 & n24028;
  assign n25378 = ~n25376 & ~n25377;
  assign n25379 = ~n25374 & ~n25378;
  assign n25380 = pi301 & n3012;
  assign n25381 = ~n24007 & ~n24014;
  assign n25382 = ~n24015 & ~n25381;
  assign n25383 = ~n25380 & ~n25382;
  assign n25384 = ~n24010 & ~n24015;
  assign n25385 = ~n24014 & ~n25384;
  assign n25386 = n25380 & ~n25385;
  assign n25387 = ~n25383 & ~n25386;
  assign n25388 = n23964 & ~n23968;
  assign n25389 = ~n23964 & n23968;
  assign n25390 = ~n25388 & ~n25389;
  assign n25391 = ~n23607 & ~n25390;
  assign n25392 = ~n23437 & ~n23441;
  assign n25393 = ~n23436 & ~n25392;
  assign n25394 = n23607 & n25390;
  assign n25395 = ~n25393 & ~n25394;
  assign n25396 = ~n25391 & ~n25395;
  assign n25397 = pi305 & n5463;
  assign n25398 = ~n23950 & ~n23957;
  assign n25399 = ~n23958 & ~n25398;
  assign n25400 = ~n25397 & ~n25399;
  assign n25401 = ~n23953 & ~n23958;
  assign n25402 = ~n23957 & ~n25401;
  assign n25403 = n25397 & ~n25402;
  assign n25404 = ~n25400 & ~n25403;
  assign n25405 = ~n23884 & ~n23895;
  assign n25406 = n23884 & n23895;
  assign n25407 = ~n23889 & ~n25406;
  assign n25408 = ~n25405 & ~n25407;
  assign n25409 = pi309 & n9517;
  assign n25410 = ~n23862 & ~n23869;
  assign n25411 = ~n23870 & ~n25410;
  assign n25412 = ~n25409 & ~n25411;
  assign n25413 = ~n23865 & ~n23870;
  assign n25414 = ~n23869 & ~n25413;
  assign n25415 = n25409 & ~n25414;
  assign n25416 = ~n25412 & ~n25415;
  assign n25417 = ~n23795 & ~n23796;
  assign n25418 = n23795 & n23796;
  assign n25419 = ~n23801 & ~n25418;
  assign n25420 = ~n25417 & ~n25419;
  assign n25421 = pi313 & n14156;
  assign n25422 = ~n23774 & ~n23781;
  assign n25423 = ~n23782 & ~n25422;
  assign n25424 = ~n25421 & ~n25423;
  assign n25425 = ~n23777 & ~n23782;
  assign n25426 = ~n23781 & ~n25425;
  assign n25427 = n25421 & ~n25426;
  assign n25428 = ~n25424 & ~n25427;
  assign n25429 = ~n23741 & ~n23742;
  assign n25430 = n23741 & n23742;
  assign n25431 = ~n23220 & ~n25430;
  assign n25432 = ~n23214 & n25431;
  assign n25433 = ~n25429 & ~n25432;
  assign n25434 = ~n23697 & n23702;
  assign n25435 = ~n23696 & ~n23702;
  assign n25436 = ~n23693 & n25435;
  assign n25437 = ~n25434 & ~n25436;
  assign n25438 = ~n23723 & ~n25437;
  assign n25439 = pi317 & n18937;
  assign n25440 = pi319 & n23069;
  assign n25441 = n23626 & ~n23631;
  assign n25442 = ~n23069 & ~n25441;
  assign n25443 = n20347 & ~n25442;
  assign n25444 = n23069 & ~n23646;
  assign n25445 = ~n25443 & ~n25444;
  assign n25446 = pi321 & ~n25445;
  assign n25447 = n20347 & n23632;
  assign n25448 = ~n25446 & ~n25447;
  assign n25449 = pi320 & ~n25448;
  assign n25450 = n23088 & n25441;
  assign n25451 = ~n25449 & ~n25450;
  assign n25452 = ~n25440 & ~n25451;
  assign n25453 = n25440 & n25451;
  assign n25454 = ~n25452 & ~n25453;
  assign n25455 = ~pi156 & ~n23060;
  assign n25456 = pi155 & n25455;
  assign n25457 = ~pi155 & pi156;
  assign n25458 = pi154 & n25457;
  assign n25459 = ~n25456 & ~n25458;
  assign n25460 = pi153 & ~n25459;
  assign n25461 = pi155 & pi156;
  assign n25462 = ~pi154 & n25461;
  assign n25463 = ~pi156 & n23060;
  assign n25464 = ~pi155 & n25463;
  assign n25465 = ~n25462 & ~n25464;
  assign n25466 = ~pi153 & ~n25465;
  assign n25467 = pi155 & ~pi156;
  assign n25468 = pi156 & ~n23060;
  assign n25469 = ~pi155 & n25468;
  assign n25470 = ~n25467 & ~n25469;
  assign n25471 = pi154 & ~n25470;
  assign n25472 = ~pi155 & ~pi156;
  assign n25473 = pi156 & n23060;
  assign n25474 = pi155 & n25473;
  assign n25475 = ~n25472 & ~n25474;
  assign n25476 = ~pi154 & ~n25475;
  assign n25477 = ~n25471 & ~n25476;
  assign n25478 = ~n25466 & n25477;
  assign n25479 = ~n25460 & n25478;
  assign n25480 = n23626 & n25479;
  assign n25481 = n1178 & n25480;
  assign n25482 = pi321 & n25479;
  assign n25483 = pi320 & n23626;
  assign n25484 = ~n25482 & ~n25483;
  assign n25485 = ~n25481 & ~n25484;
  assign n25486 = ~n25454 & ~n25485;
  assign n25487 = ~n25440 & n25451;
  assign n25488 = n25440 & ~n25451;
  assign n25489 = ~n25487 & ~n25488;
  assign n25490 = n23626 & ~n25482;
  assign n25491 = pi320 & n25490;
  assign n25492 = n25479 & ~n25483;
  assign n25493 = pi321 & n25492;
  assign n25494 = ~n25491 & ~n25493;
  assign n25495 = ~n25489 & ~n25494;
  assign n25496 = ~n25486 & ~n25495;
  assign n25497 = ~n23658 & ~n23671;
  assign n25498 = n23658 & n23671;
  assign n25499 = pi319 & ~n25498;
  assign n25500 = ~n25497 & ~n25499;
  assign n25501 = n25496 & ~n25500;
  assign n25502 = ~pi319 & ~n25497;
  assign n25503 = ~n25498 & ~n25502;
  assign n25504 = ~n25496 & ~n25503;
  assign n25505 = ~n25501 & ~n25504;
  assign n25506 = n20347 & ~n25505;
  assign n25507 = pi318 & n25506;
  assign n25508 = n20347 & ~n25498;
  assign n25509 = pi319 & n25508;
  assign n25510 = ~n25497 & ~n25509;
  assign n25511 = ~n25496 & ~n25510;
  assign n25512 = n25496 & ~n25503;
  assign n25513 = ~n25511 & ~n25512;
  assign n25514 = ~pi318 & ~n25513;
  assign n25515 = ~n23671 & ~n25496;
  assign n25516 = ~n23658 & n25515;
  assign n25517 = n25496 & ~n25497;
  assign n25518 = ~n25516 & ~n25517;
  assign n25519 = ~n20347 & ~n25518;
  assign n25520 = ~n25514 & ~n25519;
  assign n25521 = n23680 & n23688;
  assign n25522 = ~n23680 & ~n23688;
  assign n25523 = ~n23677 & ~n25522;
  assign n25524 = ~n25521 & ~n25523;
  assign n25525 = n25520 & ~n25524;
  assign n25526 = ~n25507 & n25525;
  assign n25527 = ~n25507 & n25520;
  assign n25528 = n18937 & ~n25521;
  assign n25529 = pi318 & n25528;
  assign n25530 = ~n25522 & ~n25529;
  assign n25531 = ~n25527 & ~n25530;
  assign n25532 = ~n25526 & ~n25531;
  assign n25533 = ~n25439 & ~n25532;
  assign n25534 = n25439 & n25532;
  assign n25535 = ~n25533 & ~n25534;
  assign n25536 = pi316 & n17455;
  assign n25537 = ~n23696 & n23702;
  assign n25538 = ~n25536 & ~n25537;
  assign n25539 = ~n23693 & n25538;
  assign n25540 = ~n23693 & ~n25537;
  assign n25541 = n25536 & ~n25540;
  assign n25542 = ~n25539 & ~n25541;
  assign n25543 = ~n25535 & ~n25542;
  assign n25544 = ~n25439 & n25532;
  assign n25545 = n25439 & ~n25532;
  assign n25546 = ~n25544 & ~n25545;
  assign n25547 = n25536 & ~n25537;
  assign n25548 = ~n23693 & n25547;
  assign n25549 = ~n25536 & ~n25540;
  assign n25550 = ~n25548 & ~n25549;
  assign n25551 = ~n25546 & ~n25550;
  assign n25552 = ~n25543 & ~n25551;
  assign n25553 = ~n16985 & ~n25552;
  assign n25554 = ~pi315 & ~n25552;
  assign n25555 = n16985 & n25552;
  assign n25556 = pi315 & n25555;
  assign n25557 = ~n25554 & ~n25556;
  assign n25558 = ~pi316 & ~n25557;
  assign n25559 = ~n25553 & ~n25558;
  assign n25560 = ~n25438 & ~n25559;
  assign n25561 = n16985 & n25437;
  assign n25562 = n23723 & n25552;
  assign n25563 = n25561 & n25562;
  assign n25564 = n16985 & n25438;
  assign n25565 = n23723 & ~n25437;
  assign n25566 = ~n23723 & n25437;
  assign n25567 = ~n25565 & ~n25566;
  assign n25568 = pi316 & ~n25567;
  assign n25569 = ~n25564 & ~n25568;
  assign n25570 = ~n25552 & ~n25569;
  assign n25571 = ~n25563 & ~n25570;
  assign n25572 = pi315 & ~n25571;
  assign n25573 = ~n23723 & n25552;
  assign n25574 = ~n16985 & ~n25437;
  assign n25575 = n25573 & n25574;
  assign n25576 = n23723 & ~n25552;
  assign n25577 = n25437 & n25576;
  assign n25578 = n23723 & n25437;
  assign n25579 = n16985 & ~n25578;
  assign n25580 = pi316 & n25579;
  assign n25581 = ~n25438 & ~n25580;
  assign n25582 = n25552 & ~n25581;
  assign n25583 = ~n25577 & ~n25582;
  assign n25584 = ~pi315 & ~n25583;
  assign n25585 = ~n25575 & ~n25584;
  assign n25586 = ~n25572 & n25585;
  assign n25587 = ~n25560 & n25586;
  assign n25588 = n23729 & ~n23732;
  assign n25589 = ~n23202 & n23207;
  assign n25590 = ~n23203 & ~n25589;
  assign n25591 = ~n23729 & n23732;
  assign n25592 = ~n25590 & ~n25591;
  assign n25593 = ~n25588 & ~n25592;
  assign n25594 = ~n25587 & n25593;
  assign n25595 = n25587 & ~n25593;
  assign n25596 = ~n25594 & ~n25595;
  assign n25597 = n14618 & ~n25596;
  assign n25598 = pi314 & n25597;
  assign n25599 = pi314 & n14618;
  assign n25600 = ~n25595 & ~n25599;
  assign n25601 = ~n25594 & n25600;
  assign n25602 = ~n25598 & ~n25601;
  assign n25603 = ~n25433 & ~n25602;
  assign n25604 = n25433 & ~n25601;
  assign n25605 = ~n25598 & n25604;
  assign n25606 = ~n25603 & ~n25605;
  assign n25607 = n25428 & ~n25606;
  assign n25608 = ~n25428 & n25606;
  assign n25609 = ~n25607 & ~n25608;
  assign n25610 = pi312 & n11998;
  assign n25611 = ~n10908 & ~n11998;
  assign n25612 = pi313 & ~n25611;
  assign n25613 = n23757 & ~n25612;
  assign n25614 = ~n10908 & n11998;
  assign n25615 = pi313 & ~n23757;
  assign n25616 = n25614 & n25615;
  assign n25617 = ~n25613 & ~n25616;
  assign n25618 = ~n23771 & ~n25617;
  assign n25619 = ~n11998 & n23757;
  assign n25620 = ~n23759 & ~n25619;
  assign n25621 = ~n23222 & ~n25620;
  assign n25622 = n23770 & n25621;
  assign n25623 = n10908 & ~n11998;
  assign n25624 = ~n23757 & n25623;
  assign n25625 = ~n10908 & ~n23222;
  assign n25626 = n11998 & ~n25625;
  assign n25627 = n23757 & n25626;
  assign n25628 = ~n25624 & ~n25627;
  assign n25629 = pi313 & ~n25628;
  assign n25630 = n23222 & n23781;
  assign n25631 = ~n25629 & ~n25630;
  assign n25632 = ~n23770 & ~n25631;
  assign n25633 = ~n11998 & ~n23757;
  assign n25634 = n11998 & n23757;
  assign n25635 = ~n25633 & ~n25634;
  assign n25636 = n10908 & ~n25635;
  assign n25637 = pi313 & n25636;
  assign n25638 = n23222 & n25637;
  assign n25639 = ~n25632 & ~n25638;
  assign n25640 = ~n25622 & n25639;
  assign n25641 = ~n25618 & n25640;
  assign n25642 = ~n23792 & ~n25641;
  assign n25643 = n23792 & n25641;
  assign n25644 = n23761 & ~n25643;
  assign n25645 = ~n25642 & ~n25644;
  assign n25646 = n25610 & ~n25645;
  assign n25647 = ~n23761 & ~n25642;
  assign n25648 = ~n25643 & ~n25647;
  assign n25649 = ~n25610 & ~n25648;
  assign n25650 = ~n25646 & ~n25649;
  assign n25651 = ~n25609 & ~n25650;
  assign n25652 = n25428 & n25606;
  assign n25653 = ~n25428 & ~n25606;
  assign n25654 = ~n25652 & ~n25653;
  assign n25655 = ~n25610 & ~n25645;
  assign n25656 = n25610 & ~n25648;
  assign n25657 = ~n25655 & ~n25656;
  assign n25658 = ~n25654 & ~n25657;
  assign n25659 = ~n25651 & ~n25658;
  assign n25660 = n25420 & ~n25659;
  assign n25661 = ~n25420 & n25659;
  assign n25662 = ~n25660 & ~n25661;
  assign n25663 = n10908 & ~n25662;
  assign n25664 = pi311 & n25663;
  assign n25665 = pi311 & n10908;
  assign n25666 = ~n25420 & ~n25659;
  assign n25667 = n25420 & n25659;
  assign n25668 = ~n25666 & ~n25667;
  assign n25669 = ~n25665 & ~n25668;
  assign n25670 = ~n25664 & ~n25669;
  assign n25671 = ~n9517 & ~n23812;
  assign n25672 = ~n23296 & ~n25671;
  assign n25673 = n7874 & n25672;
  assign n25674 = ~n23295 & ~n23812;
  assign n25675 = n9517 & ~n25674;
  assign n25676 = ~n25673 & ~n25675;
  assign n25677 = pi310 & ~n25676;
  assign n25678 = ~n23822 & ~n25677;
  assign n25679 = n25670 & ~n25678;
  assign n25680 = ~n25670 & n25678;
  assign n25681 = ~n25679 & ~n25680;
  assign n25682 = n9815 & ~n25681;
  assign n25683 = pi310 & n25682;
  assign n25684 = pi310 & n9815;
  assign n25685 = ~n25670 & ~n25678;
  assign n25686 = n25670 & n25678;
  assign n25687 = ~n25685 & ~n25686;
  assign n25688 = ~n25684 & ~n25687;
  assign n25689 = ~n25683 & ~n25688;
  assign n25690 = n25416 & n25689;
  assign n25691 = ~n25416 & ~n25689;
  assign n25692 = ~n25690 & ~n25691;
  assign n25693 = pi308 & n7874;
  assign n25694 = pi309 & ~n14735;
  assign n25695 = n23844 & ~n25694;
  assign n25696 = pi309 & ~n23844;
  assign n25697 = n14732 & n25696;
  assign n25698 = ~n25695 & ~n25697;
  assign n25699 = ~n23859 & ~n25698;
  assign n25700 = ~n7874 & n23844;
  assign n25701 = ~n23870 & ~n25700;
  assign n25702 = n23305 & ~n25701;
  assign n25703 = n23858 & n25702;
  assign n25704 = n14747 & ~n23844;
  assign n25705 = ~n7044 & n23305;
  assign n25706 = n7874 & ~n25705;
  assign n25707 = n23844 & n25706;
  assign n25708 = ~n25704 & ~n25707;
  assign n25709 = pi309 & ~n25708;
  assign n25710 = ~n23305 & n23845;
  assign n25711 = ~n25709 & ~n25710;
  assign n25712 = ~n23858 & ~n25711;
  assign n25713 = ~n7874 & ~n23844;
  assign n25714 = n7874 & n23844;
  assign n25715 = ~n25713 & ~n25714;
  assign n25716 = n7044 & ~n25715;
  assign n25717 = pi309 & n25716;
  assign n25718 = ~n23305 & n25717;
  assign n25719 = ~n25712 & ~n25718;
  assign n25720 = ~n25703 & n25719;
  assign n25721 = ~n25699 & n25720;
  assign n25722 = n23880 & n25721;
  assign n25723 = ~n23880 & ~n25721;
  assign n25724 = n23848 & ~n25723;
  assign n25725 = ~n25722 & ~n25724;
  assign n25726 = n25693 & ~n25725;
  assign n25727 = ~n23848 & ~n25722;
  assign n25728 = ~n25723 & ~n25727;
  assign n25729 = ~n25693 & ~n25728;
  assign n25730 = ~n25726 & ~n25729;
  assign n25731 = ~n25692 & ~n25730;
  assign n25732 = n25416 & ~n25689;
  assign n25733 = ~n25416 & n25689;
  assign n25734 = ~n25732 & ~n25733;
  assign n25735 = ~n25693 & ~n25725;
  assign n25736 = n25693 & ~n25728;
  assign n25737 = ~n25735 & ~n25736;
  assign n25738 = ~n25734 & ~n25737;
  assign n25739 = ~n25731 & ~n25738;
  assign n25740 = ~n25408 & ~n25739;
  assign n25741 = n25408 & n25739;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 = n7044 & ~n25742;
  assign n25744 = pi307 & n25743;
  assign n25745 = pi307 & n7044;
  assign n25746 = n25408 & ~n25739;
  assign n25747 = ~n25408 & n25739;
  assign n25748 = ~n25746 & ~n25747;
  assign n25749 = ~n25745 & ~n25748;
  assign n25750 = ~n25744 & ~n25749;
  assign n25751 = ~n23366 & n23920;
  assign n25752 = ~n23381 & ~n23902;
  assign n25753 = n4772 & n25752;
  assign n25754 = ~n23382 & n23900;
  assign n25755 = n5463 & ~n25754;
  assign n25756 = ~n25753 & ~n25755;
  assign n25757 = pi306 & ~n25756;
  assign n25758 = ~n25751 & ~n25757;
  assign n25759 = ~n25750 & n25758;
  assign n25760 = n25750 & ~n25758;
  assign n25761 = ~n25759 & ~n25760;
  assign n25762 = n6777 & ~n25761;
  assign n25763 = pi306 & n25762;
  assign n25764 = pi306 & n6777;
  assign n25765 = n25750 & n25758;
  assign n25766 = ~n25750 & ~n25758;
  assign n25767 = ~n25765 & ~n25766;
  assign n25768 = ~n25764 & ~n25767;
  assign n25769 = ~n25763 & ~n25768;
  assign n25770 = n25404 & n25769;
  assign n25771 = ~n25404 & ~n25769;
  assign n25772 = ~n25770 & ~n25771;
  assign n25773 = pi304 & n4772;
  assign n25774 = pi305 & n23932;
  assign n25775 = n9909 & n25774;
  assign n25776 = pi305 & ~n9912;
  assign n25777 = ~n23932 & ~n25776;
  assign n25778 = ~n25775 & ~n25777;
  assign n25779 = ~n23947 & ~n25778;
  assign n25780 = ~n4772 & ~n23932;
  assign n25781 = ~n23958 & ~n25780;
  assign n25782 = ~n23385 & ~n25781;
  assign n25783 = n23946 & n25782;
  assign n25784 = n4772 & ~n23932;
  assign n25785 = ~n4772 & n23932;
  assign n25786 = ~n25784 & ~n25785;
  assign n25787 = n4086 & ~n25786;
  assign n25788 = pi305 & n25787;
  assign n25789 = n23385 & n25788;
  assign n25790 = ~n4086 & ~n23385;
  assign n25791 = n4772 & ~n25790;
  assign n25792 = ~n23932 & n25791;
  assign n25793 = n9924 & n23932;
  assign n25794 = ~n25792 & ~n25793;
  assign n25795 = pi305 & ~n25794;
  assign n25796 = n23385 & n23933;
  assign n25797 = ~n25795 & ~n25796;
  assign n25798 = ~n23946 & ~n25797;
  assign n25799 = ~n25789 & ~n25798;
  assign n25800 = ~n25783 & n25799;
  assign n25801 = ~n25779 & n25800;
  assign n25802 = n23968 & n25801;
  assign n25803 = ~n23968 & ~n25801;
  assign n25804 = n23936 & ~n25803;
  assign n25805 = ~n25802 & ~n25804;
  assign n25806 = n25773 & ~n25805;
  assign n25807 = ~n23936 & ~n25802;
  assign n25808 = ~n25803 & ~n25807;
  assign n25809 = ~n25773 & ~n25808;
  assign n25810 = ~n25806 & ~n25809;
  assign n25811 = ~n25772 & ~n25810;
  assign n25812 = n25404 & ~n25769;
  assign n25813 = ~n25404 & n25769;
  assign n25814 = ~n25812 & ~n25813;
  assign n25815 = ~n25773 & ~n25805;
  assign n25816 = n25773 & ~n25808;
  assign n25817 = ~n25815 & ~n25816;
  assign n25818 = ~n25814 & ~n25817;
  assign n25819 = ~n25811 & ~n25818;
  assign n25820 = ~n25396 & ~n25819;
  assign n25821 = n25396 & n25819;
  assign n25822 = ~n25820 & ~n25821;
  assign n25823 = n4086 & ~n25822;
  assign n25824 = pi303 & n25823;
  assign n25825 = pi303 & n4086;
  assign n25826 = n25396 & ~n25819;
  assign n25827 = ~n25396 & n25819;
  assign n25828 = ~n25826 & ~n25827;
  assign n25829 = ~n25825 & ~n25828;
  assign n25830 = ~n25824 & ~n25829;
  assign n25831 = ~n23974 & ~n23975;
  assign n25832 = n23974 & n23975;
  assign n25833 = ~n23454 & ~n25832;
  assign n25834 = ~n23448 & n25833;
  assign n25835 = ~n25831 & ~n25834;
  assign n25836 = ~n25830 & n25835;
  assign n25837 = n25830 & ~n25835;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = n3552 & ~n25838;
  assign n25840 = pi302 & n25839;
  assign n25841 = pi302 & n3552;
  assign n25842 = n25830 & n25835;
  assign n25843 = ~n25830 & ~n25835;
  assign n25844 = ~n25842 & ~n25843;
  assign n25845 = ~n25841 & ~n25844;
  assign n25846 = ~n25840 & ~n25845;
  assign n25847 = n25387 & ~n25846;
  assign n25848 = ~n25387 & n25846;
  assign n25849 = ~n25847 & ~n25848;
  assign n25850 = pi300 & n2574;
  assign n25851 = pi301 & ~n9624;
  assign n25852 = n23990 & ~n25851;
  assign n25853 = pi301 & ~n23990;
  assign n25854 = n9627 & n25853;
  assign n25855 = ~n25852 & ~n25854;
  assign n25856 = ~n24004 & ~n25855;
  assign n25857 = ~n2574 & n23990;
  assign n25858 = ~n23992 & ~n25857;
  assign n25859 = ~n23456 & ~n25858;
  assign n25860 = n24003 & n25859;
  assign n25861 = n9636 & ~n23990;
  assign n25862 = ~n2183 & ~n23456;
  assign n25863 = n2574 & ~n25862;
  assign n25864 = n23990 & n25863;
  assign n25865 = ~n25861 & ~n25864;
  assign n25866 = pi301 & ~n25865;
  assign n25867 = n23456 & n24014;
  assign n25868 = ~n25866 & ~n25867;
  assign n25869 = ~n24003 & ~n25868;
  assign n25870 = ~n2574 & ~n23990;
  assign n25871 = n2574 & n23990;
  assign n25872 = ~n25870 & ~n25871;
  assign n25873 = n2183 & ~n25872;
  assign n25874 = pi301 & n25873;
  assign n25875 = n23456 & n25874;
  assign n25876 = ~n25869 & ~n25875;
  assign n25877 = ~n25860 & n25876;
  assign n25878 = ~n25856 & n25877;
  assign n25879 = ~n24025 & ~n25878;
  assign n25880 = n24025 & n25878;
  assign n25881 = n23994 & ~n25880;
  assign n25882 = ~n25879 & ~n25881;
  assign n25883 = n25850 & ~n25882;
  assign n25884 = ~n23994 & ~n25879;
  assign n25885 = ~n25880 & ~n25884;
  assign n25886 = ~n25850 & ~n25885;
  assign n25887 = ~n25883 & ~n25886;
  assign n25888 = ~n25849 & ~n25887;
  assign n25889 = n25387 & n25846;
  assign n25890 = ~n25387 & ~n25846;
  assign n25891 = ~n25889 & ~n25890;
  assign n25892 = ~n25850 & ~n25882;
  assign n25893 = n25850 & ~n25885;
  assign n25894 = ~n25892 & ~n25893;
  assign n25895 = ~n25891 & ~n25894;
  assign n25896 = ~n25888 & ~n25895;
  assign n25897 = n25379 & ~n25896;
  assign n25898 = ~n25379 & n25896;
  assign n25899 = ~n25897 & ~n25898;
  assign n25900 = n2183 & ~n25899;
  assign n25901 = pi299 & n25900;
  assign n25902 = pi299 & n2183;
  assign n25903 = ~n25379 & ~n25896;
  assign n25904 = n25379 & n25896;
  assign n25905 = ~n25903 & ~n25904;
  assign n25906 = ~n25902 & ~n25905;
  assign n25907 = ~n25901 & ~n25906;
  assign n25908 = ~n24032 & ~n24042;
  assign n25909 = n24032 & n24042;
  assign n25910 = ~n24033 & ~n25909;
  assign n25911 = ~n23519 & n25910;
  assign n25912 = ~n25908 & ~n25911;
  assign n25913 = n25907 & n25912;
  assign n25914 = ~n25907 & ~n25912;
  assign n25915 = ~n25913 & ~n25914;
  assign n25916 = n1840 & ~n25915;
  assign n25917 = pi298 & n25916;
  assign n25918 = pi298 & n1840;
  assign n25919 = ~n25907 & n25912;
  assign n25920 = n25907 & ~n25912;
  assign n25921 = ~n25919 & ~n25920;
  assign n25922 = ~n25918 & ~n25921;
  assign n25923 = ~n25917 & ~n25922;
  assign n25924 = n25373 & n25923;
  assign n25925 = ~n25373 & ~n25923;
  assign n25926 = ~n25924 & ~n25925;
  assign n25927 = pi296 & n1553;
  assign n25928 = n24048 & ~n24075;
  assign n25929 = ~n24060 & n25928;
  assign n25930 = ~n24048 & ~n24078;
  assign n25931 = ~n25929 & ~n25930;
  assign n25932 = ~n23583 & ~n25931;
  assign n25933 = ~n24048 & ~n24075;
  assign n25934 = ~n24060 & n25933;
  assign n25935 = n24048 & ~n24078;
  assign n25936 = ~n25934 & ~n25935;
  assign n25937 = n1553 & ~n25936;
  assign n25938 = pi297 & n25937;
  assign n25939 = ~n25932 & ~n25938;
  assign n25940 = ~n24096 & n25939;
  assign n25941 = n24096 & ~n25939;
  assign n25942 = n24061 & ~n25941;
  assign n25943 = ~n25940 & ~n25942;
  assign n25944 = n25927 & ~n25943;
  assign n25945 = ~n24061 & ~n25940;
  assign n25946 = ~n25941 & ~n25945;
  assign n25947 = ~n25927 & ~n25946;
  assign n25948 = ~n25944 & ~n25947;
  assign n25949 = ~n25926 & ~n25948;
  assign n25950 = n25373 & ~n25923;
  assign n25951 = ~n25373 & n25923;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = ~n25927 & ~n25943;
  assign n25954 = n25927 & ~n25946;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = ~n25952 & ~n25955;
  assign n25957 = ~n25949 & ~n25956;
  assign n25958 = n25364 & ~n25957;
  assign n25959 = ~n25364 & n25957;
  assign n25960 = ~n25958 & ~n25959;
  assign n25961 = ~n24117 & n25330;
  assign n25962 = pi294 & ~n1568;
  assign n25963 = ~n25961 & ~n25962;
  assign n25964 = n25961 & n25962;
  assign n25965 = ~n25963 & ~n25964;
  assign n25966 = pi293 & ~n25965;
  assign n25967 = pi128 & n25966;
  assign n25968 = pi128 & pi293;
  assign n25969 = n25961 & ~n25962;
  assign n25970 = ~n25961 & n25962;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = ~n25968 & ~n25971;
  assign n25973 = ~n25967 & ~n25972;
  assign n25974 = ~n25960 & ~n25973;
  assign n25975 = n25364 & n25957;
  assign n25976 = ~n25364 & ~n25957;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = pi293 & ~n25971;
  assign n25979 = pi128 & n25978;
  assign n25980 = ~n25965 & ~n25968;
  assign n25981 = ~n25979 & ~n25980;
  assign n25982 = ~n25977 & ~n25981;
  assign n25983 = ~n25974 & ~n25982;
  assign n25984 = n1156 & ~n25299;
  assign n25985 = pi349 & n25984;
  assign n25986 = ~n25309 & ~n25318;
  assign n25987 = ~n25985 & ~n25986;
  assign n25988 = ~n25311 & ~n25987;
  assign n25989 = ~n25310 & ~n25988;
  assign n25990 = pi258 & ~n25318;
  assign n25991 = pi128 & n25990;
  assign n25992 = pi349 & n25991;
  assign n25993 = n24146 & n24161;
  assign n25994 = ~n24146 & ~n24161;
  assign n25995 = n25264 & ~n25994;
  assign n25996 = ~n25993 & ~n25995;
  assign n25997 = ~n24146 & ~n25264;
  assign n25998 = n24146 & n25264;
  assign n25999 = ~n25997 & ~n25998;
  assign n26000 = ~n24157 & n25268;
  assign n26001 = n24161 & ~n25275;
  assign n26002 = ~n24161 & n25275;
  assign n26003 = ~n26001 & ~n26002;
  assign n26004 = ~n26000 & ~n26003;
  assign n26005 = ~n25999 & n26004;
  assign n26006 = ~n24146 & n25264;
  assign n26007 = n24146 & ~n25264;
  assign n26008 = ~n26006 & ~n26007;
  assign n26009 = ~n24161 & ~n25275;
  assign n26010 = n24161 & n25275;
  assign n26011 = ~n26009 & ~n26010;
  assign n26012 = ~n26000 & ~n26011;
  assign n26013 = ~n26008 & n26012;
  assign n26014 = n24157 & ~n25268;
  assign n26015 = ~n26013 & ~n26014;
  assign n26016 = ~n26005 & n26015;
  assign n26017 = ~n25996 & ~n26016;
  assign n26018 = n25996 & n26016;
  assign n26019 = ~n26017 & ~n26018;
  assign n26020 = pi345 & n2091;
  assign n26021 = n24181 & n25150;
  assign n26022 = ~n21965 & ~n24173;
  assign n26023 = n21965 & ~n24164;
  assign n26024 = ~n26022 & ~n26023;
  assign n26025 = ~n25152 & ~n26024;
  assign n26026 = ~n25155 & ~n26025;
  assign n26027 = n25151 & ~n26026;
  assign n26028 = n21965 & ~n24173;
  assign n26029 = ~n21965 & ~n24164;
  assign n26030 = ~n26028 & ~n26029;
  assign n26031 = ~n25155 & ~n26030;
  assign n26032 = ~n25152 & ~n26031;
  assign n26033 = ~n25151 & ~n26032;
  assign n26034 = ~n26027 & ~n26033;
  assign n26035 = ~n25149 & ~n26034;
  assign n26036 = ~n25177 & ~n26033;
  assign n26037 = ~n26027 & n26036;
  assign n26038 = ~n26035 & ~n26037;
  assign n26039 = ~n25186 & ~n26038;
  assign n26040 = ~n25177 & ~n26034;
  assign n26041 = ~n25149 & ~n26033;
  assign n26042 = ~n26027 & n26041;
  assign n26043 = ~n26040 & ~n26042;
  assign n26044 = ~n25134 & ~n26043;
  assign n26045 = ~n26039 & ~n26044;
  assign n26046 = ~n24181 & ~n25150;
  assign n26047 = n26045 & ~n26046;
  assign n26048 = ~n26021 & ~n26047;
  assign n26049 = n4596 & ~n24188;
  assign n26050 = pi341 & n26049;
  assign n26051 = ~n24181 & n25191;
  assign n26052 = n24181 & ~n25191;
  assign n26053 = ~n26051 & ~n26052;
  assign n26054 = ~n24204 & ~n26053;
  assign n26055 = n24181 & n25191;
  assign n26056 = ~n24181 & ~n25191;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = n24204 & ~n26057;
  assign n26059 = ~n26054 & ~n26058;
  assign n26060 = n24188 & ~n25197;
  assign n26061 = ~n26059 & ~n26060;
  assign n26062 = ~n26050 & ~n26061;
  assign n26063 = ~n26048 & n26062;
  assign n26064 = n26048 & ~n26062;
  assign n26065 = ~n26063 & ~n26064;
  assign n26066 = pi339 & n5732;
  assign n26067 = n24224 & n25065;
  assign n26068 = ~n25061 & ~n25085;
  assign n26069 = n25061 & n25085;
  assign n26070 = ~n26068 & ~n26069;
  assign n26071 = n11711 & ~n26070;
  assign n26072 = pi331 & n26071;
  assign n26073 = ~n25061 & n25085;
  assign n26074 = n25061 & ~n25085;
  assign n26075 = ~n26073 & ~n26074;
  assign n26076 = ~n25032 & ~n26075;
  assign n26077 = ~n26072 & ~n26076;
  assign n26078 = ~n25031 & ~n26077;
  assign n26079 = n11711 & ~n26075;
  assign n26080 = pi331 & n26079;
  assign n26081 = ~n25032 & ~n26070;
  assign n26082 = ~n26080 & ~n26081;
  assign n26083 = ~n25101 & ~n26082;
  assign n26084 = ~n26078 & ~n26083;
  assign n26085 = ~n24224 & ~n25065;
  assign n26086 = n26084 & ~n26085;
  assign n26087 = ~n26067 & ~n26086;
  assign n26088 = n9205 & ~n24231;
  assign n26089 = pi335 & n26088;
  assign n26090 = ~n24224 & n25106;
  assign n26091 = n24224 & ~n25106;
  assign n26092 = ~n26090 & ~n26091;
  assign n26093 = ~n24247 & ~n26092;
  assign n26094 = n24224 & n25106;
  assign n26095 = ~n24224 & ~n25106;
  assign n26096 = ~n26094 & ~n26095;
  assign n26097 = n24247 & ~n26096;
  assign n26098 = ~n26093 & ~n26097;
  assign n26099 = n24231 & ~n25112;
  assign n26100 = ~n26098 & ~n26099;
  assign n26101 = ~n26089 & ~n26100;
  assign n26102 = ~n26087 & n26101;
  assign n26103 = n26087 & ~n26101;
  assign n26104 = ~n26102 & ~n26103;
  assign n26105 = pi333 & n11384;
  assign n26106 = ~n24251 & ~n25003;
  assign n26107 = n24251 & n25003;
  assign n26108 = n18461 & ~n26107;
  assign n26109 = pi328 & n26108;
  assign n26110 = ~n26106 & ~n26109;
  assign n26111 = n24264 & ~n24268;
  assign n26112 = ~n24264 & n24268;
  assign n26113 = ~n24251 & n25003;
  assign n26114 = n24251 & ~n25003;
  assign n26115 = ~n26113 & ~n26114;
  assign n26116 = n18461 & ~n26115;
  assign n26117 = pi328 & n26116;
  assign n26118 = ~n26106 & ~n26107;
  assign n26119 = ~n25009 & ~n26118;
  assign n26120 = ~n26117 & ~n26119;
  assign n26121 = ~n26112 & ~n26120;
  assign n26122 = ~n26111 & ~n26121;
  assign n26123 = n26110 & n26122;
  assign n26124 = ~n26110 & ~n26122;
  assign n26125 = ~n26123 & ~n26124;
  assign n26126 = pi329 & n18461;
  assign n26127 = ~n24272 & n24982;
  assign n26128 = n24272 & ~n24982;
  assign n26129 = ~n24989 & ~n26128;
  assign n26130 = ~n26127 & ~n26129;
  assign n26131 = ~n24272 & ~n24977;
  assign n26132 = n24272 & n24977;
  assign n26133 = ~n26131 & ~n26132;
  assign n26134 = n24292 & n24981;
  assign n26135 = ~n24962 & n24982;
  assign n26136 = n24962 & ~n24982;
  assign n26137 = ~n26135 & ~n26136;
  assign n26138 = ~n26134 & ~n26137;
  assign n26139 = ~n26133 & n26138;
  assign n26140 = ~n24272 & n24977;
  assign n26141 = n24272 & ~n24977;
  assign n26142 = ~n26140 & ~n26141;
  assign n26143 = n24962 & n24982;
  assign n26144 = ~n24962 & ~n24982;
  assign n26145 = ~n26143 & ~n26144;
  assign n26146 = ~n26134 & ~n26145;
  assign n26147 = ~n26142 & n26146;
  assign n26148 = ~n24292 & ~n24981;
  assign n26149 = ~n26147 & ~n26148;
  assign n26150 = ~n26139 & n26149;
  assign n26151 = n26130 & n26150;
  assign n26152 = ~n26130 & ~n26150;
  assign n26153 = ~n26151 & ~n26152;
  assign n26154 = ~n24297 & ~n24931;
  assign n26155 = ~n24939 & ~n26154;
  assign n26156 = ~n24305 & n24942;
  assign n26157 = ~n24297 & ~n24940;
  assign n26158 = n24297 & ~n24939;
  assign n26159 = ~n24931 & n26158;
  assign n26160 = ~n26157 & ~n26159;
  assign n26161 = n24305 & ~n24942;
  assign n26162 = ~n26160 & ~n26161;
  assign n26163 = ~n26156 & ~n26162;
  assign n26164 = ~n26155 & n26163;
  assign n26165 = n26155 & ~n26163;
  assign n26166 = ~n26164 & ~n26165;
  assign n26167 = n22545 & n24912;
  assign n26168 = ~n24913 & ~n26167;
  assign n26169 = ~n22557 & ~n26168;
  assign n26170 = ~n22545 & n24907;
  assign n26171 = ~n24908 & ~n26170;
  assign n26172 = n22557 & ~n26171;
  assign n26173 = n24906 & ~n24919;
  assign n26174 = ~n26172 & ~n26173;
  assign n26175 = ~n26169 & n26174;
  assign n26176 = pi323 & n26175;
  assign n26177 = pi151 & pi263;
  assign n26178 = pi148 & pi266;
  assign n26179 = pi145 & pi269;
  assign n26180 = pi142 & pi272;
  assign n26181 = pi139 & pi275;
  assign n26182 = pi136 & pi278;
  assign n26183 = pi133 & pi281;
  assign n26184 = pi285 & ~n22092;
  assign n26185 = pi284 & n26184;
  assign n26186 = ~pi285 & n22092;
  assign n26187 = pi284 & ~n26186;
  assign n26188 = ~pi284 & ~n26184;
  assign n26189 = pi283 & ~n26188;
  assign n26190 = ~n26187 & ~n26189;
  assign n26191 = pi129 & ~n26190;
  assign n26192 = ~n26185 & ~n26191;
  assign n26193 = pi128 & ~n26192;
  assign n26194 = pi284 & ~n22092;
  assign n26195 = n22096 & n26194;
  assign n26196 = ~n26193 & ~n26195;
  assign n26197 = pi128 & pi286;
  assign n26198 = pi285 & ~n26197;
  assign n26199 = pi129 & n26198;
  assign n26200 = pi129 & pi285;
  assign n26201 = pi286 & ~n26200;
  assign n26202 = pi128 & n26201;
  assign n26203 = ~n26199 & ~n26202;
  assign n26204 = ~n26196 & ~n26203;
  assign n26205 = n26196 & n26203;
  assign n26206 = ~n26204 & ~n26205;
  assign n26207 = pi284 & ~n26206;
  assign n26208 = pi130 & n26207;
  assign n26209 = pi130 & pi284;
  assign n26210 = n26196 & ~n26203;
  assign n26211 = ~n26196 & n26203;
  assign n26212 = ~n26210 & ~n26211;
  assign n26213 = ~n26209 & ~n26212;
  assign n26214 = ~n26208 & ~n26213;
  assign n26215 = ~n24332 & ~n24358;
  assign n26216 = ~n22096 & ~n24325;
  assign n26217 = ~n24355 & ~n26216;
  assign n26218 = n24332 & ~n26217;
  assign n26219 = ~n26215 & ~n26218;
  assign n26220 = ~n22121 & n26219;
  assign n26221 = n22102 & n26220;
  assign n26222 = ~pi283 & ~n26219;
  assign n26223 = ~n24387 & ~n26222;
  assign n26224 = pi282 & n26223;
  assign n26225 = ~n24324 & ~n26219;
  assign n26226 = pi283 & ~n26225;
  assign n26227 = ~n26224 & ~n26226;
  assign n26228 = pi130 & ~n26227;
  assign n26229 = ~n26221 & ~n26228;
  assign n26230 = ~n26214 & ~n26229;
  assign n26231 = n26214 & n26229;
  assign n26232 = ~n26230 & ~n26231;
  assign n26233 = pi283 & ~n26232;
  assign n26234 = pi131 & n26233;
  assign n26235 = pi131 & pi283;
  assign n26236 = n26214 & ~n26229;
  assign n26237 = ~n26214 & n26229;
  assign n26238 = ~n26236 & ~n26237;
  assign n26239 = ~n26235 & ~n26238;
  assign n26240 = ~n26234 & ~n26239;
  assign n26241 = pi130 & ~n24387;
  assign n26242 = ~n24324 & ~n26241;
  assign n26243 = n24367 & ~n26242;
  assign n26244 = ~pi130 & ~n24324;
  assign n26245 = ~n24387 & ~n26244;
  assign n26246 = ~n24367 & ~n26245;
  assign n26247 = ~n26243 & ~n26246;
  assign n26248 = pi282 & ~n26247;
  assign n26249 = pi131 & n26248;
  assign n26250 = ~n24367 & ~n24390;
  assign n26251 = n24367 & ~n26245;
  assign n26252 = ~n26250 & ~n26251;
  assign n26253 = ~pi131 & ~n26252;
  assign n26254 = ~n22121 & ~n24367;
  assign n26255 = n22102 & n26254;
  assign n26256 = ~n24324 & n24367;
  assign n26257 = ~n26255 & ~n26256;
  assign n26258 = ~pi282 & ~n26257;
  assign n26259 = ~n26253 & ~n26258;
  assign n26260 = ~n24403 & n26259;
  assign n26261 = ~n26249 & ~n26260;
  assign n26262 = n26240 & ~n26261;
  assign n26263 = ~n26240 & n26261;
  assign n26264 = ~n26262 & ~n26263;
  assign n26265 = pi282 & ~n26264;
  assign n26266 = pi132 & n26265;
  assign n26267 = pi132 & pi282;
  assign n26268 = ~n26263 & ~n26267;
  assign n26269 = ~n26262 & n26268;
  assign n26270 = ~n26266 & ~n26269;
  assign n26271 = ~n24322 & ~n24408;
  assign n26272 = ~n24413 & ~n26271;
  assign n26273 = ~n26270 & ~n26272;
  assign n26274 = ~n26269 & ~n26271;
  assign n26275 = ~n26266 & n26274;
  assign n26276 = ~n24413 & n26275;
  assign n26277 = ~n26273 & ~n26276;
  assign n26278 = ~n26183 & n26277;
  assign n26279 = n26183 & ~n26277;
  assign n26280 = ~n26278 & ~n26279;
  assign n26281 = pi280 & ~n24418;
  assign n26282 = pi133 & n26281;
  assign n26283 = pi134 & pi280;
  assign n26284 = ~n24311 & ~n24417;
  assign n26285 = ~n24415 & n26284;
  assign n26286 = ~n24442 & ~n26285;
  assign n26287 = ~n26283 & ~n26286;
  assign n26288 = ~n26282 & n26287;
  assign n26289 = ~n26282 & ~n26286;
  assign n26290 = n26283 & ~n26289;
  assign n26291 = ~n26288 & ~n26290;
  assign n26292 = ~n26280 & ~n26291;
  assign n26293 = ~n26183 & ~n26277;
  assign n26294 = n26183 & n26277;
  assign n26295 = ~n26293 & ~n26294;
  assign n26296 = n26283 & ~n26286;
  assign n26297 = ~n26282 & n26296;
  assign n26298 = ~n26283 & ~n26289;
  assign n26299 = ~n26297 & ~n26298;
  assign n26300 = ~n26295 & ~n26299;
  assign n26301 = ~n26292 & ~n26300;
  assign n26302 = n24458 & ~n24475;
  assign n26303 = ~n24458 & n24475;
  assign n26304 = ~n24466 & ~n26303;
  assign n26305 = n24457 & n26304;
  assign n26306 = ~n26302 & ~n26305;
  assign n26307 = n26301 & n26306;
  assign n26308 = ~n26301 & ~n26306;
  assign n26309 = ~n26307 & ~n26308;
  assign n26310 = pi135 & pi279;
  assign n26311 = n24490 & ~n24495;
  assign n26312 = ~n24496 & ~n26311;
  assign n26313 = n26310 & ~n26312;
  assign n26314 = ~n24490 & ~n24496;
  assign n26315 = ~n24495 & ~n26314;
  assign n26316 = ~n26310 & ~n26315;
  assign n26317 = ~n26313 & ~n26316;
  assign n26318 = ~n26309 & ~n26317;
  assign n26319 = n26301 & ~n26306;
  assign n26320 = ~n26301 & n26306;
  assign n26321 = ~n26319 & ~n26320;
  assign n26322 = ~n26310 & ~n26312;
  assign n26323 = n26310 & ~n26315;
  assign n26324 = ~n26322 & ~n26323;
  assign n26325 = ~n26321 & ~n26324;
  assign n26326 = ~n26318 & ~n26325;
  assign n26327 = ~n26182 & n26326;
  assign n26328 = n26182 & ~n26326;
  assign n26329 = ~n26327 & ~n26328;
  assign n26330 = pi137 & pi277;
  assign n26331 = pi278 & ~n24488;
  assign n26332 = pi135 & n26331;
  assign n26333 = ~n24490 & ~n24497;
  assign n26334 = ~n26332 & ~n26333;
  assign n26335 = ~n24506 & n26334;
  assign n26336 = n24506 & ~n26334;
  assign n26337 = n24489 & ~n26336;
  assign n26338 = ~n26335 & ~n26337;
  assign n26339 = n26330 & ~n26338;
  assign n26340 = ~n24489 & ~n26335;
  assign n26341 = ~n26336 & ~n26340;
  assign n26342 = ~n26330 & ~n26341;
  assign n26343 = ~n26339 & ~n26342;
  assign n26344 = ~n26329 & ~n26343;
  assign n26345 = ~n26182 & ~n26326;
  assign n26346 = n26182 & n26326;
  assign n26347 = ~n26345 & ~n26346;
  assign n26348 = ~n26330 & ~n26338;
  assign n26349 = n26330 & ~n26341;
  assign n26350 = ~n26348 & ~n26349;
  assign n26351 = ~n26347 & ~n26350;
  assign n26352 = ~n26344 & ~n26351;
  assign n26353 = n24510 & ~n24535;
  assign n26354 = ~n24510 & n24535;
  assign n26355 = ~n24526 & ~n26354;
  assign n26356 = ~n26353 & ~n26355;
  assign n26357 = n26352 & ~n26356;
  assign n26358 = ~n26352 & n26356;
  assign n26359 = ~n26357 & ~n26358;
  assign n26360 = pi138 & pi276;
  assign n26361 = n24549 & ~n24555;
  assign n26362 = ~n24554 & ~n26361;
  assign n26363 = n26360 & ~n26362;
  assign n26364 = ~n24549 & ~n24554;
  assign n26365 = ~n24555 & ~n26364;
  assign n26366 = ~n26360 & ~n26365;
  assign n26367 = ~n26363 & ~n26366;
  assign n26368 = ~n26359 & ~n26367;
  assign n26369 = n26352 & n26356;
  assign n26370 = ~n26352 & ~n26356;
  assign n26371 = ~n26369 & ~n26370;
  assign n26372 = ~n26360 & ~n26362;
  assign n26373 = n26360 & ~n26365;
  assign n26374 = ~n26372 & ~n26373;
  assign n26375 = ~n26371 & ~n26374;
  assign n26376 = ~n26368 & ~n26375;
  assign n26377 = ~n26181 & ~n26376;
  assign n26378 = n26181 & n26376;
  assign n26379 = ~n26377 & ~n26378;
  assign n26380 = pi275 & ~n24556;
  assign n26381 = pi138 & n26380;
  assign n26382 = ~n24547 & ~n24549;
  assign n26383 = ~n24548 & ~n26382;
  assign n26384 = ~n26381 & n26383;
  assign n26385 = pi140 & pi274;
  assign n26386 = ~n26381 & ~n26382;
  assign n26387 = pi274 & ~n26386;
  assign n26388 = pi139 & n26387;
  assign n26389 = n24566 & ~n26388;
  assign n26390 = n26385 & ~n26389;
  assign n26391 = ~n26384 & n26390;
  assign n26392 = ~n26384 & ~n26389;
  assign n26393 = ~n26385 & ~n26392;
  assign n26394 = ~n26391 & ~n26393;
  assign n26395 = ~n26379 & ~n26394;
  assign n26396 = ~n26181 & n26376;
  assign n26397 = n26181 & ~n26376;
  assign n26398 = ~n26396 & ~n26397;
  assign n26399 = ~n26385 & ~n26389;
  assign n26400 = ~n26384 & n26399;
  assign n26401 = n26385 & ~n26392;
  assign n26402 = ~n26400 & ~n26401;
  assign n26403 = ~n26398 & ~n26402;
  assign n26404 = ~n26395 & ~n26403;
  assign n26405 = ~n24569 & ~n24570;
  assign n26406 = n24569 & n24570;
  assign n26407 = ~n24589 & ~n26406;
  assign n26408 = ~n26405 & ~n26407;
  assign n26409 = n26404 & n26408;
  assign n26410 = ~n26404 & ~n26408;
  assign n26411 = ~n26409 & ~n26410;
  assign n26412 = pi141 & pi273;
  assign n26413 = n24609 & ~n24615;
  assign n26414 = ~n24614 & ~n26413;
  assign n26415 = n26412 & ~n26414;
  assign n26416 = ~n24609 & ~n24614;
  assign n26417 = ~n24615 & ~n26416;
  assign n26418 = ~n26412 & ~n26417;
  assign n26419 = ~n26415 & ~n26418;
  assign n26420 = ~n26411 & ~n26419;
  assign n26421 = n26404 & ~n26408;
  assign n26422 = ~n26404 & n26408;
  assign n26423 = ~n26421 & ~n26422;
  assign n26424 = ~n26412 & ~n26414;
  assign n26425 = n26412 & ~n26417;
  assign n26426 = ~n26424 & ~n26425;
  assign n26427 = ~n26423 & ~n26426;
  assign n26428 = ~n26420 & ~n26427;
  assign n26429 = ~n26180 & ~n26428;
  assign n26430 = n26180 & n26428;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = pi272 & ~n24616;
  assign n26433 = pi141 & n26432;
  assign n26434 = ~n24607 & ~n24609;
  assign n26435 = ~n24608 & ~n26434;
  assign n26436 = ~n26433 & n26435;
  assign n26437 = pi143 & pi271;
  assign n26438 = ~n26433 & ~n26434;
  assign n26439 = pi271 & ~n26438;
  assign n26440 = pi142 & n26439;
  assign n26441 = n24626 & ~n26440;
  assign n26442 = n26437 & ~n26441;
  assign n26443 = ~n26436 & n26442;
  assign n26444 = ~n26436 & ~n26441;
  assign n26445 = ~n26437 & ~n26444;
  assign n26446 = ~n26443 & ~n26445;
  assign n26447 = ~n26431 & ~n26446;
  assign n26448 = ~n26180 & n26428;
  assign n26449 = n26180 & ~n26428;
  assign n26450 = ~n26448 & ~n26449;
  assign n26451 = ~n26437 & ~n26441;
  assign n26452 = ~n26436 & n26451;
  assign n26453 = n26437 & ~n26444;
  assign n26454 = ~n26452 & ~n26453;
  assign n26455 = ~n26450 & ~n26454;
  assign n26456 = ~n26447 & ~n26455;
  assign n26457 = ~n24630 & ~n24655;
  assign n26458 = n24630 & n24655;
  assign n26459 = ~n24649 & ~n26458;
  assign n26460 = ~n26457 & ~n26459;
  assign n26461 = n26456 & ~n26460;
  assign n26462 = ~n26456 & n26460;
  assign n26463 = ~n26461 & ~n26462;
  assign n26464 = pi144 & pi270;
  assign n26465 = n24669 & ~n24674;
  assign n26466 = ~n24675 & ~n26465;
  assign n26467 = n26464 & ~n26466;
  assign n26468 = ~n24669 & ~n24675;
  assign n26469 = ~n24674 & ~n26468;
  assign n26470 = ~n26464 & ~n26469;
  assign n26471 = ~n26467 & ~n26470;
  assign n26472 = ~n26463 & ~n26471;
  assign n26473 = n26456 & n26460;
  assign n26474 = ~n26456 & ~n26460;
  assign n26475 = ~n26473 & ~n26474;
  assign n26476 = ~n26464 & ~n26466;
  assign n26477 = n26464 & ~n26469;
  assign n26478 = ~n26476 & ~n26477;
  assign n26479 = ~n26475 & ~n26478;
  assign n26480 = ~n26472 & ~n26479;
  assign n26481 = ~n26179 & n26480;
  assign n26482 = n26179 & ~n26480;
  assign n26483 = ~n26481 & ~n26482;
  assign n26484 = pi269 & ~n24676;
  assign n26485 = pi144 & n26484;
  assign n26486 = ~n24667 & ~n24669;
  assign n26487 = ~n26485 & ~n26486;
  assign n26488 = pi268 & ~n26487;
  assign n26489 = pi145 & n26488;
  assign n26490 = pi146 & pi268;
  assign n26491 = ~n24668 & ~n26486;
  assign n26492 = ~n26485 & n26491;
  assign n26493 = ~n24685 & ~n26492;
  assign n26494 = ~n26490 & ~n26493;
  assign n26495 = ~n26489 & n26494;
  assign n26496 = ~n26489 & ~n26493;
  assign n26497 = n26490 & ~n26496;
  assign n26498 = ~n26495 & ~n26497;
  assign n26499 = ~n26483 & ~n26498;
  assign n26500 = ~n26179 & ~n26480;
  assign n26501 = n26179 & n26480;
  assign n26502 = ~n26500 & ~n26501;
  assign n26503 = n26490 & ~n26493;
  assign n26504 = ~n26489 & n26503;
  assign n26505 = ~n26490 & ~n26496;
  assign n26506 = ~n26504 & ~n26505;
  assign n26507 = ~n26502 & ~n26506;
  assign n26508 = ~n26499 & ~n26507;
  assign n26509 = ~n24689 & ~n24714;
  assign n26510 = n24689 & n24714;
  assign n26511 = ~n24708 & ~n26510;
  assign n26512 = ~n26509 & ~n26511;
  assign n26513 = n26508 & ~n26512;
  assign n26514 = ~n26508 & n26512;
  assign n26515 = ~n26513 & ~n26514;
  assign n26516 = pi147 & pi267;
  assign n26517 = n24728 & ~n24733;
  assign n26518 = ~n24734 & ~n26517;
  assign n26519 = n26516 & ~n26518;
  assign n26520 = ~n24728 & ~n24734;
  assign n26521 = ~n24733 & ~n26520;
  assign n26522 = ~n26516 & ~n26521;
  assign n26523 = ~n26519 & ~n26522;
  assign n26524 = ~n26515 & ~n26523;
  assign n26525 = n26508 & n26512;
  assign n26526 = ~n26508 & ~n26512;
  assign n26527 = ~n26525 & ~n26526;
  assign n26528 = ~n26516 & ~n26518;
  assign n26529 = n26516 & ~n26521;
  assign n26530 = ~n26528 & ~n26529;
  assign n26531 = ~n26527 & ~n26530;
  assign n26532 = ~n26524 & ~n26531;
  assign n26533 = ~n26178 & n26532;
  assign n26534 = n26178 & ~n26532;
  assign n26535 = ~n26533 & ~n26534;
  assign n26536 = pi266 & ~n24735;
  assign n26537 = pi147 & n26536;
  assign n26538 = ~n24726 & ~n24728;
  assign n26539 = ~n26537 & ~n26538;
  assign n26540 = pi265 & ~n26539;
  assign n26541 = pi148 & n26540;
  assign n26542 = pi149 & pi265;
  assign n26543 = ~n24727 & ~n26538;
  assign n26544 = ~n26537 & n26543;
  assign n26545 = ~n24744 & ~n26544;
  assign n26546 = ~n26542 & ~n26545;
  assign n26547 = ~n26541 & n26546;
  assign n26548 = ~n26541 & ~n26545;
  assign n26549 = n26542 & ~n26548;
  assign n26550 = ~n26547 & ~n26549;
  assign n26551 = ~n26535 & ~n26550;
  assign n26552 = ~n26178 & ~n26532;
  assign n26553 = n26178 & n26532;
  assign n26554 = ~n26552 & ~n26553;
  assign n26555 = n26542 & ~n26545;
  assign n26556 = ~n26541 & n26555;
  assign n26557 = ~n26542 & ~n26548;
  assign n26558 = ~n26556 & ~n26557;
  assign n26559 = ~n26554 & ~n26558;
  assign n26560 = ~n26551 & ~n26559;
  assign n26561 = n24748 & ~n24773;
  assign n26562 = ~n24748 & n24773;
  assign n26563 = ~n24764 & ~n26562;
  assign n26564 = ~n26561 & ~n26563;
  assign n26565 = n26560 & n26564;
  assign n26566 = ~n26560 & ~n26564;
  assign n26567 = ~n26565 & ~n26566;
  assign n26568 = pi150 & pi264;
  assign n26569 = n24787 & ~n24793;
  assign n26570 = ~n24792 & ~n26569;
  assign n26571 = n26568 & ~n26570;
  assign n26572 = ~n24787 & ~n24792;
  assign n26573 = ~n24793 & ~n26572;
  assign n26574 = ~n26568 & ~n26573;
  assign n26575 = ~n26571 & ~n26574;
  assign n26576 = ~n26567 & ~n26575;
  assign n26577 = n26560 & ~n26564;
  assign n26578 = ~n26560 & n26564;
  assign n26579 = ~n26577 & ~n26578;
  assign n26580 = ~n26568 & ~n26570;
  assign n26581 = n26568 & ~n26573;
  assign n26582 = ~n26580 & ~n26581;
  assign n26583 = ~n26579 & ~n26582;
  assign n26584 = ~n26576 & ~n26583;
  assign n26585 = ~n26177 & n26584;
  assign n26586 = n26177 & ~n26584;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = pi263 & ~n24794;
  assign n26589 = pi150 & n26588;
  assign n26590 = ~n24785 & ~n24787;
  assign n26591 = ~n26589 & ~n26590;
  assign n26592 = pi262 & ~n26591;
  assign n26593 = pi151 & n26592;
  assign n26594 = pi152 & pi262;
  assign n26595 = ~n24786 & ~n26590;
  assign n26596 = ~n26589 & n26595;
  assign n26597 = ~n24812 & ~n26596;
  assign n26598 = ~n26594 & ~n26597;
  assign n26599 = ~n26593 & n26598;
  assign n26600 = ~n26593 & ~n26597;
  assign n26601 = n26594 & ~n26600;
  assign n26602 = ~n26599 & ~n26601;
  assign n26603 = ~n26587 & ~n26602;
  assign n26604 = ~n26177 & ~n26584;
  assign n26605 = n26177 & n26584;
  assign n26606 = ~n26604 & ~n26605;
  assign n26607 = n26594 & ~n26597;
  assign n26608 = ~n26593 & n26607;
  assign n26609 = ~n26594 & ~n26600;
  assign n26610 = ~n26608 & ~n26609;
  assign n26611 = ~n26606 & ~n26610;
  assign n26612 = ~n26603 & ~n26611;
  assign n26613 = n24816 & ~n24857;
  assign n26614 = ~n24816 & n24857;
  assign n26615 = ~n24848 & ~n26614;
  assign n26616 = ~n26613 & ~n26615;
  assign n26617 = n26612 & ~n26616;
  assign n26618 = ~n26612 & n26616;
  assign n26619 = ~n26617 & ~n26618;
  assign n26620 = pi153 & pi261;
  assign n26621 = n24872 & ~n24900;
  assign n26622 = ~n24899 & ~n26621;
  assign n26623 = n26620 & ~n26622;
  assign n26624 = ~n24872 & ~n24899;
  assign n26625 = ~n24900 & ~n26624;
  assign n26626 = ~n26620 & ~n26625;
  assign n26627 = ~n26623 & ~n26626;
  assign n26628 = ~n26619 & ~n26627;
  assign n26629 = n26612 & n26616;
  assign n26630 = ~n26612 & ~n26616;
  assign n26631 = ~n26629 & ~n26630;
  assign n26632 = ~n26620 & ~n26622;
  assign n26633 = n26620 & ~n26625;
  assign n26634 = ~n26632 & ~n26633;
  assign n26635 = ~n26631 & ~n26634;
  assign n26636 = ~n26628 & ~n26635;
  assign n26637 = n24871 & n24884;
  assign n26638 = n24872 & ~n24901;
  assign n26639 = ~n24870 & ~n24872;
  assign n26640 = ~n26638 & ~n26639;
  assign n26641 = ~n24871 & ~n24884;
  assign n26642 = ~n26640 & ~n26641;
  assign n26643 = ~n26637 & ~n26642;
  assign n26644 = n26636 & ~n26643;
  assign n26645 = ~n26636 & n26643;
  assign n26646 = ~n26644 & ~n26645;
  assign n26647 = pi155 & pi259;
  assign n26648 = pi154 & pi260;
  assign n26649 = ~n26647 & ~n26648;
  assign n26650 = n26647 & n26648;
  assign n26651 = ~n26649 & ~n26650;
  assign n26652 = ~n24875 & n24884;
  assign n26653 = ~n24884 & ~n24892;
  assign n26654 = ~n26652 & ~n26653;
  assign n26655 = ~n24901 & ~n26654;
  assign n26656 = n24884 & ~n24892;
  assign n26657 = ~n24875 & ~n24884;
  assign n26658 = ~n26656 & ~n26657;
  assign n26659 = ~n24870 & ~n26658;
  assign n26660 = ~n26655 & ~n26659;
  assign n26661 = n24885 & ~n26660;
  assign n26662 = pi156 & pi258;
  assign n26663 = n26661 & n26662;
  assign n26664 = ~n26661 & ~n26662;
  assign n26665 = ~n26663 & ~n26664;
  assign n26666 = ~n26651 & ~n26665;
  assign n26667 = n26647 & ~n26648;
  assign n26668 = ~n26647 & n26648;
  assign n26669 = ~n26667 & ~n26668;
  assign n26670 = ~n26661 & n26662;
  assign n26671 = n26661 & ~n26662;
  assign n26672 = ~n26670 & ~n26671;
  assign n26673 = ~n26669 & ~n26672;
  assign n26674 = ~n26666 & ~n26673;
  assign n26675 = ~n26646 & ~n26674;
  assign n26676 = n26636 & n26643;
  assign n26677 = ~n26636 & ~n26643;
  assign n26678 = ~n26676 & ~n26677;
  assign n26679 = ~n26665 & ~n26669;
  assign n26680 = ~n26651 & ~n26672;
  assign n26681 = ~n26679 & ~n26680;
  assign n26682 = ~n26678 & ~n26681;
  assign n26683 = ~n26675 & ~n26682;
  assign n26684 = ~n22545 & ~n24913;
  assign n26685 = n22545 & ~n24912;
  assign n26686 = ~n22557 & ~n26685;
  assign n26687 = ~n26684 & ~n26686;
  assign n26688 = n26683 & n26687;
  assign n26689 = ~n26683 & ~n26687;
  assign n26690 = ~n26688 & ~n26689;
  assign n26691 = ~n24906 & ~n26690;
  assign n26692 = n26683 & ~n26687;
  assign n26693 = ~n26683 & n26687;
  assign n26694 = ~n26692 & ~n26693;
  assign n26695 = n24906 & ~n26694;
  assign n26696 = ~n26691 & ~n26695;
  assign n26697 = pi322 & ~n26696;
  assign n26698 = ~n26176 & ~n26697;
  assign n26699 = n26175 & ~n26696;
  assign n26700 = pi323 & n26699;
  assign n26701 = pi322 & n26700;
  assign n26702 = ~n26698 & ~n26701;
  assign n26703 = pi325 & n21479;
  assign n26704 = ~n22557 & ~n24926;
  assign n26705 = n22557 & ~n24919;
  assign n26706 = ~n26704 & ~n26705;
  assign n26707 = pi324 & n26706;
  assign n26708 = n26703 & n26707;
  assign n26709 = ~n26703 & ~n26707;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = ~n26702 & ~n26710;
  assign n26712 = ~n26703 & n26707;
  assign n26713 = n26703 & ~n26707;
  assign n26714 = ~n26712 & ~n26713;
  assign n26715 = ~n26701 & ~n26714;
  assign n26716 = ~n26698 & n26715;
  assign n26717 = ~n26711 & ~n26716;
  assign n26718 = ~n26166 & ~n26717;
  assign n26719 = ~n26155 & ~n26163;
  assign n26720 = n26155 & n26163;
  assign n26721 = ~n26719 & ~n26720;
  assign n26722 = ~n26702 & ~n26714;
  assign n26723 = ~n26701 & ~n26710;
  assign n26724 = ~n26698 & n26723;
  assign n26725 = ~n26722 & ~n26724;
  assign n26726 = ~n26721 & ~n26725;
  assign n26727 = ~n26718 & ~n26726;
  assign n26728 = n24941 & ~n24977;
  assign n26729 = ~n24939 & ~n24942;
  assign n26730 = ~n24931 & n26729;
  assign n26731 = n21479 & ~n24940;
  assign n26732 = pi324 & n26731;
  assign n26733 = ~n26730 & ~n26732;
  assign n26734 = ~n24956 & ~n26733;
  assign n26735 = ~n24940 & ~n24942;
  assign n26736 = n24940 & n24942;
  assign n26737 = ~n26735 & ~n26736;
  assign n26738 = ~n24308 & ~n26737;
  assign n26739 = ~n26734 & ~n26738;
  assign n26740 = ~n24941 & n24977;
  assign n26741 = ~n26739 & ~n26740;
  assign n26742 = ~n26728 & ~n26741;
  assign n26743 = n26727 & n26742;
  assign n26744 = ~n26727 & ~n26742;
  assign n26745 = ~n26743 & ~n26744;
  assign n26746 = pi327 & n19557;
  assign n26747 = pi326 & n19970;
  assign n26748 = n26746 & n26747;
  assign n26749 = ~n26746 & ~n26747;
  assign n26750 = ~n26748 & ~n26749;
  assign n26751 = ~n26745 & ~n26750;
  assign n26752 = ~n26727 & n26742;
  assign n26753 = n26727 & ~n26742;
  assign n26754 = ~n26752 & ~n26753;
  assign n26755 = ~n26746 & n26747;
  assign n26756 = n26746 & ~n26747;
  assign n26757 = ~n26755 & ~n26756;
  assign n26758 = ~n26754 & ~n26757;
  assign n26759 = ~n26751 & ~n26758;
  assign n26760 = ~n26153 & ~n26759;
  assign n26761 = n26130 & ~n26150;
  assign n26762 = ~n26130 & n26150;
  assign n26763 = ~n26761 & ~n26762;
  assign n26764 = ~n26750 & ~n26754;
  assign n26765 = ~n26745 & ~n26757;
  assign n26766 = ~n26764 & ~n26765;
  assign n26767 = ~n26763 & ~n26766;
  assign n26768 = ~n26760 & ~n26767;
  assign n26769 = ~n26126 & n26768;
  assign n26770 = n26126 & ~n26768;
  assign n26771 = ~n26769 & ~n26770;
  assign n26772 = n19539 & ~n26771;
  assign n26773 = pi328 & n26772;
  assign n26774 = pi328 & n19539;
  assign n26775 = n26126 & n26768;
  assign n26776 = ~n26126 & ~n26768;
  assign n26777 = ~n26775 & ~n26776;
  assign n26778 = ~n26774 & ~n26777;
  assign n26779 = ~n26773 & ~n26778;
  assign n26780 = ~n26125 & ~n26779;
  assign n26781 = n26110 & ~n26122;
  assign n26782 = ~n26110 & n26122;
  assign n26783 = ~n26781 & ~n26782;
  assign n26784 = n19539 & ~n26777;
  assign n26785 = pi328 & n26784;
  assign n26786 = ~n26771 & ~n26774;
  assign n26787 = ~n26785 & ~n26786;
  assign n26788 = ~n26783 & ~n26787;
  assign n26789 = ~n26780 & ~n26788;
  assign n26790 = ~n25028 & n25032;
  assign n26791 = n25028 & ~n25032;
  assign n26792 = n11711 & ~n25049;
  assign n26793 = ~n25050 & ~n26792;
  assign n26794 = n12917 & ~n26793;
  assign n26795 = pi330 & n26794;
  assign n26796 = ~n12917 & ~n26792;
  assign n26797 = pi330 & ~n26796;
  assign n26798 = ~n25050 & ~n26797;
  assign n26799 = ~n26795 & ~n26798;
  assign n26800 = n25024 & ~n26799;
  assign n26801 = ~n25024 & n26799;
  assign n26802 = ~n26800 & ~n26801;
  assign n26803 = ~n26791 & ~n26802;
  assign n26804 = ~n26790 & ~n26803;
  assign n26805 = n26789 & n26804;
  assign n26806 = ~n26789 & ~n26804;
  assign n26807 = ~n26805 & ~n26806;
  assign n26808 = pi331 & n12917;
  assign n26809 = n25024 & ~n26798;
  assign n26810 = ~n26795 & ~n26809;
  assign n26811 = n13762 & n26810;
  assign n26812 = pi330 & n26811;
  assign n26813 = pi330 & n13762;
  assign n26814 = ~n26810 & ~n26813;
  assign n26815 = ~n26812 & ~n26814;
  assign n26816 = ~n26808 & n26815;
  assign n26817 = n26808 & ~n26815;
  assign n26818 = ~n26816 & ~n26817;
  assign n26819 = pi332 & n11711;
  assign n26820 = n22004 & ~n24207;
  assign n26821 = ~n22004 & ~n24216;
  assign n26822 = ~n26820 & ~n26821;
  assign n26823 = ~n25067 & ~n26822;
  assign n26824 = ~n25070 & ~n26823;
  assign n26825 = n25066 & ~n26824;
  assign n26826 = ~n25064 & ~n26825;
  assign n26827 = ~n25101 & n26826;
  assign n26828 = ~n25066 & n26824;
  assign n26829 = ~n25092 & ~n26825;
  assign n26830 = ~n25031 & n26829;
  assign n26831 = ~n26828 & ~n26830;
  assign n26832 = ~n26827 & n26831;
  assign n26833 = n26819 & ~n26832;
  assign n26834 = ~n26819 & n26832;
  assign n26835 = ~n26833 & ~n26834;
  assign n26836 = ~n26818 & ~n26835;
  assign n26837 = n26808 & n26815;
  assign n26838 = ~n26808 & ~n26815;
  assign n26839 = ~n26837 & ~n26838;
  assign n26840 = ~n26819 & ~n26832;
  assign n26841 = n26819 & n26832;
  assign n26842 = ~n26840 & ~n26841;
  assign n26843 = ~n26839 & ~n26842;
  assign n26844 = ~n26836 & ~n26843;
  assign n26845 = ~n26807 & ~n26844;
  assign n26846 = n26789 & ~n26804;
  assign n26847 = ~n26789 & n26804;
  assign n26848 = ~n26846 & ~n26847;
  assign n26849 = ~n26835 & ~n26839;
  assign n26850 = ~n26818 & ~n26842;
  assign n26851 = ~n26849 & ~n26850;
  assign n26852 = ~n26848 & ~n26851;
  assign n26853 = ~n26845 & ~n26852;
  assign n26854 = ~n26105 & n26853;
  assign n26855 = n26105 & ~n26853;
  assign n26856 = ~n26854 & ~n26855;
  assign n26857 = pi335 & n10561;
  assign n26858 = n9205 & ~n24235;
  assign n26859 = pi334 & n26858;
  assign n26860 = ~n24236 & ~n26859;
  assign n26861 = ~pi334 & ~n26860;
  assign n26862 = ~n24244 & n26860;
  assign n26863 = ~n11366 & ~n26862;
  assign n26864 = ~n26861 & ~n26863;
  assign n26865 = ~n26096 & ~n26864;
  assign n26866 = ~n11366 & ~n26860;
  assign n26867 = n10561 & n26866;
  assign n26868 = ~n10561 & n26860;
  assign n26869 = n10561 & ~n26860;
  assign n26870 = ~n26092 & ~n26869;
  assign n26871 = ~n26868 & ~n26870;
  assign n26872 = n11366 & ~n26871;
  assign n26873 = ~n26867 & ~n26872;
  assign n26874 = pi334 & ~n26873;
  assign n26875 = ~n26865 & ~n26874;
  assign n26876 = n26857 & ~n26875;
  assign n26877 = ~n26857 & n26875;
  assign n26878 = ~n26876 & ~n26877;
  assign n26879 = ~n26856 & ~n26878;
  assign n26880 = n26105 & n26853;
  assign n26881 = ~n26105 & ~n26853;
  assign n26882 = ~n26880 & ~n26881;
  assign n26883 = ~n26857 & ~n26875;
  assign n26884 = n26857 & n26875;
  assign n26885 = ~n26883 & ~n26884;
  assign n26886 = ~n26882 & ~n26885;
  assign n26887 = ~n26879 & ~n26886;
  assign n26888 = ~n26104 & ~n26887;
  assign n26889 = ~n26087 & ~n26101;
  assign n26890 = n26087 & n26101;
  assign n26891 = ~n26889 & ~n26890;
  assign n26892 = ~n26878 & ~n26882;
  assign n26893 = ~n26856 & ~n26885;
  assign n26894 = ~n26892 & ~n26893;
  assign n26895 = ~n26891 & ~n26894;
  assign n26896 = ~n26888 & ~n26895;
  assign n26897 = ~n25131 & n25135;
  assign n26898 = ~n25127 & ~n25146;
  assign n26899 = n25127 & n25146;
  assign n26900 = ~n26898 & ~n26899;
  assign n26901 = n25131 & ~n25135;
  assign n26902 = ~n26900 & ~n26901;
  assign n26903 = ~n26897 & ~n26902;
  assign n26904 = n26896 & n26903;
  assign n26905 = ~n26896 & ~n26903;
  assign n26906 = ~n26904 & ~n26905;
  assign n26907 = pi337 & n6556;
  assign n26908 = ~n25127 & ~n25141;
  assign n26909 = n25127 & n25141;
  assign n26910 = ~n6556 & ~n26909;
  assign n26911 = ~n26908 & ~n26910;
  assign n26912 = n9205 & ~n26911;
  assign n26913 = ~n9205 & ~n26908;
  assign n26914 = n6556 & n26913;
  assign n26915 = ~n26912 & ~n26914;
  assign n26916 = pi336 & ~n26915;
  assign n26917 = pi336 & n9205;
  assign n26918 = n25127 & ~n26917;
  assign n26919 = n25141 & n26918;
  assign n26920 = ~n26916 & ~n26919;
  assign n26921 = ~n26907 & n26920;
  assign n26922 = n26907 & ~n26920;
  assign n26923 = ~n26921 & ~n26922;
  assign n26924 = pi338 & n5973;
  assign n26925 = ~n25149 & ~n25186;
  assign n26926 = ~n25134 & ~n25177;
  assign n26927 = ~n26033 & ~n26926;
  assign n26928 = ~n26925 & n26927;
  assign n26929 = ~n26027 & ~n26928;
  assign n26930 = n26924 & n26929;
  assign n26931 = ~n26924 & ~n26929;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = ~n26923 & ~n26932;
  assign n26934 = n26907 & n26920;
  assign n26935 = ~n26907 & ~n26920;
  assign n26936 = ~n26934 & ~n26935;
  assign n26937 = ~n26924 & n26929;
  assign n26938 = n26924 & ~n26929;
  assign n26939 = ~n26937 & ~n26938;
  assign n26940 = ~n26936 & ~n26939;
  assign n26941 = ~n26933 & ~n26940;
  assign n26942 = ~n26906 & ~n26941;
  assign n26943 = n26896 & ~n26903;
  assign n26944 = ~n26896 & n26903;
  assign n26945 = ~n26943 & ~n26944;
  assign n26946 = ~n26932 & ~n26936;
  assign n26947 = ~n26923 & ~n26939;
  assign n26948 = ~n26946 & ~n26947;
  assign n26949 = ~n26945 & ~n26948;
  assign n26950 = ~n26942 & ~n26949;
  assign n26951 = ~n26066 & n26950;
  assign n26952 = n26066 & ~n26950;
  assign n26953 = ~n26951 & ~n26952;
  assign n26954 = pi341 & n5257;
  assign n26955 = n4596 & ~n24192;
  assign n26956 = pi340 & n26955;
  assign n26957 = ~n24193 & ~n26956;
  assign n26958 = ~pi340 & ~n26957;
  assign n26959 = ~n24201 & n26957;
  assign n26960 = ~n5714 & ~n26959;
  assign n26961 = ~n26958 & ~n26960;
  assign n26962 = ~n26057 & ~n26961;
  assign n26963 = ~n5714 & ~n26957;
  assign n26964 = n5257 & n26963;
  assign n26965 = ~n5257 & n26957;
  assign n26966 = n5257 & ~n26957;
  assign n26967 = ~n26053 & ~n26966;
  assign n26968 = ~n26965 & ~n26967;
  assign n26969 = n5714 & ~n26968;
  assign n26970 = ~n26964 & ~n26969;
  assign n26971 = pi340 & ~n26970;
  assign n26972 = ~n26962 & ~n26971;
  assign n26973 = n26954 & ~n26972;
  assign n26974 = ~n26954 & n26972;
  assign n26975 = ~n26973 & ~n26974;
  assign n26976 = ~n26953 & ~n26975;
  assign n26977 = n26066 & n26950;
  assign n26978 = ~n26066 & ~n26950;
  assign n26979 = ~n26977 & ~n26978;
  assign n26980 = ~n26954 & ~n26972;
  assign n26981 = n26954 & n26972;
  assign n26982 = ~n26980 & ~n26981;
  assign n26983 = ~n26979 & ~n26982;
  assign n26984 = ~n26976 & ~n26983;
  assign n26985 = ~n26065 & ~n26984;
  assign n26986 = ~n26048 & ~n26062;
  assign n26987 = n26048 & n26062;
  assign n26988 = ~n26986 & ~n26987;
  assign n26989 = ~n26975 & ~n26979;
  assign n26990 = ~n26953 & ~n26982;
  assign n26991 = ~n26989 & ~n26990;
  assign n26992 = ~n26988 & ~n26991;
  assign n26993 = ~n26985 & ~n26992;
  assign n26994 = ~n25216 & n25220;
  assign n26995 = ~n25212 & ~n25231;
  assign n26996 = n25212 & n25231;
  assign n26997 = ~n26995 & ~n26996;
  assign n26998 = n25216 & ~n25220;
  assign n26999 = ~n26997 & ~n26998;
  assign n27000 = ~n26994 & ~n26999;
  assign n27001 = n26993 & n27000;
  assign n27002 = ~n26993 & ~n27000;
  assign n27003 = ~n27001 & ~n27002;
  assign n27004 = pi343 & n2887;
  assign n27005 = ~n25212 & ~n25226;
  assign n27006 = n25212 & n25226;
  assign n27007 = ~n2887 & ~n27006;
  assign n27008 = ~n27005 & ~n27007;
  assign n27009 = n4596 & ~n27008;
  assign n27010 = ~n4596 & ~n27005;
  assign n27011 = n2887 & n27010;
  assign n27012 = ~n27009 & ~n27011;
  assign n27013 = pi342 & ~n27012;
  assign n27014 = pi342 & n4596;
  assign n27015 = n25212 & ~n27014;
  assign n27016 = n25226 & n27015;
  assign n27017 = ~n27013 & ~n27016;
  assign n27018 = ~n27004 & n27017;
  assign n27019 = n27004 & ~n27017;
  assign n27020 = ~n27018 & ~n27019;
  assign n27021 = pi344 & n2464;
  assign n27022 = ~n25234 & ~n25252;
  assign n27023 = ~n25259 & n27022;
  assign n27024 = ~n25250 & ~n25252;
  assign n27025 = ~n25219 & n27024;
  assign n27026 = ~n25251 & ~n27025;
  assign n27027 = ~n27023 & n27026;
  assign n27028 = n27021 & ~n27027;
  assign n27029 = ~n27021 & n27027;
  assign n27030 = ~n27028 & ~n27029;
  assign n27031 = ~n27020 & ~n27030;
  assign n27032 = n27004 & n27017;
  assign n27033 = ~n27004 & ~n27017;
  assign n27034 = ~n27032 & ~n27033;
  assign n27035 = ~n27021 & ~n27027;
  assign n27036 = n27021 & n27027;
  assign n27037 = ~n27035 & ~n27036;
  assign n27038 = ~n27034 & ~n27037;
  assign n27039 = ~n27031 & ~n27038;
  assign n27040 = ~n27003 & ~n27039;
  assign n27041 = n26993 & ~n27000;
  assign n27042 = ~n26993 & n27000;
  assign n27043 = ~n27041 & ~n27042;
  assign n27044 = ~n27030 & ~n27034;
  assign n27045 = ~n27020 & ~n27037;
  assign n27046 = ~n27044 & ~n27045;
  assign n27047 = ~n27043 & ~n27046;
  assign n27048 = ~n27040 & ~n27047;
  assign n27049 = ~n26020 & n27048;
  assign n27050 = n26020 & ~n27048;
  assign n27051 = ~n27049 & ~n27050;
  assign n27052 = pi347 & n1442;
  assign n27053 = ~n25269 & ~n25273;
  assign n27054 = ~n24148 & n27053;
  assign n27055 = pi346 & n1729;
  assign n27056 = n24161 & ~n27055;
  assign n27057 = ~n27054 & n27056;
  assign n27058 = n1442 & ~n25270;
  assign n27059 = pi346 & n27058;
  assign n27060 = ~n24161 & n27055;
  assign n27061 = ~n27059 & n27060;
  assign n27062 = ~n27057 & ~n27061;
  assign n27063 = ~n25999 & ~n27062;
  assign n27064 = n24161 & n27055;
  assign n27065 = ~n27059 & n27064;
  assign n27066 = ~n24161 & ~n27055;
  assign n27067 = ~n27054 & n27066;
  assign n27068 = ~n27065 & ~n27067;
  assign n27069 = ~n26008 & ~n27068;
  assign n27070 = ~n27055 & n27059;
  assign n27071 = n27054 & n27055;
  assign n27072 = ~n27059 & n27071;
  assign n27073 = ~n27070 & ~n27072;
  assign n27074 = ~n27069 & n27073;
  assign n27075 = ~n27063 & n27074;
  assign n27076 = n27052 & ~n27075;
  assign n27077 = ~n27052 & n27075;
  assign n27078 = ~n27076 & ~n27077;
  assign n27079 = ~n27051 & ~n27078;
  assign n27080 = n26020 & n27048;
  assign n27081 = ~n26020 & ~n27048;
  assign n27082 = ~n27080 & ~n27081;
  assign n27083 = ~n27052 & ~n27075;
  assign n27084 = n27052 & n27075;
  assign n27085 = ~n27083 & ~n27084;
  assign n27086 = ~n27082 & ~n27085;
  assign n27087 = ~n27079 & ~n27086;
  assign n27088 = ~n26019 & ~n27087;
  assign n27089 = ~n25996 & n26016;
  assign n27090 = n25996 & ~n26016;
  assign n27091 = ~n27089 & ~n27090;
  assign n27092 = ~n27078 & ~n27082;
  assign n27093 = ~n27051 & ~n27085;
  assign n27094 = ~n27092 & ~n27093;
  assign n27095 = ~n27091 & ~n27094;
  assign n27096 = ~n27088 & ~n27095;
  assign n27097 = n25992 & ~n27096;
  assign n27098 = ~n25992 & n27096;
  assign n27099 = ~n27097 & ~n27098;
  assign n27100 = n24122 & n25296;
  assign n27101 = ~n24122 & ~n25296;
  assign n27102 = ~n1154 & ~n27101;
  assign n27103 = ~n27100 & ~n27102;
  assign n27104 = ~n1256 & ~n27103;
  assign n27105 = pi348 & n27104;
  assign n27106 = ~n1154 & n25296;
  assign n27107 = n1256 & ~n27106;
  assign n27108 = pi348 & ~n27107;
  assign n27109 = n1154 & ~n25296;
  assign n27110 = n24122 & ~n27109;
  assign n27111 = ~n27108 & ~n27110;
  assign n27112 = ~n27105 & ~n27111;
  assign n27113 = ~n1154 & ~n27112;
  assign n27114 = pi349 & n27113;
  assign n27115 = pi349 & ~n1154;
  assign n27116 = ~n27111 & ~n27115;
  assign n27117 = ~n27105 & n27116;
  assign n27118 = ~n27114 & ~n27117;
  assign n27119 = ~n27099 & ~n27118;
  assign n27120 = n25992 & n27096;
  assign n27121 = ~n25992 & ~n27096;
  assign n27122 = ~n27120 & ~n27121;
  assign n27123 = ~n27112 & ~n27115;
  assign n27124 = n27112 & n27115;
  assign n27125 = ~n27123 & ~n27124;
  assign n27126 = ~n27122 & ~n27125;
  assign n27127 = ~n27119 & ~n27126;
  assign n27128 = pi286 & ~n27127;
  assign n27129 = ~pi286 & n27127;
  assign n27130 = ~n27128 & ~n27129;
  assign n27131 = pi258 & ~n27130;
  assign n27132 = pi128 & n27131;
  assign n27133 = pi350 & n27132;
  assign n27134 = pi286 & n27127;
  assign n27135 = ~pi286 & ~n27127;
  assign n27136 = ~n27134 & ~n27135;
  assign n27137 = pi350 & n1156;
  assign n27138 = ~n27136 & ~n27137;
  assign n27139 = ~n27133 & ~n27138;
  assign n27140 = ~n25989 & ~n27139;
  assign n27141 = n25989 & n27139;
  assign n27142 = ~n27140 & ~n27141;
  assign n27143 = ~n25983 & ~n27142;
  assign n27144 = ~n25989 & n27139;
  assign n27145 = n25989 & ~n27139;
  assign n27146 = ~n27144 & ~n27145;
  assign n27147 = n25983 & ~n27146;
  assign n27148 = ~n27143 & ~n27147;
  assign n27149 = ~n25324 & ~n25346;
  assign n27150 = n25324 & n25346;
  assign n27151 = n24117 & ~n25330;
  assign n27152 = ~n25961 & ~n27151;
  assign n27153 = ~n27150 & ~n27152;
  assign n27154 = ~n27149 & ~n27153;
  assign n27155 = n27148 & n27154;
  assign n27156 = ~n27148 & ~n27154;
  assign n27157 = ~n27155 & ~n27156;
  assign n27158 = ~n831 & ~n27157;
  assign n27159 = ~n25356 & ~n27158;
  assign n27160 = pi161 & ~n27159;
  assign n27161 = ~n25355 & ~n27160;
  assign po221 = ~pi160 & n27161;
  assign n27163 = ~pi093 & ~pi161;
  assign n27164 = ~pi287 & n831;
  assign n27165 = ~n25965 & ~n25977;
  assign n27166 = ~n25960 & ~n25971;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = pi293 & ~n27167;
  assign n27169 = pi128 & n27168;
  assign n27170 = ~pi128 & pi293;
  assign n27171 = ~n27169 & ~n27170;
  assign n27172 = pi129 & ~n27171;
  assign n27173 = pi293 & ~n27169;
  assign n27174 = n1567 & n27173;
  assign n27175 = ~n27172 & ~n27174;
  assign n27176 = ~n25367 & ~n25923;
  assign n27177 = pi301 & n3552;
  assign n27178 = pi305 & n6777;
  assign n27179 = pi309 & n9815;
  assign n27180 = pi313 & n14618;
  assign n27181 = ~n25540 & ~n25544;
  assign n27182 = ~n25545 & ~n27181;
  assign n27183 = pi154 & pi156;
  assign n27184 = ~n23615 & ~n27183;
  assign n27185 = pi153 & ~n27184;
  assign n27186 = ~pi155 & ~n25468;
  assign n27187 = pi154 & ~n27186;
  assign n27188 = ~n25461 & ~n27187;
  assign n27189 = ~n27185 & n27188;
  assign n27190 = pi157 & n27189;
  assign n27191 = ~pi157 & ~n27189;
  assign n27192 = ~n27190 & ~n27191;
  assign n27193 = pi156 & ~n27192;
  assign n27194 = pi157 & ~n27189;
  assign n27195 = ~pi157 & n27189;
  assign n27196 = ~n27194 & ~n27195;
  assign n27197 = ~pi156 & ~n27196;
  assign n27198 = ~n27193 & ~n27197;
  assign n27199 = ~n25451 & n25479;
  assign n27200 = ~pi320 & ~n27199;
  assign n27201 = ~n23626 & ~n25479;
  assign n27202 = n23626 & n25451;
  assign n27203 = pi320 & n27199;
  assign n27204 = ~n27202 & ~n27203;
  assign n27205 = ~n27201 & n27204;
  assign n27206 = ~n27200 & n27205;
  assign n27207 = n27198 & ~n27206;
  assign n27208 = ~n25451 & ~n27198;
  assign n27209 = ~pi320 & n25479;
  assign n27210 = n27208 & n27209;
  assign n27211 = ~n27207 & ~n27210;
  assign n27212 = pi321 & ~n27211;
  assign n27213 = n25451 & ~n27198;
  assign n27214 = ~n23626 & n27213;
  assign n27215 = n23626 & ~n25451;
  assign n27216 = ~pi321 & ~n27215;
  assign n27217 = ~n27214 & ~n27216;
  assign n27218 = n25479 & ~n27217;
  assign n27219 = pi321 & n27198;
  assign n27220 = ~n25451 & ~n27219;
  assign n27221 = ~n25479 & n27220;
  assign n27222 = n23626 & n27221;
  assign n27223 = ~n27218 & ~n27222;
  assign n27224 = pi320 & ~n27223;
  assign n27225 = ~n27212 & ~n27224;
  assign n27226 = pi319 & n23626;
  assign n27227 = ~n27225 & ~n27226;
  assign n27228 = n23626 & n27225;
  assign n27229 = pi319 & n27228;
  assign n27230 = ~n27227 & ~n27229;
  assign n27231 = ~n25451 & ~n25483;
  assign n27232 = pi320 & n27202;
  assign n27233 = ~n27231 & ~n27232;
  assign n27234 = ~n25482 & ~n27233;
  assign n27235 = n25451 & ~n25483;
  assign n27236 = pi320 & n27215;
  assign n27237 = ~n27235 & ~n27236;
  assign n27238 = n25479 & ~n27237;
  assign n27239 = pi321 & n27238;
  assign n27240 = ~n27234 & ~n27239;
  assign n27241 = ~n23671 & ~n27240;
  assign n27242 = ~n23658 & n27241;
  assign n27243 = ~n23069 & n27240;
  assign n27244 = ~n25498 & ~n27243;
  assign n27245 = n20347 & n27244;
  assign n27246 = ~n25497 & n27240;
  assign n27247 = n23069 & ~n27246;
  assign n27248 = ~n27245 & ~n27247;
  assign n27249 = pi319 & ~n27248;
  assign n27250 = ~n27242 & ~n27249;
  assign n27251 = ~n27230 & ~n27250;
  assign n27252 = n27230 & n27250;
  assign n27253 = ~n27251 & ~n27252;
  assign n27254 = n23069 & ~n27253;
  assign n27255 = pi318 & n27254;
  assign n27256 = pi318 & n23069;
  assign n27257 = n27230 & ~n27250;
  assign n27258 = ~n27230 & n27250;
  assign n27259 = ~n27257 & ~n27258;
  assign n27260 = ~n27256 & ~n27259;
  assign n27261 = ~n27255 & ~n27260;
  assign n27262 = ~n25507 & ~n25522;
  assign n27263 = ~n25529 & n27262;
  assign n27264 = n25520 & ~n27263;
  assign n27265 = ~n27261 & ~n27264;
  assign n27266 = n27261 & n27264;
  assign n27267 = ~n27265 & ~n27266;
  assign n27268 = n20347 & ~n27267;
  assign n27269 = pi317 & n27268;
  assign n27270 = pi317 & n20347;
  assign n27271 = ~n27266 & ~n27270;
  assign n27272 = ~n27265 & n27271;
  assign n27273 = ~n27269 & ~n27272;
  assign n27274 = ~n27182 & ~n27273;
  assign n27275 = n27182 & ~n27272;
  assign n27276 = ~n27269 & n27275;
  assign n27277 = ~n27274 & ~n27276;
  assign n27278 = ~n25532 & ~n25537;
  assign n27279 = ~n23693 & n27278;
  assign n27280 = n25532 & ~n25540;
  assign n27281 = ~n27279 & ~n27280;
  assign n27282 = ~n25439 & ~n27281;
  assign n27283 = n25532 & ~n25537;
  assign n27284 = ~n23693 & n27283;
  assign n27285 = ~n25532 & ~n25540;
  assign n27286 = ~n27284 & ~n27285;
  assign n27287 = n18937 & ~n27286;
  assign n27288 = pi317 & n27287;
  assign n27289 = ~n27282 & ~n27288;
  assign n27290 = ~n23723 & ~n27289;
  assign n27291 = ~n25437 & n27290;
  assign n27292 = ~n17455 & n27289;
  assign n27293 = ~n25578 & ~n27292;
  assign n27294 = n16985 & n27293;
  assign n27295 = ~n25438 & n27289;
  assign n27296 = n17455 & ~n27295;
  assign n27297 = ~n27294 & ~n27296;
  assign n27298 = pi316 & ~n27297;
  assign n27299 = ~n27291 & ~n27298;
  assign n27300 = n27277 & ~n27299;
  assign n27301 = ~n27277 & n27299;
  assign n27302 = ~n27300 & ~n27301;
  assign n27303 = pi316 & n18937;
  assign n27304 = pi315 & n17455;
  assign n27305 = ~n27303 & ~n27304;
  assign n27306 = n27303 & n27304;
  assign n27307 = ~n27305 & ~n27306;
  assign n27308 = ~n27302 & ~n27307;
  assign n27309 = ~n27277 & ~n27299;
  assign n27310 = n27277 & n27299;
  assign n27311 = ~n27309 & ~n27310;
  assign n27312 = n18937 & ~n27304;
  assign n27313 = pi316 & n27312;
  assign n27314 = n17455 & ~n27303;
  assign n27315 = pi315 & n27314;
  assign n27316 = ~n27313 & ~n27315;
  assign n27317 = ~n27311 & ~n27316;
  assign n27318 = ~n27308 & ~n27317;
  assign n27319 = ~n23703 & ~n25438;
  assign n27320 = ~n25578 & ~n27319;
  assign n27321 = ~n25552 & ~n27320;
  assign n27322 = ~n25582 & ~n27321;
  assign n27323 = ~n25593 & ~n27322;
  assign n27324 = n25593 & n27322;
  assign n27325 = n16985 & ~n27324;
  assign n27326 = pi315 & n27325;
  assign n27327 = ~n27323 & ~n27326;
  assign n27328 = n27318 & n27327;
  assign n27329 = ~n27318 & ~n27327;
  assign n27330 = ~n27328 & ~n27329;
  assign n27331 = pi314 & n16985;
  assign n27332 = ~n25604 & ~n27331;
  assign n27333 = ~n25598 & n27332;
  assign n27334 = ~n25598 & ~n25604;
  assign n27335 = n27331 & ~n27334;
  assign n27336 = ~n27333 & ~n27335;
  assign n27337 = ~n27330 & ~n27336;
  assign n27338 = n27318 & ~n27327;
  assign n27339 = ~n27318 & n27327;
  assign n27340 = ~n27338 & ~n27339;
  assign n27341 = ~n25604 & n27331;
  assign n27342 = ~n25598 & n27341;
  assign n27343 = ~n27331 & ~n27334;
  assign n27344 = ~n27342 & ~n27343;
  assign n27345 = ~n27340 & ~n27344;
  assign n27346 = ~n27337 & ~n27345;
  assign n27347 = ~n27180 & n27346;
  assign n27348 = n27180 & ~n27346;
  assign n27349 = ~n27347 & ~n27348;
  assign n27350 = pi312 & n14156;
  assign n27351 = n23222 & ~n23781;
  assign n27352 = n10908 & ~n25633;
  assign n27353 = pi313 & n27352;
  assign n27354 = ~n27351 & ~n27353;
  assign n27355 = ~n23770 & ~n27354;
  assign n27356 = n23222 & n27352;
  assign n27357 = ~n25634 & ~n27356;
  assign n27358 = pi313 & ~n27357;
  assign n27359 = ~n27355 & ~n27358;
  assign n27360 = n25606 & ~n27359;
  assign n27361 = ~n25606 & n27359;
  assign n27362 = n25421 & ~n27361;
  assign n27363 = ~n27360 & ~n27362;
  assign n27364 = n27350 & ~n27363;
  assign n27365 = ~n25421 & ~n27360;
  assign n27366 = ~n27361 & ~n27365;
  assign n27367 = ~n27350 & ~n27366;
  assign n27368 = ~n27364 & ~n27367;
  assign n27369 = ~n27349 & ~n27368;
  assign n27370 = ~n27180 & ~n27346;
  assign n27371 = n27180 & n27346;
  assign n27372 = ~n27370 & ~n27371;
  assign n27373 = ~n27350 & ~n27363;
  assign n27374 = n27350 & ~n27366;
  assign n27375 = ~n27373 & ~n27374;
  assign n27376 = ~n27372 & ~n27375;
  assign n27377 = ~n27369 & ~n27376;
  assign n27378 = n25610 & ~n25654;
  assign n27379 = ~n25610 & n25654;
  assign n27380 = ~n25645 & ~n27379;
  assign n27381 = ~n27378 & ~n27380;
  assign n27382 = n27377 & n27381;
  assign n27383 = ~n27377 & ~n27381;
  assign n27384 = ~n27382 & ~n27383;
  assign n27385 = pi311 & n11998;
  assign n27386 = n25665 & ~n25666;
  assign n27387 = ~n25667 & ~n27386;
  assign n27388 = n27385 & ~n27387;
  assign n27389 = ~n25665 & ~n25667;
  assign n27390 = ~n25666 & ~n27389;
  assign n27391 = ~n27385 & ~n27390;
  assign n27392 = ~n27388 & ~n27391;
  assign n27393 = ~n27384 & ~n27392;
  assign n27394 = n27377 & ~n27381;
  assign n27395 = ~n27377 & n27381;
  assign n27396 = ~n27394 & ~n27395;
  assign n27397 = ~n27385 & ~n27387;
  assign n27398 = n27385 & ~n27390;
  assign n27399 = ~n27397 & ~n27398;
  assign n27400 = ~n27396 & ~n27399;
  assign n27401 = ~n27393 & ~n27400;
  assign n27402 = ~pi310 & n27401;
  assign n27403 = ~n10908 & n27401;
  assign n27404 = n10908 & ~n27401;
  assign n27405 = pi310 & n27404;
  assign n27406 = ~n27403 & ~n27405;
  assign n27407 = ~n9815 & ~n27406;
  assign n27408 = ~n27402 & ~n27407;
  assign n27409 = ~n25679 & ~n27408;
  assign n27410 = n25678 & ~n27406;
  assign n27411 = n9815 & ~n25678;
  assign n27412 = n10908 & n27401;
  assign n27413 = n27411 & n27412;
  assign n27414 = ~n27410 & ~n27413;
  assign n27415 = ~n25670 & ~n27414;
  assign n27416 = ~n25678 & n27412;
  assign n27417 = ~n10908 & ~n27401;
  assign n27418 = n9815 & n27417;
  assign n27419 = ~n27416 & ~n27418;
  assign n27420 = pi310 & ~n27419;
  assign n27421 = pi310 & n10908;
  assign n27422 = ~n27401 & ~n27421;
  assign n27423 = ~n25678 & n27422;
  assign n27424 = n9815 & n25678;
  assign n27425 = n27412 & n27424;
  assign n27426 = ~n27423 & ~n27425;
  assign n27427 = ~n27420 & n27426;
  assign n27428 = n25670 & ~n27427;
  assign n27429 = ~n25678 & n27417;
  assign n27430 = n25684 & n27429;
  assign n27431 = ~n27428 & ~n27430;
  assign n27432 = ~n27415 & n27431;
  assign n27433 = ~n27409 & n27432;
  assign n27434 = ~n27179 & ~n27433;
  assign n27435 = n27179 & n27433;
  assign n27436 = ~n27434 & ~n27435;
  assign n27437 = pi308 & n9517;
  assign n27438 = n7044 & ~n25700;
  assign n27439 = pi309 & n27438;
  assign n27440 = ~n23305 & ~n23869;
  assign n27441 = ~n27439 & ~n27440;
  assign n27442 = ~n23858 & ~n27441;
  assign n27443 = n7874 & ~n23844;
  assign n27444 = ~n23305 & n27438;
  assign n27445 = ~n27443 & ~n27444;
  assign n27446 = pi309 & ~n27445;
  assign n27447 = ~n27442 & ~n27446;
  assign n27448 = ~n25689 & ~n27447;
  assign n27449 = n25689 & n27447;
  assign n27450 = n25409 & ~n27449;
  assign n27451 = ~n27448 & ~n27450;
  assign n27452 = n27437 & ~n27451;
  assign n27453 = ~n25409 & ~n27448;
  assign n27454 = ~n27449 & ~n27453;
  assign n27455 = ~n27437 & ~n27454;
  assign n27456 = ~n27452 & ~n27455;
  assign n27457 = ~n27436 & ~n27456;
  assign n27458 = ~n27179 & n27433;
  assign n27459 = n27179 & ~n27433;
  assign n27460 = ~n27458 & ~n27459;
  assign n27461 = ~n27437 & ~n27451;
  assign n27462 = n27437 & ~n27454;
  assign n27463 = ~n27461 & ~n27462;
  assign n27464 = ~n27460 & ~n27463;
  assign n27465 = ~n27457 & ~n27464;
  assign n27466 = ~n25692 & ~n25693;
  assign n27467 = n25692 & n25693;
  assign n27468 = ~n25728 & ~n27467;
  assign n27469 = ~n27466 & ~n27468;
  assign n27470 = n27465 & n27469;
  assign n27471 = ~n27465 & ~n27469;
  assign n27472 = ~n27470 & ~n27471;
  assign n27473 = pi307 & n7874;
  assign n27474 = ~n25740 & n25745;
  assign n27475 = ~n25741 & ~n27474;
  assign n27476 = n27473 & ~n27475;
  assign n27477 = ~n25741 & ~n25745;
  assign n27478 = ~n25740 & ~n27477;
  assign n27479 = ~n27473 & ~n27478;
  assign n27480 = ~n27476 & ~n27479;
  assign n27481 = ~n27472 & ~n27480;
  assign n27482 = n27465 & ~n27469;
  assign n27483 = ~n27465 & n27469;
  assign n27484 = ~n27482 & ~n27483;
  assign n27485 = ~n27473 & ~n27475;
  assign n27486 = n27473 & ~n27478;
  assign n27487 = ~n27485 & ~n27486;
  assign n27488 = ~n27484 & ~n27487;
  assign n27489 = ~n27481 & ~n27488;
  assign n27490 = ~pi306 & n27489;
  assign n27491 = ~n7044 & n27489;
  assign n27492 = n7044 & ~n27489;
  assign n27493 = pi306 & n27492;
  assign n27494 = ~n27491 & ~n27493;
  assign n27495 = ~n6777 & ~n27494;
  assign n27496 = ~n27490 & ~n27495;
  assign n27497 = ~n25766 & ~n27496;
  assign n27498 = n6777 & ~n25758;
  assign n27499 = n7044 & n27489;
  assign n27500 = n27498 & n27499;
  assign n27501 = n25758 & ~n27494;
  assign n27502 = ~n27500 & ~n27501;
  assign n27503 = n25750 & ~n27502;
  assign n27504 = ~n25758 & n27499;
  assign n27505 = ~n7044 & ~n27489;
  assign n27506 = n6777 & n27505;
  assign n27507 = ~n27504 & ~n27506;
  assign n27508 = pi306 & ~n27507;
  assign n27509 = n6777 & n25758;
  assign n27510 = n27499 & n27509;
  assign n27511 = pi306 & n7044;
  assign n27512 = ~n27489 & ~n27511;
  assign n27513 = ~n25758 & n27512;
  assign n27514 = ~n27510 & ~n27513;
  assign n27515 = ~n27508 & n27514;
  assign n27516 = ~n25750 & ~n27515;
  assign n27517 = ~n25758 & n27505;
  assign n27518 = n25764 & n27517;
  assign n27519 = ~n27516 & ~n27518;
  assign n27520 = ~n27503 & n27519;
  assign n27521 = ~n27497 & n27520;
  assign n27522 = ~n27178 & n27521;
  assign n27523 = n27178 & ~n27521;
  assign n27524 = ~n27522 & ~n27523;
  assign n27525 = pi304 & n5463;
  assign n27526 = n23385 & ~n23957;
  assign n27527 = n4086 & ~n25780;
  assign n27528 = pi305 & n27527;
  assign n27529 = ~n27526 & ~n27528;
  assign n27530 = ~n23946 & ~n27529;
  assign n27531 = n4772 & n23932;
  assign n27532 = n23385 & n27527;
  assign n27533 = ~n27531 & ~n27532;
  assign n27534 = pi305 & ~n27533;
  assign n27535 = ~n27530 & ~n27534;
  assign n27536 = n25769 & ~n27535;
  assign n27537 = ~n25769 & n27535;
  assign n27538 = n25397 & ~n27537;
  assign n27539 = ~n27536 & ~n27538;
  assign n27540 = n27525 & ~n27539;
  assign n27541 = ~n25397 & ~n27536;
  assign n27542 = ~n27537 & ~n27541;
  assign n27543 = ~n27525 & ~n27542;
  assign n27544 = ~n27540 & ~n27543;
  assign n27545 = ~n27524 & ~n27544;
  assign n27546 = ~n27178 & ~n27521;
  assign n27547 = n27178 & n27521;
  assign n27548 = ~n27546 & ~n27547;
  assign n27549 = ~n27525 & ~n27539;
  assign n27550 = n27525 & ~n27542;
  assign n27551 = ~n27549 & ~n27550;
  assign n27552 = ~n27548 & ~n27551;
  assign n27553 = ~n27545 & ~n27552;
  assign n27554 = ~n25773 & ~n25814;
  assign n27555 = n25773 & n25814;
  assign n27556 = ~n25808 & ~n27555;
  assign n27557 = ~n27554 & ~n27556;
  assign n27558 = n27553 & ~n27557;
  assign n27559 = ~n27553 & n27557;
  assign n27560 = ~n27558 & ~n27559;
  assign n27561 = pi303 & n4772;
  assign n27562 = n25825 & ~n25827;
  assign n27563 = ~n25826 & ~n27562;
  assign n27564 = n27561 & ~n27563;
  assign n27565 = ~n25825 & ~n25826;
  assign n27566 = ~n25827 & ~n27565;
  assign n27567 = ~n27561 & ~n27566;
  assign n27568 = ~n27564 & ~n27567;
  assign n27569 = ~n27560 & ~n27568;
  assign n27570 = n27553 & n27557;
  assign n27571 = ~n27553 & ~n27557;
  assign n27572 = ~n27570 & ~n27571;
  assign n27573 = ~n27561 & ~n27563;
  assign n27574 = n27561 & ~n27566;
  assign n27575 = ~n27573 & ~n27574;
  assign n27576 = ~n27572 & ~n27575;
  assign n27577 = ~n27569 & ~n27576;
  assign n27578 = ~pi302 & ~n27577;
  assign n27579 = ~n4086 & ~n27577;
  assign n27580 = n4086 & n27577;
  assign n27581 = pi302 & n27580;
  assign n27582 = ~n27579 & ~n27581;
  assign n27583 = ~n3552 & ~n27582;
  assign n27584 = ~n27578 & ~n27583;
  assign n27585 = ~n25842 & ~n27584;
  assign n27586 = ~n25838 & ~n27577;
  assign n27587 = n3552 & n27586;
  assign n27588 = ~n25835 & n27577;
  assign n27589 = ~n25830 & n27588;
  assign n27590 = n25835 & ~n27577;
  assign n27591 = n25830 & n27590;
  assign n27592 = ~n27589 & ~n27591;
  assign n27593 = pi302 & ~n27592;
  assign n27594 = ~n27587 & ~n27593;
  assign n27595 = n4086 & ~n27594;
  assign n27596 = ~n25835 & ~n27577;
  assign n27597 = ~n25830 & n27596;
  assign n27598 = n3552 & ~n25843;
  assign n27599 = pi302 & n27598;
  assign n27600 = ~n25842 & ~n27599;
  assign n27601 = n27577 & ~n27600;
  assign n27602 = ~n27597 & ~n27601;
  assign n27603 = ~n4086 & ~n27602;
  assign n27604 = n25835 & n27577;
  assign n27605 = ~pi302 & n25830;
  assign n27606 = n27604 & n27605;
  assign n27607 = ~n27603 & ~n27606;
  assign n27608 = ~n27595 & n27607;
  assign n27609 = ~n27585 & n27608;
  assign n27610 = ~n27177 & n27609;
  assign n27611 = n27177 & ~n27609;
  assign n27612 = ~n27610 & ~n27611;
  assign n27613 = pi300 & n3012;
  assign n27614 = n23456 & ~n24014;
  assign n27615 = n2183 & ~n25870;
  assign n27616 = pi301 & n27615;
  assign n27617 = ~n27614 & ~n27616;
  assign n27618 = ~n24003 & ~n27617;
  assign n27619 = n23456 & n27615;
  assign n27620 = ~n25871 & ~n27619;
  assign n27621 = pi301 & ~n27620;
  assign n27622 = ~n27618 & ~n27621;
  assign n27623 = n25846 & ~n27622;
  assign n27624 = ~n25846 & n27622;
  assign n27625 = n25380 & ~n27624;
  assign n27626 = ~n27623 & ~n27625;
  assign n27627 = n27613 & ~n27626;
  assign n27628 = ~n25380 & ~n27623;
  assign n27629 = ~n27624 & ~n27628;
  assign n27630 = ~n27613 & ~n27629;
  assign n27631 = ~n27627 & ~n27630;
  assign n27632 = ~n27612 & ~n27631;
  assign n27633 = ~n27177 & ~n27609;
  assign n27634 = n27177 & n27609;
  assign n27635 = ~n27633 & ~n27634;
  assign n27636 = ~n27613 & ~n27626;
  assign n27637 = n27613 & ~n27629;
  assign n27638 = ~n27636 & ~n27637;
  assign n27639 = ~n27635 & ~n27638;
  assign n27640 = ~n27632 & ~n27639;
  assign n27641 = n25850 & ~n25891;
  assign n27642 = ~n25850 & n25891;
  assign n27643 = ~n25882 & ~n27642;
  assign n27644 = ~n27641 & ~n27643;
  assign n27645 = n27640 & n27644;
  assign n27646 = ~n27640 & ~n27644;
  assign n27647 = ~n27645 & ~n27646;
  assign n27648 = pi299 & n2574;
  assign n27649 = n25902 & ~n25903;
  assign n27650 = ~n25904 & ~n27649;
  assign n27651 = n27648 & ~n27650;
  assign n27652 = ~n25902 & ~n25904;
  assign n27653 = ~n25903 & ~n27652;
  assign n27654 = ~n27648 & ~n27653;
  assign n27655 = ~n27651 & ~n27654;
  assign n27656 = ~n27647 & ~n27655;
  assign n27657 = n27640 & ~n27644;
  assign n27658 = ~n27640 & n27644;
  assign n27659 = ~n27657 & ~n27658;
  assign n27660 = ~n27648 & ~n27650;
  assign n27661 = n27648 & ~n27653;
  assign n27662 = ~n27660 & ~n27661;
  assign n27663 = ~n27659 & ~n27662;
  assign n27664 = ~n27656 & ~n27663;
  assign n27665 = ~pi298 & n27664;
  assign n27666 = ~n2183 & n27664;
  assign n27667 = n2183 & ~n27664;
  assign n27668 = pi298 & n27667;
  assign n27669 = ~n27666 & ~n27668;
  assign n27670 = ~n1840 & ~n27669;
  assign n27671 = ~n27665 & ~n27670;
  assign n27672 = ~n25913 & ~n27671;
  assign n27673 = n25912 & n27664;
  assign n27674 = n25907 & n27673;
  assign n27675 = ~n25912 & ~n27664;
  assign n27676 = ~n25907 & n27675;
  assign n27677 = ~n27674 & ~n27676;
  assign n27678 = pi298 & ~n27677;
  assign n27679 = ~n25921 & n27664;
  assign n27680 = n1840 & n27679;
  assign n27681 = ~n27678 & ~n27680;
  assign n27682 = n2183 & ~n27681;
  assign n27683 = n25912 & ~n27664;
  assign n27684 = ~pi298 & n25907;
  assign n27685 = n27683 & n27684;
  assign n27686 = ~n25912 & n27664;
  assign n27687 = ~n25907 & n27686;
  assign n27688 = n1840 & ~n25914;
  assign n27689 = pi298 & n27688;
  assign n27690 = ~n25913 & ~n27689;
  assign n27691 = ~n27664 & ~n27690;
  assign n27692 = ~n27687 & ~n27691;
  assign n27693 = ~n2183 & ~n27692;
  assign n27694 = ~n27685 & ~n27693;
  assign n27695 = ~n27682 & n27694;
  assign n27696 = ~n27672 & n27695;
  assign n27697 = pi297 & ~n6883;
  assign n27698 = n27696 & ~n27697;
  assign n27699 = pi297 & ~n27696;
  assign n27700 = n6886 & n27699;
  assign n27701 = ~n27698 & ~n27700;
  assign n27702 = ~n27176 & ~n27701;
  assign n27703 = ~n1840 & n27696;
  assign n27704 = pi297 & n1840;
  assign n27705 = ~n27696 & n27704;
  assign n27706 = ~n27703 & ~n27705;
  assign n27707 = n25923 & ~n27706;
  assign n27708 = n25367 & n27707;
  assign n27709 = n6897 & ~n27696;
  assign n27710 = ~n1533 & n25923;
  assign n27711 = n1840 & ~n27710;
  assign n27712 = n27696 & n27711;
  assign n27713 = ~n27709 & ~n27712;
  assign n27714 = pi297 & ~n27713;
  assign n27715 = ~n27696 & ~n27704;
  assign n27716 = ~n25923 & n27715;
  assign n27717 = ~n27714 & ~n27716;
  assign n27718 = ~n25367 & ~n27717;
  assign n27719 = ~n1840 & ~n27696;
  assign n27720 = n1840 & n27696;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = n1533 & ~n27721;
  assign n27723 = pi297 & n27722;
  assign n27724 = ~n25923 & n27723;
  assign n27725 = ~n27718 & ~n27724;
  assign n27726 = ~n27708 & n27725;
  assign n27727 = ~n27702 & n27726;
  assign n27728 = ~n25926 & ~n25927;
  assign n27729 = n25926 & n25927;
  assign n27730 = ~n25946 & ~n27729;
  assign n27731 = ~n27728 & ~n27730;
  assign n27732 = n27727 & ~n27731;
  assign n27733 = ~n27727 & n27731;
  assign n27734 = ~n27732 & ~n27733;
  assign n27735 = n1533 & ~n27734;
  assign n27736 = pi296 & n27735;
  assign n27737 = pi296 & n1533;
  assign n27738 = ~n27727 & ~n27731;
  assign n27739 = n27727 & n27731;
  assign n27740 = ~n27738 & ~n27739;
  assign n27741 = ~n27737 & ~n27740;
  assign n27742 = ~n27736 & ~n27741;
  assign n27743 = ~n24117 & n25962;
  assign n27744 = n25330 & n27743;
  assign n27745 = ~n25963 & ~n25977;
  assign n27746 = ~n27744 & ~n27745;
  assign n27747 = n27742 & ~n27746;
  assign n27748 = ~n27742 & n27746;
  assign n27749 = ~n27747 & ~n27748;
  assign n27750 = n25362 & ~n25957;
  assign n27751 = ~n25362 & n25957;
  assign n27752 = ~n1515 & ~n27751;
  assign n27753 = ~n27750 & ~n27752;
  assign n27754 = n1553 & ~n27753;
  assign n27755 = ~n1553 & ~n27750;
  assign n27756 = n1515 & n27755;
  assign n27757 = ~n27754 & ~n27756;
  assign n27758 = pi295 & ~n27757;
  assign n27759 = pi295 & n1553;
  assign n27760 = n25957 & ~n27759;
  assign n27761 = ~n25362 & n27760;
  assign n27762 = ~n27758 & ~n27761;
  assign n27763 = pi294 & n1515;
  assign n27764 = n27762 & ~n27763;
  assign n27765 = n1515 & ~n27762;
  assign n27766 = pi294 & n27765;
  assign n27767 = ~n27764 & ~n27766;
  assign n27768 = ~n27749 & ~n27767;
  assign n27769 = ~n27742 & ~n27746;
  assign n27770 = n27742 & n27746;
  assign n27771 = ~n27769 & ~n27770;
  assign n27772 = ~n27762 & ~n27763;
  assign n27773 = n1515 & n27762;
  assign n27774 = pi294 & n27773;
  assign n27775 = ~n27772 & ~n27774;
  assign n27776 = ~n27771 & ~n27775;
  assign n27777 = ~n27768 & ~n27776;
  assign n27778 = ~n27175 & n27777;
  assign n27779 = n27175 & ~n27777;
  assign n27780 = ~n27778 & ~n27779;
  assign n27781 = pi292 & ~n27780;
  assign n27782 = pi128 & n27781;
  assign n27783 = pi128 & pi292;
  assign n27784 = n27175 & n27777;
  assign n27785 = ~n27175 & ~n27777;
  assign n27786 = ~n27784 & ~n27785;
  assign n27787 = ~n27783 & ~n27786;
  assign n27788 = ~n27782 & ~n27787;
  assign n27789 = n1156 & n27127;
  assign n27790 = ~n1154 & ~n27789;
  assign n27791 = n1154 & n27127;
  assign n27792 = n1156 & n27791;
  assign n27793 = ~n27790 & ~n27792;
  assign n27794 = pi350 & ~n27793;
  assign n27795 = n25996 & ~n27048;
  assign n27796 = ~n25996 & n27048;
  assign n27797 = ~n27795 & ~n27796;
  assign n27798 = n26016 & n27052;
  assign n27799 = n26020 & ~n27075;
  assign n27800 = ~n26020 & n27075;
  assign n27801 = ~n27799 & ~n27800;
  assign n27802 = ~n27798 & ~n27801;
  assign n27803 = ~n27797 & n27802;
  assign n27804 = n25996 & n27048;
  assign n27805 = ~n25996 & ~n27048;
  assign n27806 = ~n27804 & ~n27805;
  assign n27807 = ~n26020 & ~n27075;
  assign n27808 = n26020 & n27075;
  assign n27809 = ~n27807 & ~n27808;
  assign n27810 = ~n27798 & ~n27809;
  assign n27811 = ~n27806 & n27810;
  assign n27812 = ~n26016 & ~n27052;
  assign n27813 = ~n27811 & ~n27812;
  assign n27814 = ~n27803 & n27813;
  assign n27815 = ~n1154 & n25992;
  assign n27816 = pi349 & n27815;
  assign n27817 = ~n25992 & ~n27115;
  assign n27818 = ~n27096 & ~n27111;
  assign n27819 = ~n27105 & n27818;
  assign n27820 = n27096 & ~n27112;
  assign n27821 = ~n27819 & ~n27820;
  assign n27822 = ~n27817 & ~n27821;
  assign n27823 = ~n27816 & ~n27822;
  assign n27824 = n27814 & n27823;
  assign n27825 = ~n27814 & ~n27823;
  assign n27826 = ~n27824 & ~n27825;
  assign n27827 = n27096 & ~n27111;
  assign n27828 = ~n27105 & ~n27827;
  assign n27829 = n1442 & n27828;
  assign n27830 = pi348 & n27829;
  assign n27831 = pi348 & n1442;
  assign n27832 = ~n27828 & ~n27831;
  assign n27833 = ~n27830 & ~n27832;
  assign n27834 = ~n26048 & n26950;
  assign n27835 = n26048 & ~n26950;
  assign n27836 = ~n27834 & ~n27835;
  assign n27837 = ~n26062 & n26954;
  assign n27838 = n26066 & ~n26972;
  assign n27839 = ~n26066 & n26972;
  assign n27840 = ~n27838 & ~n27839;
  assign n27841 = ~n27837 & ~n27840;
  assign n27842 = ~n27836 & n27841;
  assign n27843 = n26048 & n26950;
  assign n27844 = ~n26048 & ~n26950;
  assign n27845 = ~n27843 & ~n27844;
  assign n27846 = ~n26066 & ~n26972;
  assign n27847 = n26066 & n26972;
  assign n27848 = ~n27846 & ~n27847;
  assign n27849 = ~n27837 & ~n27848;
  assign n27850 = ~n27845 & n27849;
  assign n27851 = n26062 & ~n26954;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = ~n27842 & n27852;
  assign n27854 = ~n27000 & n27004;
  assign n27855 = n27000 & ~n27004;
  assign n27856 = n2887 & ~n27005;
  assign n27857 = ~n27006 & ~n27856;
  assign n27858 = n4596 & ~n27857;
  assign n27859 = pi342 & n27858;
  assign n27860 = ~n4596 & ~n27856;
  assign n27861 = pi342 & ~n27860;
  assign n27862 = ~n27006 & ~n27861;
  assign n27863 = ~n27859 & ~n27862;
  assign n27864 = n26993 & ~n27863;
  assign n27865 = ~n26993 & n27863;
  assign n27866 = ~n27864 & ~n27865;
  assign n27867 = ~n27855 & ~n27866;
  assign n27868 = ~n27854 & ~n27867;
  assign n27869 = n27853 & n27868;
  assign n27870 = ~n27853 & ~n27868;
  assign n27871 = ~n27869 & ~n27870;
  assign n27872 = pi341 & n5714;
  assign n27873 = ~n26087 & n26853;
  assign n27874 = n26087 & ~n26853;
  assign n27875 = ~n27873 & ~n27874;
  assign n27876 = ~n26101 & n26857;
  assign n27877 = n26105 & ~n26875;
  assign n27878 = ~n26105 & n26875;
  assign n27879 = ~n27877 & ~n27878;
  assign n27880 = ~n27876 & ~n27879;
  assign n27881 = ~n27875 & n27880;
  assign n27882 = n26087 & n26853;
  assign n27883 = ~n26087 & ~n26853;
  assign n27884 = ~n27882 & ~n27883;
  assign n27885 = ~n26105 & ~n26875;
  assign n27886 = n26105 & n26875;
  assign n27887 = ~n27885 & ~n27886;
  assign n27888 = ~n27876 & ~n27887;
  assign n27889 = ~n27884 & n27888;
  assign n27890 = n26101 & ~n26857;
  assign n27891 = ~n27889 & ~n27890;
  assign n27892 = ~n27881 & n27891;
  assign n27893 = ~n26903 & n26907;
  assign n27894 = n26903 & ~n26907;
  assign n27895 = n6556 & ~n26908;
  assign n27896 = ~n26909 & ~n27895;
  assign n27897 = n9205 & ~n27896;
  assign n27898 = pi336 & n27897;
  assign n27899 = ~n9205 & ~n27895;
  assign n27900 = pi336 & ~n27899;
  assign n27901 = ~n26909 & ~n27900;
  assign n27902 = ~n27898 & ~n27901;
  assign n27903 = n26896 & ~n27902;
  assign n27904 = ~n26896 & n27902;
  assign n27905 = ~n27903 & ~n27904;
  assign n27906 = ~n27894 & ~n27905;
  assign n27907 = ~n27893 & ~n27906;
  assign n27908 = n27892 & n27907;
  assign n27909 = ~n27892 & ~n27907;
  assign n27910 = ~n27908 & ~n27909;
  assign n27911 = pi335 & n11366;
  assign n27912 = ~n26122 & ~n26126;
  assign n27913 = n26122 & n26126;
  assign n27914 = ~n26110 & n26768;
  assign n27915 = n26110 & ~n26768;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = n19539 & ~n27916;
  assign n27918 = pi328 & n27917;
  assign n27919 = ~n26110 & ~n26768;
  assign n27920 = n26110 & n26768;
  assign n27921 = ~n27919 & ~n27920;
  assign n27922 = ~n26774 & ~n27921;
  assign n27923 = ~n27918 & ~n27922;
  assign n27924 = ~n27913 & ~n27923;
  assign n27925 = ~n27912 & ~n27924;
  assign n27926 = ~n26804 & n26808;
  assign n27927 = ~n26789 & ~n26815;
  assign n27928 = n26789 & n26815;
  assign n27929 = ~n27927 & ~n27928;
  assign n27930 = n26804 & ~n26808;
  assign n27931 = ~n27929 & ~n27930;
  assign n27932 = ~n27926 & ~n27931;
  assign n27933 = n27925 & n27932;
  assign n27934 = ~n27925 & ~n27932;
  assign n27935 = ~n27933 & ~n27934;
  assign n27936 = ~n26789 & n26810;
  assign n27937 = n26789 & ~n26810;
  assign n27938 = ~n13762 & ~n27937;
  assign n27939 = ~n27936 & ~n27938;
  assign n27940 = n18461 & ~n27939;
  assign n27941 = ~n18461 & ~n27936;
  assign n27942 = n13762 & n27941;
  assign n27943 = ~n27940 & ~n27942;
  assign n27944 = pi330 & ~n27943;
  assign n27945 = pi330 & n18461;
  assign n27946 = n26789 & ~n27945;
  assign n27947 = ~n26810 & n27946;
  assign n27948 = ~n27944 & ~n27947;
  assign n27949 = ~n26130 & ~n26742;
  assign n27950 = n26130 & n26742;
  assign n27951 = ~n27949 & ~n27950;
  assign n27952 = n26150 & n26746;
  assign n27953 = ~n26727 & n26747;
  assign n27954 = n26727 & ~n26747;
  assign n27955 = ~n27953 & ~n27954;
  assign n27956 = ~n27952 & ~n27955;
  assign n27957 = ~n27951 & n27956;
  assign n27958 = ~n26130 & n26742;
  assign n27959 = n26130 & ~n26742;
  assign n27960 = ~n27958 & ~n27959;
  assign n27961 = n26727 & n26747;
  assign n27962 = ~n26727 & ~n26747;
  assign n27963 = ~n27961 & ~n27962;
  assign n27964 = ~n27952 & ~n27963;
  assign n27965 = ~n27960 & n27964;
  assign n27966 = ~n26150 & ~n26746;
  assign n27967 = ~n27965 & ~n27966;
  assign n27968 = ~n27957 & n27967;
  assign n27969 = n19539 & ~n27920;
  assign n27970 = pi328 & n27969;
  assign n27971 = ~n27919 & ~n27970;
  assign n27972 = n27968 & ~n27971;
  assign n27973 = ~n27968 & n27971;
  assign n27974 = ~n27972 & ~n27973;
  assign n27975 = pi327 & n19970;
  assign n27976 = n26703 & ~n26742;
  assign n27977 = ~n26155 & ~n26702;
  assign n27978 = n26155 & ~n26701;
  assign n27979 = ~n26698 & n27978;
  assign n27980 = ~n27977 & ~n27979;
  assign n27981 = ~n26707 & ~n27980;
  assign n27982 = n26155 & ~n26702;
  assign n27983 = ~n26155 & ~n26701;
  assign n27984 = ~n26698 & n27983;
  assign n27985 = ~n27982 & ~n27984;
  assign n27986 = n26706 & ~n27985;
  assign n27987 = pi324 & n27986;
  assign n27988 = ~n27981 & ~n27987;
  assign n27989 = n26163 & ~n27988;
  assign n27990 = ~n26163 & n27988;
  assign n27991 = ~n27989 & ~n27990;
  assign n27992 = ~n26703 & n26742;
  assign n27993 = ~n27991 & ~n27992;
  assign n27994 = ~n27976 & ~n27993;
  assign n27995 = ~n26130 & n26747;
  assign n27996 = n26130 & ~n26747;
  assign n27997 = ~n26754 & ~n27996;
  assign n27998 = ~n27995 & ~n27997;
  assign n27999 = n27994 & ~n27998;
  assign n28000 = ~n27994 & n27998;
  assign n28001 = ~n27999 & ~n28000;
  assign n28002 = pi324 & n26175;
  assign n28003 = ~n26155 & ~n26698;
  assign n28004 = ~n26701 & ~n28003;
  assign n28005 = ~n28002 & ~n28004;
  assign n28006 = n28002 & n28004;
  assign n28007 = ~n28005 & ~n28006;
  assign n28008 = ~n24906 & ~n26694;
  assign n28009 = n24906 & ~n26690;
  assign n28010 = ~n28008 & ~n28009;
  assign n28011 = pi323 & n28010;
  assign n28012 = ~n26643 & n26648;
  assign n28013 = n26643 & ~n26648;
  assign n28014 = ~n26636 & ~n28013;
  assign n28015 = ~n28012 & ~n28014;
  assign n28016 = n26647 & n26661;
  assign n28017 = n26648 & ~n26678;
  assign n28018 = ~n26646 & ~n26648;
  assign n28019 = ~n28017 & ~n28018;
  assign n28020 = ~n26647 & ~n26661;
  assign n28021 = ~n28019 & ~n28020;
  assign n28022 = ~n28016 & ~n28021;
  assign n28023 = n28015 & ~n28022;
  assign n28024 = ~n28015 & n28022;
  assign n28025 = ~n28023 & ~n28024;
  assign n28026 = n26277 & ~n26286;
  assign n28027 = ~n26282 & n28026;
  assign n28028 = ~n26277 & ~n26289;
  assign n28029 = ~n28027 & ~n28028;
  assign n28030 = ~n26183 & ~n28029;
  assign n28031 = ~n26277 & ~n26286;
  assign n28032 = ~n26282 & n28031;
  assign n28033 = n26277 & ~n26289;
  assign n28034 = ~n28032 & ~n28033;
  assign n28035 = pi281 & ~n28034;
  assign n28036 = pi133 & n28035;
  assign n28037 = ~n28030 & ~n28036;
  assign n28038 = ~n26306 & ~n28037;
  assign n28039 = pi133 & pi282;
  assign n28040 = pi132 & pi283;
  assign n28041 = pi131 & pi284;
  assign n28042 = ~n26196 & n26197;
  assign n28043 = pi129 & pi286;
  assign n28044 = pi287 & ~n28043;
  assign n28045 = pi128 & n28044;
  assign n28046 = pi128 & pi287;
  assign n28047 = pi286 & ~n28046;
  assign n28048 = pi129 & n28047;
  assign n28049 = ~n28045 & ~n28048;
  assign n28050 = ~pi285 & ~n28049;
  assign n28051 = ~pi130 & ~n28049;
  assign n28052 = pi285 & n28049;
  assign n28053 = pi130 & n28052;
  assign n28054 = ~n28051 & ~n28053;
  assign n28055 = ~pi129 & ~n28054;
  assign n28056 = ~n28050 & ~n28055;
  assign n28057 = ~n28042 & ~n28056;
  assign n28058 = n26196 & n26197;
  assign n28059 = ~n26196 & ~n26197;
  assign n28060 = ~n28058 & ~n28059;
  assign n28061 = pi129 & ~n28060;
  assign n28062 = pi285 & n28042;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = ~n28049 & ~n28063;
  assign n28065 = pi285 & n26196;
  assign n28066 = ~n26197 & n28049;
  assign n28067 = n28065 & n28066;
  assign n28068 = ~n28064 & ~n28067;
  assign n28069 = pi130 & ~n28068;
  assign n28070 = ~n26197 & ~n28049;
  assign n28071 = n26196 & n28070;
  assign n28072 = n26196 & ~n26197;
  assign n28073 = pi285 & ~n28072;
  assign n28074 = pi129 & n28073;
  assign n28075 = ~n28042 & ~n28074;
  assign n28076 = n28049 & ~n28075;
  assign n28077 = ~n28071 & ~n28076;
  assign n28078 = ~pi130 & ~n28077;
  assign n28079 = n26197 & n28049;
  assign n28080 = ~pi285 & ~n26196;
  assign n28081 = n28079 & n28080;
  assign n28082 = ~n28078 & ~n28081;
  assign n28083 = ~n28069 & n28082;
  assign n28084 = ~n28057 & n28083;
  assign n28085 = ~n28041 & n28084;
  assign n28086 = n28041 & ~n28084;
  assign n28087 = ~n28085 & ~n28086;
  assign n28088 = n26209 & ~n26229;
  assign n28089 = ~n26209 & n26229;
  assign n28090 = ~n26212 & ~n28089;
  assign n28091 = ~n28088 & ~n28090;
  assign n28092 = ~n28087 & ~n28091;
  assign n28093 = ~n28041 & ~n28084;
  assign n28094 = n28041 & n28084;
  assign n28095 = ~n28093 & ~n28094;
  assign n28096 = ~n26206 & ~n28088;
  assign n28097 = ~n28089 & ~n28096;
  assign n28098 = ~n28095 & ~n28097;
  assign n28099 = ~n28092 & ~n28098;
  assign n28100 = ~n28040 & n28099;
  assign n28101 = n28040 & ~n28099;
  assign n28102 = ~n28100 & ~n28101;
  assign n28103 = n26235 & ~n26261;
  assign n28104 = ~n26235 & n26261;
  assign n28105 = ~n26238 & ~n28104;
  assign n28106 = ~n28103 & ~n28105;
  assign n28107 = ~n28102 & ~n28106;
  assign n28108 = ~n28040 & ~n28099;
  assign n28109 = n28040 & n28099;
  assign n28110 = ~n28108 & ~n28109;
  assign n28111 = ~n26232 & ~n28103;
  assign n28112 = ~n28104 & ~n28111;
  assign n28113 = ~n28110 & ~n28112;
  assign n28114 = ~n28107 & ~n28113;
  assign n28115 = ~n28039 & ~n28114;
  assign n28116 = n28039 & n28114;
  assign n28117 = ~n28115 & ~n28116;
  assign n28118 = ~n26266 & ~n26272;
  assign n28119 = ~n26269 & ~n28118;
  assign n28120 = ~n28117 & ~n28119;
  assign n28121 = ~n28039 & n28114;
  assign n28122 = n28039 & ~n28114;
  assign n28123 = ~n28121 & ~n28122;
  assign n28124 = ~n28118 & ~n28123;
  assign n28125 = ~n26269 & n28124;
  assign n28126 = ~n28120 & ~n28125;
  assign n28127 = ~n26289 & ~n26293;
  assign n28128 = ~n26294 & ~n28127;
  assign n28129 = n28126 & ~n28128;
  assign n28130 = ~n26286 & ~n26294;
  assign n28131 = ~n26282 & n28130;
  assign n28132 = ~n26293 & ~n28131;
  assign n28133 = ~n28126 & ~n28132;
  assign n28134 = ~n28129 & ~n28133;
  assign n28135 = ~pi134 & n28134;
  assign n28136 = ~pi281 & n28134;
  assign n28137 = pi281 & ~n28134;
  assign n28138 = pi134 & n28137;
  assign n28139 = ~n28136 & ~n28138;
  assign n28140 = ~pi280 & ~n28139;
  assign n28141 = ~n28135 & ~n28140;
  assign n28142 = ~n28038 & ~n28141;
  assign n28143 = ~n26306 & n28134;
  assign n28144 = ~n28037 & n28143;
  assign n28145 = n26306 & ~n28134;
  assign n28146 = n28037 & n28145;
  assign n28147 = ~n28144 & ~n28146;
  assign n28148 = pi134 & ~n28147;
  assign n28149 = ~n26306 & n28037;
  assign n28150 = n26306 & ~n28037;
  assign n28151 = ~n28149 & ~n28150;
  assign n28152 = n28134 & ~n28151;
  assign n28153 = pi280 & n28152;
  assign n28154 = ~n28148 & ~n28153;
  assign n28155 = pi281 & ~n28154;
  assign n28156 = ~pi134 & ~n28037;
  assign n28157 = ~n26306 & ~n28134;
  assign n28158 = n28156 & n28157;
  assign n28159 = n26306 & n28134;
  assign n28160 = n28037 & n28159;
  assign n28161 = n26306 & n28037;
  assign n28162 = pi280 & ~n28161;
  assign n28163 = pi134 & n28162;
  assign n28164 = ~n28038 & ~n28163;
  assign n28165 = ~n28134 & ~n28164;
  assign n28166 = ~n28160 & ~n28165;
  assign n28167 = ~pi281 & ~n28166;
  assign n28168 = ~n28158 & ~n28167;
  assign n28169 = ~n28155 & n28168;
  assign n28170 = ~n28142 & n28169;
  assign n28171 = ~n26309 & ~n26310;
  assign n28172 = n26309 & n26310;
  assign n28173 = ~n26315 & ~n28172;
  assign n28174 = ~n28171 & ~n28173;
  assign n28175 = ~n28170 & n28174;
  assign n28176 = n28170 & ~n28174;
  assign n28177 = ~n28175 & ~n28176;
  assign n28178 = pi136 & pi279;
  assign n28179 = pi135 & pi280;
  assign n28180 = n28178 & n28179;
  assign n28181 = ~n28178 & ~n28179;
  assign n28182 = ~n28180 & ~n28181;
  assign n28183 = ~n28177 & ~n28182;
  assign n28184 = n28170 & n28174;
  assign n28185 = ~n28170 & ~n28174;
  assign n28186 = ~n28184 & ~n28185;
  assign n28187 = pi279 & ~n28179;
  assign n28188 = pi136 & n28187;
  assign n28189 = pi280 & ~n28178;
  assign n28190 = pi135 & n28189;
  assign n28191 = ~n28188 & ~n28190;
  assign n28192 = ~n28186 & ~n28191;
  assign n28193 = ~n28183 & ~n28192;
  assign n28194 = pi278 & n26326;
  assign n28195 = ~pi278 & ~n26326;
  assign n28196 = pi277 & ~n28195;
  assign n28197 = ~n24506 & n28196;
  assign n28198 = ~n28194 & ~n28197;
  assign n28199 = pi136 & ~n28198;
  assign n28200 = pi136 & n28196;
  assign n28201 = ~n24506 & ~n26345;
  assign n28202 = ~n28200 & ~n28201;
  assign n28203 = n26334 & ~n28202;
  assign n28204 = ~n28199 & ~n28203;
  assign n28205 = n28193 & n28204;
  assign n28206 = ~n28193 & ~n28204;
  assign n28207 = ~n28205 & ~n28206;
  assign n28208 = pi137 & pi278;
  assign n28209 = ~pi277 & ~pi278;
  assign n28210 = pi136 & ~n28209;
  assign n28211 = n26326 & ~n28210;
  assign n28212 = ~pi277 & pi278;
  assign n28213 = pi136 & ~n26326;
  assign n28214 = n28212 & n28213;
  assign n28215 = ~n28211 & ~n28214;
  assign n28216 = ~n26335 & ~n28215;
  assign n28217 = ~pi278 & n26326;
  assign n28218 = ~n26328 & ~n28217;
  assign n28219 = n24506 & ~n28218;
  assign n28220 = ~n26334 & n28219;
  assign n28221 = ~n28194 & ~n28195;
  assign n28222 = pi277 & ~n28221;
  assign n28223 = pi136 & n28222;
  assign n28224 = ~n24506 & n28223;
  assign n28225 = pi277 & ~pi278;
  assign n28226 = ~n26326 & n28225;
  assign n28227 = ~pi277 & n24506;
  assign n28228 = pi278 & ~n28227;
  assign n28229 = n26326 & n28228;
  assign n28230 = ~n28226 & ~n28229;
  assign n28231 = pi136 & ~n28230;
  assign n28232 = ~n24506 & n26345;
  assign n28233 = ~n28231 & ~n28232;
  assign n28234 = n26334 & ~n28233;
  assign n28235 = ~n28224 & ~n28234;
  assign n28236 = ~n28220 & n28235;
  assign n28237 = ~n28216 & n28236;
  assign n28238 = ~n26356 & ~n28237;
  assign n28239 = n26356 & n28237;
  assign n28240 = n26330 & ~n28239;
  assign n28241 = ~n28238 & ~n28240;
  assign n28242 = n28208 & ~n28241;
  assign n28243 = ~n26330 & ~n28238;
  assign n28244 = ~n28239 & ~n28243;
  assign n28245 = ~n28208 & ~n28244;
  assign n28246 = ~n28242 & ~n28245;
  assign n28247 = ~n28207 & ~n28246;
  assign n28248 = n28193 & ~n28204;
  assign n28249 = ~n28193 & n28204;
  assign n28250 = ~n28248 & ~n28249;
  assign n28251 = ~n28208 & ~n28241;
  assign n28252 = n28208 & ~n28244;
  assign n28253 = ~n28251 & ~n28252;
  assign n28254 = ~n28250 & ~n28253;
  assign n28255 = ~n28247 & ~n28254;
  assign n28256 = ~n26360 & ~n26371;
  assign n28257 = n26360 & n26371;
  assign n28258 = ~n26365 & ~n28257;
  assign n28259 = ~n28256 & ~n28258;
  assign n28260 = ~n28255 & n28259;
  assign n28261 = n28255 & ~n28259;
  assign n28262 = ~n28260 & ~n28261;
  assign n28263 = pi139 & pi276;
  assign n28264 = pi138 & pi277;
  assign n28265 = n28263 & n28264;
  assign n28266 = ~n28263 & ~n28264;
  assign n28267 = ~n28265 & ~n28266;
  assign n28268 = ~n28262 & ~n28267;
  assign n28269 = n28255 & n28259;
  assign n28270 = ~n28255 & ~n28259;
  assign n28271 = ~n28269 & ~n28270;
  assign n28272 = pi276 & ~n28264;
  assign n28273 = pi139 & n28272;
  assign n28274 = pi277 & ~n28263;
  assign n28275 = pi138 & n28274;
  assign n28276 = ~n28273 & ~n28275;
  assign n28277 = ~n28271 & ~n28276;
  assign n28278 = ~n28268 & ~n28277;
  assign n28279 = ~n26389 & ~n26396;
  assign n28280 = ~n26384 & n28279;
  assign n28281 = ~n26397 & ~n28280;
  assign n28282 = n28278 & n28281;
  assign n28283 = ~n28278 & ~n28281;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = pi140 & pi275;
  assign n28286 = ~n26376 & ~n26389;
  assign n28287 = ~n26384 & n28286;
  assign n28288 = n26376 & ~n26392;
  assign n28289 = ~n28287 & ~n28288;
  assign n28290 = ~n26181 & ~n28289;
  assign n28291 = n26376 & ~n26389;
  assign n28292 = ~n26384 & n28291;
  assign n28293 = ~n26376 & ~n26392;
  assign n28294 = ~n28292 & ~n28293;
  assign n28295 = pi275 & ~n28294;
  assign n28296 = pi139 & n28295;
  assign n28297 = ~n28290 & ~n28296;
  assign n28298 = n26408 & n28297;
  assign n28299 = ~n26408 & ~n28297;
  assign n28300 = n26385 & ~n28299;
  assign n28301 = ~n28298 & ~n28300;
  assign n28302 = n28285 & ~n28301;
  assign n28303 = ~n26385 & ~n28298;
  assign n28304 = ~n28299 & ~n28303;
  assign n28305 = ~n28285 & ~n28304;
  assign n28306 = ~n28302 & ~n28305;
  assign n28307 = ~n28284 & ~n28306;
  assign n28308 = n28278 & ~n28281;
  assign n28309 = ~n28278 & n28281;
  assign n28310 = ~n28308 & ~n28309;
  assign n28311 = ~n28285 & ~n28301;
  assign n28312 = n28285 & ~n28304;
  assign n28313 = ~n28311 & ~n28312;
  assign n28314 = ~n28310 & ~n28313;
  assign n28315 = ~n28307 & ~n28314;
  assign n28316 = ~n26412 & ~n26423;
  assign n28317 = n26412 & n26423;
  assign n28318 = ~n26417 & ~n28317;
  assign n28319 = ~n28316 & ~n28318;
  assign n28320 = ~n28315 & n28319;
  assign n28321 = n28315 & ~n28319;
  assign n28322 = ~n28320 & ~n28321;
  assign n28323 = pi142 & pi273;
  assign n28324 = pi141 & pi274;
  assign n28325 = n28323 & n28324;
  assign n28326 = ~n28323 & ~n28324;
  assign n28327 = ~n28325 & ~n28326;
  assign n28328 = ~n28322 & ~n28327;
  assign n28329 = n28315 & n28319;
  assign n28330 = ~n28315 & ~n28319;
  assign n28331 = ~n28329 & ~n28330;
  assign n28332 = pi273 & ~n28324;
  assign n28333 = pi142 & n28332;
  assign n28334 = pi274 & ~n28323;
  assign n28335 = pi141 & n28334;
  assign n28336 = ~n28333 & ~n28335;
  assign n28337 = ~n28331 & ~n28336;
  assign n28338 = ~n28328 & ~n28337;
  assign n28339 = ~n26441 & ~n26448;
  assign n28340 = ~n26436 & n28339;
  assign n28341 = ~n26449 & ~n28340;
  assign n28342 = n28338 & ~n28341;
  assign n28343 = ~n28338 & n28341;
  assign n28344 = ~n28342 & ~n28343;
  assign n28345 = pi143 & pi272;
  assign n28346 = ~n26428 & ~n26441;
  assign n28347 = ~n26436 & n28346;
  assign n28348 = n26428 & ~n26444;
  assign n28349 = ~n28347 & ~n28348;
  assign n28350 = ~n26180 & ~n28349;
  assign n28351 = n26428 & ~n26441;
  assign n28352 = ~n26436 & n28351;
  assign n28353 = ~n26428 & ~n26444;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = pi272 & ~n28354;
  assign n28356 = pi142 & n28355;
  assign n28357 = ~n28350 & ~n28356;
  assign n28358 = n26460 & n28357;
  assign n28359 = ~n26460 & ~n28357;
  assign n28360 = n26437 & ~n28359;
  assign n28361 = ~n28358 & ~n28360;
  assign n28362 = n28345 & ~n28361;
  assign n28363 = ~n26437 & ~n28358;
  assign n28364 = ~n28359 & ~n28363;
  assign n28365 = ~n28345 & ~n28364;
  assign n28366 = ~n28362 & ~n28365;
  assign n28367 = ~n28344 & ~n28366;
  assign n28368 = n28338 & n28341;
  assign n28369 = ~n28338 & ~n28341;
  assign n28370 = ~n28368 & ~n28369;
  assign n28371 = ~n28345 & ~n28361;
  assign n28372 = n28345 & ~n28364;
  assign n28373 = ~n28371 & ~n28372;
  assign n28374 = ~n28370 & ~n28373;
  assign n28375 = ~n28367 & ~n28374;
  assign n28376 = n26464 & ~n26475;
  assign n28377 = ~n26464 & n26475;
  assign n28378 = ~n26466 & ~n28377;
  assign n28379 = ~n28376 & ~n28378;
  assign n28380 = ~n28375 & n28379;
  assign n28381 = n28375 & ~n28379;
  assign n28382 = ~n28380 & ~n28381;
  assign n28383 = pi145 & pi270;
  assign n28384 = pi144 & pi271;
  assign n28385 = n28383 & n28384;
  assign n28386 = ~n28383 & ~n28384;
  assign n28387 = ~n28385 & ~n28386;
  assign n28388 = ~n28382 & ~n28387;
  assign n28389 = n28375 & n28379;
  assign n28390 = ~n28375 & ~n28379;
  assign n28391 = ~n28389 & ~n28390;
  assign n28392 = pi270 & ~n28384;
  assign n28393 = pi145 & n28392;
  assign n28394 = pi271 & ~n28383;
  assign n28395 = pi144 & n28394;
  assign n28396 = ~n28393 & ~n28395;
  assign n28397 = ~n28391 & ~n28396;
  assign n28398 = ~n28388 & ~n28397;
  assign n28399 = ~n26496 & ~n26500;
  assign n28400 = ~n26501 & ~n28399;
  assign n28401 = n28398 & ~n28400;
  assign n28402 = ~n28398 & n28400;
  assign n28403 = ~n28401 & ~n28402;
  assign n28404 = pi146 & pi269;
  assign n28405 = ~n26480 & ~n26493;
  assign n28406 = ~n26489 & n28405;
  assign n28407 = n26480 & ~n26496;
  assign n28408 = ~n28406 & ~n28407;
  assign n28409 = ~n26179 & ~n28408;
  assign n28410 = n26480 & ~n26493;
  assign n28411 = ~n26489 & n28410;
  assign n28412 = ~n26480 & ~n26496;
  assign n28413 = ~n28411 & ~n28412;
  assign n28414 = pi269 & ~n28413;
  assign n28415 = pi145 & n28414;
  assign n28416 = ~n28409 & ~n28415;
  assign n28417 = n26512 & n28416;
  assign n28418 = ~n26512 & ~n28416;
  assign n28419 = n26490 & ~n28418;
  assign n28420 = ~n28417 & ~n28419;
  assign n28421 = n28404 & ~n28420;
  assign n28422 = ~n26490 & ~n28417;
  assign n28423 = ~n28418 & ~n28422;
  assign n28424 = ~n28404 & ~n28423;
  assign n28425 = ~n28421 & ~n28424;
  assign n28426 = ~n28403 & ~n28425;
  assign n28427 = n28398 & n28400;
  assign n28428 = ~n28398 & ~n28400;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 = ~n28404 & ~n28420;
  assign n28431 = n28404 & ~n28423;
  assign n28432 = ~n28430 & ~n28431;
  assign n28433 = ~n28429 & ~n28432;
  assign n28434 = ~n28426 & ~n28433;
  assign n28435 = n26516 & ~n26527;
  assign n28436 = ~n26516 & n26527;
  assign n28437 = ~n26518 & ~n28436;
  assign n28438 = ~n28435 & ~n28437;
  assign n28439 = ~n28434 & n28438;
  assign n28440 = n28434 & ~n28438;
  assign n28441 = ~n28439 & ~n28440;
  assign n28442 = pi148 & pi267;
  assign n28443 = pi147 & pi268;
  assign n28444 = n28442 & n28443;
  assign n28445 = ~n28442 & ~n28443;
  assign n28446 = ~n28444 & ~n28445;
  assign n28447 = ~n28441 & ~n28446;
  assign n28448 = n28434 & n28438;
  assign n28449 = ~n28434 & ~n28438;
  assign n28450 = ~n28448 & ~n28449;
  assign n28451 = pi267 & ~n28443;
  assign n28452 = pi148 & n28451;
  assign n28453 = pi268 & ~n28442;
  assign n28454 = pi147 & n28453;
  assign n28455 = ~n28452 & ~n28454;
  assign n28456 = ~n28450 & ~n28455;
  assign n28457 = ~n28447 & ~n28456;
  assign n28458 = ~n26548 & ~n26552;
  assign n28459 = ~n26553 & ~n28458;
  assign n28460 = n28457 & n28459;
  assign n28461 = ~n28457 & ~n28459;
  assign n28462 = ~n28460 & ~n28461;
  assign n28463 = pi149 & pi266;
  assign n28464 = n26532 & ~n26545;
  assign n28465 = ~n26541 & n28464;
  assign n28466 = ~n26532 & ~n26548;
  assign n28467 = ~n28465 & ~n28466;
  assign n28468 = ~n26178 & ~n28467;
  assign n28469 = ~n26532 & ~n26545;
  assign n28470 = ~n26541 & n28469;
  assign n28471 = n26532 & ~n26548;
  assign n28472 = ~n28470 & ~n28471;
  assign n28473 = pi266 & ~n28472;
  assign n28474 = pi148 & n28473;
  assign n28475 = ~n28468 & ~n28474;
  assign n28476 = ~n26564 & ~n28475;
  assign n28477 = n26564 & n28475;
  assign n28478 = n26542 & ~n28477;
  assign n28479 = ~n28476 & ~n28478;
  assign n28480 = n28463 & ~n28479;
  assign n28481 = ~n26542 & ~n28476;
  assign n28482 = ~n28477 & ~n28481;
  assign n28483 = ~n28463 & ~n28482;
  assign n28484 = ~n28480 & ~n28483;
  assign n28485 = ~n28462 & ~n28484;
  assign n28486 = n28457 & ~n28459;
  assign n28487 = ~n28457 & n28459;
  assign n28488 = ~n28486 & ~n28487;
  assign n28489 = ~n28463 & ~n28479;
  assign n28490 = n28463 & ~n28482;
  assign n28491 = ~n28489 & ~n28490;
  assign n28492 = ~n28488 & ~n28491;
  assign n28493 = ~n28485 & ~n28492;
  assign n28494 = ~n26567 & ~n26568;
  assign n28495 = n26567 & n26568;
  assign n28496 = ~n26573 & ~n28495;
  assign n28497 = ~n28494 & ~n28496;
  assign n28498 = ~n28493 & n28497;
  assign n28499 = n28493 & ~n28497;
  assign n28500 = ~n28498 & ~n28499;
  assign n28501 = pi151 & pi264;
  assign n28502 = pi150 & pi265;
  assign n28503 = n28501 & n28502;
  assign n28504 = ~n28501 & ~n28502;
  assign n28505 = ~n28503 & ~n28504;
  assign n28506 = ~n28500 & ~n28505;
  assign n28507 = n28493 & n28497;
  assign n28508 = ~n28493 & ~n28497;
  assign n28509 = ~n28507 & ~n28508;
  assign n28510 = pi264 & ~n28502;
  assign n28511 = pi151 & n28510;
  assign n28512 = pi265 & ~n28501;
  assign n28513 = pi150 & n28512;
  assign n28514 = ~n28511 & ~n28513;
  assign n28515 = ~n28509 & ~n28514;
  assign n28516 = ~n28506 & ~n28515;
  assign n28517 = ~n26600 & ~n26604;
  assign n28518 = ~n26605 & ~n28517;
  assign n28519 = n28516 & n28518;
  assign n28520 = ~n28516 & ~n28518;
  assign n28521 = ~n28519 & ~n28520;
  assign n28522 = pi152 & pi263;
  assign n28523 = n26584 & ~n26597;
  assign n28524 = ~n26593 & n28523;
  assign n28525 = ~n26584 & ~n26600;
  assign n28526 = ~n28524 & ~n28525;
  assign n28527 = ~n26177 & ~n28526;
  assign n28528 = ~n26584 & ~n26597;
  assign n28529 = ~n26593 & n28528;
  assign n28530 = n26584 & ~n26600;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = pi263 & ~n28531;
  assign n28533 = pi151 & n28532;
  assign n28534 = ~n28527 & ~n28533;
  assign n28535 = ~n26616 & ~n28534;
  assign n28536 = n26616 & n28534;
  assign n28537 = n26594 & ~n28536;
  assign n28538 = ~n28535 & ~n28537;
  assign n28539 = n28522 & ~n28538;
  assign n28540 = ~n26594 & ~n28535;
  assign n28541 = ~n28536 & ~n28540;
  assign n28542 = ~n28522 & ~n28541;
  assign n28543 = ~n28539 & ~n28542;
  assign n28544 = ~n28521 & ~n28543;
  assign n28545 = n28516 & ~n28518;
  assign n28546 = ~n28516 & n28518;
  assign n28547 = ~n28545 & ~n28546;
  assign n28548 = ~n28522 & ~n28538;
  assign n28549 = n28522 & ~n28541;
  assign n28550 = ~n28548 & ~n28549;
  assign n28551 = ~n28547 & ~n28550;
  assign n28552 = ~n28544 & ~n28551;
  assign n28553 = ~n26620 & ~n26631;
  assign n28554 = n26620 & n26631;
  assign n28555 = ~n26625 & ~n28554;
  assign n28556 = ~n28553 & ~n28555;
  assign n28557 = n28552 & n28556;
  assign n28558 = ~n28552 & ~n28556;
  assign n28559 = ~n28557 & ~n28558;
  assign n28560 = pi262 & ~n28559;
  assign n28561 = pi153 & n28560;
  assign n28562 = pi153 & pi262;
  assign n28563 = ~n28552 & n28556;
  assign n28564 = n28552 & ~n28556;
  assign n28565 = ~n28563 & ~n28564;
  assign n28566 = ~n28562 & ~n28565;
  assign n28567 = ~n28561 & ~n28566;
  assign n28568 = pi261 & ~n28567;
  assign n28569 = pi154 & n28568;
  assign n28570 = pi154 & pi261;
  assign n28571 = ~n28566 & ~n28570;
  assign n28572 = ~n28561 & n28571;
  assign n28573 = ~n28569 & ~n28572;
  assign n28574 = pi260 & ~n28573;
  assign n28575 = pi155 & n28574;
  assign n28576 = pi155 & pi260;
  assign n28577 = ~n28572 & ~n28576;
  assign n28578 = ~n28569 & n28577;
  assign n28579 = ~n28575 & ~n28578;
  assign n28580 = ~n28025 & ~n28579;
  assign n28581 = n28015 & n28022;
  assign n28582 = ~n28015 & ~n28022;
  assign n28583 = ~n28581 & ~n28582;
  assign n28584 = ~n28573 & ~n28576;
  assign n28585 = n28573 & n28576;
  assign n28586 = ~n28584 & ~n28585;
  assign n28587 = ~n28583 & ~n28586;
  assign n28588 = ~n28580 & ~n28587;
  assign n28589 = ~n24906 & ~n26688;
  assign n28590 = ~n26689 & ~n28589;
  assign n28591 = n28588 & n28590;
  assign n28592 = ~n28588 & ~n28590;
  assign n28593 = ~n28591 & ~n28592;
  assign n28594 = ~n26651 & n26661;
  assign n28595 = ~n26661 & ~n26669;
  assign n28596 = ~n28594 & ~n28595;
  assign n28597 = ~n26678 & ~n28596;
  assign n28598 = n26661 & ~n26669;
  assign n28599 = ~n26651 & ~n26661;
  assign n28600 = ~n28598 & ~n28599;
  assign n28601 = ~n26646 & ~n28600;
  assign n28602 = ~n28597 & ~n28601;
  assign n28603 = n26662 & ~n28602;
  assign n28604 = ~pi259 & n28603;
  assign n28605 = pi259 & ~n28603;
  assign n28606 = pi156 & n28605;
  assign n28607 = ~n28604 & ~n28606;
  assign n28608 = n26683 & n28607;
  assign n28609 = ~n26683 & ~n28607;
  assign n28610 = ~n28608 & ~n28609;
  assign n28611 = pi258 & ~n28610;
  assign n28612 = pi157 & n28611;
  assign n28613 = pi157 & pi258;
  assign n28614 = ~n26683 & n28607;
  assign n28615 = n26683 & ~n28607;
  assign n28616 = ~n28614 & ~n28615;
  assign n28617 = ~n28613 & ~n28616;
  assign n28618 = ~n28612 & ~n28617;
  assign n28619 = ~n28593 & ~n28618;
  assign n28620 = n28588 & ~n28590;
  assign n28621 = ~n28588 & n28590;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = pi258 & ~n28616;
  assign n28624 = pi157 & n28623;
  assign n28625 = ~n28610 & ~n28613;
  assign n28626 = ~n28624 & ~n28625;
  assign n28627 = ~n28622 & ~n28626;
  assign n28628 = ~n28619 & ~n28627;
  assign n28629 = pi322 & n28628;
  assign n28630 = ~n28011 & ~n28629;
  assign n28631 = n28010 & n28628;
  assign n28632 = n1445 & n28631;
  assign n28633 = ~n28630 & ~n28632;
  assign n28634 = ~n28007 & ~n28633;
  assign n28635 = ~n28002 & n28004;
  assign n28636 = n28002 & ~n28004;
  assign n28637 = ~n28635 & ~n28636;
  assign n28638 = ~n28011 & n28628;
  assign n28639 = pi322 & n28638;
  assign n28640 = n28010 & ~n28629;
  assign n28641 = pi323 & n28640;
  assign n28642 = ~n28639 & ~n28641;
  assign n28643 = ~n28637 & ~n28642;
  assign n28644 = ~n28634 & ~n28643;
  assign n28645 = ~n26163 & n26707;
  assign n28646 = n26163 & ~n26707;
  assign n28647 = ~n27980 & ~n28646;
  assign n28648 = ~n28645 & ~n28647;
  assign n28649 = n28644 & ~n28648;
  assign n28650 = ~n28644 & n28648;
  assign n28651 = ~n28649 & ~n28650;
  assign n28652 = pi326 & n21479;
  assign n28653 = pi325 & n26706;
  assign n28654 = n28652 & n28653;
  assign n28655 = ~n28652 & ~n28653;
  assign n28656 = ~n28654 & ~n28655;
  assign n28657 = ~n28651 & ~n28656;
  assign n28658 = ~n28644 & ~n28648;
  assign n28659 = n28644 & n28648;
  assign n28660 = ~n28658 & ~n28659;
  assign n28661 = ~n28652 & n28653;
  assign n28662 = n28652 & ~n28653;
  assign n28663 = ~n28661 & ~n28662;
  assign n28664 = ~n28660 & ~n28663;
  assign n28665 = ~n28657 & ~n28664;
  assign n28666 = ~n28001 & ~n28665;
  assign n28667 = n27994 & n27998;
  assign n28668 = ~n27994 & ~n27998;
  assign n28669 = ~n28667 & ~n28668;
  assign n28670 = ~n28656 & ~n28660;
  assign n28671 = ~n28651 & ~n28663;
  assign n28672 = ~n28670 & ~n28671;
  assign n28673 = ~n28669 & ~n28672;
  assign n28674 = ~n28666 & ~n28673;
  assign n28675 = ~n27975 & n28674;
  assign n28676 = n27975 & ~n28674;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = pi329 & n19539;
  assign n28679 = pi328 & n19557;
  assign n28680 = n28678 & n28679;
  assign n28681 = ~n28678 & ~n28679;
  assign n28682 = ~n28680 & ~n28681;
  assign n28683 = ~n28677 & ~n28682;
  assign n28684 = n27975 & n28674;
  assign n28685 = ~n27975 & ~n28674;
  assign n28686 = ~n28684 & ~n28685;
  assign n28687 = ~n28678 & n28679;
  assign n28688 = n28678 & ~n28679;
  assign n28689 = ~n28687 & ~n28688;
  assign n28690 = ~n28686 & ~n28689;
  assign n28691 = ~n28683 & ~n28690;
  assign n28692 = ~n27974 & ~n28691;
  assign n28693 = n27968 & n27971;
  assign n28694 = ~n27968 & ~n27971;
  assign n28695 = ~n28693 & ~n28694;
  assign n28696 = ~n28682 & ~n28686;
  assign n28697 = ~n28677 & ~n28689;
  assign n28698 = ~n28696 & ~n28697;
  assign n28699 = ~n28695 & ~n28698;
  assign n28700 = ~n28692 & ~n28699;
  assign n28701 = ~n27948 & ~n28700;
  assign n28702 = n27948 & n28700;
  assign n28703 = ~n28701 & ~n28702;
  assign n28704 = n13762 & ~n28703;
  assign n28705 = pi331 & n28704;
  assign n28706 = pi331 & n13762;
  assign n28707 = n27948 & ~n28700;
  assign n28708 = ~n27948 & n28700;
  assign n28709 = ~n28707 & ~n28708;
  assign n28710 = ~n28706 & ~n28709;
  assign n28711 = ~n28705 & ~n28710;
  assign n28712 = ~n27935 & ~n28711;
  assign n28713 = ~n27925 & n27932;
  assign n28714 = n27925 & ~n27932;
  assign n28715 = ~n28713 & ~n28714;
  assign n28716 = n13762 & ~n28709;
  assign n28717 = pi331 & n28716;
  assign n28718 = ~n28703 & ~n28706;
  assign n28719 = ~n28717 & ~n28718;
  assign n28720 = ~n28715 & ~n28719;
  assign n28721 = ~n28712 & ~n28720;
  assign n28722 = ~n26087 & n26105;
  assign n28723 = n26087 & ~n26105;
  assign n28724 = n26853 & ~n28723;
  assign n28725 = ~n28722 & ~n28724;
  assign n28726 = n28721 & n28725;
  assign n28727 = ~n28721 & ~n28725;
  assign n28728 = ~n28726 & ~n28727;
  assign n28729 = pi333 & n11711;
  assign n28730 = ~n26818 & ~n26841;
  assign n28731 = ~n26848 & n28730;
  assign n28732 = ~n26839 & ~n26841;
  assign n28733 = ~n26807 & n28732;
  assign n28734 = ~n26840 & ~n28733;
  assign n28735 = ~n28731 & n28734;
  assign n28736 = pi332 & n12917;
  assign n28737 = n28735 & ~n28736;
  assign n28738 = n12917 & ~n28735;
  assign n28739 = pi332 & n28738;
  assign n28740 = ~n28737 & ~n28739;
  assign n28741 = ~n28729 & n28740;
  assign n28742 = n28729 & ~n28740;
  assign n28743 = ~n28741 & ~n28742;
  assign n28744 = pi334 & n11384;
  assign n28745 = pi334 & n26869;
  assign n28746 = ~n26096 & ~n26862;
  assign n28747 = ~n28745 & ~n28746;
  assign n28748 = n11366 & ~n28747;
  assign n28749 = pi334 & n28748;
  assign n28750 = n26105 & ~n27875;
  assign n28751 = ~n26105 & ~n27884;
  assign n28752 = ~n28750 & ~n28751;
  assign n28753 = pi334 & n11366;
  assign n28754 = n28747 & ~n28753;
  assign n28755 = ~n28752 & ~n28754;
  assign n28756 = ~n28749 & ~n28755;
  assign n28757 = n28744 & n28756;
  assign n28758 = ~n28744 & ~n28756;
  assign n28759 = ~n28757 & ~n28758;
  assign n28760 = ~n28743 & ~n28759;
  assign n28761 = n28729 & n28740;
  assign n28762 = ~n28729 & ~n28740;
  assign n28763 = ~n28761 & ~n28762;
  assign n28764 = ~n28744 & n28756;
  assign n28765 = n28744 & ~n28756;
  assign n28766 = ~n28764 & ~n28765;
  assign n28767 = ~n28763 & ~n28766;
  assign n28768 = ~n28760 & ~n28767;
  assign n28769 = ~n28728 & ~n28768;
  assign n28770 = n28721 & ~n28725;
  assign n28771 = ~n28721 & n28725;
  assign n28772 = ~n28770 & ~n28771;
  assign n28773 = ~n28759 & ~n28763;
  assign n28774 = ~n28743 & ~n28766;
  assign n28775 = ~n28773 & ~n28774;
  assign n28776 = ~n28772 & ~n28775;
  assign n28777 = ~n28769 & ~n28776;
  assign n28778 = ~n27911 & n28777;
  assign n28779 = n27911 & ~n28777;
  assign n28780 = ~n28778 & ~n28779;
  assign n28781 = pi337 & n9205;
  assign n28782 = pi336 & n10561;
  assign n28783 = n26896 & ~n27901;
  assign n28784 = ~n27898 & ~n28783;
  assign n28785 = ~n28782 & ~n28784;
  assign n28786 = n10561 & ~n28783;
  assign n28787 = pi336 & n28786;
  assign n28788 = ~n27898 & n28787;
  assign n28789 = ~n28785 & ~n28788;
  assign n28790 = n28781 & ~n28789;
  assign n28791 = ~n28781 & n28789;
  assign n28792 = ~n28790 & ~n28791;
  assign n28793 = ~n28780 & ~n28792;
  assign n28794 = n27911 & n28777;
  assign n28795 = ~n27911 & ~n28777;
  assign n28796 = ~n28794 & ~n28795;
  assign n28797 = ~n28781 & ~n28789;
  assign n28798 = n28781 & n28789;
  assign n28799 = ~n28797 & ~n28798;
  assign n28800 = ~n28796 & ~n28799;
  assign n28801 = ~n28793 & ~n28800;
  assign n28802 = ~n27910 & ~n28801;
  assign n28803 = n27892 & ~n27907;
  assign n28804 = ~n27892 & n27907;
  assign n28805 = ~n28803 & ~n28804;
  assign n28806 = ~n28792 & ~n28796;
  assign n28807 = ~n28780 & ~n28799;
  assign n28808 = ~n28806 & ~n28807;
  assign n28809 = ~n28805 & ~n28808;
  assign n28810 = ~n28802 & ~n28809;
  assign n28811 = ~n26048 & n26066;
  assign n28812 = n26048 & ~n26066;
  assign n28813 = n26950 & ~n28812;
  assign n28814 = ~n28811 & ~n28813;
  assign n28815 = n28810 & n28814;
  assign n28816 = ~n28810 & ~n28814;
  assign n28817 = ~n28815 & ~n28816;
  assign n28818 = pi339 & n5973;
  assign n28819 = ~n26923 & ~n26938;
  assign n28820 = ~n26945 & n28819;
  assign n28821 = ~n26936 & ~n26938;
  assign n28822 = ~n26906 & n28821;
  assign n28823 = ~n26937 & ~n28822;
  assign n28824 = ~n28820 & n28823;
  assign n28825 = pi338 & n6556;
  assign n28826 = n28824 & ~n28825;
  assign n28827 = n6556 & ~n28824;
  assign n28828 = pi338 & n28827;
  assign n28829 = ~n28826 & ~n28828;
  assign n28830 = ~n28818 & n28829;
  assign n28831 = n28818 & ~n28829;
  assign n28832 = ~n28830 & ~n28831;
  assign n28833 = pi340 & n5732;
  assign n28834 = pi340 & n26966;
  assign n28835 = ~n26057 & ~n26959;
  assign n28836 = ~n28834 & ~n28835;
  assign n28837 = n5714 & ~n28836;
  assign n28838 = pi340 & n28837;
  assign n28839 = n26066 & ~n27836;
  assign n28840 = ~n26066 & ~n27845;
  assign n28841 = ~n28839 & ~n28840;
  assign n28842 = pi340 & n5714;
  assign n28843 = n28836 & ~n28842;
  assign n28844 = ~n28841 & ~n28843;
  assign n28845 = ~n28838 & ~n28844;
  assign n28846 = n28833 & n28845;
  assign n28847 = ~n28833 & ~n28845;
  assign n28848 = ~n28846 & ~n28847;
  assign n28849 = ~n28832 & ~n28848;
  assign n28850 = n28818 & n28829;
  assign n28851 = ~n28818 & ~n28829;
  assign n28852 = ~n28850 & ~n28851;
  assign n28853 = ~n28833 & n28845;
  assign n28854 = n28833 & ~n28845;
  assign n28855 = ~n28853 & ~n28854;
  assign n28856 = ~n28852 & ~n28855;
  assign n28857 = ~n28849 & ~n28856;
  assign n28858 = ~n28817 & ~n28857;
  assign n28859 = n28810 & ~n28814;
  assign n28860 = ~n28810 & n28814;
  assign n28861 = ~n28859 & ~n28860;
  assign n28862 = ~n28848 & ~n28852;
  assign n28863 = ~n28832 & ~n28855;
  assign n28864 = ~n28862 & ~n28863;
  assign n28865 = ~n28861 & ~n28864;
  assign n28866 = ~n28858 & ~n28865;
  assign n28867 = ~n27872 & n28866;
  assign n28868 = n27872 & ~n28866;
  assign n28869 = ~n28867 & ~n28868;
  assign n28870 = pi343 & n4596;
  assign n28871 = pi342 & n5257;
  assign n28872 = n26993 & ~n27862;
  assign n28873 = ~n27859 & ~n28872;
  assign n28874 = ~n28871 & ~n28873;
  assign n28875 = n5257 & ~n28872;
  assign n28876 = pi342 & n28875;
  assign n28877 = ~n27859 & n28876;
  assign n28878 = ~n28874 & ~n28877;
  assign n28879 = n28870 & ~n28878;
  assign n28880 = ~n28870 & n28878;
  assign n28881 = ~n28879 & ~n28880;
  assign n28882 = ~n28869 & ~n28881;
  assign n28883 = n27872 & n28866;
  assign n28884 = ~n27872 & ~n28866;
  assign n28885 = ~n28883 & ~n28884;
  assign n28886 = ~n28870 & ~n28878;
  assign n28887 = n28870 & n28878;
  assign n28888 = ~n28886 & ~n28887;
  assign n28889 = ~n28885 & ~n28888;
  assign n28890 = ~n28882 & ~n28889;
  assign n28891 = ~n27871 & ~n28890;
  assign n28892 = n27853 & ~n27868;
  assign n28893 = ~n27853 & n27868;
  assign n28894 = ~n28892 & ~n28893;
  assign n28895 = ~n28881 & ~n28885;
  assign n28896 = ~n28869 & ~n28888;
  assign n28897 = ~n28895 & ~n28896;
  assign n28898 = ~n28894 & ~n28897;
  assign n28899 = ~n28891 & ~n28898;
  assign n28900 = ~n25996 & n26020;
  assign n28901 = n25996 & ~n26020;
  assign n28902 = n27048 & ~n28901;
  assign n28903 = ~n28900 & ~n28902;
  assign n28904 = n28899 & n28903;
  assign n28905 = ~n28899 & ~n28903;
  assign n28906 = ~n28904 & ~n28905;
  assign n28907 = pi345 & n2464;
  assign n28908 = ~n27020 & ~n27036;
  assign n28909 = ~n27043 & n28908;
  assign n28910 = ~n27034 & ~n27036;
  assign n28911 = ~n27003 & n28910;
  assign n28912 = ~n27035 & ~n28911;
  assign n28913 = ~n28909 & n28912;
  assign n28914 = pi344 & n2887;
  assign n28915 = n28913 & ~n28914;
  assign n28916 = n2887 & ~n28913;
  assign n28917 = pi344 & n28916;
  assign n28918 = ~n28915 & ~n28917;
  assign n28919 = ~n28907 & n28918;
  assign n28920 = n28907 & ~n28918;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = pi347 & n1729;
  assign n28923 = pi346 & n2091;
  assign n28924 = n1729 & ~n26008;
  assign n28925 = pi345 & n28924;
  assign n28926 = ~n24161 & ~n25999;
  assign n28927 = ~n27054 & ~n28926;
  assign n28928 = ~n28925 & n28927;
  assign n28929 = ~n27059 & ~n28928;
  assign n28930 = ~n27055 & n28929;
  assign n28931 = ~n28923 & ~n28930;
  assign n28932 = n26020 & n28931;
  assign n28933 = n27055 & ~n28929;
  assign n28934 = n28923 & ~n28933;
  assign n28935 = ~n26020 & n28934;
  assign n28936 = ~n28932 & ~n28935;
  assign n28937 = ~n27797 & ~n28936;
  assign n28938 = n26020 & n28934;
  assign n28939 = ~n26020 & n28931;
  assign n28940 = ~n28938 & ~n28939;
  assign n28941 = ~n27806 & ~n28940;
  assign n28942 = ~n28923 & ~n28929;
  assign n28943 = n27055 & n28942;
  assign n28944 = n28923 & n28929;
  assign n28945 = ~n27055 & n28944;
  assign n28946 = ~n28943 & ~n28945;
  assign n28947 = ~n28941 & n28946;
  assign n28948 = ~n28937 & n28947;
  assign n28949 = n28922 & ~n28948;
  assign n28950 = ~n28922 & n28948;
  assign n28951 = ~n28949 & ~n28950;
  assign n28952 = ~n28921 & ~n28951;
  assign n28953 = n28907 & n28918;
  assign n28954 = ~n28907 & ~n28918;
  assign n28955 = ~n28953 & ~n28954;
  assign n28956 = ~n28922 & ~n28948;
  assign n28957 = n28922 & n28948;
  assign n28958 = ~n28956 & ~n28957;
  assign n28959 = ~n28955 & ~n28958;
  assign n28960 = ~n28952 & ~n28959;
  assign n28961 = ~n28906 & ~n28960;
  assign n28962 = n28899 & ~n28903;
  assign n28963 = ~n28899 & n28903;
  assign n28964 = ~n28962 & ~n28963;
  assign n28965 = ~n28951 & ~n28955;
  assign n28966 = ~n28921 & ~n28958;
  assign n28967 = ~n28965 & ~n28966;
  assign n28968 = ~n28964 & ~n28967;
  assign n28969 = ~n28961 & ~n28968;
  assign n28970 = n27833 & n28969;
  assign n28971 = ~n27833 & ~n28969;
  assign n28972 = ~n28970 & ~n28971;
  assign n28973 = ~n1256 & ~n28972;
  assign n28974 = pi349 & n28973;
  assign n28975 = pi349 & ~n1256;
  assign n28976 = ~n27833 & n28969;
  assign n28977 = n27833 & ~n28969;
  assign n28978 = ~n28976 & ~n28977;
  assign n28979 = ~n28975 & ~n28978;
  assign n28980 = ~n28974 & ~n28979;
  assign n28981 = ~n27826 & ~n28980;
  assign n28982 = n27814 & ~n27823;
  assign n28983 = ~n27814 & n27823;
  assign n28984 = ~n28982 & ~n28983;
  assign n28985 = ~n1256 & ~n28978;
  assign n28986 = pi349 & n28985;
  assign n28987 = ~n28972 & ~n28975;
  assign n28988 = ~n28986 & ~n28987;
  assign n28989 = ~n28984 & ~n28988;
  assign n28990 = ~n28981 & ~n28989;
  assign n28991 = ~n27794 & ~n28990;
  assign n28992 = n27794 & n28990;
  assign n28993 = ~n28991 & ~n28992;
  assign n28994 = ~pi286 & ~n25989;
  assign n28995 = pi286 & n25989;
  assign n28996 = n27127 & ~n27137;
  assign n28997 = pi350 & ~n27127;
  assign n28998 = n1156 & n28997;
  assign n28999 = ~n28996 & ~n28998;
  assign n29000 = ~n28995 & ~n28999;
  assign n29001 = ~n28994 & ~n29000;
  assign n29002 = ~pi287 & n29001;
  assign n29003 = pi287 & ~n29001;
  assign n29004 = ~n29002 & ~n29003;
  assign n29005 = n1156 & ~n29004;
  assign n29006 = pi351 & n29005;
  assign n29007 = pi351 & n1156;
  assign n29008 = ~pi287 & ~n29001;
  assign n29009 = pi287 & n29001;
  assign n29010 = ~n29008 & ~n29009;
  assign n29011 = ~n29007 & ~n29010;
  assign n29012 = ~n29006 & ~n29011;
  assign n29013 = ~n28993 & ~n29012;
  assign n29014 = ~n27794 & n28990;
  assign n29015 = n27794 & ~n28990;
  assign n29016 = ~n29014 & ~n29015;
  assign n29017 = n1156 & ~n29010;
  assign n29018 = pi351 & n29017;
  assign n29019 = ~n29004 & ~n29007;
  assign n29020 = ~n29018 & ~n29019;
  assign n29021 = ~n29016 & ~n29020;
  assign n29022 = ~n29013 & ~n29021;
  assign n29023 = ~n27788 & ~n29022;
  assign n29024 = n27788 & n29022;
  assign n29025 = ~n29023 & ~n29024;
  assign n29026 = n25983 & ~n27154;
  assign n29027 = ~n25983 & n27154;
  assign n29028 = ~n27142 & ~n29027;
  assign n29029 = ~n29026 & ~n29028;
  assign n29030 = n29025 & n29029;
  assign n29031 = ~n29025 & ~n29029;
  assign n29032 = ~n29030 & ~n29031;
  assign n29033 = ~n831 & ~n29032;
  assign n29034 = ~n27164 & ~n29033;
  assign n29035 = pi161 & ~n29034;
  assign n29036 = ~n27163 & ~n29035;
  assign po222 = ~pi160 & n29036;
  assign n29038 = pi094 & ~pi161;
  assign n29039 = n27789 & n28990;
  assign n29040 = ~n27789 & ~n28990;
  assign n29041 = ~n1154 & ~n29040;
  assign n29042 = ~n29039 & ~n29041;
  assign n29043 = n1256 & ~n29042;
  assign n29044 = n1154 & ~n28990;
  assign n29045 = ~n1154 & n28990;
  assign n29046 = ~n27789 & ~n29045;
  assign n29047 = ~n29044 & ~n29046;
  assign n29048 = ~n1256 & ~n29047;
  assign n29049 = ~n29043 & ~n29048;
  assign n29050 = pi350 & ~n29049;
  assign n29051 = n27814 & n28922;
  assign n29052 = ~n28918 & ~n28948;
  assign n29053 = n28918 & n28948;
  assign n29054 = ~n29052 & ~n29053;
  assign n29055 = n2464 & ~n29054;
  assign n29056 = pi345 & n29055;
  assign n29057 = ~n28918 & n28948;
  assign n29058 = n28918 & ~n28948;
  assign n29059 = ~n29057 & ~n29058;
  assign n29060 = ~n28907 & ~n29059;
  assign n29061 = ~n29056 & ~n29060;
  assign n29062 = ~n28906 & ~n29061;
  assign n29063 = n2464 & ~n29059;
  assign n29064 = pi345 & n29063;
  assign n29065 = ~n28907 & ~n29054;
  assign n29066 = ~n29064 & ~n29065;
  assign n29067 = ~n28964 & ~n29066;
  assign n29068 = ~n29062 & ~n29067;
  assign n29069 = ~n27814 & ~n28922;
  assign n29070 = n29068 & ~n29069;
  assign n29071 = ~n29051 & ~n29070;
  assign n29072 = ~n27814 & n28969;
  assign n29073 = n27814 & ~n28969;
  assign n29074 = ~n29072 & ~n29073;
  assign n29075 = ~n27833 & ~n29074;
  assign n29076 = n27814 & n28969;
  assign n29077 = ~n27814 & ~n28969;
  assign n29078 = ~n29076 & ~n29077;
  assign n29079 = n27833 & ~n29078;
  assign n29080 = ~n29075 & ~n29079;
  assign n29081 = n27823 & ~n28975;
  assign n29082 = ~n29080 & ~n29081;
  assign n29083 = ~n1256 & ~n27823;
  assign n29084 = pi349 & n29083;
  assign n29085 = ~n29082 & ~n29084;
  assign n29086 = ~n29071 & n29085;
  assign n29087 = n29071 & ~n29085;
  assign n29088 = ~n29086 & ~n29087;
  assign n29089 = pi347 & n2091;
  assign n29090 = n27853 & n27872;
  assign n29091 = ~n27853 & ~n27872;
  assign n29092 = n28866 & ~n29091;
  assign n29093 = ~n29090 & ~n29092;
  assign n29094 = ~n27853 & n28866;
  assign n29095 = n27853 & ~n28866;
  assign n29096 = ~n29094 & ~n29095;
  assign n29097 = n27872 & ~n28878;
  assign n29098 = ~n27872 & n28878;
  assign n29099 = ~n29097 & ~n29098;
  assign n29100 = n27868 & ~n28870;
  assign n29101 = ~n29099 & ~n29100;
  assign n29102 = ~n29096 & n29101;
  assign n29103 = ~n27868 & n28870;
  assign n29104 = ~n27853 & ~n28866;
  assign n29105 = n27853 & n28866;
  assign n29106 = ~n29104 & ~n29105;
  assign n29107 = ~n27872 & ~n28878;
  assign n29108 = n27872 & n28878;
  assign n29109 = ~n29107 & ~n29108;
  assign n29110 = ~n29100 & ~n29109;
  assign n29111 = ~n29106 & n29110;
  assign n29112 = ~n29103 & ~n29111;
  assign n29113 = ~n29102 & n29112;
  assign n29114 = ~n29093 & n29113;
  assign n29115 = n29093 & ~n29113;
  assign n29116 = ~n29114 & ~n29115;
  assign n29117 = pi341 & n5732;
  assign n29118 = n27892 & n27911;
  assign n29119 = ~n27892 & ~n27911;
  assign n29120 = n28777 & ~n29119;
  assign n29121 = ~n29118 & ~n29120;
  assign n29122 = ~n27892 & n28777;
  assign n29123 = n27892 & ~n28777;
  assign n29124 = ~n29122 & ~n29123;
  assign n29125 = n27911 & ~n28789;
  assign n29126 = ~n27911 & n28789;
  assign n29127 = ~n29125 & ~n29126;
  assign n29128 = n27907 & ~n28781;
  assign n29129 = ~n29127 & ~n29128;
  assign n29130 = ~n29124 & n29129;
  assign n29131 = ~n27907 & n28781;
  assign n29132 = ~n27892 & ~n28777;
  assign n29133 = n27892 & n28777;
  assign n29134 = ~n29132 & ~n29133;
  assign n29135 = ~n27911 & ~n28789;
  assign n29136 = n27911 & n28789;
  assign n29137 = ~n29135 & ~n29136;
  assign n29138 = ~n29128 & ~n29137;
  assign n29139 = ~n29134 & n29138;
  assign n29140 = ~n29131 & ~n29139;
  assign n29141 = ~n29130 & n29140;
  assign n29142 = ~n29121 & n29141;
  assign n29143 = n29121 & ~n29141;
  assign n29144 = ~n29142 & ~n29143;
  assign n29145 = pi335 & n11384;
  assign n29146 = n27925 & n28678;
  assign n29147 = n19557 & ~n28677;
  assign n29148 = pi328 & n29147;
  assign n29149 = ~n28679 & ~n28686;
  assign n29150 = ~n29148 & ~n29149;
  assign n29151 = ~n27974 & ~n29150;
  assign n29152 = n19557 & ~n28686;
  assign n29153 = pi328 & n29152;
  assign n29154 = ~n28677 & ~n28679;
  assign n29155 = ~n29153 & ~n29154;
  assign n29156 = ~n28695 & ~n29155;
  assign n29157 = ~n29151 & ~n29156;
  assign n29158 = ~n27925 & ~n28678;
  assign n29159 = n29157 & ~n29158;
  assign n29160 = ~n29146 & ~n29159;
  assign n29161 = ~n27932 & n28706;
  assign n29162 = n27925 & ~n28700;
  assign n29163 = ~n27925 & n28700;
  assign n29164 = ~n29162 & ~n29163;
  assign n29165 = ~n27948 & ~n29164;
  assign n29166 = n27925 & n28700;
  assign n29167 = ~n27925 & ~n28700;
  assign n29168 = ~n29166 & ~n29167;
  assign n29169 = n27948 & ~n29168;
  assign n29170 = ~n29165 & ~n29169;
  assign n29171 = n27932 & ~n28706;
  assign n29172 = ~n29170 & ~n29171;
  assign n29173 = ~n29161 & ~n29172;
  assign n29174 = ~n29160 & n29173;
  assign n29175 = n29160 & ~n29173;
  assign n29176 = ~n29174 & ~n29175;
  assign n29177 = pi330 & n19539;
  assign n29178 = n13762 & ~n27936;
  assign n29179 = ~n27937 & ~n29178;
  assign n29180 = n18461 & ~n29179;
  assign n29181 = pi330 & n29180;
  assign n29182 = ~n18461 & ~n29178;
  assign n29183 = pi330 & ~n29182;
  assign n29184 = ~n27937 & ~n29183;
  assign n29185 = ~n29168 & ~n29184;
  assign n29186 = ~n29181 & ~n29185;
  assign n29187 = ~n29177 & ~n29186;
  assign n29188 = n29164 & ~n29184;
  assign n29189 = n19539 & ~n29188;
  assign n29190 = pi330 & n29189;
  assign n29191 = ~n29181 & n29190;
  assign n29192 = ~n29187 & ~n29191;
  assign n29193 = n27968 & n27975;
  assign n29194 = ~n27968 & ~n27975;
  assign n29195 = n28674 & ~n29194;
  assign n29196 = ~n29193 & ~n29195;
  assign n29197 = ~n27971 & n28679;
  assign n29198 = ~n27968 & ~n28674;
  assign n29199 = n27968 & n28674;
  assign n29200 = ~n29198 & ~n29199;
  assign n29201 = n27975 & ~n29200;
  assign n29202 = n27968 & ~n28674;
  assign n29203 = ~n27968 & n28674;
  assign n29204 = ~n29202 & ~n29203;
  assign n29205 = ~n27975 & ~n29204;
  assign n29206 = ~n29201 & ~n29205;
  assign n29207 = n27971 & ~n28679;
  assign n29208 = ~n29206 & ~n29207;
  assign n29209 = ~n29197 & ~n29208;
  assign n29210 = ~n29196 & n29209;
  assign n29211 = n29196 & ~n29209;
  assign n29212 = ~n29210 & ~n29211;
  assign n29213 = pi327 & n21479;
  assign n29214 = ~n27994 & n28653;
  assign n29215 = n27994 & ~n28653;
  assign n29216 = ~n28651 & ~n29215;
  assign n29217 = ~n29214 & ~n29216;
  assign n29218 = ~n27994 & n28648;
  assign n29219 = n27994 & ~n28648;
  assign n29220 = ~n29218 & ~n29219;
  assign n29221 = ~n28644 & n28653;
  assign n29222 = n28644 & ~n28653;
  assign n29223 = ~n29221 & ~n29222;
  assign n29224 = n27998 & ~n28652;
  assign n29225 = ~n29223 & ~n29224;
  assign n29226 = ~n29220 & n29225;
  assign n29227 = ~n27998 & n28652;
  assign n29228 = ~n27994 & ~n28648;
  assign n29229 = n27994 & n28648;
  assign n29230 = ~n29228 & ~n29229;
  assign n29231 = n28644 & n28653;
  assign n29232 = ~n28644 & ~n28653;
  assign n29233 = ~n29231 & ~n29232;
  assign n29234 = ~n29224 & ~n29233;
  assign n29235 = ~n29230 & n29234;
  assign n29236 = ~n29227 & ~n29235;
  assign n29237 = ~n29226 & n29236;
  assign n29238 = n29217 & n29237;
  assign n29239 = ~n29217 & ~n29237;
  assign n29240 = ~n29238 & ~n29239;
  assign n29241 = pi324 & n28010;
  assign n29242 = ~n28004 & n28010;
  assign n29243 = pi323 & n29242;
  assign n29244 = n28004 & ~n28011;
  assign n29245 = n28628 & ~n29244;
  assign n29246 = pi322 & n29245;
  assign n29247 = ~n29243 & ~n29246;
  assign n29248 = ~n29241 & ~n29247;
  assign n29249 = n29241 & n29247;
  assign n29250 = ~n29248 & ~n29249;
  assign n29251 = pi323 & n28628;
  assign n29252 = pi154 & pi262;
  assign n29253 = pi151 & pi265;
  assign n29254 = pi148 & pi268;
  assign n29255 = pi145 & pi271;
  assign n29256 = pi142 & pi274;
  assign n29257 = pi139 & pi277;
  assign n29258 = pi136 & pi280;
  assign n29259 = pi134 & pi282;
  assign n29260 = n28114 & n28119;
  assign n29261 = ~n28114 & ~n28119;
  assign n29262 = ~n29260 & ~n29261;
  assign n29263 = pi282 & ~n29262;
  assign n29264 = pi133 & n29263;
  assign n29265 = pi133 & pi283;
  assign n29266 = pi131 & pi285;
  assign n29267 = pi287 & ~n26196;
  assign n29268 = pi286 & n29267;
  assign n29269 = ~pi287 & n26196;
  assign n29270 = pi286 & ~n29269;
  assign n29271 = ~pi286 & ~n29267;
  assign n29272 = pi285 & ~n29271;
  assign n29273 = ~n29270 & ~n29272;
  assign n29274 = pi129 & ~n29273;
  assign n29275 = ~n29268 & ~n29274;
  assign n29276 = pi128 & ~n29275;
  assign n29277 = pi286 & ~n26196;
  assign n29278 = n26200 & n29277;
  assign n29279 = ~n29276 & ~n29278;
  assign n29280 = pi129 & pi287;
  assign n29281 = pi288 & ~n29280;
  assign n29282 = pi128 & n29281;
  assign n29283 = pi128 & pi288;
  assign n29284 = pi287 & ~n29283;
  assign n29285 = pi129 & n29284;
  assign n29286 = ~n29282 & ~n29285;
  assign n29287 = n29279 & n29286;
  assign n29288 = ~n29279 & ~n29286;
  assign n29289 = ~n29287 & ~n29288;
  assign n29290 = pi286 & ~n29289;
  assign n29291 = pi130 & n29290;
  assign n29292 = pi130 & pi286;
  assign n29293 = ~n29279 & n29286;
  assign n29294 = n29279 & ~n29286;
  assign n29295 = ~n29293 & ~n29294;
  assign n29296 = ~n29292 & ~n29295;
  assign n29297 = ~n29291 & ~n29296;
  assign n29298 = ~n28049 & ~n28075;
  assign n29299 = ~n26200 & ~n28042;
  assign n29300 = ~n28072 & ~n29299;
  assign n29301 = n28049 & ~n29300;
  assign n29302 = ~n29298 & ~n29301;
  assign n29303 = ~n28091 & n29302;
  assign n29304 = n28091 & ~n29302;
  assign n29305 = pi285 & ~n29304;
  assign n29306 = pi130 & n29305;
  assign n29307 = ~n29303 & ~n29306;
  assign n29308 = ~n29297 & ~n29307;
  assign n29309 = pi130 & pi285;
  assign n29310 = ~n29303 & ~n29309;
  assign n29311 = ~n29304 & ~n29310;
  assign n29312 = n29297 & ~n29311;
  assign n29313 = ~n29308 & ~n29312;
  assign n29314 = ~n29266 & n29313;
  assign n29315 = n29266 & ~n29313;
  assign n29316 = ~n29314 & ~n29315;
  assign n29317 = pi132 & pi284;
  assign n29318 = ~n28084 & ~n28091;
  assign n29319 = n28084 & n28091;
  assign n29320 = ~n29318 & ~n29319;
  assign n29321 = ~n28106 & n29320;
  assign n29322 = n28106 & ~n29320;
  assign n29323 = n28041 & ~n29322;
  assign n29324 = ~n29321 & ~n29323;
  assign n29325 = n29317 & ~n29324;
  assign n29326 = ~n28041 & ~n29321;
  assign n29327 = ~n29322 & ~n29326;
  assign n29328 = ~n29317 & ~n29327;
  assign n29329 = ~n29325 & ~n29328;
  assign n29330 = ~n29316 & ~n29329;
  assign n29331 = ~n29266 & ~n29313;
  assign n29332 = n29266 & n29313;
  assign n29333 = ~n29331 & ~n29332;
  assign n29334 = ~n29317 & ~n29324;
  assign n29335 = n29317 & ~n29327;
  assign n29336 = ~n29334 & ~n29335;
  assign n29337 = ~n29333 & ~n29336;
  assign n29338 = ~n29330 & ~n29337;
  assign n29339 = ~n29265 & n29338;
  assign n29340 = n29265 & ~n29338;
  assign n29341 = ~n29339 & ~n29340;
  assign n29342 = n28040 & n28119;
  assign n29343 = ~n28099 & n28106;
  assign n29344 = n28099 & ~n28106;
  assign n29345 = ~n29343 & ~n29344;
  assign n29346 = ~n28040 & ~n28119;
  assign n29347 = ~n29345 & ~n29346;
  assign n29348 = ~n29342 & ~n29347;
  assign n29349 = ~n29341 & ~n29348;
  assign n29350 = ~n29265 & ~n29338;
  assign n29351 = n29265 & n29338;
  assign n29352 = ~n29350 & ~n29351;
  assign n29353 = ~n28099 & ~n28106;
  assign n29354 = n28099 & n28106;
  assign n29355 = ~n29353 & ~n29354;
  assign n29356 = ~n29342 & ~n29355;
  assign n29357 = ~n29346 & ~n29356;
  assign n29358 = ~n29352 & ~n29357;
  assign n29359 = ~n29349 & ~n29358;
  assign n29360 = ~n28039 & n29262;
  assign n29361 = ~n28128 & ~n29360;
  assign n29362 = ~n29359 & ~n29361;
  assign n29363 = ~n29264 & n29362;
  assign n29364 = ~n29264 & ~n29361;
  assign n29365 = n29359 & ~n29364;
  assign n29366 = ~n29363 & ~n29365;
  assign n29367 = ~n29259 & ~n29366;
  assign n29368 = n29359 & ~n29361;
  assign n29369 = ~n29264 & n29368;
  assign n29370 = ~n29359 & ~n29364;
  assign n29371 = ~n29369 & ~n29370;
  assign n29372 = pi282 & ~n29371;
  assign n29373 = pi134 & n29372;
  assign n29374 = ~n29367 & ~n29373;
  assign n29375 = ~n28037 & n28157;
  assign n29376 = ~n28136 & ~n28161;
  assign n29377 = pi280 & n29376;
  assign n29378 = ~n28038 & n28134;
  assign n29379 = pi281 & ~n29378;
  assign n29380 = ~n29377 & ~n29379;
  assign n29381 = pi134 & ~n29380;
  assign n29382 = ~n29375 & ~n29381;
  assign n29383 = n29374 & n29382;
  assign n29384 = ~n29374 & ~n29382;
  assign n29385 = ~n29383 & ~n29384;
  assign n29386 = pi135 & pi281;
  assign n29387 = n28179 & ~n28185;
  assign n29388 = ~n28184 & ~n29387;
  assign n29389 = n29386 & ~n29388;
  assign n29390 = ~n28179 & ~n28184;
  assign n29391 = ~n28185 & ~n29390;
  assign n29392 = ~n29386 & ~n29391;
  assign n29393 = ~n29389 & ~n29392;
  assign n29394 = ~n29385 & ~n29393;
  assign n29395 = n29374 & ~n29382;
  assign n29396 = ~n29374 & n29382;
  assign n29397 = ~n29395 & ~n29396;
  assign n29398 = ~n29386 & ~n29388;
  assign n29399 = n29386 & ~n29391;
  assign n29400 = ~n29398 & ~n29399;
  assign n29401 = ~n29397 & ~n29400;
  assign n29402 = ~n29394 & ~n29401;
  assign n29403 = ~n29258 & n29402;
  assign n29404 = n29258 & ~n29402;
  assign n29405 = ~n29403 & ~n29404;
  assign n29406 = pi280 & ~n28186;
  assign n29407 = pi135 & n29406;
  assign n29408 = ~n28177 & ~n28179;
  assign n29409 = ~n29407 & ~n29408;
  assign n29410 = pi279 & ~n29409;
  assign n29411 = pi136 & n29410;
  assign n29412 = pi137 & pi279;
  assign n29413 = ~n28178 & ~n29408;
  assign n29414 = ~n29407 & n29413;
  assign n29415 = ~n28204 & ~n29414;
  assign n29416 = ~n29412 & ~n29415;
  assign n29417 = ~n29411 & n29416;
  assign n29418 = ~n29411 & ~n29415;
  assign n29419 = n29412 & ~n29418;
  assign n29420 = ~n29417 & ~n29419;
  assign n29421 = ~n29405 & ~n29420;
  assign n29422 = ~n29258 & ~n29402;
  assign n29423 = n29258 & n29402;
  assign n29424 = ~n29422 & ~n29423;
  assign n29425 = n29412 & ~n29415;
  assign n29426 = ~n29411 & n29425;
  assign n29427 = ~n29412 & ~n29418;
  assign n29428 = ~n29426 & ~n29427;
  assign n29429 = ~n29424 & ~n29428;
  assign n29430 = ~n29421 & ~n29429;
  assign n29431 = n28208 & ~n28250;
  assign n29432 = ~n28208 & n28250;
  assign n29433 = ~n28241 & ~n29432;
  assign n29434 = ~n29431 & ~n29433;
  assign n29435 = n29430 & ~n29434;
  assign n29436 = ~n29430 & n29434;
  assign n29437 = ~n29435 & ~n29436;
  assign n29438 = pi138 & pi278;
  assign n29439 = n28264 & ~n28270;
  assign n29440 = ~n28269 & ~n29439;
  assign n29441 = n29438 & ~n29440;
  assign n29442 = ~n28264 & ~n28269;
  assign n29443 = ~n28270 & ~n29442;
  assign n29444 = ~n29438 & ~n29443;
  assign n29445 = ~n29441 & ~n29444;
  assign n29446 = ~n29437 & ~n29445;
  assign n29447 = n29430 & n29434;
  assign n29448 = ~n29430 & ~n29434;
  assign n29449 = ~n29447 & ~n29448;
  assign n29450 = ~n29438 & ~n29440;
  assign n29451 = n29438 & ~n29443;
  assign n29452 = ~n29450 & ~n29451;
  assign n29453 = ~n29449 & ~n29452;
  assign n29454 = ~n29446 & ~n29453;
  assign n29455 = ~n29257 & ~n29454;
  assign n29456 = n29257 & n29454;
  assign n29457 = ~n29455 & ~n29456;
  assign n29458 = pi277 & ~n28271;
  assign n29459 = pi138 & n29458;
  assign n29460 = ~n28262 & ~n28264;
  assign n29461 = ~n28263 & ~n29460;
  assign n29462 = ~n29459 & n29461;
  assign n29463 = pi140 & pi276;
  assign n29464 = ~n29459 & ~n29460;
  assign n29465 = pi276 & ~n29464;
  assign n29466 = pi139 & n29465;
  assign n29467 = n28281 & ~n29466;
  assign n29468 = n29463 & ~n29467;
  assign n29469 = ~n29462 & n29468;
  assign n29470 = ~n29462 & ~n29467;
  assign n29471 = ~n29463 & ~n29470;
  assign n29472 = ~n29469 & ~n29471;
  assign n29473 = ~n29457 & ~n29472;
  assign n29474 = ~n29257 & n29454;
  assign n29475 = n29257 & ~n29454;
  assign n29476 = ~n29474 & ~n29475;
  assign n29477 = ~n29463 & ~n29467;
  assign n29478 = ~n29462 & n29477;
  assign n29479 = n29463 & ~n29470;
  assign n29480 = ~n29478 & ~n29479;
  assign n29481 = ~n29476 & ~n29480;
  assign n29482 = ~n29473 & ~n29481;
  assign n29483 = ~n28284 & ~n28285;
  assign n29484 = n28284 & n28285;
  assign n29485 = ~n28304 & ~n29484;
  assign n29486 = ~n29483 & ~n29485;
  assign n29487 = n29482 & n29486;
  assign n29488 = ~n29482 & ~n29486;
  assign n29489 = ~n29487 & ~n29488;
  assign n29490 = pi141 & pi275;
  assign n29491 = n28324 & ~n28330;
  assign n29492 = ~n28329 & ~n29491;
  assign n29493 = n29490 & ~n29492;
  assign n29494 = ~n28324 & ~n28329;
  assign n29495 = ~n28330 & ~n29494;
  assign n29496 = ~n29490 & ~n29495;
  assign n29497 = ~n29493 & ~n29496;
  assign n29498 = ~n29489 & ~n29497;
  assign n29499 = n29482 & ~n29486;
  assign n29500 = ~n29482 & n29486;
  assign n29501 = ~n29499 & ~n29500;
  assign n29502 = ~n29490 & ~n29492;
  assign n29503 = n29490 & ~n29495;
  assign n29504 = ~n29502 & ~n29503;
  assign n29505 = ~n29501 & ~n29504;
  assign n29506 = ~n29498 & ~n29505;
  assign n29507 = ~n29256 & ~n29506;
  assign n29508 = n29256 & n29506;
  assign n29509 = ~n29507 & ~n29508;
  assign n29510 = pi274 & ~n28331;
  assign n29511 = pi141 & n29510;
  assign n29512 = ~n28322 & ~n28324;
  assign n29513 = ~n28323 & ~n29512;
  assign n29514 = ~n29511 & n29513;
  assign n29515 = pi143 & pi273;
  assign n29516 = ~n29511 & ~n29512;
  assign n29517 = pi273 & ~n29516;
  assign n29518 = pi142 & n29517;
  assign n29519 = n28341 & ~n29518;
  assign n29520 = n29515 & ~n29519;
  assign n29521 = ~n29514 & n29520;
  assign n29522 = ~n29514 & ~n29519;
  assign n29523 = ~n29515 & ~n29522;
  assign n29524 = ~n29521 & ~n29523;
  assign n29525 = ~n29509 & ~n29524;
  assign n29526 = ~n29256 & n29506;
  assign n29527 = n29256 & ~n29506;
  assign n29528 = ~n29526 & ~n29527;
  assign n29529 = ~n29515 & ~n29519;
  assign n29530 = ~n29514 & n29529;
  assign n29531 = n29515 & ~n29522;
  assign n29532 = ~n29530 & ~n29531;
  assign n29533 = ~n29528 & ~n29532;
  assign n29534 = ~n29525 & ~n29533;
  assign n29535 = ~n28345 & ~n28370;
  assign n29536 = n28345 & n28370;
  assign n29537 = ~n28364 & ~n29536;
  assign n29538 = ~n29535 & ~n29537;
  assign n29539 = n29534 & ~n29538;
  assign n29540 = ~n29534 & n29538;
  assign n29541 = ~n29539 & ~n29540;
  assign n29542 = pi144 & pi272;
  assign n29543 = n28384 & ~n28389;
  assign n29544 = ~n28390 & ~n29543;
  assign n29545 = n29542 & ~n29544;
  assign n29546 = ~n28384 & ~n28390;
  assign n29547 = ~n28389 & ~n29546;
  assign n29548 = ~n29542 & ~n29547;
  assign n29549 = ~n29545 & ~n29548;
  assign n29550 = ~n29541 & ~n29549;
  assign n29551 = n29534 & n29538;
  assign n29552 = ~n29534 & ~n29538;
  assign n29553 = ~n29551 & ~n29552;
  assign n29554 = ~n29542 & ~n29544;
  assign n29555 = n29542 & ~n29547;
  assign n29556 = ~n29554 & ~n29555;
  assign n29557 = ~n29553 & ~n29556;
  assign n29558 = ~n29550 & ~n29557;
  assign n29559 = ~n29255 & n29558;
  assign n29560 = n29255 & ~n29558;
  assign n29561 = ~n29559 & ~n29560;
  assign n29562 = pi271 & ~n28391;
  assign n29563 = pi144 & n29562;
  assign n29564 = ~n28382 & ~n28384;
  assign n29565 = ~n29563 & ~n29564;
  assign n29566 = pi270 & ~n29565;
  assign n29567 = pi145 & n29566;
  assign n29568 = pi146 & pi270;
  assign n29569 = ~n28383 & ~n29564;
  assign n29570 = ~n29563 & n29569;
  assign n29571 = ~n28400 & ~n29570;
  assign n29572 = ~n29568 & ~n29571;
  assign n29573 = ~n29567 & n29572;
  assign n29574 = ~n29567 & ~n29571;
  assign n29575 = n29568 & ~n29574;
  assign n29576 = ~n29573 & ~n29575;
  assign n29577 = ~n29561 & ~n29576;
  assign n29578 = ~n29255 & ~n29558;
  assign n29579 = n29255 & n29558;
  assign n29580 = ~n29578 & ~n29579;
  assign n29581 = n29568 & ~n29571;
  assign n29582 = ~n29567 & n29581;
  assign n29583 = ~n29568 & ~n29574;
  assign n29584 = ~n29582 & ~n29583;
  assign n29585 = ~n29580 & ~n29584;
  assign n29586 = ~n29577 & ~n29585;
  assign n29587 = ~n28404 & ~n28429;
  assign n29588 = n28404 & n28429;
  assign n29589 = ~n28423 & ~n29588;
  assign n29590 = ~n29587 & ~n29589;
  assign n29591 = n29586 & ~n29590;
  assign n29592 = ~n29586 & n29590;
  assign n29593 = ~n29591 & ~n29592;
  assign n29594 = pi147 & pi269;
  assign n29595 = n28443 & ~n28448;
  assign n29596 = ~n28449 & ~n29595;
  assign n29597 = n29594 & ~n29596;
  assign n29598 = ~n28443 & ~n28449;
  assign n29599 = ~n28448 & ~n29598;
  assign n29600 = ~n29594 & ~n29599;
  assign n29601 = ~n29597 & ~n29600;
  assign n29602 = ~n29593 & ~n29601;
  assign n29603 = n29586 & n29590;
  assign n29604 = ~n29586 & ~n29590;
  assign n29605 = ~n29603 & ~n29604;
  assign n29606 = ~n29594 & ~n29596;
  assign n29607 = n29594 & ~n29599;
  assign n29608 = ~n29606 & ~n29607;
  assign n29609 = ~n29605 & ~n29608;
  assign n29610 = ~n29602 & ~n29609;
  assign n29611 = ~n29254 & n29610;
  assign n29612 = n29254 & ~n29610;
  assign n29613 = ~n29611 & ~n29612;
  assign n29614 = pi268 & ~n28450;
  assign n29615 = pi147 & n29614;
  assign n29616 = ~n28441 & ~n28443;
  assign n29617 = ~n29615 & ~n29616;
  assign n29618 = pi267 & ~n29617;
  assign n29619 = pi148 & n29618;
  assign n29620 = pi149 & pi267;
  assign n29621 = ~n28442 & ~n29616;
  assign n29622 = ~n29615 & n29621;
  assign n29623 = ~n28459 & ~n29622;
  assign n29624 = ~n29620 & ~n29623;
  assign n29625 = ~n29619 & n29624;
  assign n29626 = ~n29619 & ~n29623;
  assign n29627 = n29620 & ~n29626;
  assign n29628 = ~n29625 & ~n29627;
  assign n29629 = ~n29613 & ~n29628;
  assign n29630 = ~n29254 & ~n29610;
  assign n29631 = n29254 & n29610;
  assign n29632 = ~n29630 & ~n29631;
  assign n29633 = n29620 & ~n29623;
  assign n29634 = ~n29619 & n29633;
  assign n29635 = ~n29620 & ~n29626;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = ~n29632 & ~n29636;
  assign n29638 = ~n29629 & ~n29637;
  assign n29639 = n28463 & ~n28488;
  assign n29640 = ~n28463 & n28488;
  assign n29641 = ~n28479 & ~n29640;
  assign n29642 = ~n29639 & ~n29641;
  assign n29643 = n29638 & n29642;
  assign n29644 = ~n29638 & ~n29642;
  assign n29645 = ~n29643 & ~n29644;
  assign n29646 = pi150 & pi266;
  assign n29647 = n28502 & ~n28508;
  assign n29648 = ~n28507 & ~n29647;
  assign n29649 = n29646 & ~n29648;
  assign n29650 = ~n28502 & ~n28507;
  assign n29651 = ~n28508 & ~n29650;
  assign n29652 = ~n29646 & ~n29651;
  assign n29653 = ~n29649 & ~n29652;
  assign n29654 = ~n29645 & ~n29653;
  assign n29655 = n29638 & ~n29642;
  assign n29656 = ~n29638 & n29642;
  assign n29657 = ~n29655 & ~n29656;
  assign n29658 = ~n29646 & ~n29648;
  assign n29659 = n29646 & ~n29651;
  assign n29660 = ~n29658 & ~n29659;
  assign n29661 = ~n29657 & ~n29660;
  assign n29662 = ~n29654 & ~n29661;
  assign n29663 = ~n29253 & n29662;
  assign n29664 = n29253 & ~n29662;
  assign n29665 = ~n29663 & ~n29664;
  assign n29666 = pi265 & ~n28509;
  assign n29667 = pi150 & n29666;
  assign n29668 = ~n28500 & ~n28502;
  assign n29669 = ~n29667 & ~n29668;
  assign n29670 = pi264 & ~n29669;
  assign n29671 = pi151 & n29670;
  assign n29672 = pi152 & pi264;
  assign n29673 = ~n28501 & ~n29668;
  assign n29674 = ~n29667 & n29673;
  assign n29675 = ~n28518 & ~n29674;
  assign n29676 = ~n29672 & ~n29675;
  assign n29677 = ~n29671 & n29676;
  assign n29678 = ~n29671 & ~n29675;
  assign n29679 = n29672 & ~n29678;
  assign n29680 = ~n29677 & ~n29679;
  assign n29681 = ~n29665 & ~n29680;
  assign n29682 = ~n29253 & ~n29662;
  assign n29683 = n29253 & n29662;
  assign n29684 = ~n29682 & ~n29683;
  assign n29685 = n29672 & ~n29675;
  assign n29686 = ~n29671 & n29685;
  assign n29687 = ~n29672 & ~n29678;
  assign n29688 = ~n29686 & ~n29687;
  assign n29689 = ~n29684 & ~n29688;
  assign n29690 = ~n29681 & ~n29689;
  assign n29691 = n28522 & ~n28547;
  assign n29692 = ~n28522 & n28547;
  assign n29693 = ~n28538 & ~n29692;
  assign n29694 = ~n29691 & ~n29693;
  assign n29695 = n29690 & ~n29694;
  assign n29696 = ~n29690 & n29694;
  assign n29697 = ~n29695 & ~n29696;
  assign n29698 = pi153 & pi263;
  assign n29699 = ~n28558 & n28562;
  assign n29700 = ~n28557 & ~n29699;
  assign n29701 = n29698 & ~n29700;
  assign n29702 = ~n28557 & ~n28562;
  assign n29703 = ~n28558 & ~n29702;
  assign n29704 = ~n29698 & ~n29703;
  assign n29705 = ~n29701 & ~n29704;
  assign n29706 = ~n29697 & ~n29705;
  assign n29707 = n29690 & n29694;
  assign n29708 = ~n29690 & ~n29694;
  assign n29709 = ~n29707 & ~n29708;
  assign n29710 = ~n29698 & ~n29700;
  assign n29711 = n29698 & ~n29703;
  assign n29712 = ~n29710 & ~n29711;
  assign n29713 = ~n29709 & ~n29712;
  assign n29714 = ~n29706 & ~n29713;
  assign n29715 = ~n29252 & ~n29714;
  assign n29716 = n29252 & n29714;
  assign n29717 = ~n29715 & ~n29716;
  assign n29718 = pi155 & pi261;
  assign n29719 = n28015 & ~n28569;
  assign n29720 = n29718 & ~n29719;
  assign n29721 = ~n28572 & n29720;
  assign n29722 = ~n28572 & ~n29719;
  assign n29723 = ~n29718 & ~n29722;
  assign n29724 = ~n29721 & ~n29723;
  assign n29725 = ~n29717 & ~n29724;
  assign n29726 = ~n29252 & n29714;
  assign n29727 = n29252 & ~n29714;
  assign n29728 = ~n29726 & ~n29727;
  assign n29729 = ~n29718 & ~n29719;
  assign n29730 = ~n28572 & n29729;
  assign n29731 = n29718 & ~n29722;
  assign n29732 = ~n29730 & ~n29731;
  assign n29733 = ~n29728 & ~n29732;
  assign n29734 = ~n29725 & ~n29733;
  assign n29735 = pi260 & ~n28022;
  assign n29736 = pi155 & n29735;
  assign n29737 = n28022 & ~n28576;
  assign n29738 = n28015 & ~n28572;
  assign n29739 = ~n28569 & n29738;
  assign n29740 = ~n28015 & ~n28573;
  assign n29741 = ~n29739 & ~n29740;
  assign n29742 = ~n29737 & ~n29741;
  assign n29743 = ~n29736 & ~n29742;
  assign n29744 = n29734 & n29743;
  assign n29745 = ~n29734 & ~n29743;
  assign n29746 = ~n29744 & ~n29745;
  assign n29747 = pi156 & pi259;
  assign n29748 = ~n28603 & ~n29747;
  assign n29749 = pi156 & pi260;
  assign n29750 = pi259 & n28603;
  assign n29751 = ~n28588 & ~n29750;
  assign n29752 = ~n29749 & ~n29751;
  assign n29753 = ~n29748 & n29752;
  assign n29754 = ~n29748 & ~n29751;
  assign n29755 = n29749 & ~n29754;
  assign n29756 = ~n29753 & ~n29755;
  assign n29757 = ~n29746 & ~n29756;
  assign n29758 = n29734 & ~n29743;
  assign n29759 = ~n29734 & n29743;
  assign n29760 = ~n29758 & ~n29759;
  assign n29761 = n29749 & ~n29751;
  assign n29762 = ~n29748 & n29761;
  assign n29763 = ~n29749 & ~n29754;
  assign n29764 = ~n29762 & ~n29763;
  assign n29765 = ~n29760 & ~n29764;
  assign n29766 = ~n29757 & ~n29765;
  assign n29767 = ~n26683 & ~n28590;
  assign n29768 = n26683 & n28590;
  assign n29769 = ~n28588 & n28607;
  assign n29770 = n28588 & ~n28607;
  assign n29771 = ~n29769 & ~n29770;
  assign n29772 = pi258 & ~n29771;
  assign n29773 = pi157 & n29772;
  assign n29774 = ~n28588 & ~n28607;
  assign n29775 = n28588 & n28607;
  assign n29776 = ~n29774 & ~n29775;
  assign n29777 = ~n28613 & ~n29776;
  assign n29778 = ~n29773 & ~n29777;
  assign n29779 = ~n29768 & ~n29778;
  assign n29780 = ~n29767 & ~n29779;
  assign n29781 = n29766 & n29780;
  assign n29782 = ~n29766 & ~n29780;
  assign n29783 = ~n29781 & ~n29782;
  assign n29784 = pi158 & pi258;
  assign n29785 = pi157 & pi259;
  assign n29786 = ~n29784 & ~n29785;
  assign n29787 = n29784 & n29785;
  assign n29788 = ~n29786 & ~n29787;
  assign n29789 = ~n29748 & ~n29750;
  assign n29790 = ~n28588 & n29789;
  assign n29791 = n28588 & ~n29789;
  assign n29792 = ~n29790 & ~n29791;
  assign n29793 = pi258 & ~n29792;
  assign n29794 = pi157 & n29793;
  assign n29795 = ~n28613 & ~n29792;
  assign n29796 = ~n28588 & ~n29789;
  assign n29797 = n28588 & n29789;
  assign n29798 = ~n29796 & ~n29797;
  assign n29799 = pi258 & ~n29798;
  assign n29800 = pi157 & n29799;
  assign n29801 = ~n29795 & ~n29800;
  assign n29802 = n29794 & ~n29801;
  assign n29803 = ~n29794 & n29801;
  assign n29804 = ~n29802 & ~n29803;
  assign n29805 = ~n29788 & ~n29804;
  assign n29806 = n29784 & ~n29785;
  assign n29807 = ~n29784 & n29785;
  assign n29808 = ~n29806 & ~n29807;
  assign n29809 = ~n29794 & ~n29801;
  assign n29810 = n29794 & n29801;
  assign n29811 = ~n29809 & ~n29810;
  assign n29812 = ~n29808 & ~n29811;
  assign n29813 = ~n29805 & ~n29812;
  assign n29814 = ~n29783 & ~n29813;
  assign n29815 = n29766 & ~n29780;
  assign n29816 = ~n29766 & n29780;
  assign n29817 = ~n29815 & ~n29816;
  assign n29818 = ~n29804 & ~n29808;
  assign n29819 = ~n29788 & ~n29811;
  assign n29820 = ~n29818 & ~n29819;
  assign n29821 = ~n29817 & ~n29820;
  assign n29822 = ~n29814 & ~n29821;
  assign n29823 = pi322 & n29822;
  assign n29824 = ~n29251 & ~n29823;
  assign n29825 = n28628 & n29822;
  assign n29826 = n1445 & n29825;
  assign n29827 = ~n29824 & ~n29826;
  assign n29828 = ~n29250 & ~n29827;
  assign n29829 = ~n29241 & n29247;
  assign n29830 = n29241 & ~n29247;
  assign n29831 = ~n29829 & ~n29830;
  assign n29832 = ~n29251 & n29822;
  assign n29833 = pi322 & n29832;
  assign n29834 = n28628 & ~n29823;
  assign n29835 = pi323 & n29834;
  assign n29836 = ~n29833 & ~n29835;
  assign n29837 = ~n29831 & ~n29836;
  assign n29838 = ~n29828 & ~n29837;
  assign n29839 = n28002 & ~n28648;
  assign n29840 = ~n28004 & ~n28629;
  assign n29841 = n28004 & n28628;
  assign n29842 = pi322 & n29841;
  assign n29843 = ~n29840 & ~n29842;
  assign n29844 = ~n28011 & ~n29843;
  assign n29845 = n28004 & ~n28629;
  assign n29846 = ~n28004 & n28628;
  assign n29847 = pi322 & n29846;
  assign n29848 = ~n29845 & ~n29847;
  assign n29849 = n28010 & ~n29848;
  assign n29850 = pi323 & n29849;
  assign n29851 = ~n29844 & ~n29850;
  assign n29852 = ~n28002 & n28648;
  assign n29853 = ~n29851 & ~n29852;
  assign n29854 = ~n29839 & ~n29853;
  assign n29855 = n29838 & ~n29854;
  assign n29856 = ~n29838 & n29854;
  assign n29857 = ~n29855 & ~n29856;
  assign n29858 = pi326 & n26706;
  assign n29859 = pi325 & n26175;
  assign n29860 = n29858 & n29859;
  assign n29861 = ~n29858 & ~n29859;
  assign n29862 = ~n29860 & ~n29861;
  assign n29863 = ~n29857 & ~n29862;
  assign n29864 = ~n29838 & ~n29854;
  assign n29865 = n29838 & n29854;
  assign n29866 = ~n29864 & ~n29865;
  assign n29867 = ~n29858 & n29859;
  assign n29868 = n29858 & ~n29859;
  assign n29869 = ~n29867 & ~n29868;
  assign n29870 = ~n29866 & ~n29869;
  assign n29871 = ~n29863 & ~n29870;
  assign n29872 = ~n29240 & ~n29871;
  assign n29873 = n29217 & ~n29237;
  assign n29874 = ~n29217 & n29237;
  assign n29875 = ~n29873 & ~n29874;
  assign n29876 = ~n29862 & ~n29866;
  assign n29877 = ~n29857 & ~n29869;
  assign n29878 = ~n29876 & ~n29877;
  assign n29879 = ~n29875 & ~n29878;
  assign n29880 = ~n29872 & ~n29879;
  assign n29881 = ~n29213 & n29880;
  assign n29882 = n29213 & ~n29880;
  assign n29883 = ~n29881 & ~n29882;
  assign n29884 = pi329 & n19557;
  assign n29885 = pi328 & n19970;
  assign n29886 = n29884 & n29885;
  assign n29887 = ~n29884 & ~n29885;
  assign n29888 = ~n29886 & ~n29887;
  assign n29889 = ~n29883 & ~n29888;
  assign n29890 = n29213 & n29880;
  assign n29891 = ~n29213 & ~n29880;
  assign n29892 = ~n29890 & ~n29891;
  assign n29893 = ~n29884 & n29885;
  assign n29894 = n29884 & ~n29885;
  assign n29895 = ~n29893 & ~n29894;
  assign n29896 = ~n29892 & ~n29895;
  assign n29897 = ~n29889 & ~n29896;
  assign n29898 = ~n29212 & ~n29897;
  assign n29899 = ~n29196 & ~n29209;
  assign n29900 = n29196 & n29209;
  assign n29901 = ~n29899 & ~n29900;
  assign n29902 = ~n29888 & ~n29892;
  assign n29903 = ~n29883 & ~n29895;
  assign n29904 = ~n29902 & ~n29903;
  assign n29905 = ~n29901 & ~n29904;
  assign n29906 = ~n29898 & ~n29905;
  assign n29907 = ~n29192 & ~n29906;
  assign n29908 = n29192 & n29906;
  assign n29909 = ~n29907 & ~n29908;
  assign n29910 = n18461 & ~n29909;
  assign n29911 = pi331 & n29910;
  assign n29912 = pi331 & n18461;
  assign n29913 = n29192 & ~n29906;
  assign n29914 = ~n29192 & n29906;
  assign n29915 = ~n29913 & ~n29914;
  assign n29916 = ~n29912 & ~n29915;
  assign n29917 = ~n29911 & ~n29916;
  assign n29918 = ~n29176 & ~n29917;
  assign n29919 = n29160 & n29173;
  assign n29920 = ~n29160 & ~n29173;
  assign n29921 = ~n29919 & ~n29920;
  assign n29922 = n18461 & ~n29915;
  assign n29923 = pi331 & n29922;
  assign n29924 = ~n29909 & ~n29912;
  assign n29925 = ~n29923 & ~n29924;
  assign n29926 = ~n29921 & ~n29925;
  assign n29927 = ~n29918 & ~n29926;
  assign n29928 = ~n28725 & n28729;
  assign n29929 = ~n28721 & ~n28740;
  assign n29930 = n28721 & n28740;
  assign n29931 = ~n29929 & ~n29930;
  assign n29932 = n28725 & ~n28729;
  assign n29933 = ~n29931 & ~n29932;
  assign n29934 = ~n29928 & ~n29933;
  assign n29935 = n29927 & n29934;
  assign n29936 = ~n29927 & ~n29934;
  assign n29937 = ~n29935 & ~n29936;
  assign n29938 = pi333 & n12917;
  assign n29939 = ~n28721 & ~n28735;
  assign n29940 = n28721 & n28735;
  assign n29941 = ~n12917 & ~n29940;
  assign n29942 = ~n29939 & ~n29941;
  assign n29943 = n13762 & ~n29942;
  assign n29944 = ~n13762 & ~n29939;
  assign n29945 = n12917 & n29944;
  assign n29946 = ~n29943 & ~n29945;
  assign n29947 = pi332 & ~n29946;
  assign n29948 = pi332 & n13762;
  assign n29949 = n28721 & ~n29948;
  assign n29950 = n28735 & n29949;
  assign n29951 = ~n29947 & ~n29950;
  assign n29952 = ~n29938 & n29951;
  assign n29953 = n29938 & ~n29951;
  assign n29954 = ~n29952 & ~n29953;
  assign n29955 = pi334 & n11711;
  assign n29956 = ~n28743 & ~n28765;
  assign n29957 = ~n28772 & n29956;
  assign n29958 = ~n28763 & ~n28765;
  assign n29959 = ~n28728 & n29958;
  assign n29960 = ~n28764 & ~n29959;
  assign n29961 = ~n29957 & n29960;
  assign n29962 = n29955 & ~n29961;
  assign n29963 = ~n29955 & n29961;
  assign n29964 = ~n29962 & ~n29963;
  assign n29965 = ~n29954 & ~n29964;
  assign n29966 = n29938 & n29951;
  assign n29967 = ~n29938 & ~n29951;
  assign n29968 = ~n29966 & ~n29967;
  assign n29969 = ~n29955 & ~n29961;
  assign n29970 = n29955 & n29961;
  assign n29971 = ~n29969 & ~n29970;
  assign n29972 = ~n29968 & ~n29971;
  assign n29973 = ~n29965 & ~n29972;
  assign n29974 = ~n29937 & ~n29973;
  assign n29975 = n29927 & ~n29934;
  assign n29976 = ~n29927 & n29934;
  assign n29977 = ~n29975 & ~n29976;
  assign n29978 = ~n29964 & ~n29968;
  assign n29979 = ~n29954 & ~n29971;
  assign n29980 = ~n29978 & ~n29979;
  assign n29981 = ~n29977 & ~n29980;
  assign n29982 = ~n29974 & ~n29981;
  assign n29983 = ~n29145 & n29982;
  assign n29984 = n29145 & ~n29982;
  assign n29985 = ~n29983 & ~n29984;
  assign n29986 = pi337 & n10561;
  assign n29987 = pi336 & n11366;
  assign n29988 = ~n28782 & n28784;
  assign n29989 = ~n29987 & ~n29988;
  assign n29990 = n27911 & n29989;
  assign n29991 = n28782 & ~n28784;
  assign n29992 = n29987 & ~n29991;
  assign n29993 = ~n27911 & n29992;
  assign n29994 = ~n29990 & ~n29993;
  assign n29995 = ~n29134 & ~n29994;
  assign n29996 = n27911 & n29992;
  assign n29997 = ~n27911 & n29989;
  assign n29998 = ~n29996 & ~n29997;
  assign n29999 = ~n29124 & ~n29998;
  assign n30000 = ~n28784 & ~n29987;
  assign n30001 = n28782 & n30000;
  assign n30002 = n28784 & n29987;
  assign n30003 = ~n28782 & n30002;
  assign n30004 = ~n30001 & ~n30003;
  assign n30005 = ~n29999 & n30004;
  assign n30006 = ~n29995 & n30005;
  assign n30007 = n29986 & ~n30006;
  assign n30008 = ~n29986 & n30006;
  assign n30009 = ~n30007 & ~n30008;
  assign n30010 = ~n29985 & ~n30009;
  assign n30011 = n29145 & n29982;
  assign n30012 = ~n29145 & ~n29982;
  assign n30013 = ~n30011 & ~n30012;
  assign n30014 = ~n29986 & ~n30006;
  assign n30015 = n29986 & n30006;
  assign n30016 = ~n30014 & ~n30015;
  assign n30017 = ~n30013 & ~n30016;
  assign n30018 = ~n30010 & ~n30017;
  assign n30019 = ~n29144 & ~n30018;
  assign n30020 = ~n29121 & ~n29141;
  assign n30021 = n29121 & n29141;
  assign n30022 = ~n30020 & ~n30021;
  assign n30023 = ~n30009 & ~n30013;
  assign n30024 = ~n29985 & ~n30016;
  assign n30025 = ~n30023 & ~n30024;
  assign n30026 = ~n30022 & ~n30025;
  assign n30027 = ~n30019 & ~n30026;
  assign n30028 = ~n28814 & n28818;
  assign n30029 = ~n28810 & ~n28829;
  assign n30030 = n28810 & n28829;
  assign n30031 = ~n30029 & ~n30030;
  assign n30032 = n28814 & ~n28818;
  assign n30033 = ~n30031 & ~n30032;
  assign n30034 = ~n30028 & ~n30033;
  assign n30035 = n30027 & n30034;
  assign n30036 = ~n30027 & ~n30034;
  assign n30037 = ~n30035 & ~n30036;
  assign n30038 = pi339 & n6556;
  assign n30039 = ~n28810 & ~n28824;
  assign n30040 = n28810 & n28824;
  assign n30041 = ~n6556 & ~n30040;
  assign n30042 = ~n30039 & ~n30041;
  assign n30043 = n9205 & ~n30042;
  assign n30044 = ~n9205 & ~n30039;
  assign n30045 = n6556 & n30044;
  assign n30046 = ~n30043 & ~n30045;
  assign n30047 = pi338 & ~n30046;
  assign n30048 = pi338 & n9205;
  assign n30049 = n28810 & ~n30048;
  assign n30050 = n28824 & n30049;
  assign n30051 = ~n30047 & ~n30050;
  assign n30052 = ~n30038 & n30051;
  assign n30053 = n30038 & ~n30051;
  assign n30054 = ~n30052 & ~n30053;
  assign n30055 = pi340 & n5973;
  assign n30056 = ~n28832 & ~n28854;
  assign n30057 = ~n28861 & n30056;
  assign n30058 = ~n28852 & ~n28854;
  assign n30059 = ~n28817 & n30058;
  assign n30060 = ~n28853 & ~n30059;
  assign n30061 = ~n30057 & n30060;
  assign n30062 = n30055 & ~n30061;
  assign n30063 = ~n30055 & n30061;
  assign n30064 = ~n30062 & ~n30063;
  assign n30065 = ~n30054 & ~n30064;
  assign n30066 = n30038 & n30051;
  assign n30067 = ~n30038 & ~n30051;
  assign n30068 = ~n30066 & ~n30067;
  assign n30069 = ~n30055 & ~n30061;
  assign n30070 = n30055 & n30061;
  assign n30071 = ~n30069 & ~n30070;
  assign n30072 = ~n30068 & ~n30071;
  assign n30073 = ~n30065 & ~n30072;
  assign n30074 = ~n30037 & ~n30073;
  assign n30075 = n30027 & ~n30034;
  assign n30076 = ~n30027 & n30034;
  assign n30077 = ~n30075 & ~n30076;
  assign n30078 = ~n30064 & ~n30068;
  assign n30079 = ~n30054 & ~n30071;
  assign n30080 = ~n30078 & ~n30079;
  assign n30081 = ~n30077 & ~n30080;
  assign n30082 = ~n30074 & ~n30081;
  assign n30083 = ~n29117 & n30082;
  assign n30084 = n29117 & ~n30082;
  assign n30085 = ~n30083 & ~n30084;
  assign n30086 = pi343 & n5257;
  assign n30087 = pi342 & n5714;
  assign n30088 = ~n28871 & n28873;
  assign n30089 = ~n30087 & ~n30088;
  assign n30090 = n27872 & n30089;
  assign n30091 = n28871 & ~n28873;
  assign n30092 = n30087 & ~n30091;
  assign n30093 = ~n27872 & n30092;
  assign n30094 = ~n30090 & ~n30093;
  assign n30095 = ~n29106 & ~n30094;
  assign n30096 = n27872 & n30092;
  assign n30097 = ~n27872 & n30089;
  assign n30098 = ~n30096 & ~n30097;
  assign n30099 = ~n29096 & ~n30098;
  assign n30100 = ~n28873 & ~n30087;
  assign n30101 = n28871 & n30100;
  assign n30102 = n28873 & n30087;
  assign n30103 = ~n28871 & n30102;
  assign n30104 = ~n30101 & ~n30103;
  assign n30105 = ~n30099 & n30104;
  assign n30106 = ~n30095 & n30105;
  assign n30107 = n30086 & ~n30106;
  assign n30108 = ~n30086 & n30106;
  assign n30109 = ~n30107 & ~n30108;
  assign n30110 = ~n30085 & ~n30109;
  assign n30111 = n29117 & n30082;
  assign n30112 = ~n29117 & ~n30082;
  assign n30113 = ~n30111 & ~n30112;
  assign n30114 = ~n30086 & ~n30106;
  assign n30115 = n30086 & n30106;
  assign n30116 = ~n30114 & ~n30115;
  assign n30117 = ~n30113 & ~n30116;
  assign n30118 = ~n30110 & ~n30117;
  assign n30119 = ~n29116 & ~n30118;
  assign n30120 = ~n29093 & ~n29113;
  assign n30121 = n29093 & n29113;
  assign n30122 = ~n30120 & ~n30121;
  assign n30123 = ~n30109 & ~n30113;
  assign n30124 = ~n30085 & ~n30116;
  assign n30125 = ~n30123 & ~n30124;
  assign n30126 = ~n30122 & ~n30125;
  assign n30127 = ~n30119 & ~n30126;
  assign n30128 = ~n28903 & n28907;
  assign n30129 = ~n28899 & ~n28918;
  assign n30130 = n28899 & n28918;
  assign n30131 = ~n30129 & ~n30130;
  assign n30132 = n28903 & ~n28907;
  assign n30133 = ~n30131 & ~n30132;
  assign n30134 = ~n30128 & ~n30133;
  assign n30135 = n30127 & n30134;
  assign n30136 = ~n30127 & ~n30134;
  assign n30137 = ~n30135 & ~n30136;
  assign n30138 = pi345 & n2887;
  assign n30139 = ~n28899 & ~n28913;
  assign n30140 = n28899 & n28913;
  assign n30141 = ~n2887 & ~n30140;
  assign n30142 = ~n30139 & ~n30141;
  assign n30143 = n4596 & ~n30142;
  assign n30144 = ~n4596 & ~n30139;
  assign n30145 = n2887 & n30144;
  assign n30146 = ~n30143 & ~n30145;
  assign n30147 = pi344 & ~n30146;
  assign n30148 = pi344 & n4596;
  assign n30149 = n28899 & ~n30148;
  assign n30150 = n28913 & n30149;
  assign n30151 = ~n30147 & ~n30150;
  assign n30152 = ~n30138 & n30151;
  assign n30153 = n30138 & ~n30151;
  assign n30154 = ~n30152 & ~n30153;
  assign n30155 = pi346 & n2464;
  assign n30156 = n26020 & ~n27797;
  assign n30157 = ~n26020 & ~n27806;
  assign n30158 = ~n30156 & ~n30157;
  assign n30159 = ~n28930 & ~n30158;
  assign n30160 = ~n28933 & ~n30159;
  assign n30161 = n28923 & ~n30160;
  assign n30162 = ~n28921 & ~n30161;
  assign n30163 = ~n28964 & n30162;
  assign n30164 = ~n28923 & n30160;
  assign n30165 = ~n28955 & ~n30161;
  assign n30166 = ~n28906 & n30165;
  assign n30167 = ~n30164 & ~n30166;
  assign n30168 = ~n30163 & n30167;
  assign n30169 = n30155 & ~n30168;
  assign n30170 = ~n30155 & n30168;
  assign n30171 = ~n30169 & ~n30170;
  assign n30172 = ~n30154 & ~n30171;
  assign n30173 = n30138 & n30151;
  assign n30174 = ~n30138 & ~n30151;
  assign n30175 = ~n30173 & ~n30174;
  assign n30176 = ~n30155 & ~n30168;
  assign n30177 = n30155 & n30168;
  assign n30178 = ~n30176 & ~n30177;
  assign n30179 = ~n30175 & ~n30178;
  assign n30180 = ~n30172 & ~n30179;
  assign n30181 = ~n30137 & ~n30180;
  assign n30182 = n30127 & ~n30134;
  assign n30183 = ~n30127 & n30134;
  assign n30184 = ~n30182 & ~n30183;
  assign n30185 = ~n30171 & ~n30175;
  assign n30186 = ~n30154 & ~n30178;
  assign n30187 = ~n30185 & ~n30186;
  assign n30188 = ~n30184 & ~n30187;
  assign n30189 = ~n30181 & ~n30188;
  assign n30190 = ~n29089 & n30189;
  assign n30191 = n29089 & ~n30189;
  assign n30192 = ~n30190 & ~n30191;
  assign n30193 = pi349 & n1442;
  assign n30194 = ~pi348 & ~n27828;
  assign n30195 = n27828 & ~n27831;
  assign n30196 = ~n1729 & ~n30195;
  assign n30197 = ~n30194 & ~n30196;
  assign n30198 = ~n29078 & ~n30197;
  assign n30199 = ~n1729 & ~n27828;
  assign n30200 = n1442 & n30199;
  assign n30201 = ~n1442 & n27828;
  assign n30202 = n1442 & ~n27828;
  assign n30203 = ~n29074 & ~n30202;
  assign n30204 = ~n30201 & ~n30203;
  assign n30205 = n1729 & ~n30204;
  assign n30206 = ~n30200 & ~n30205;
  assign n30207 = pi348 & ~n30206;
  assign n30208 = ~n30198 & ~n30207;
  assign n30209 = n30193 & ~n30208;
  assign n30210 = ~n30193 & n30208;
  assign n30211 = ~n30209 & ~n30210;
  assign n30212 = ~n30192 & ~n30211;
  assign n30213 = n29089 & n30189;
  assign n30214 = ~n29089 & ~n30189;
  assign n30215 = ~n30213 & ~n30214;
  assign n30216 = ~n30193 & ~n30208;
  assign n30217 = n30193 & n30208;
  assign n30218 = ~n30216 & ~n30217;
  assign n30219 = ~n30215 & ~n30218;
  assign n30220 = ~n30212 & ~n30219;
  assign n30221 = ~n29088 & ~n30220;
  assign n30222 = ~n29071 & ~n29085;
  assign n30223 = n29071 & n29085;
  assign n30224 = ~n30222 & ~n30223;
  assign n30225 = ~n30211 & ~n30215;
  assign n30226 = ~n30192 & ~n30218;
  assign n30227 = ~n30225 & ~n30226;
  assign n30228 = ~n30224 & ~n30227;
  assign n30229 = ~n30221 & ~n30228;
  assign n30230 = ~n29050 & ~n30229;
  assign n30231 = n29050 & n30229;
  assign n30232 = ~n30230 & ~n30231;
  assign n30233 = pi258 & ~n29016;
  assign n30234 = pi128 & n30233;
  assign n30235 = pi351 & n30234;
  assign n30236 = pi351 & ~n1154;
  assign n30237 = ~n30235 & ~n30236;
  assign n30238 = n30235 & n30236;
  assign n30239 = ~n30237 & ~n30238;
  assign n30240 = n1156 & ~n30239;
  assign n30241 = pi352 & n30240;
  assign n30242 = pi352 & n1156;
  assign n30243 = n30235 & ~n30236;
  assign n30244 = ~n30235 & n30236;
  assign n30245 = ~n30243 & ~n30244;
  assign n30246 = ~n30242 & ~n30245;
  assign n30247 = ~n30241 & ~n30246;
  assign n30248 = ~n30232 & ~n30247;
  assign n30249 = ~n29050 & n30229;
  assign n30250 = n29050 & ~n30229;
  assign n30251 = ~n30249 & ~n30250;
  assign n30252 = n1156 & ~n30245;
  assign n30253 = pi352 & n30252;
  assign n30254 = ~n30239 & ~n30242;
  assign n30255 = ~n30253 & ~n30254;
  assign n30256 = ~n30251 & ~n30255;
  assign n30257 = ~n30248 & ~n30256;
  assign n30258 = ~n29022 & ~n29029;
  assign n30259 = n29022 & n29029;
  assign n30260 = n27788 & ~n30259;
  assign n30261 = ~n30258 & ~n30260;
  assign n30262 = n30257 & n30261;
  assign n30263 = ~n30257 & ~n30261;
  assign n30264 = ~n30262 & ~n30263;
  assign n30265 = pi130 & pi293;
  assign n30266 = ~pi129 & ~n30265;
  assign n30267 = pi293 & ~n12284;
  assign n30268 = ~n1514 & n30267;
  assign n30269 = n27777 & ~n30268;
  assign n30270 = ~n30266 & ~n30269;
  assign n30271 = n27169 & ~n30270;
  assign n30272 = ~pi130 & n27777;
  assign n30273 = ~pi129 & n30272;
  assign n30274 = pi130 & ~n27777;
  assign n30275 = pi129 & n30274;
  assign n30276 = ~n30273 & ~n30275;
  assign n30277 = pi128 & ~n30276;
  assign n30278 = ~n27169 & n27777;
  assign n30279 = pi130 & n30278;
  assign n30280 = ~pi130 & ~n27777;
  assign n30281 = pi129 & n30280;
  assign n30282 = ~n30279 & ~n30281;
  assign n30283 = ~pi128 & ~n30282;
  assign n30284 = pi129 & n27777;
  assign n30285 = ~pi129 & ~n27777;
  assign n30286 = ~n30284 & ~n30285;
  assign n30287 = ~n27169 & ~n30286;
  assign n30288 = pi130 & n30287;
  assign n30289 = ~n30283 & ~n30288;
  assign n30290 = ~n30277 & n30289;
  assign n30291 = pi293 & ~n30290;
  assign n30292 = ~n30271 & ~n30291;
  assign n30293 = n25357 & n25957;
  assign n30294 = ~n25357 & ~n25957;
  assign n30295 = ~n25362 & ~n30294;
  assign n30296 = ~n30293 & ~n30295;
  assign n30297 = n27742 & ~n30296;
  assign n30298 = pi297 & n2183;
  assign n30299 = n27696 & ~n27704;
  assign n30300 = n25367 & n25923;
  assign n30301 = n25365 & ~n30300;
  assign n30302 = ~n27176 & ~n30301;
  assign n30303 = ~n30299 & ~n30302;
  assign n30304 = ~n27705 & ~n30303;
  assign n30305 = ~n30298 & ~n30304;
  assign n30306 = ~n25365 & ~n27176;
  assign n30307 = ~n30300 & ~n30306;
  assign n30308 = ~n27705 & ~n30307;
  assign n30309 = ~n30299 & ~n30308;
  assign n30310 = n30298 & ~n30309;
  assign n30311 = ~n30305 & ~n30310;
  assign n30312 = n27525 & n27557;
  assign n30313 = pi305 & n27521;
  assign n30314 = n17127 & n30313;
  assign n30315 = pi305 & ~n17124;
  assign n30316 = ~n27521 & ~n30315;
  assign n30317 = ~n30314 & ~n30316;
  assign n30318 = ~n27536 & ~n30317;
  assign n30319 = ~n6777 & ~n27521;
  assign n30320 = ~n27547 & ~n30319;
  assign n30321 = ~n25769 & ~n30320;
  assign n30322 = n27535 & n30321;
  assign n30323 = n6777 & ~n27521;
  assign n30324 = ~n6777 & n27521;
  assign n30325 = ~n30323 & ~n30324;
  assign n30326 = n5463 & ~n30325;
  assign n30327 = pi305 & n30326;
  assign n30328 = n25769 & n30327;
  assign n30329 = ~n5463 & ~n25769;
  assign n30330 = n6777 & ~n30329;
  assign n30331 = ~n27521 & n30330;
  assign n30332 = n17136 & n27521;
  assign n30333 = ~n30331 & ~n30332;
  assign n30334 = pi305 & ~n30333;
  assign n30335 = n25769 & n27522;
  assign n30336 = ~n30334 & ~n30335;
  assign n30337 = ~n27535 & ~n30336;
  assign n30338 = ~n30328 & ~n30337;
  assign n30339 = ~n30322 & n30338;
  assign n30340 = ~n30318 & n30339;
  assign n30341 = ~n27525 & ~n27557;
  assign n30342 = n30340 & ~n30341;
  assign n30343 = ~n30312 & ~n30342;
  assign n30344 = n25830 & n27604;
  assign n30345 = ~n25843 & ~n27579;
  assign n30346 = n3552 & n30345;
  assign n30347 = ~n25842 & ~n27577;
  assign n30348 = n4086 & ~n30347;
  assign n30349 = ~n30346 & ~n30348;
  assign n30350 = pi302 & ~n30349;
  assign n30351 = ~n30344 & ~n30350;
  assign n30352 = ~n30343 & n30351;
  assign n30353 = n30343 & ~n30351;
  assign n30354 = ~n30352 & ~n30353;
  assign n30355 = ~n25819 & n25825;
  assign n30356 = n25819 & ~n25825;
  assign n30357 = n25396 & ~n30356;
  assign n30358 = ~n30355 & ~n30357;
  assign n30359 = n27561 & ~n30358;
  assign n30360 = ~n27561 & n30358;
  assign n30361 = ~n27572 & ~n30360;
  assign n30362 = ~n30359 & ~n30361;
  assign n30363 = pi303 & n5463;
  assign n30364 = ~n30362 & ~n30363;
  assign n30365 = n5463 & n30362;
  assign n30366 = pi303 & n30365;
  assign n30367 = ~n30364 & ~n30366;
  assign n30368 = n25769 & ~n27546;
  assign n30369 = n5463 & ~n30319;
  assign n30370 = pi305 & n30369;
  assign n30371 = ~n30368 & ~n30370;
  assign n30372 = ~n27535 & ~n30371;
  assign n30373 = n6777 & n27521;
  assign n30374 = n25769 & n30369;
  assign n30375 = ~n30373 & ~n30374;
  assign n30376 = pi305 & ~n30375;
  assign n30377 = ~n30372 & ~n30376;
  assign n30378 = n27437 & n27469;
  assign n30379 = n25409 & ~n25689;
  assign n30380 = ~n25409 & n25689;
  assign n30381 = ~n27447 & ~n30380;
  assign n30382 = ~n30379 & ~n30381;
  assign n30383 = ~n27433 & ~n30382;
  assign n30384 = n27433 & n30382;
  assign n30385 = ~n30383 & ~n30384;
  assign n30386 = n27179 & ~n30385;
  assign n30387 = ~n27433 & n30382;
  assign n30388 = n27433 & ~n30382;
  assign n30389 = ~n30387 & ~n30388;
  assign n30390 = ~n27179 & ~n30389;
  assign n30391 = ~n30386 & ~n30390;
  assign n30392 = ~n27437 & ~n27469;
  assign n30393 = ~n30391 & ~n30392;
  assign n30394 = ~n30378 & ~n30393;
  assign n30395 = ~n25758 & ~n27489;
  assign n30396 = ~n25750 & n30395;
  assign n30397 = ~n25765 & ~n27491;
  assign n30398 = n6777 & n30397;
  assign n30399 = ~n25766 & n27489;
  assign n30400 = n7044 & ~n30399;
  assign n30401 = ~n30398 & ~n30400;
  assign n30402 = pi306 & ~n30401;
  assign n30403 = ~n30396 & ~n30402;
  assign n30404 = ~n30394 & n30403;
  assign n30405 = n30394 & ~n30403;
  assign n30406 = ~n30404 & ~n30405;
  assign n30407 = n25739 & n25745;
  assign n30408 = ~n25739 & ~n25745;
  assign n30409 = n25408 & ~n30408;
  assign n30410 = ~n30407 & ~n30409;
  assign n30411 = n27473 & ~n30410;
  assign n30412 = ~n27473 & n30410;
  assign n30413 = ~n27472 & ~n30412;
  assign n30414 = ~n30411 & ~n30413;
  assign n30415 = pi307 & n9517;
  assign n30416 = ~n30414 & ~n30415;
  assign n30417 = n9517 & n30414;
  assign n30418 = pi307 & n30417;
  assign n30419 = ~n30416 & ~n30418;
  assign n30420 = n25659 & n25665;
  assign n30421 = ~n25659 & ~n25665;
  assign n30422 = n25420 & ~n30421;
  assign n30423 = ~n30420 & ~n30422;
  assign n30424 = n27384 & ~n30423;
  assign n30425 = n25606 & ~n27370;
  assign n30426 = ~n14618 & ~n27346;
  assign n30427 = n14156 & ~n30426;
  assign n30428 = pi313 & n30427;
  assign n30429 = ~n30425 & ~n30428;
  assign n30430 = ~n27359 & ~n30429;
  assign n30431 = n14618 & n27346;
  assign n30432 = n25606 & n30427;
  assign n30433 = ~n30431 & ~n30432;
  assign n30434 = pi313 & ~n30433;
  assign n30435 = ~n30430 & ~n30434;
  assign n30436 = pi313 & n16985;
  assign n30437 = ~n30435 & ~n30436;
  assign n30438 = n16985 & n30435;
  assign n30439 = pi313 & n30438;
  assign n30440 = ~n30437 & ~n30439;
  assign n30441 = n27304 & ~n27327;
  assign n30442 = ~n27304 & n27327;
  assign n30443 = n18937 & ~n27311;
  assign n30444 = pi316 & n30443;
  assign n30445 = ~n27302 & ~n27303;
  assign n30446 = ~n30444 & ~n30445;
  assign n30447 = ~n30442 & ~n30446;
  assign n30448 = ~n30441 & ~n30447;
  assign n30449 = ~n27330 & ~n27331;
  assign n30450 = n27330 & n27331;
  assign n30451 = ~n25604 & ~n30450;
  assign n30452 = ~n25598 & n30451;
  assign n30453 = ~n30449 & ~n30452;
  assign n30454 = n30448 & ~n30453;
  assign n30455 = ~n30448 & n30453;
  assign n30456 = ~n30454 & ~n30455;
  assign n30457 = pi316 & n20347;
  assign n30458 = pi320 & n27198;
  assign n30459 = ~pi156 & n27190;
  assign n30460 = pi156 & n27191;
  assign n30461 = ~n30459 & ~n30460;
  assign n30462 = pi158 & n30461;
  assign n30463 = ~pi158 & ~n30461;
  assign n30464 = ~n30462 & ~n30463;
  assign n30465 = ~n30458 & ~n30464;
  assign n30466 = pi321 & n30465;
  assign n30467 = pi158 & ~n30461;
  assign n30468 = ~pi158 & n30461;
  assign n30469 = ~n30467 & ~n30468;
  assign n30470 = pi321 & n30469;
  assign n30471 = n27198 & ~n30470;
  assign n30472 = pi320 & n30471;
  assign n30473 = ~n30466 & ~n30472;
  assign n30474 = pi319 & n25479;
  assign n30475 = n30473 & ~n30474;
  assign n30476 = n25479 & ~n30473;
  assign n30477 = pi319 & n30476;
  assign n30478 = ~n30475 & ~n30477;
  assign n30479 = ~n25451 & n27198;
  assign n30480 = ~n25479 & ~n30479;
  assign n30481 = n23626 & ~n30480;
  assign n30482 = n25479 & ~n27213;
  assign n30483 = ~n30481 & ~n30482;
  assign n30484 = pi321 & ~n30483;
  assign n30485 = n23626 & n27199;
  assign n30486 = ~n30484 & ~n30485;
  assign n30487 = pi320 & ~n30486;
  assign n30488 = n25482 & n30479;
  assign n30489 = ~n30487 & ~n30488;
  assign n30490 = ~n27225 & ~n27250;
  assign n30491 = n27225 & n27250;
  assign n30492 = n23626 & ~n30491;
  assign n30493 = pi319 & n30492;
  assign n30494 = ~n30490 & ~n30493;
  assign n30495 = n30489 & n30494;
  assign n30496 = ~n30489 & ~n30494;
  assign n30497 = ~n30495 & ~n30496;
  assign n30498 = ~n30478 & ~n30497;
  assign n30499 = ~n30489 & n30494;
  assign n30500 = n30489 & ~n30494;
  assign n30501 = ~n30499 & ~n30500;
  assign n30502 = ~n30473 & ~n30474;
  assign n30503 = n25479 & n30473;
  assign n30504 = pi319 & n30503;
  assign n30505 = ~n30502 & ~n30504;
  assign n30506 = ~n30501 & ~n30505;
  assign n30507 = ~n30498 & ~n30506;
  assign n30508 = pi318 & n23626;
  assign n30509 = n30507 & ~n30508;
  assign n30510 = n23626 & ~n30507;
  assign n30511 = pi318 & n30510;
  assign n30512 = ~n30509 & ~n30511;
  assign n30513 = ~n27256 & ~n27264;
  assign n30514 = ~n27259 & ~n30513;
  assign n30515 = n23069 & n27264;
  assign n30516 = pi318 & n30515;
  assign n30517 = ~n30514 & ~n30516;
  assign n30518 = ~n30512 & ~n30517;
  assign n30519 = n30512 & n30517;
  assign n30520 = ~n30518 & ~n30519;
  assign n30521 = n23069 & ~n30520;
  assign n30522 = pi317 & n30521;
  assign n30523 = pi317 & n23069;
  assign n30524 = n30512 & ~n30517;
  assign n30525 = ~n30512 & n30517;
  assign n30526 = ~n30524 & ~n30525;
  assign n30527 = ~n30523 & ~n30526;
  assign n30528 = ~n30522 & ~n30527;
  assign n30529 = ~n27182 & ~n27272;
  assign n30530 = ~n30528 & ~n30529;
  assign n30531 = ~n27269 & n30530;
  assign n30532 = ~n27269 & ~n30529;
  assign n30533 = n30528 & ~n30532;
  assign n30534 = ~n30531 & ~n30533;
  assign n30535 = ~n30457 & ~n30534;
  assign n30536 = n30528 & ~n30529;
  assign n30537 = ~n27269 & n30536;
  assign n30538 = ~n30528 & ~n30532;
  assign n30539 = ~n30537 & ~n30538;
  assign n30540 = n20347 & ~n30539;
  assign n30541 = pi316 & n30540;
  assign n30542 = ~n30535 & ~n30541;
  assign n30543 = n18937 & ~n27310;
  assign n30544 = pi316 & n30543;
  assign n30545 = ~n27309 & ~n30544;
  assign n30546 = n30542 & n30545;
  assign n30547 = ~n30542 & ~n30545;
  assign n30548 = ~n30546 & ~n30547;
  assign n30549 = n18937 & ~n30548;
  assign n30550 = pi315 & n30549;
  assign n30551 = pi315 & n18937;
  assign n30552 = ~n30542 & n30545;
  assign n30553 = n30542 & ~n30545;
  assign n30554 = ~n30552 & ~n30553;
  assign n30555 = ~n30551 & ~n30554;
  assign n30556 = ~n30550 & ~n30555;
  assign n30557 = pi314 & n17455;
  assign n30558 = n30556 & ~n30557;
  assign n30559 = n17455 & ~n30556;
  assign n30560 = pi314 & n30559;
  assign n30561 = ~n30558 & ~n30560;
  assign n30562 = ~n30456 & ~n30561;
  assign n30563 = ~n30448 & ~n30453;
  assign n30564 = n30448 & n30453;
  assign n30565 = ~n30563 & ~n30564;
  assign n30566 = ~n30556 & ~n30557;
  assign n30567 = n17455 & n30556;
  assign n30568 = pi314 & n30567;
  assign n30569 = ~n30566 & ~n30568;
  assign n30570 = ~n30565 & ~n30569;
  assign n30571 = ~n30562 & ~n30570;
  assign n30572 = n30440 & ~n30571;
  assign n30573 = ~n30440 & n30571;
  assign n30574 = ~n30572 & ~n30573;
  assign n30575 = pi312 & n14618;
  assign n30576 = ~n14156 & ~n14618;
  assign n30577 = pi313 & ~n30576;
  assign n30578 = n27346 & ~n30577;
  assign n30579 = ~n14156 & n14618;
  assign n30580 = pi313 & ~n27346;
  assign n30581 = n30579 & n30580;
  assign n30582 = ~n30578 & ~n30581;
  assign n30583 = ~n27360 & ~n30582;
  assign n30584 = ~n14618 & n27346;
  assign n30585 = ~n27348 & ~n30584;
  assign n30586 = ~n25606 & ~n30585;
  assign n30587 = n27359 & n30586;
  assign n30588 = n14156 & ~n14618;
  assign n30589 = ~n27346 & n30588;
  assign n30590 = ~n14156 & ~n25606;
  assign n30591 = n14618 & ~n30590;
  assign n30592 = n27346 & n30591;
  assign n30593 = ~n30589 & ~n30592;
  assign n30594 = pi313 & ~n30593;
  assign n30595 = n25606 & n27370;
  assign n30596 = ~n30594 & ~n30595;
  assign n30597 = ~n27359 & ~n30596;
  assign n30598 = ~n30426 & ~n30431;
  assign n30599 = n14156 & ~n30598;
  assign n30600 = pi313 & n30599;
  assign n30601 = n25606 & n30600;
  assign n30602 = ~n30597 & ~n30601;
  assign n30603 = ~n30587 & n30602;
  assign n30604 = ~n30583 & n30603;
  assign n30605 = ~n27381 & ~n30604;
  assign n30606 = n27381 & n30604;
  assign n30607 = n27350 & ~n30606;
  assign n30608 = ~n30605 & ~n30607;
  assign n30609 = n30575 & ~n30608;
  assign n30610 = ~n27350 & ~n30605;
  assign n30611 = ~n30606 & ~n30610;
  assign n30612 = ~n30575 & ~n30611;
  assign n30613 = ~n30609 & ~n30612;
  assign n30614 = ~n30574 & ~n30613;
  assign n30615 = n30440 & n30571;
  assign n30616 = ~n30440 & ~n30571;
  assign n30617 = ~n30615 & ~n30616;
  assign n30618 = ~n30575 & ~n30608;
  assign n30619 = n30575 & ~n30611;
  assign n30620 = ~n30618 & ~n30619;
  assign n30621 = ~n30617 & ~n30620;
  assign n30622 = ~n30614 & ~n30621;
  assign n30623 = ~n11998 & ~n14156;
  assign n30624 = pi311 & ~n30623;
  assign n30625 = ~n30622 & ~n30624;
  assign n30626 = ~n11998 & n30622;
  assign n30627 = pi311 & n14156;
  assign n30628 = n30626 & n30627;
  assign n30629 = ~n30625 & ~n30628;
  assign n30630 = ~n30424 & ~n30629;
  assign n30631 = n27384 & n30423;
  assign n30632 = ~n27384 & ~n30423;
  assign n30633 = ~n30631 & ~n30632;
  assign n30634 = n11998 & ~n30633;
  assign n30635 = ~n30622 & n30634;
  assign n30636 = ~n27384 & n30622;
  assign n30637 = n30423 & n30636;
  assign n30638 = n27384 & ~n30622;
  assign n30639 = ~n30423 & n30638;
  assign n30640 = ~n30637 & ~n30639;
  assign n30641 = pi311 & ~n30640;
  assign n30642 = ~n30635 & ~n30641;
  assign n30643 = n14156 & ~n30642;
  assign n30644 = ~n27384 & ~n30622;
  assign n30645 = n30423 & n30644;
  assign n30646 = ~n27384 & n30423;
  assign n30647 = n11998 & ~n30646;
  assign n30648 = pi311 & n30647;
  assign n30649 = ~n30424 & ~n30648;
  assign n30650 = n30622 & ~n30649;
  assign n30651 = ~n30645 & ~n30650;
  assign n30652 = ~n14156 & ~n30651;
  assign n30653 = ~pi311 & ~n30423;
  assign n30654 = n27384 & n30622;
  assign n30655 = n30653 & n30654;
  assign n30656 = ~n30652 & ~n30655;
  assign n30657 = ~n30643 & n30656;
  assign n30658 = ~n30630 & n30657;
  assign n30659 = ~n25678 & n27401;
  assign n30660 = n25670 & n30659;
  assign n30661 = ~n25680 & ~n27417;
  assign n30662 = n9815 & n30661;
  assign n30663 = ~n25679 & ~n27401;
  assign n30664 = n10908 & ~n30663;
  assign n30665 = ~n30662 & ~n30664;
  assign n30666 = pi310 & ~n30665;
  assign n30667 = ~n30660 & ~n30666;
  assign n30668 = n30658 & ~n30667;
  assign n30669 = ~n30658 & n30667;
  assign n30670 = ~n30668 & ~n30669;
  assign n30671 = n11998 & ~n30670;
  assign n30672 = pi310 & n30671;
  assign n30673 = pi310 & n11998;
  assign n30674 = ~n30658 & ~n30667;
  assign n30675 = n30658 & n30667;
  assign n30676 = ~n30674 & ~n30675;
  assign n30677 = ~n30673 & ~n30676;
  assign n30678 = ~n30672 & ~n30677;
  assign n30679 = ~pi309 & n30678;
  assign n30680 = ~n10908 & n30678;
  assign n30681 = n10908 & ~n30678;
  assign n30682 = pi309 & n30681;
  assign n30683 = ~n30680 & ~n30682;
  assign n30684 = ~n9815 & ~n30683;
  assign n30685 = ~n30679 & ~n30684;
  assign n30686 = ~n30383 & ~n30685;
  assign n30687 = ~n27433 & n30678;
  assign n30688 = ~n30382 & n30687;
  assign n30689 = n27433 & ~n30678;
  assign n30690 = n30382 & n30689;
  assign n30691 = ~n30688 & ~n30690;
  assign n30692 = pi309 & ~n30691;
  assign n30693 = ~n30389 & n30678;
  assign n30694 = n9815 & n30693;
  assign n30695 = ~n30692 & ~n30694;
  assign n30696 = n10908 & ~n30695;
  assign n30697 = n27433 & n30678;
  assign n30698 = n30382 & n30697;
  assign n30699 = n9815 & ~n30384;
  assign n30700 = pi309 & n30699;
  assign n30701 = ~n30383 & ~n30700;
  assign n30702 = ~n30678 & ~n30701;
  assign n30703 = ~n30698 & ~n30702;
  assign n30704 = ~n10908 & ~n30703;
  assign n30705 = ~n27433 & ~n30678;
  assign n30706 = ~pi309 & ~n30382;
  assign n30707 = n30705 & n30706;
  assign n30708 = ~n30704 & ~n30707;
  assign n30709 = ~n30696 & n30708;
  assign n30710 = ~n30686 & n30709;
  assign n30711 = pi308 & n9815;
  assign n30712 = n30710 & ~n30711;
  assign n30713 = n9815 & ~n30710;
  assign n30714 = pi308 & n30713;
  assign n30715 = ~n30712 & ~n30714;
  assign n30716 = n30419 & n30715;
  assign n30717 = ~n30419 & ~n30715;
  assign n30718 = ~n30716 & ~n30717;
  assign n30719 = n7874 & ~n30718;
  assign n30720 = pi306 & n30719;
  assign n30721 = pi306 & n7874;
  assign n30722 = ~n30419 & n30715;
  assign n30723 = n30419 & ~n30715;
  assign n30724 = ~n30722 & ~n30723;
  assign n30725 = ~n30721 & ~n30724;
  assign n30726 = ~n30720 & ~n30725;
  assign n30727 = ~n30406 & ~n30726;
  assign n30728 = ~n30394 & ~n30403;
  assign n30729 = n30394 & n30403;
  assign n30730 = ~n30728 & ~n30729;
  assign n30731 = n7874 & ~n30724;
  assign n30732 = pi306 & n30731;
  assign n30733 = ~n30718 & ~n30721;
  assign n30734 = ~n30732 & ~n30733;
  assign n30735 = ~n30730 & ~n30734;
  assign n30736 = ~n30727 & ~n30735;
  assign n30737 = ~n30377 & ~n30736;
  assign n30738 = n30377 & n30736;
  assign n30739 = ~n30737 & ~n30738;
  assign n30740 = n7044 & ~n30739;
  assign n30741 = pi305 & n30740;
  assign n30742 = pi305 & n7044;
  assign n30743 = n30377 & ~n30736;
  assign n30744 = ~n30377 & n30736;
  assign n30745 = ~n30743 & ~n30744;
  assign n30746 = ~n30742 & ~n30745;
  assign n30747 = ~n30741 & ~n30746;
  assign n30748 = pi304 & n6777;
  assign n30749 = ~n30747 & n30748;
  assign n30750 = n30747 & ~n30748;
  assign n30751 = ~n30749 & ~n30750;
  assign n30752 = n30367 & n30751;
  assign n30753 = ~n30367 & ~n30751;
  assign n30754 = ~n30752 & ~n30753;
  assign n30755 = n4772 & ~n30754;
  assign n30756 = pi302 & n30755;
  assign n30757 = pi302 & n4772;
  assign n30758 = ~n30367 & n30751;
  assign n30759 = n30367 & ~n30751;
  assign n30760 = ~n30758 & ~n30759;
  assign n30761 = ~n30757 & ~n30760;
  assign n30762 = ~n30756 & ~n30761;
  assign n30763 = ~n30354 & ~n30762;
  assign n30764 = ~n30343 & ~n30351;
  assign n30765 = n30343 & n30351;
  assign n30766 = ~n30764 & ~n30765;
  assign n30767 = n4772 & ~n30760;
  assign n30768 = pi302 & n30767;
  assign n30769 = ~n30754 & ~n30757;
  assign n30770 = ~n30768 & ~n30769;
  assign n30771 = ~n30766 & ~n30770;
  assign n30772 = ~n30763 & ~n30771;
  assign n30773 = n27613 & ~n27644;
  assign n30774 = pi301 & ~n11042;
  assign n30775 = n27609 & ~n30774;
  assign n30776 = pi301 & ~n27609;
  assign n30777 = n11045 & n30776;
  assign n30778 = ~n30775 & ~n30777;
  assign n30779 = ~n27623 & ~n30778;
  assign n30780 = ~n3552 & n27609;
  assign n30781 = ~n27611 & ~n30780;
  assign n30782 = ~n25846 & ~n30781;
  assign n30783 = n27622 & n30782;
  assign n30784 = n11054 & ~n27609;
  assign n30785 = ~n3012 & ~n25846;
  assign n30786 = n3552 & ~n30785;
  assign n30787 = n27609 & n30786;
  assign n30788 = ~n30784 & ~n30787;
  assign n30789 = pi301 & ~n30788;
  assign n30790 = n25846 & n27633;
  assign n30791 = ~n30789 & ~n30790;
  assign n30792 = ~n27622 & ~n30791;
  assign n30793 = ~n3552 & ~n27609;
  assign n30794 = n3552 & n27609;
  assign n30795 = ~n30793 & ~n30794;
  assign n30796 = n3012 & ~n30795;
  assign n30797 = pi301 & n30796;
  assign n30798 = n25846 & n30797;
  assign n30799 = ~n30792 & ~n30798;
  assign n30800 = ~n30783 & n30799;
  assign n30801 = ~n30779 & n30800;
  assign n30802 = ~n27613 & n27644;
  assign n30803 = ~n30801 & ~n30802;
  assign n30804 = ~n30773 & ~n30803;
  assign n30805 = ~n30772 & n30804;
  assign n30806 = n30772 & ~n30804;
  assign n30807 = ~n30805 & ~n30806;
  assign n30808 = n25846 & ~n27633;
  assign n30809 = n3012 & ~n30793;
  assign n30810 = pi301 & n30809;
  assign n30811 = ~n30808 & ~n30810;
  assign n30812 = ~n27622 & ~n30811;
  assign n30813 = n25846 & n30809;
  assign n30814 = ~n30794 & ~n30813;
  assign n30815 = pi301 & ~n30814;
  assign n30816 = ~n30812 & ~n30815;
  assign n30817 = pi301 & n4086;
  assign n30818 = ~n30816 & ~n30817;
  assign n30819 = n4086 & n30816;
  assign n30820 = pi301 & n30819;
  assign n30821 = ~n30818 & ~n30820;
  assign n30822 = pi300 & n3552;
  assign n30823 = ~n30821 & n30822;
  assign n30824 = n30821 & ~n30822;
  assign n30825 = ~n30823 & ~n30824;
  assign n30826 = ~n30807 & ~n30825;
  assign n30827 = ~n30772 & ~n30804;
  assign n30828 = n30772 & n30804;
  assign n30829 = ~n30827 & ~n30828;
  assign n30830 = ~n30821 & ~n30822;
  assign n30831 = n30821 & n30822;
  assign n30832 = ~n30830 & ~n30831;
  assign n30833 = ~n30829 & ~n30832;
  assign n30834 = ~n30826 & ~n30833;
  assign n30835 = ~n2183 & ~n27664;
  assign n30836 = ~n25914 & ~n30835;
  assign n30837 = n1840 & n30836;
  assign n30838 = ~n25913 & ~n27664;
  assign n30839 = n2183 & ~n30838;
  assign n30840 = ~n30837 & ~n30839;
  assign n30841 = pi298 & ~n30840;
  assign n30842 = ~n27674 & ~n30841;
  assign n30843 = n30834 & n30842;
  assign n30844 = ~n30834 & ~n30842;
  assign n30845 = ~n30843 & ~n30844;
  assign n30846 = pi299 & n3012;
  assign n30847 = ~n27647 & ~n27648;
  assign n30848 = n27647 & n27648;
  assign n30849 = ~n27653 & ~n30848;
  assign n30850 = ~n30847 & ~n30849;
  assign n30851 = ~n30846 & n30850;
  assign n30852 = n30846 & ~n30850;
  assign n30853 = ~n30851 & ~n30852;
  assign n30854 = n2574 & ~n30853;
  assign n30855 = pi298 & n30854;
  assign n30856 = pi298 & n2574;
  assign n30857 = n30846 & n30850;
  assign n30858 = ~n30846 & ~n30850;
  assign n30859 = ~n30857 & ~n30858;
  assign n30860 = ~n30856 & ~n30859;
  assign n30861 = ~n30855 & ~n30860;
  assign n30862 = ~n30845 & ~n30861;
  assign n30863 = n30834 & ~n30842;
  assign n30864 = ~n30834 & n30842;
  assign n30865 = ~n30863 & ~n30864;
  assign n30866 = n2574 & ~n30859;
  assign n30867 = pi298 & n30866;
  assign n30868 = ~n30853 & ~n30856;
  assign n30869 = ~n30867 & ~n30868;
  assign n30870 = ~n30865 & ~n30869;
  assign n30871 = ~n30862 & ~n30870;
  assign n30872 = n30311 & n30871;
  assign n30873 = ~n30311 & ~n30871;
  assign n30874 = ~n30872 & ~n30873;
  assign n30875 = pi296 & n1840;
  assign n30876 = n27737 & ~n27738;
  assign n30877 = ~n27739 & ~n30876;
  assign n30878 = n30875 & ~n30877;
  assign n30879 = ~n27737 & ~n27739;
  assign n30880 = ~n27738 & ~n30879;
  assign n30881 = ~n30875 & ~n30880;
  assign n30882 = ~n30878 & ~n30881;
  assign n30883 = ~n30874 & ~n30882;
  assign n30884 = n30311 & ~n30871;
  assign n30885 = ~n30311 & n30871;
  assign n30886 = ~n30884 & ~n30885;
  assign n30887 = ~n30875 & ~n30877;
  assign n30888 = n30875 & ~n30880;
  assign n30889 = ~n30887 & ~n30888;
  assign n30890 = ~n30886 & ~n30889;
  assign n30891 = ~n30883 & ~n30890;
  assign n30892 = ~pi295 & n30891;
  assign n30893 = ~n1533 & n30891;
  assign n30894 = n1533 & ~n30891;
  assign n30895 = pi295 & n30894;
  assign n30896 = ~n30893 & ~n30895;
  assign n30897 = ~n1553 & ~n30896;
  assign n30898 = ~n30892 & ~n30897;
  assign n30899 = ~n30297 & ~n30898;
  assign n30900 = n27742 & n30891;
  assign n30901 = ~n30296 & n30900;
  assign n30902 = ~n27742 & ~n30891;
  assign n30903 = n30296 & n30902;
  assign n30904 = ~n30901 & ~n30903;
  assign n30905 = pi295 & ~n30904;
  assign n30906 = ~n27742 & ~n30296;
  assign n30907 = n27742 & n30296;
  assign n30908 = ~n30906 & ~n30907;
  assign n30909 = n30891 & ~n30908;
  assign n30910 = n1553 & n30909;
  assign n30911 = ~n30905 & ~n30910;
  assign n30912 = n1533 & ~n30911;
  assign n30913 = n27742 & ~n30891;
  assign n30914 = ~pi295 & ~n30296;
  assign n30915 = n30913 & n30914;
  assign n30916 = ~n27742 & n30891;
  assign n30917 = n30296 & n30916;
  assign n30918 = ~n27742 & n30296;
  assign n30919 = n1553 & ~n30918;
  assign n30920 = pi295 & n30919;
  assign n30921 = ~n30297 & ~n30920;
  assign n30922 = ~n30891 & ~n30921;
  assign n30923 = ~n30917 & ~n30922;
  assign n30924 = ~n1533 & ~n30923;
  assign n30925 = ~n30915 & ~n30924;
  assign n30926 = ~n30912 & n30925;
  assign n30927 = ~n30899 & n30926;
  assign n30928 = n27742 & n27762;
  assign n30929 = ~n27742 & ~n27762;
  assign n30930 = ~n30928 & ~n30929;
  assign n30931 = n27746 & ~n27763;
  assign n30932 = ~n30930 & ~n30931;
  assign n30933 = n1515 & ~n27746;
  assign n30934 = pi294 & n30933;
  assign n30935 = ~n30932 & ~n30934;
  assign n30936 = ~n30927 & n30935;
  assign n30937 = n30927 & ~n30935;
  assign n30938 = ~n30936 & ~n30937;
  assign n30939 = n1553 & ~n30938;
  assign n30940 = pi294 & n30939;
  assign n30941 = pi294 & n1553;
  assign n30942 = n30927 & n30935;
  assign n30943 = ~n30927 & ~n30935;
  assign n30944 = ~n30942 & ~n30943;
  assign n30945 = ~n30941 & ~n30944;
  assign n30946 = ~n30940 & ~n30945;
  assign n30947 = n30292 & ~n30946;
  assign n30948 = ~n30292 & n30946;
  assign n30949 = ~n30947 & ~n30948;
  assign n30950 = pi292 & ~n27786;
  assign n30951 = pi128 & n30950;
  assign n30952 = pi292 & ~n1568;
  assign n30953 = ~n30951 & ~n30952;
  assign n30954 = n30951 & n30952;
  assign n30955 = ~n30953 & ~n30954;
  assign n30956 = pi291 & ~n30955;
  assign n30957 = pi128 & n30956;
  assign n30958 = pi128 & pi291;
  assign n30959 = n30951 & ~n30952;
  assign n30960 = ~n30951 & n30952;
  assign n30961 = ~n30959 & ~n30960;
  assign n30962 = ~n30958 & ~n30961;
  assign n30963 = ~n30957 & ~n30962;
  assign n30964 = ~n30949 & ~n30963;
  assign n30965 = n30292 & n30946;
  assign n30966 = ~n30292 & ~n30946;
  assign n30967 = ~n30965 & ~n30966;
  assign n30968 = pi291 & ~n30961;
  assign n30969 = pi128 & n30968;
  assign n30970 = ~n30955 & ~n30958;
  assign n30971 = ~n30969 & ~n30970;
  assign n30972 = ~n30967 & ~n30971;
  assign n30973 = ~n30964 & ~n30972;
  assign n30974 = n1156 & ~n28993;
  assign n30975 = pi351 & n30974;
  assign n30976 = ~n29007 & ~n29016;
  assign n30977 = ~n30975 & ~n30976;
  assign n30978 = ~n29009 & ~n30977;
  assign n30979 = ~n29008 & ~n30978;
  assign n30980 = n30973 & n30979;
  assign n30981 = ~n30973 & ~n30979;
  assign n30982 = ~n30980 & ~n30981;
  assign n30983 = pi288 & ~n30982;
  assign n30984 = ~n30973 & n30979;
  assign n30985 = n30973 & ~n30979;
  assign n30986 = ~n30984 & ~n30985;
  assign n30987 = ~pi288 & ~n30986;
  assign n30988 = ~n30983 & ~n30987;
  assign n30989 = ~n30264 & ~n30988;
  assign n30990 = n30257 & ~n30261;
  assign n30991 = ~n30257 & n30261;
  assign n30992 = ~n30990 & ~n30991;
  assign n30993 = pi288 & ~n30986;
  assign n30994 = ~pi288 & ~n30982;
  assign n30995 = ~n30993 & ~n30994;
  assign n30996 = ~n30992 & ~n30995;
  assign n30997 = ~n30989 & ~n30996;
  assign n30998 = ~n831 & ~n30997;
  assign n30999 = ~pi288 & n831;
  assign n31000 = ~n30998 & ~n30999;
  assign n31001 = pi161 & n31000;
  assign n31002 = ~n29038 & ~n31001;
  assign po223 = ~pi160 & ~n31002;
  assign n31004 = pi095 & ~pi161;
  assign n31005 = ~pi289 & n831;
  assign n31006 = pi161 & ~n31005;
  assign n31007 = n1335 & n30272;
  assign n31008 = ~pi129 & n27169;
  assign n31009 = pi129 & ~n27169;
  assign n31010 = n27777 & ~n31009;
  assign n31011 = pi128 & n31010;
  assign n31012 = ~n31008 & ~n31011;
  assign n31013 = pi130 & ~n31012;
  assign n31014 = ~n31007 & ~n31013;
  assign n31015 = pi293 & ~n31014;
  assign n31016 = pi290 & ~pi291;
  assign n31017 = ~pi290 & pi291;
  assign n31018 = ~pi129 & n31017;
  assign n31019 = ~n31016 & ~n31018;
  assign n31020 = pi128 & ~n31019;
  assign n31021 = pi128 & ~pi290;
  assign n31022 = pi291 & ~n31021;
  assign n31023 = pi129 & n31022;
  assign n31024 = ~n31020 & ~n31023;
  assign n31025 = ~n30948 & ~n31024;
  assign n31026 = pi129 & pi291;
  assign n31027 = ~pi128 & ~n31026;
  assign n31028 = pi291 & ~n1175;
  assign n31029 = ~pi290 & ~n31028;
  assign n31030 = pi290 & pi291;
  assign n31031 = ~pi129 & n31030;
  assign n31032 = ~n31029 & ~n31031;
  assign n31033 = ~n31027 & n31032;
  assign n31034 = n30946 & ~n31033;
  assign n31035 = ~n30292 & n31034;
  assign n31036 = ~n31025 & ~n31035;
  assign n31037 = n31015 & ~n31036;
  assign n31038 = ~n31015 & n31036;
  assign n31039 = n1515 & n31038;
  assign n31040 = ~n31037 & ~n31039;
  assign n31041 = pi292 & ~n31040;
  assign n31042 = ~n31015 & ~n31036;
  assign n31043 = ~n1515 & n31042;
  assign n31044 = n31015 & n31036;
  assign n31045 = ~n31042 & ~n31044;
  assign n31046 = ~pi292 & ~n31045;
  assign n31047 = ~n31043 & ~n31046;
  assign n31048 = ~n31041 & n31047;
  assign n31049 = pi352 & ~n1154;
  assign n31050 = ~n1256 & ~n31049;
  assign n31051 = pi351 & n31050;
  assign n31052 = pi351 & ~n1256;
  assign n31053 = ~n1154 & ~n31052;
  assign n31054 = pi352 & n31053;
  assign n31055 = ~n31051 & ~n31054;
  assign n31056 = ~n30955 & ~n30967;
  assign n31057 = ~n30949 & ~n30961;
  assign n31058 = ~n31056 & ~n31057;
  assign n31059 = pi291 & ~n31058;
  assign n31060 = pi128 & n31059;
  assign n31061 = ~n1533 & ~n30891;
  assign n31062 = ~n30918 & ~n31061;
  assign n31063 = n1553 & n31062;
  assign n31064 = ~n30297 & ~n30891;
  assign n31065 = n1533 & ~n31064;
  assign n31066 = ~n31063 & ~n31065;
  assign n31067 = pi295 & ~n31066;
  assign n31068 = ~n30901 & ~n31067;
  assign n31069 = pi296 & n2183;
  assign n31070 = n1840 & ~n31069;
  assign n31071 = pi295 & n31070;
  assign n31072 = pi295 & n1840;
  assign n31073 = n2183 & ~n31072;
  assign n31074 = pi296 & n31073;
  assign n31075 = ~n31071 & ~n31074;
  assign n31076 = n31068 & n31075;
  assign n31077 = ~n31068 & ~n31075;
  assign n31078 = ~n31076 & ~n31077;
  assign n31079 = n31060 & ~n31078;
  assign n31080 = n31068 & ~n31075;
  assign n31081 = ~n31068 & n31075;
  assign n31082 = ~n31080 & ~n31081;
  assign n31083 = ~n31060 & ~n31082;
  assign n31084 = ~n31079 & ~n31083;
  assign n31085 = ~n30874 & ~n30875;
  assign n31086 = n30874 & n30875;
  assign n31087 = ~n30880 & ~n31086;
  assign n31088 = ~n31085 & ~n31087;
  assign n31089 = pi297 & n2574;
  assign n31090 = n31088 & ~n31089;
  assign n31091 = n2574 & ~n31088;
  assign n31092 = pi297 & n31091;
  assign n31093 = ~n31090 & ~n31092;
  assign n31094 = n30834 & n30846;
  assign n31095 = ~n30834 & ~n30846;
  assign n31096 = n30850 & ~n31095;
  assign n31097 = ~n31094 & ~n31096;
  assign n31098 = n30772 & n30821;
  assign n31099 = ~n30772 & ~n30821;
  assign n31100 = ~n31098 & ~n31099;
  assign n31101 = n30804 & ~n30822;
  assign n31102 = ~n31100 & ~n31101;
  assign n31103 = n3552 & ~n30804;
  assign n31104 = pi300 & n31103;
  assign n31105 = ~n31102 & ~n31104;
  assign n31106 = pi304 & n7044;
  assign n31107 = n31105 & ~n31106;
  assign n31108 = n7044 & ~n31105;
  assign n31109 = pi304 & n31108;
  assign n31110 = ~n31107 & ~n31109;
  assign n31111 = n5463 & ~n30362;
  assign n31112 = pi303 & n31111;
  assign n31113 = n30343 & ~n30751;
  assign n31114 = ~n30343 & n30751;
  assign n31115 = ~n31113 & ~n31114;
  assign n31116 = n30362 & ~n30363;
  assign n31117 = ~n31115 & ~n31116;
  assign n31118 = ~n31112 & ~n31117;
  assign n31119 = ~n30343 & n30747;
  assign n31120 = n30343 & ~n30747;
  assign n31121 = n30748 & ~n31120;
  assign n31122 = ~n31119 & ~n31121;
  assign n31123 = n9517 & ~n30414;
  assign n31124 = pi307 & n31123;
  assign n31125 = n30394 & ~n30715;
  assign n31126 = ~n30394 & n30715;
  assign n31127 = ~n31125 & ~n31126;
  assign n31128 = n30414 & ~n30415;
  assign n31129 = ~n31127 & ~n31128;
  assign n31130 = ~n31124 & ~n31129;
  assign n31131 = n30394 & ~n30710;
  assign n31132 = ~n30394 & n30710;
  assign n31133 = ~n30711 & ~n31132;
  assign n31134 = ~n31131 & ~n31133;
  assign n31135 = n11998 & ~n31134;
  assign n31136 = pi309 & n31135;
  assign n31137 = pi309 & n11998;
  assign n31138 = n9815 & ~n31131;
  assign n31139 = pi308 & n31138;
  assign n31140 = ~n31132 & ~n31139;
  assign n31141 = ~n31137 & ~n31140;
  assign n31142 = ~n31136 & ~n31141;
  assign n31143 = pi312 & n16985;
  assign n31144 = n31142 & ~n31143;
  assign n31145 = n16985 & ~n31142;
  assign n31146 = pi312 & n31145;
  assign n31147 = ~n31144 & ~n31146;
  assign n31148 = ~n30423 & n30654;
  assign n31149 = n30622 & n30647;
  assign n31150 = n11998 & n27384;
  assign n31151 = ~n30622 & ~n31150;
  assign n31152 = ~n11998 & ~n27384;
  assign n31153 = ~n30423 & ~n31152;
  assign n31154 = n31151 & ~n31153;
  assign n31155 = n14156 & ~n31154;
  assign n31156 = ~n31149 & ~n31155;
  assign n31157 = pi311 & ~n31156;
  assign n31158 = ~n31148 & ~n31157;
  assign n31159 = n25479 & ~n30494;
  assign n31160 = pi319 & n31159;
  assign n31161 = n30473 & ~n30489;
  assign n31162 = ~n30473 & n30489;
  assign n31163 = ~n31161 & ~n31162;
  assign n31164 = ~n30474 & n30494;
  assign n31165 = ~n31163 & ~n31164;
  assign n31166 = ~n31160 & ~n31165;
  assign n31167 = n30507 & ~n30517;
  assign n31168 = ~n30507 & n30517;
  assign n31169 = n23626 & ~n31168;
  assign n31170 = pi318 & n31169;
  assign n31171 = ~n31167 & ~n31170;
  assign n31172 = ~n31166 & ~n31171;
  assign n31173 = n31166 & n31171;
  assign n31174 = ~n31172 & ~n31173;
  assign n31175 = n30534 & n30545;
  assign n31176 = ~n30534 & ~n30545;
  assign n31177 = ~n20347 & ~n31176;
  assign n31178 = ~n31175 & ~n31177;
  assign n31179 = n23069 & ~n31178;
  assign n31180 = ~n23069 & ~n31175;
  assign n31181 = n20347 & n31180;
  assign n31182 = ~n31179 & ~n31181;
  assign n31183 = pi316 & ~n31182;
  assign n31184 = pi316 & n23069;
  assign n31185 = ~n30545 & ~n31184;
  assign n31186 = ~n30534 & n31185;
  assign n31187 = ~n31183 & ~n31186;
  assign n31188 = n30575 & ~n30617;
  assign n31189 = ~n30575 & n30617;
  assign n31190 = ~n30608 & ~n31189;
  assign n31191 = ~n31188 & ~n31190;
  assign n31192 = n31187 & n31191;
  assign n31193 = ~n31187 & ~n31191;
  assign n31194 = ~n31192 & ~n31193;
  assign n31195 = n17455 & ~n31194;
  assign n31196 = pi313 & n31195;
  assign n31197 = pi313 & n17455;
  assign n31198 = ~n31187 & n31191;
  assign n31199 = n31187 & ~n31191;
  assign n31200 = ~n31198 & ~n31199;
  assign n31201 = ~n31197 & ~n31200;
  assign n31202 = ~n31196 & ~n31201;
  assign n31203 = ~n31174 & ~n31202;
  assign n31204 = ~n31166 & n31171;
  assign n31205 = n31166 & ~n31171;
  assign n31206 = ~n31204 & ~n31205;
  assign n31207 = n17455 & ~n31200;
  assign n31208 = pi313 & n31207;
  assign n31209 = ~n31194 & ~n31197;
  assign n31210 = ~n31208 & ~n31209;
  assign n31211 = ~n31206 & ~n31210;
  assign n31212 = ~n31203 & ~n31211;
  assign n31213 = n31158 & ~n31212;
  assign n31214 = ~n31158 & n31212;
  assign n31215 = ~n31213 & ~n31214;
  assign n31216 = ~n31147 & ~n31215;
  assign n31217 = ~n31158 & ~n31212;
  assign n31218 = n31158 & n31212;
  assign n31219 = ~n31217 & ~n31218;
  assign n31220 = ~n31142 & ~n31143;
  assign n31221 = n16985 & n31142;
  assign n31222 = pi312 & n31221;
  assign n31223 = ~n31220 & ~n31222;
  assign n31224 = ~n31219 & ~n31223;
  assign n31225 = ~n31216 & ~n31224;
  assign n31226 = ~n31130 & n31225;
  assign n31227 = n31130 & ~n31225;
  assign n31228 = ~n31226 & ~n31227;
  assign n31229 = pi308 & n10908;
  assign n31230 = pi307 & n9815;
  assign n31231 = ~n31229 & ~n31230;
  assign n31232 = n9815 & n10908;
  assign n31233 = pi307 & pi308;
  assign n31234 = n31232 & n31233;
  assign n31235 = ~n31231 & ~n31234;
  assign n31236 = ~n31228 & ~n31235;
  assign n31237 = ~n31130 & ~n31225;
  assign n31238 = n31130 & n31225;
  assign n31239 = ~n31237 & ~n31238;
  assign n31240 = n9815 & ~n31229;
  assign n31241 = pi307 & n31240;
  assign n31242 = n10908 & ~n31230;
  assign n31243 = pi308 & n31242;
  assign n31244 = ~n31241 & ~n31243;
  assign n31245 = ~n31239 & ~n31244;
  assign n31246 = ~n31236 & ~n31245;
  assign n31247 = pi305 & n7874;
  assign n31248 = ~n31246 & ~n31247;
  assign n31249 = n7874 & n31246;
  assign n31250 = pi305 & n31249;
  assign n31251 = ~n31248 & ~n31250;
  assign n31252 = ~n31122 & ~n31251;
  assign n31253 = ~n30748 & ~n31119;
  assign n31254 = ~n31120 & ~n31253;
  assign n31255 = n31246 & ~n31247;
  assign n31256 = n7874 & ~n31246;
  assign n31257 = pi305 & n31256;
  assign n31258 = ~n31255 & ~n31257;
  assign n31259 = ~n31254 & ~n31258;
  assign n31260 = ~n31252 & ~n31259;
  assign n31261 = n31118 & ~n31260;
  assign n31262 = ~n31118 & n31260;
  assign n31263 = ~n31261 & ~n31262;
  assign n31264 = ~n31110 & ~n31263;
  assign n31265 = ~n31118 & ~n31260;
  assign n31266 = n31118 & n31260;
  assign n31267 = ~n31265 & ~n31266;
  assign n31268 = ~n31105 & ~n31106;
  assign n31269 = n7044 & n31105;
  assign n31270 = pi304 & n31269;
  assign n31271 = ~n31268 & ~n31270;
  assign n31272 = ~n31267 & ~n31271;
  assign n31273 = ~n31264 & ~n31272;
  assign n31274 = pi300 & n4086;
  assign n31275 = n31273 & ~n31274;
  assign n31276 = n4086 & ~n31273;
  assign n31277 = pi300 & n31276;
  assign n31278 = ~n31275 & ~n31277;
  assign n31279 = n31097 & ~n31278;
  assign n31280 = ~n31097 & n31278;
  assign n31281 = ~n31279 & ~n31280;
  assign n31282 = ~n31093 & ~n31281;
  assign n31283 = ~n31097 & ~n31278;
  assign n31284 = n31097 & n31278;
  assign n31285 = ~n31283 & ~n31284;
  assign n31286 = ~n31088 & ~n31089;
  assign n31287 = n2574 & n31088;
  assign n31288 = pi297 & n31287;
  assign n31289 = ~n31286 & ~n31288;
  assign n31290 = ~n31285 & ~n31289;
  assign n31291 = ~n31282 & ~n31290;
  assign n31292 = ~n30834 & n30850;
  assign n31293 = n30834 & ~n30850;
  assign n31294 = ~n31292 & ~n31293;
  assign n31295 = ~n30846 & ~n31294;
  assign n31296 = ~n30834 & ~n30850;
  assign n31297 = n30834 & n30850;
  assign n31298 = ~n31296 & ~n31297;
  assign n31299 = n30846 & ~n31298;
  assign n31300 = ~n31295 & ~n31299;
  assign n31301 = n30842 & ~n30856;
  assign n31302 = ~n31300 & ~n31301;
  assign n31303 = n2574 & ~n30842;
  assign n31304 = pi298 & n31303;
  assign n31305 = ~n31302 & ~n31304;
  assign n31306 = pi302 & n5463;
  assign n31307 = n4772 & ~n30351;
  assign n31308 = pi302 & n31307;
  assign n31309 = n30343 & n30751;
  assign n31310 = ~n30343 & ~n30751;
  assign n31311 = ~n31309 & ~n31310;
  assign n31312 = ~n30367 & ~n31311;
  assign n31313 = n30367 & ~n31115;
  assign n31314 = ~n31312 & ~n31313;
  assign n31315 = n30351 & ~n30757;
  assign n31316 = ~n31314 & ~n31315;
  assign n31317 = ~n31308 & ~n31316;
  assign n31318 = n30742 & ~n30743;
  assign n31319 = ~n30744 & ~n31318;
  assign n31320 = n30394 & n30715;
  assign n31321 = ~n30394 & ~n30715;
  assign n31322 = ~n31320 & ~n31321;
  assign n31323 = ~n30419 & ~n31322;
  assign n31324 = n30419 & ~n31127;
  assign n31325 = ~n31323 & ~n31324;
  assign n31326 = n30403 & ~n30721;
  assign n31327 = ~n31325 & ~n31326;
  assign n31328 = n7874 & ~n30403;
  assign n31329 = pi306 & n31328;
  assign n31330 = ~n31327 & ~n31329;
  assign n31331 = pi310 & n14156;
  assign n31332 = n31330 & ~n31331;
  assign n31333 = n14156 & ~n31330;
  assign n31334 = pi310 & n31333;
  assign n31335 = ~n31332 & ~n31334;
  assign n31336 = ~n30382 & n30705;
  assign n31337 = ~n30384 & ~n30680;
  assign n31338 = n9815 & n31337;
  assign n31339 = ~n30383 & n30678;
  assign n31340 = n10908 & ~n31339;
  assign n31341 = ~n31338 & ~n31340;
  assign n31342 = pi309 & ~n31341;
  assign n31343 = ~n31336 & ~n31342;
  assign n31344 = n11998 & ~n30669;
  assign n31345 = pi310 & n31344;
  assign n31346 = ~n30668 & ~n31345;
  assign n31347 = pi311 & n14618;
  assign n31348 = ~n31346 & ~n31347;
  assign n31349 = n14618 & n31346;
  assign n31350 = pi311 & n31349;
  assign n31351 = ~n31348 & ~n31350;
  assign n31352 = ~n30435 & n30571;
  assign n31353 = n30435 & ~n30571;
  assign n31354 = n16985 & ~n31353;
  assign n31355 = pi313 & n31354;
  assign n31356 = ~n31352 & ~n31355;
  assign n31357 = pi314 & n18937;
  assign n31358 = ~n30532 & ~n31357;
  assign n31359 = ~n30528 & n31358;
  assign n31360 = n18937 & ~n30538;
  assign n31361 = pi314 & n31360;
  assign n31362 = ~n31359 & ~n31361;
  assign n31363 = n30448 & ~n30556;
  assign n31364 = ~n30448 & n30556;
  assign n31365 = ~n31363 & ~n31364;
  assign n31366 = ~n30453 & ~n30557;
  assign n31367 = ~n31365 & ~n31366;
  assign n31368 = n17455 & n30453;
  assign n31369 = pi314 & n31368;
  assign n31370 = ~n31367 & ~n31369;
  assign n31371 = ~n31362 & ~n31370;
  assign n31372 = n31362 & n31370;
  assign n31373 = ~n31371 & ~n31372;
  assign n31374 = ~n30448 & n30551;
  assign n31375 = n30448 & ~n30551;
  assign n31376 = ~n30554 & ~n31375;
  assign n31377 = ~n31374 & ~n31376;
  assign n31378 = ~n31373 & ~n31377;
  assign n31379 = ~n31362 & n31370;
  assign n31380 = n31362 & ~n31370;
  assign n31381 = ~n31379 & ~n31380;
  assign n31382 = ~n30548 & ~n31374;
  assign n31383 = ~n31375 & ~n31382;
  assign n31384 = ~n31381 & ~n31383;
  assign n31385 = ~n31378 & ~n31384;
  assign n31386 = pi319 & n27198;
  assign n31387 = ~pi158 & ~pi159;
  assign n31388 = pi157 & n31387;
  assign n31389 = pi159 & ~n27189;
  assign n31390 = pi158 & n31389;
  assign n31391 = ~n31388 & ~n31390;
  assign n31392 = pi156 & ~n31391;
  assign n31393 = pi158 & ~pi159;
  assign n31394 = ~pi157 & n31393;
  assign n31395 = pi159 & n27189;
  assign n31396 = ~pi158 & n31395;
  assign n31397 = ~n31394 & ~n31396;
  assign n31398 = ~pi156 & ~n31397;
  assign n31399 = pi158 & pi159;
  assign n31400 = ~pi159 & ~n27189;
  assign n31401 = ~pi158 & n31400;
  assign n31402 = ~n31399 & ~n31401;
  assign n31403 = pi157 & ~n31402;
  assign n31404 = ~pi158 & pi159;
  assign n31405 = ~pi159 & n27189;
  assign n31406 = pi158 & n31405;
  assign n31407 = ~n31404 & ~n31406;
  assign n31408 = ~pi157 & ~n31407;
  assign n31409 = ~n31403 & ~n31408;
  assign n31410 = ~n31398 & n31409;
  assign n31411 = ~n31392 & n31410;
  assign n31412 = pi321 & ~n31411;
  assign n31413 = pi317 & n23626;
  assign n31414 = n31412 & ~n31413;
  assign n31415 = n23626 & ~n31412;
  assign n31416 = pi317 & n31415;
  assign n31417 = ~n31414 & ~n31416;
  assign n31418 = ~n31386 & ~n31417;
  assign n31419 = ~n31412 & ~n31413;
  assign n31420 = n23626 & n31412;
  assign n31421 = pi317 & n31420;
  assign n31422 = ~n31419 & ~n31421;
  assign n31423 = n27198 & ~n31422;
  assign n31424 = pi319 & n31423;
  assign n31425 = ~n31418 & ~n31424;
  assign n31426 = ~n30458 & n30489;
  assign n31427 = ~n30464 & ~n31426;
  assign n31428 = pi321 & n31427;
  assign n31429 = n27198 & ~n30489;
  assign n31430 = pi320 & n31429;
  assign n31431 = ~n31428 & ~n31430;
  assign n31432 = n31425 & n31431;
  assign n31433 = ~n31425 & ~n31431;
  assign n31434 = ~n31432 & ~n31433;
  assign n31435 = n23069 & ~n30526;
  assign n31436 = pi317 & n31435;
  assign n31437 = pi320 & ~n30464;
  assign n31438 = ~n31436 & ~n31437;
  assign n31439 = n31436 & n31437;
  assign n31440 = ~n31438 & ~n31439;
  assign n31441 = n25479 & ~n31440;
  assign n31442 = pi318 & n31441;
  assign n31443 = pi318 & n25479;
  assign n31444 = n31436 & ~n31437;
  assign n31445 = ~n31436 & n31437;
  assign n31446 = ~n31444 & ~n31445;
  assign n31447 = ~n31443 & ~n31446;
  assign n31448 = ~n31442 & ~n31447;
  assign n31449 = ~n31434 & ~n31448;
  assign n31450 = n31425 & ~n31431;
  assign n31451 = ~n31425 & n31431;
  assign n31452 = ~n31450 & ~n31451;
  assign n31453 = n25479 & ~n31446;
  assign n31454 = pi318 & n31453;
  assign n31455 = ~n31440 & ~n31443;
  assign n31456 = ~n31454 & ~n31455;
  assign n31457 = ~n31452 & ~n31456;
  assign n31458 = ~n31449 & ~n31457;
  assign n31459 = ~n31385 & n31458;
  assign n31460 = n31385 & ~n31458;
  assign n31461 = ~n31459 & ~n31460;
  assign n31462 = n20347 & ~n31461;
  assign n31463 = pi315 & n31462;
  assign n31464 = pi315 & n20347;
  assign n31465 = n31385 & n31458;
  assign n31466 = ~n31385 & ~n31458;
  assign n31467 = ~n31465 & ~n31466;
  assign n31468 = ~n31464 & ~n31467;
  assign n31469 = ~n31463 & ~n31468;
  assign n31470 = n31356 & ~n31469;
  assign n31471 = ~n31356 & n31469;
  assign n31472 = ~n31470 & ~n31471;
  assign n31473 = ~n31351 & ~n31472;
  assign n31474 = ~n31356 & ~n31469;
  assign n31475 = n31356 & n31469;
  assign n31476 = ~n31474 & ~n31475;
  assign n31477 = n31346 & ~n31347;
  assign n31478 = n14618 & ~n31346;
  assign n31479 = pi311 & n31478;
  assign n31480 = ~n31477 & ~n31479;
  assign n31481 = ~n31476 & ~n31480;
  assign n31482 = ~n31473 & ~n31481;
  assign n31483 = n31343 & ~n31482;
  assign n31484 = ~n31343 & n31482;
  assign n31485 = ~n31483 & ~n31484;
  assign n31486 = ~n31335 & ~n31485;
  assign n31487 = ~n31343 & ~n31482;
  assign n31488 = n31343 & n31482;
  assign n31489 = ~n31487 & ~n31488;
  assign n31490 = ~n31330 & ~n31331;
  assign n31491 = n14156 & n31330;
  assign n31492 = pi310 & n31491;
  assign n31493 = ~n31490 & ~n31492;
  assign n31494 = ~n31489 & ~n31493;
  assign n31495 = ~n31486 & ~n31494;
  assign n31496 = pi306 & n9517;
  assign n31497 = ~n31495 & ~n31496;
  assign n31498 = n9517 & n31495;
  assign n31499 = pi306 & n31498;
  assign n31500 = ~n31497 & ~n31499;
  assign n31501 = ~n31319 & ~n31500;
  assign n31502 = ~n30742 & ~n30744;
  assign n31503 = ~n30743 & ~n31502;
  assign n31504 = n31495 & ~n31496;
  assign n31505 = n9517 & ~n31495;
  assign n31506 = pi306 & n31505;
  assign n31507 = ~n31504 & ~n31506;
  assign n31508 = ~n31503 & ~n31507;
  assign n31509 = ~n31501 & ~n31508;
  assign n31510 = ~n31317 & n31509;
  assign n31511 = n31317 & ~n31509;
  assign n31512 = ~n31510 & ~n31511;
  assign n31513 = n6777 & ~n31512;
  assign n31514 = pi303 & n31513;
  assign n31515 = pi303 & n6777;
  assign n31516 = n31317 & n31509;
  assign n31517 = ~n31317 & ~n31509;
  assign n31518 = ~n31516 & ~n31517;
  assign n31519 = ~n31515 & ~n31518;
  assign n31520 = ~n31514 & ~n31519;
  assign n31521 = pi301 & n4772;
  assign n31522 = ~n31520 & ~n31521;
  assign n31523 = n4772 & n31520;
  assign n31524 = pi301 & n31523;
  assign n31525 = ~n31522 & ~n31524;
  assign n31526 = ~n31306 & ~n31525;
  assign n31527 = n31520 & ~n31521;
  assign n31528 = n4772 & ~n31520;
  assign n31529 = pi301 & n31528;
  assign n31530 = ~n31527 & ~n31529;
  assign n31531 = n5463 & ~n31530;
  assign n31532 = pi302 & n31531;
  assign n31533 = ~n31526 & ~n31532;
  assign n31534 = n30772 & ~n30816;
  assign n31535 = ~n30772 & n30816;
  assign n31536 = n4086 & ~n31535;
  assign n31537 = pi301 & n31536;
  assign n31538 = ~n31534 & ~n31537;
  assign n31539 = n31533 & ~n31538;
  assign n31540 = ~n30817 & ~n31534;
  assign n31541 = ~n31535 & ~n31540;
  assign n31542 = ~n31533 & ~n31541;
  assign n31543 = ~n31539 & ~n31542;
  assign n31544 = ~n31305 & n31543;
  assign n31545 = n31305 & ~n31543;
  assign n31546 = ~n31544 & ~n31545;
  assign n31547 = n3552 & ~n31546;
  assign n31548 = pi299 & n31547;
  assign n31549 = pi299 & n3552;
  assign n31550 = n31305 & n31543;
  assign n31551 = ~n31305 & ~n31543;
  assign n31552 = ~n31550 & ~n31551;
  assign n31553 = ~n31549 & ~n31552;
  assign n31554 = ~n31548 & ~n31553;
  assign n31555 = pi298 & n3012;
  assign n31556 = ~n31554 & ~n31555;
  assign n31557 = n3012 & n31554;
  assign n31558 = pi298 & n31557;
  assign n31559 = ~n31556 & ~n31558;
  assign n31560 = n1533 & ~n27703;
  assign n31561 = pi297 & n31560;
  assign n31562 = ~n25923 & ~n30299;
  assign n31563 = ~n31561 & ~n31562;
  assign n31564 = ~n25367 & ~n31563;
  assign n31565 = n1840 & ~n27696;
  assign n31566 = ~n25923 & n31560;
  assign n31567 = ~n31565 & ~n31566;
  assign n31568 = pi297 & ~n31567;
  assign n31569 = ~n31564 & ~n31568;
  assign n31570 = ~n30871 & ~n31569;
  assign n31571 = n30871 & n31569;
  assign n31572 = n30298 & ~n31571;
  assign n31573 = ~n31570 & ~n31572;
  assign n31574 = ~n31559 & ~n31573;
  assign n31575 = n31554 & ~n31555;
  assign n31576 = n3012 & ~n31554;
  assign n31577 = pi298 & n31576;
  assign n31578 = ~n31575 & ~n31577;
  assign n31579 = ~n30298 & ~n31570;
  assign n31580 = ~n31571 & ~n31579;
  assign n31581 = ~n31578 & ~n31580;
  assign n31582 = ~n31574 & ~n31581;
  assign n31583 = n1553 & ~n30942;
  assign n31584 = pi294 & n31583;
  assign n31585 = ~n30943 & ~n31584;
  assign n31586 = ~n31582 & ~n31585;
  assign n31587 = ~n30941 & ~n30943;
  assign n31588 = ~n30942 & ~n31587;
  assign n31589 = n31582 & ~n31588;
  assign n31590 = ~n31586 & ~n31589;
  assign n31591 = ~n31291 & ~n31590;
  assign n31592 = n31291 & n31590;
  assign n31593 = ~n31591 & ~n31592;
  assign n31594 = ~n31084 & ~n31593;
  assign n31595 = n31291 & ~n31590;
  assign n31596 = ~n31291 & n31590;
  assign n31597 = ~n31595 & ~n31596;
  assign n31598 = n31060 & ~n31082;
  assign n31599 = ~n31060 & ~n31078;
  assign n31600 = ~n31598 & ~n31599;
  assign n31601 = ~n31597 & ~n31600;
  assign n31602 = ~n31594 & ~n31601;
  assign n31603 = n31055 & ~n31602;
  assign n31604 = ~n31055 & n31602;
  assign n31605 = ~n31603 & ~n31604;
  assign n31606 = n30257 & n30979;
  assign n31607 = ~n30257 & ~n30979;
  assign n31608 = pi288 & ~n31607;
  assign n31609 = ~n31606 & ~n31608;
  assign n31610 = ~n31605 & ~n31609;
  assign n31611 = ~n31055 & ~n31602;
  assign n31612 = n31055 & n31602;
  assign n31613 = ~n31611 & ~n31612;
  assign n31614 = ~pi288 & ~n31606;
  assign n31615 = ~n31607 & ~n31614;
  assign n31616 = ~n31613 & ~n31615;
  assign n31617 = ~n31610 & ~n31616;
  assign n31618 = ~n1256 & ~n29042;
  assign n31619 = pi350 & n31618;
  assign n31620 = n1256 & ~n29039;
  assign n31621 = ~n29041 & n31620;
  assign n31622 = pi350 & ~n31621;
  assign n31623 = n30229 & n31622;
  assign n31624 = pi258 & ~n31623;
  assign n31625 = pi128 & n31624;
  assign n31626 = ~n31619 & n31625;
  assign n31627 = pi353 & n31626;
  assign n31628 = pi353 & n1156;
  assign n31629 = ~n31619 & ~n31623;
  assign n31630 = ~n31628 & ~n31629;
  assign n31631 = ~n31627 & ~n31630;
  assign n31632 = n29071 & n30189;
  assign n31633 = ~n29071 & ~n30189;
  assign n31634 = ~n31632 & ~n31633;
  assign n31635 = n29089 & ~n30208;
  assign n31636 = ~n29089 & n30208;
  assign n31637 = ~n31635 & ~n31636;
  assign n31638 = n29085 & ~n30193;
  assign n31639 = ~n31637 & ~n31638;
  assign n31640 = ~n31634 & n31639;
  assign n31641 = ~n29085 & n30193;
  assign n31642 = n29071 & ~n30189;
  assign n31643 = ~n29071 & n30189;
  assign n31644 = ~n31642 & ~n31643;
  assign n31645 = ~n29089 & ~n30208;
  assign n31646 = n29089 & n30208;
  assign n31647 = ~n31645 & ~n31646;
  assign n31648 = ~n31638 & ~n31647;
  assign n31649 = ~n31644 & n31648;
  assign n31650 = ~n31641 & ~n31649;
  assign n31651 = ~n31640 & n31650;
  assign n31652 = ~n30154 & ~n30177;
  assign n31653 = ~n30184 & n31652;
  assign n31654 = ~n30175 & ~n30177;
  assign n31655 = ~n30137 & n31654;
  assign n31656 = ~n30176 & ~n31655;
  assign n31657 = ~n31653 & n31656;
  assign n31658 = pi345 & n4596;
  assign n31659 = n31657 & ~n31658;
  assign n31660 = n4596 & ~n31657;
  assign n31661 = pi345 & n31660;
  assign n31662 = ~n31659 & ~n31661;
  assign n31663 = n30134 & ~n30138;
  assign n31664 = ~n30134 & n30138;
  assign n31665 = ~n30127 & n30151;
  assign n31666 = n30127 & ~n30151;
  assign n31667 = ~n31665 & ~n31666;
  assign n31668 = ~n31664 & ~n31667;
  assign n31669 = ~n31663 & ~n31668;
  assign n31670 = n5257 & ~n31669;
  assign n31671 = pi344 & n31670;
  assign n31672 = pi344 & n5257;
  assign n31673 = ~n30127 & ~n30151;
  assign n31674 = n30127 & n30151;
  assign n31675 = ~n31673 & ~n31674;
  assign n31676 = ~n31672 & ~n31675;
  assign n31677 = ~n31663 & n31676;
  assign n31678 = ~n30134 & ~n31672;
  assign n31679 = n30138 & n31678;
  assign n31680 = ~n31677 & ~n31679;
  assign n31681 = ~n31671 & n31680;
  assign n31682 = ~n29093 & n30082;
  assign n31683 = n29093 & ~n30082;
  assign n31684 = ~n31682 & ~n31683;
  assign n31685 = n29117 & ~n31684;
  assign n31686 = ~n29093 & ~n30082;
  assign n31687 = n29093 & n30082;
  assign n31688 = ~n31686 & ~n31687;
  assign n31689 = ~n29117 & ~n31688;
  assign n31690 = ~n31685 & ~n31689;
  assign n31691 = n27872 & ~n29106;
  assign n31692 = ~n27872 & ~n29096;
  assign n31693 = ~n31691 & ~n31692;
  assign n31694 = ~n30088 & ~n31693;
  assign n31695 = ~n30091 & ~n31694;
  assign n31696 = ~n30087 & n31695;
  assign n31697 = ~n31690 & ~n31696;
  assign n31698 = n30087 & ~n31695;
  assign n31699 = ~n31697 & ~n31698;
  assign n31700 = n29117 & ~n31683;
  assign n31701 = ~n31682 & ~n31700;
  assign n31702 = n29121 & n29982;
  assign n31703 = ~n29121 & ~n29982;
  assign n31704 = ~n31702 & ~n31703;
  assign n31705 = n29145 & ~n30006;
  assign n31706 = ~n29145 & n30006;
  assign n31707 = ~n31705 & ~n31706;
  assign n31708 = n29141 & ~n29986;
  assign n31709 = ~n31707 & ~n31708;
  assign n31710 = ~n31704 & n31709;
  assign n31711 = ~n29141 & n29986;
  assign n31712 = n29121 & ~n29982;
  assign n31713 = ~n29121 & n29982;
  assign n31714 = ~n31712 & ~n31713;
  assign n31715 = ~n29145 & ~n30006;
  assign n31716 = n29145 & n30006;
  assign n31717 = ~n31715 & ~n31716;
  assign n31718 = ~n31708 & ~n31717;
  assign n31719 = ~n31714 & n31718;
  assign n31720 = ~n31711 & ~n31719;
  assign n31721 = ~n31710 & n31720;
  assign n31722 = ~n29954 & ~n29970;
  assign n31723 = ~n29977 & n31722;
  assign n31724 = ~n29968 & ~n29970;
  assign n31725 = ~n29937 & n31724;
  assign n31726 = ~n29969 & ~n31725;
  assign n31727 = ~n31723 & n31726;
  assign n31728 = pi333 & n13762;
  assign n31729 = n31727 & ~n31728;
  assign n31730 = n13762 & ~n31727;
  assign n31731 = pi333 & n31730;
  assign n31732 = ~n31729 & ~n31731;
  assign n31733 = n29934 & ~n29938;
  assign n31734 = ~n29934 & n29938;
  assign n31735 = ~n29927 & n29951;
  assign n31736 = n29927 & ~n29951;
  assign n31737 = ~n31735 & ~n31736;
  assign n31738 = ~n31734 & ~n31737;
  assign n31739 = ~n31733 & ~n31738;
  assign n31740 = n18461 & ~n31739;
  assign n31741 = pi332 & n31740;
  assign n31742 = pi332 & n18461;
  assign n31743 = ~n29927 & ~n29951;
  assign n31744 = n29927 & n29951;
  assign n31745 = ~n31743 & ~n31744;
  assign n31746 = ~n31742 & ~n31745;
  assign n31747 = ~n31733 & n31746;
  assign n31748 = ~n29934 & ~n31742;
  assign n31749 = n29938 & n31748;
  assign n31750 = ~n31747 & ~n31749;
  assign n31751 = ~n31741 & n31750;
  assign n31752 = n29196 & n29880;
  assign n31753 = n21479 & ~n31752;
  assign n31754 = ~n26706 & n31753;
  assign n31755 = ~n21479 & n29196;
  assign n31756 = n21479 & ~n29196;
  assign n31757 = n29880 & ~n31756;
  assign n31758 = ~n31755 & ~n31757;
  assign n31759 = n26706 & ~n31758;
  assign n31760 = ~n31754 & ~n31759;
  assign n31761 = pi327 & ~n31760;
  assign n31762 = pi327 & n26706;
  assign n31763 = ~n29196 & ~n31762;
  assign n31764 = ~n29880 & n31763;
  assign n31765 = ~n31761 & ~n31764;
  assign n31766 = ~n29160 & ~n29906;
  assign n31767 = n29160 & n29906;
  assign n31768 = ~n31766 & ~n31767;
  assign n31769 = ~n29217 & n29859;
  assign n31770 = n29217 & ~n29859;
  assign n31771 = ~n29857 & ~n31770;
  assign n31772 = ~n31769 & ~n31771;
  assign n31773 = n29173 & ~n29912;
  assign n31774 = ~n31772 & ~n31773;
  assign n31775 = ~n29192 & n31774;
  assign n31776 = ~n29173 & n29912;
  assign n31777 = n31772 & ~n31776;
  assign n31778 = n29192 & n31777;
  assign n31779 = ~n31775 & ~n31778;
  assign n31780 = ~n31768 & ~n31779;
  assign n31781 = ~n29160 & n29906;
  assign n31782 = n29160 & ~n29906;
  assign n31783 = ~n31781 & ~n31782;
  assign n31784 = ~n29192 & n31777;
  assign n31785 = n29192 & n31774;
  assign n31786 = ~n31784 & ~n31785;
  assign n31787 = ~n31783 & ~n31786;
  assign n31788 = ~n29173 & ~n31772;
  assign n31789 = n29912 & n31788;
  assign n31790 = n29173 & n31772;
  assign n31791 = ~n29912 & n31790;
  assign n31792 = ~n31789 & ~n31791;
  assign n31793 = ~n31787 & n31792;
  assign n31794 = ~n31780 & n31793;
  assign n31795 = n31765 & n31794;
  assign n31796 = ~n31765 & ~n31794;
  assign n31797 = ~n31795 & ~n31796;
  assign n31798 = ~n29181 & ~n29188;
  assign n31799 = n29177 & ~n31798;
  assign n31800 = ~n29177 & n31798;
  assign n31801 = ~n31783 & ~n31800;
  assign n31802 = ~n31799 & ~n31801;
  assign n31803 = ~n31797 & ~n31802;
  assign n31804 = n31765 & ~n31794;
  assign n31805 = ~n31765 & n31794;
  assign n31806 = ~n31804 & ~n31805;
  assign n31807 = ~n31768 & ~n31799;
  assign n31808 = ~n31800 & ~n31807;
  assign n31809 = ~n31806 & ~n31808;
  assign n31810 = ~n31803 & ~n31809;
  assign n31811 = ~n31751 & ~n31810;
  assign n31812 = n31751 & n31810;
  assign n31813 = ~n31811 & ~n31812;
  assign n31814 = ~n31732 & ~n31813;
  assign n31815 = n31751 & ~n31810;
  assign n31816 = ~n31751 & n31810;
  assign n31817 = ~n31815 & ~n31816;
  assign n31818 = ~n31727 & ~n31728;
  assign n31819 = n13762 & n31727;
  assign n31820 = pi333 & n31819;
  assign n31821 = ~n31818 & ~n31820;
  assign n31822 = ~n31817 & ~n31821;
  assign n31823 = ~n31814 & ~n31822;
  assign n31824 = n31721 & ~n31823;
  assign n31825 = ~n31721 & n31823;
  assign n31826 = ~n31824 & ~n31825;
  assign n31827 = n6556 & ~n30039;
  assign n31828 = ~n30040 & ~n31827;
  assign n31829 = n9205 & ~n31828;
  assign n31830 = pi338 & n31829;
  assign n31831 = pi337 & n11366;
  assign n31832 = ~n9205 & ~n31827;
  assign n31833 = pi338 & ~n31832;
  assign n31834 = ~n30040 & ~n31833;
  assign n31835 = n30027 & ~n31834;
  assign n31836 = ~n31831 & ~n31835;
  assign n31837 = ~n31830 & n31836;
  assign n31838 = ~n31830 & ~n31835;
  assign n31839 = n31831 & ~n31838;
  assign n31840 = ~n31837 & ~n31839;
  assign n31841 = ~n31826 & ~n31840;
  assign n31842 = n31721 & n31823;
  assign n31843 = ~n31721 & ~n31823;
  assign n31844 = ~n31842 & ~n31843;
  assign n31845 = n31831 & ~n31835;
  assign n31846 = ~n31830 & n31845;
  assign n31847 = ~n31831 & ~n31838;
  assign n31848 = ~n31846 & ~n31847;
  assign n31849 = ~n31844 & ~n31848;
  assign n31850 = ~n31841 & ~n31849;
  assign n31851 = pi340 & n6556;
  assign n31852 = ~n31850 & ~n31851;
  assign n31853 = n6556 & n31850;
  assign n31854 = pi340 & n31853;
  assign n31855 = ~n31852 & ~n31854;
  assign n31856 = ~n31701 & ~n31855;
  assign n31857 = ~n29117 & ~n31682;
  assign n31858 = ~n31683 & ~n31857;
  assign n31859 = n31850 & ~n31851;
  assign n31860 = n6556 & ~n31850;
  assign n31861 = pi340 & n31860;
  assign n31862 = ~n31859 & ~n31861;
  assign n31863 = ~n31858 & ~n31862;
  assign n31864 = ~n31856 & ~n31863;
  assign n31865 = ~n31699 & n31864;
  assign n31866 = n31699 & ~n31864;
  assign n31867 = ~n31865 & ~n31866;
  assign n31868 = pi341 & n5973;
  assign n31869 = pi342 & n5732;
  assign n31870 = ~n31868 & ~n31869;
  assign n31871 = pi341 & pi342;
  assign n31872 = n5976 & n31871;
  assign n31873 = ~n31870 & ~n31872;
  assign n31874 = ~n31867 & ~n31873;
  assign n31875 = ~n31699 & ~n31864;
  assign n31876 = n31699 & n31864;
  assign n31877 = ~n31875 & ~n31876;
  assign n31878 = n5973 & ~n31869;
  assign n31879 = pi341 & n31878;
  assign n31880 = n5732 & ~n31868;
  assign n31881 = pi342 & n31880;
  assign n31882 = ~n31879 & ~n31881;
  assign n31883 = ~n31877 & ~n31882;
  assign n31884 = ~n31874 & ~n31883;
  assign n31885 = ~n31681 & ~n31884;
  assign n31886 = n31681 & n31884;
  assign n31887 = ~n31885 & ~n31886;
  assign n31888 = ~n31662 & ~n31887;
  assign n31889 = n31681 & ~n31884;
  assign n31890 = ~n31681 & n31884;
  assign n31891 = ~n31889 & ~n31890;
  assign n31892 = ~n31657 & ~n31658;
  assign n31893 = n4596 & n31657;
  assign n31894 = pi345 & n31893;
  assign n31895 = ~n31892 & ~n31894;
  assign n31896 = ~n31891 & ~n31895;
  assign n31897 = ~n31888 & ~n31896;
  assign n31898 = pi348 & n30202;
  assign n31899 = ~n29078 & ~n30195;
  assign n31900 = ~n31898 & ~n31899;
  assign n31901 = n1729 & ~n31900;
  assign n31902 = pi348 & n31901;
  assign n31903 = n29089 & ~n31644;
  assign n31904 = ~n29089 & ~n31634;
  assign n31905 = ~n31903 & ~n31904;
  assign n31906 = pi348 & n1729;
  assign n31907 = n31900 & ~n31906;
  assign n31908 = ~n31905 & ~n31907;
  assign n31909 = ~n31902 & ~n31908;
  assign n31910 = ~n31897 & n31909;
  assign n31911 = n31897 & ~n31909;
  assign n31912 = ~n31910 & ~n31911;
  assign n31913 = ~n31651 & ~n31912;
  assign n31914 = ~n31897 & ~n31909;
  assign n31915 = n31897 & n31909;
  assign n31916 = ~n31914 & ~n31915;
  assign n31917 = n31651 & ~n31916;
  assign n31918 = ~n31913 & ~n31917;
  assign n31919 = pi348 & n2091;
  assign n31920 = n2464 & ~n31919;
  assign n31921 = pi347 & n31920;
  assign n31922 = pi347 & n2464;
  assign n31923 = n2091 & ~n31922;
  assign n31924 = pi348 & n31923;
  assign n31925 = ~n31921 & ~n31924;
  assign n31926 = n29089 & ~n31642;
  assign n31927 = ~n31643 & ~n31926;
  assign n31928 = n29117 & ~n30106;
  assign n31929 = ~n29117 & n30106;
  assign n31930 = ~n31928 & ~n31929;
  assign n31931 = n29113 & ~n30086;
  assign n31932 = ~n31930 & ~n31931;
  assign n31933 = ~n31688 & n31932;
  assign n31934 = ~n29113 & n30086;
  assign n31935 = ~n29117 & ~n30106;
  assign n31936 = n29117 & n30106;
  assign n31937 = ~n31935 & ~n31936;
  assign n31938 = ~n31931 & ~n31937;
  assign n31939 = ~n31684 & n31938;
  assign n31940 = ~n31934 & ~n31939;
  assign n31941 = ~n31933 & n31940;
  assign n31942 = ~n30054 & ~n30070;
  assign n31943 = ~n30077 & n31942;
  assign n31944 = ~n30068 & ~n30070;
  assign n31945 = ~n30037 & n31944;
  assign n31946 = ~n30069 & ~n31945;
  assign n31947 = ~n31943 & n31946;
  assign n31948 = pi339 & n9205;
  assign n31949 = n31947 & ~n31948;
  assign n31950 = n9205 & ~n31947;
  assign n31951 = pi339 & n31950;
  assign n31952 = ~n31949 & ~n31951;
  assign n31953 = n30034 & ~n30038;
  assign n31954 = ~n30034 & n30038;
  assign n31955 = ~n30027 & n30051;
  assign n31956 = n30027 & ~n30051;
  assign n31957 = ~n31955 & ~n31956;
  assign n31958 = ~n31954 & ~n31957;
  assign n31959 = ~n31953 & ~n31958;
  assign n31960 = n10561 & ~n31959;
  assign n31961 = pi338 & n31960;
  assign n31962 = pi338 & n10561;
  assign n31963 = ~n30027 & ~n30051;
  assign n31964 = n30027 & n30051;
  assign n31965 = ~n31963 & ~n31964;
  assign n31966 = ~n31962 & ~n31965;
  assign n31967 = ~n31953 & n31966;
  assign n31968 = ~n30034 & ~n31962;
  assign n31969 = n30038 & n31968;
  assign n31970 = ~n31967 & ~n31969;
  assign n31971 = ~n31961 & n31970;
  assign n31972 = ~n29145 & ~n31713;
  assign n31973 = ~n31712 & ~n31972;
  assign n31974 = n12917 & ~n31973;
  assign n31975 = pi334 & n31974;
  assign n31976 = pi334 & n12917;
  assign n31977 = ~n29121 & n29145;
  assign n31978 = n29121 & ~n29145;
  assign n31979 = n29982 & ~n31978;
  assign n31980 = ~n31977 & ~n31979;
  assign n31981 = ~n31976 & ~n31980;
  assign n31982 = ~n31975 & ~n31981;
  assign n31983 = n28721 & n29927;
  assign n31984 = n28735 & n31983;
  assign n31985 = ~n13762 & ~n29927;
  assign n31986 = ~n29939 & ~n31985;
  assign n31987 = n12917 & n31986;
  assign n31988 = ~n29927 & ~n29940;
  assign n31989 = n13762 & ~n31988;
  assign n31990 = ~n31987 & ~n31989;
  assign n31991 = pi332 & ~n31990;
  assign n31992 = ~n31984 & ~n31991;
  assign n31993 = pi331 & n19539;
  assign n31994 = ~n31992 & ~n31993;
  assign n31995 = n19539 & n31992;
  assign n31996 = pi331 & n31995;
  assign n31997 = ~n31994 & ~n31996;
  assign n31998 = ~n29247 & ~n29823;
  assign n31999 = n29247 & n29822;
  assign n32000 = pi322 & n31999;
  assign n32001 = ~n31998 & ~n32000;
  assign n32002 = ~n29251 & ~n32001;
  assign n32003 = n29247 & ~n29823;
  assign n32004 = ~n29247 & n29822;
  assign n32005 = pi322 & n32004;
  assign n32006 = ~n32003 & ~n32005;
  assign n32007 = n28628 & ~n32006;
  assign n32008 = pi323 & n32007;
  assign n32009 = ~n32002 & ~n32008;
  assign n32010 = n29854 & n32009;
  assign n32011 = ~pi325 & ~n32010;
  assign n32012 = pi324 & n32011;
  assign n32013 = ~n29854 & ~n32009;
  assign n32014 = ~pi324 & ~n32013;
  assign n32015 = ~n32010 & ~n32014;
  assign n32016 = pi325 & ~n32015;
  assign n32017 = ~n32012 & ~n32016;
  assign n32018 = n28010 & ~n32017;
  assign n32019 = pi325 & n28010;
  assign n32020 = ~n29854 & ~n32019;
  assign n32021 = ~n32009 & n32020;
  assign n32022 = ~n32018 & ~n32021;
  assign n32023 = pi330 & n19557;
  assign n32024 = n32022 & ~n32023;
  assign n32025 = n19557 & ~n32022;
  assign n32026 = pi330 & n32025;
  assign n32027 = ~n32024 & ~n32026;
  assign n32028 = ~n29160 & ~n29209;
  assign n32029 = n29884 & n32028;
  assign n32030 = ~n29196 & ~n29880;
  assign n32031 = ~n31752 & ~n32030;
  assign n32032 = n21479 & ~n32031;
  assign n32033 = pi327 & n32032;
  assign n32034 = n29196 & ~n29880;
  assign n32035 = ~n29196 & n29880;
  assign n32036 = ~n32034 & ~n32035;
  assign n32037 = ~n29213 & ~n32036;
  assign n32038 = ~n32033 & ~n32037;
  assign n32039 = ~n29160 & n29884;
  assign n32040 = n29160 & ~n29884;
  assign n32041 = ~n29209 & ~n32040;
  assign n32042 = ~n32039 & ~n32041;
  assign n32043 = ~n32038 & ~n32042;
  assign n32044 = ~n32029 & ~n32043;
  assign n32045 = n29885 & ~n32044;
  assign n32046 = n29160 & n29209;
  assign n32047 = n32038 & n32046;
  assign n32048 = ~n32028 & n32038;
  assign n32049 = ~n32046 & ~n32048;
  assign n32050 = ~n29885 & ~n32049;
  assign n32051 = ~n32047 & ~n32050;
  assign n32052 = ~n29884 & ~n32051;
  assign n32053 = ~n29885 & n32038;
  assign n32054 = n32046 & n32053;
  assign n32055 = ~n29209 & ~n32038;
  assign n32056 = n32039 & n32055;
  assign n32057 = ~n32054 & ~n32056;
  assign n32058 = ~n32052 & n32057;
  assign n32059 = ~n32045 & n32058;
  assign n32060 = n28628 & ~n29247;
  assign n32061 = pi323 & n32060;
  assign n32062 = n29247 & ~n29251;
  assign n32063 = n29822 & ~n32062;
  assign n32064 = pi322 & n32063;
  assign n32065 = ~n32061 & ~n32064;
  assign n32066 = n29785 & n29794;
  assign n32067 = ~n29785 & ~n29794;
  assign n32068 = ~n32066 & ~n32067;
  assign n32069 = ~n29714 & n29722;
  assign n32070 = n29714 & ~n29722;
  assign n32071 = n29252 & ~n32070;
  assign n32072 = ~n32069 & ~n32071;
  assign n32073 = n29254 & ~n29626;
  assign n32074 = ~n29254 & n29626;
  assign n32075 = n29610 & ~n32074;
  assign n32076 = ~n32073 & ~n32075;
  assign n32077 = pi139 & pi278;
  assign n32078 = pi137 & pi280;
  assign n32079 = pi133 & pi284;
  assign n32080 = pi286 & ~n29307;
  assign n32081 = pi130 & n32080;
  assign n32082 = ~n29292 & n29307;
  assign n32083 = ~n29295 & ~n32082;
  assign n32084 = ~n32081 & ~n32083;
  assign n32085 = n32079 & ~n32084;
  assign n32086 = ~n29289 & n29307;
  assign n32087 = ~n29287 & ~n29307;
  assign n32088 = ~n29288 & n32087;
  assign n32089 = ~n29292 & ~n32088;
  assign n32090 = ~n32086 & ~n32089;
  assign n32091 = ~n32079 & ~n32090;
  assign n32092 = ~n32085 & ~n32091;
  assign n32093 = pi282 & n32092;
  assign n32094 = pi135 & n32093;
  assign n32095 = pi135 & pi282;
  assign n32096 = ~n32092 & ~n32095;
  assign n32097 = ~n32094 & ~n32096;
  assign n32098 = ~n32078 & ~n32097;
  assign n32099 = pi282 & ~n32092;
  assign n32100 = pi135 & n32099;
  assign n32101 = n32092 & ~n32095;
  assign n32102 = ~n32100 & ~n32101;
  assign n32103 = pi280 & ~n32102;
  assign n32104 = pi137 & n32103;
  assign n32105 = ~n32098 & ~n32104;
  assign n32106 = ~n32077 & n32105;
  assign n32107 = n32077 & ~n32105;
  assign n32108 = ~n32106 & ~n32107;
  assign n32109 = n29256 & n29522;
  assign n32110 = ~n29256 & ~n29522;
  assign n32111 = ~n29506 & ~n32110;
  assign n32112 = ~n32109 & ~n32111;
  assign n32113 = n29463 & n29486;
  assign n32114 = ~n29454 & n29470;
  assign n32115 = n29454 & ~n29470;
  assign n32116 = ~n32114 & ~n32115;
  assign n32117 = n29257 & ~n32116;
  assign n32118 = ~n29454 & ~n29470;
  assign n32119 = n29454 & n29470;
  assign n32120 = ~n32118 & ~n32119;
  assign n32121 = ~n29257 & ~n32120;
  assign n32122 = ~n32117 & ~n32121;
  assign n32123 = ~n29463 & ~n29486;
  assign n32124 = ~n32122 & ~n32123;
  assign n32125 = ~n32113 & ~n32124;
  assign n32126 = n32112 & ~n32125;
  assign n32127 = ~n32112 & n32125;
  assign n32128 = ~n32126 & ~n32127;
  assign n32129 = pi271 & ~n32128;
  assign n32130 = pi146 & n32129;
  assign n32131 = pi146 & pi271;
  assign n32132 = ~n32112 & ~n32125;
  assign n32133 = n32112 & n32125;
  assign n32134 = ~n32132 & ~n32133;
  assign n32135 = ~n32131 & ~n32134;
  assign n32136 = ~n32130 & ~n32135;
  assign n32137 = ~n32108 & ~n32136;
  assign n32138 = ~n32077 & ~n32105;
  assign n32139 = n32077 & n32105;
  assign n32140 = ~n32138 & ~n32139;
  assign n32141 = pi271 & ~n32134;
  assign n32142 = pi146 & n32141;
  assign n32143 = ~n32128 & ~n32131;
  assign n32144 = ~n32142 & ~n32143;
  assign n32145 = ~n32140 & ~n32144;
  assign n32146 = ~n32137 & ~n32145;
  assign n32147 = ~n32076 & n32146;
  assign n32148 = n32076 & ~n32146;
  assign n32149 = ~n32147 & ~n32148;
  assign n32150 = pi148 & pi150;
  assign n32151 = pi267 & pi269;
  assign n32152 = n32150 & n32151;
  assign n32153 = pi150 & pi267;
  assign n32154 = pi148 & pi269;
  assign n32155 = ~n32153 & ~n32154;
  assign n32156 = ~n32152 & ~n32155;
  assign n32157 = ~n32149 & ~n32156;
  assign n32158 = ~n32076 & ~n32146;
  assign n32159 = n32076 & n32146;
  assign n32160 = ~n32158 & ~n32159;
  assign n32161 = pi269 & ~n32153;
  assign n32162 = pi148 & n32161;
  assign n32163 = pi267 & ~n32154;
  assign n32164 = pi150 & n32163;
  assign n32165 = ~n32162 & ~n32164;
  assign n32166 = ~n32160 & ~n32165;
  assign n32167 = ~n32157 & ~n32166;
  assign n32168 = n29253 & ~n29678;
  assign n32169 = ~n29253 & n29678;
  assign n32170 = n29662 & ~n32169;
  assign n32171 = ~n32168 & ~n32170;
  assign n32172 = n32167 & ~n32171;
  assign n32173 = ~n29662 & n29678;
  assign n32174 = n29662 & ~n29678;
  assign n32175 = ~n29253 & ~n32174;
  assign n32176 = ~n32173 & ~n32175;
  assign n32177 = ~n32167 & ~n32176;
  assign n32178 = ~n32172 & ~n32177;
  assign n32179 = pi157 & pi260;
  assign n32180 = n32178 & ~n32179;
  assign n32181 = pi260 & ~n32178;
  assign n32182 = pi157 & n32181;
  assign n32183 = ~n32180 & ~n32182;
  assign n32184 = ~n32072 & ~n32183;
  assign n32185 = ~n29252 & ~n32069;
  assign n32186 = ~n32070 & ~n32185;
  assign n32187 = ~n32178 & ~n32179;
  assign n32188 = pi260 & n32178;
  assign n32189 = pi157 & n32188;
  assign n32190 = ~n32187 & ~n32189;
  assign n32191 = ~n32186 & ~n32190;
  assign n32192 = ~n32184 & ~n32191;
  assign n32193 = n29766 & n32192;
  assign n32194 = ~n29766 & ~n32192;
  assign n32195 = n29784 & n32194;
  assign n32196 = ~n32193 & ~n32195;
  assign n32197 = ~n32068 & ~n32196;
  assign n32198 = ~n29784 & n32192;
  assign n32199 = n29785 & ~n29794;
  assign n32200 = ~n29785 & n29794;
  assign n32201 = ~n32199 & ~n32200;
  assign n32202 = ~n29766 & n32192;
  assign n32203 = n29766 & ~n32192;
  assign n32204 = n29784 & n32203;
  assign n32205 = ~n32202 & ~n32204;
  assign n32206 = ~n32201 & ~n32205;
  assign n32207 = ~n32198 & ~n32206;
  assign n32208 = ~n32197 & n32207;
  assign n32209 = n29718 & ~n29743;
  assign n32210 = ~n32069 & ~n32070;
  assign n32211 = n29252 & ~n32210;
  assign n32212 = ~n29714 & ~n29722;
  assign n32213 = n29714 & n29722;
  assign n32214 = ~n32212 & ~n32213;
  assign n32215 = ~n29252 & ~n32214;
  assign n32216 = ~n32211 & ~n32215;
  assign n32217 = ~n29718 & n29743;
  assign n32218 = ~n32216 & ~n32217;
  assign n32219 = ~n32209 & ~n32218;
  assign n32220 = ~n29610 & n29626;
  assign n32221 = n29610 & ~n29626;
  assign n32222 = ~n32220 & ~n32221;
  assign n32223 = pi268 & ~n32222;
  assign n32224 = pi148 & n32223;
  assign n32225 = n29610 & n29626;
  assign n32226 = ~n29610 & ~n29626;
  assign n32227 = ~n32225 & ~n32226;
  assign n32228 = ~n29254 & ~n32227;
  assign n32229 = ~n32224 & ~n32228;
  assign n32230 = ~n29642 & ~n32229;
  assign n32231 = n29642 & n32229;
  assign n32232 = n29620 & ~n32231;
  assign n32233 = ~n32230 & ~n32232;
  assign n32234 = n29515 & n29538;
  assign n32235 = ~n29506 & n29522;
  assign n32236 = n29506 & ~n29522;
  assign n32237 = ~n32235 & ~n32236;
  assign n32238 = n29256 & ~n32237;
  assign n32239 = ~n29506 & ~n29522;
  assign n32240 = n29506 & n29522;
  assign n32241 = ~n32239 & ~n32240;
  assign n32242 = ~n29256 & ~n32241;
  assign n32243 = ~n32238 & ~n32242;
  assign n32244 = ~n29515 & ~n29538;
  assign n32245 = ~n32243 & ~n32244;
  assign n32246 = ~n32234 & ~n32245;
  assign n32247 = n29412 & ~n29434;
  assign n32248 = ~n29402 & n29418;
  assign n32249 = n29402 & ~n29418;
  assign n32250 = ~n32248 & ~n32249;
  assign n32251 = n29258 & ~n32250;
  assign n32252 = ~n29402 & ~n29418;
  assign n32253 = n29402 & n29418;
  assign n32254 = ~n32252 & ~n32253;
  assign n32255 = ~n29258 & ~n32254;
  assign n32256 = ~n32251 & ~n32255;
  assign n32257 = ~n29412 & n29434;
  assign n32258 = ~n32256 & ~n32257;
  assign n32259 = ~n32247 & ~n32258;
  assign n32260 = pi287 & ~n29279;
  assign n32261 = pi129 & n32260;
  assign n32262 = n29279 & ~n29280;
  assign n32263 = pi288 & ~n32262;
  assign n32264 = pi128 & n32263;
  assign n32265 = ~n32261 & ~n32264;
  assign n32266 = n28041 & ~n28106;
  assign n32267 = ~n28041 & n28106;
  assign n32268 = n29320 & ~n32267;
  assign n32269 = ~n32266 & ~n32268;
  assign n32270 = n29266 & ~n32269;
  assign n32271 = ~n29266 & n32269;
  assign n32272 = n29313 & ~n32271;
  assign n32273 = ~n32270 & ~n32272;
  assign n32274 = ~n32265 & n32273;
  assign n32275 = n32265 & ~n32273;
  assign n32276 = ~n32274 & ~n32275;
  assign n32277 = n29265 & ~n29364;
  assign n32278 = n29338 & ~n29348;
  assign n32279 = ~n29338 & n29348;
  assign n32280 = ~n32278 & ~n32279;
  assign n32281 = ~n29265 & n29364;
  assign n32282 = ~n32280 & ~n32281;
  assign n32283 = ~n32277 & ~n32282;
  assign n32284 = pi286 & n32283;
  assign n32285 = pi131 & n32284;
  assign n32286 = pi131 & pi286;
  assign n32287 = ~n32283 & ~n32286;
  assign n32288 = ~n32285 & ~n32287;
  assign n32289 = ~n32276 & ~n32288;
  assign n32290 = n32265 & n32273;
  assign n32291 = ~n32265 & ~n32273;
  assign n32292 = ~n32290 & ~n32291;
  assign n32293 = n32283 & ~n32286;
  assign n32294 = pi286 & ~n32283;
  assign n32295 = pi131 & n32294;
  assign n32296 = ~n32293 & ~n32295;
  assign n32297 = ~n32292 & ~n32296;
  assign n32298 = ~n32289 & ~n32297;
  assign n32299 = n28174 & n28179;
  assign n32300 = ~n28174 & ~n28179;
  assign n32301 = n28170 & ~n32300;
  assign n32302 = ~n32299 & ~n32301;
  assign n32303 = n29386 & ~n32302;
  assign n32304 = ~n29386 & n32302;
  assign n32305 = ~n29397 & ~n32304;
  assign n32306 = ~n32303 & ~n32305;
  assign n32307 = n32298 & ~n32306;
  assign n32308 = ~n29385 & ~n32303;
  assign n32309 = ~n32304 & ~n32308;
  assign n32310 = ~n32298 & ~n32309;
  assign n32311 = ~n32307 & ~n32310;
  assign n32312 = n32259 & n32311;
  assign n32313 = ~n32259 & ~n32311;
  assign n32314 = ~n32312 & ~n32313;
  assign n32315 = pi141 & pi143;
  assign n32316 = pi274 & pi276;
  assign n32317 = n32315 & n32316;
  assign n32318 = pi143 & pi274;
  assign n32319 = pi141 & pi276;
  assign n32320 = ~n32318 & ~n32319;
  assign n32321 = ~n32317 & ~n32320;
  assign n32322 = ~n32314 & ~n32321;
  assign n32323 = n32259 & ~n32311;
  assign n32324 = ~n32259 & n32311;
  assign n32325 = ~n32323 & ~n32324;
  assign n32326 = pi276 & ~n32318;
  assign n32327 = pi141 & n32326;
  assign n32328 = pi274 & ~n32319;
  assign n32329 = pi143 & n32328;
  assign n32330 = ~n32327 & ~n32329;
  assign n32331 = ~n32325 & ~n32330;
  assign n32332 = ~n32322 & ~n32331;
  assign n32333 = n32246 & ~n32332;
  assign n32334 = ~n32246 & n32332;
  assign n32335 = ~n32333 & ~n32334;
  assign n32336 = n29568 & n29590;
  assign n32337 = ~n29558 & n29574;
  assign n32338 = n29558 & ~n29574;
  assign n32339 = ~n32337 & ~n32338;
  assign n32340 = n29255 & ~n32339;
  assign n32341 = ~n29558 & ~n29574;
  assign n32342 = n29558 & n29574;
  assign n32343 = ~n32341 & ~n32342;
  assign n32344 = ~n29255 & ~n32343;
  assign n32345 = ~n32340 & ~n32344;
  assign n32346 = ~n29568 & ~n29590;
  assign n32347 = ~n32345 & ~n32346;
  assign n32348 = ~n32336 & ~n32347;
  assign n32349 = pi272 & n32348;
  assign n32350 = pi145 & n32349;
  assign n32351 = pi145 & pi272;
  assign n32352 = ~n32348 & ~n32351;
  assign n32353 = ~n32350 & ~n32352;
  assign n32354 = ~n32335 & ~n32353;
  assign n32355 = ~n32246 & ~n32332;
  assign n32356 = n32246 & n32332;
  assign n32357 = ~n32355 & ~n32356;
  assign n32358 = n32348 & ~n32351;
  assign n32359 = pi272 & ~n32348;
  assign n32360 = pi145 & n32359;
  assign n32361 = ~n32358 & ~n32360;
  assign n32362 = ~n32357 & ~n32361;
  assign n32363 = ~n32354 & ~n32362;
  assign n32364 = pi152 & pi265;
  assign n32365 = n32363 & ~n32364;
  assign n32366 = pi265 & ~n32363;
  assign n32367 = pi152 & n32366;
  assign n32368 = ~n32365 & ~n32367;
  assign n32369 = ~n32233 & ~n32368;
  assign n32370 = ~n29620 & ~n32230;
  assign n32371 = ~n32231 & ~n32370;
  assign n32372 = ~n32363 & ~n32364;
  assign n32373 = pi265 & n32363;
  assign n32374 = pi152 & n32373;
  assign n32375 = ~n32372 & ~n32374;
  assign n32376 = ~n32371 & ~n32375;
  assign n32377 = ~n32369 & ~n32376;
  assign n32378 = ~n32219 & ~n32377;
  assign n32379 = n32219 & n32377;
  assign n32380 = ~n32378 & ~n32379;
  assign n32381 = n28556 & n28562;
  assign n32382 = ~n28556 & ~n28562;
  assign n32383 = n28552 & ~n32382;
  assign n32384 = ~n32381 & ~n32383;
  assign n32385 = n29698 & ~n32384;
  assign n32386 = ~n29698 & n32384;
  assign n32387 = ~n29697 & ~n32386;
  assign n32388 = ~n32385 & ~n32387;
  assign n32389 = n29255 & ~n29574;
  assign n32390 = ~n29255 & n29574;
  assign n32391 = n29558 & ~n32390;
  assign n32392 = ~n32389 & ~n32391;
  assign n32393 = n29257 & n29470;
  assign n32394 = ~n29257 & ~n29470;
  assign n32395 = ~n29454 & ~n32394;
  assign n32396 = ~n32393 & ~n32395;
  assign n32397 = n29313 & n32269;
  assign n32398 = ~n29313 & ~n32269;
  assign n32399 = ~n32397 & ~n32398;
  assign n32400 = pi285 & ~n32399;
  assign n32401 = pi131 & n32400;
  assign n32402 = ~n29313 & n32269;
  assign n32403 = n29313 & ~n32269;
  assign n32404 = ~n32402 & ~n32403;
  assign n32405 = ~n29266 & ~n32404;
  assign n32406 = ~n32401 & ~n32405;
  assign n32407 = n29348 & ~n32406;
  assign n32408 = ~n29348 & n32406;
  assign n32409 = ~n29317 & ~n32408;
  assign n32410 = ~n32407 & ~n32409;
  assign n32411 = pi287 & ~n32410;
  assign n32412 = pi130 & n32411;
  assign n32413 = pi130 & pi287;
  assign n32414 = n29317 & ~n29348;
  assign n32415 = ~n29317 & n29348;
  assign n32416 = n32406 & ~n32415;
  assign n32417 = ~n32414 & ~n32416;
  assign n32418 = ~n32413 & ~n32417;
  assign n32419 = ~n32412 & ~n32418;
  assign n32420 = pi282 & ~n29382;
  assign n32421 = pi134 & n32420;
  assign n32422 = ~n29359 & n29364;
  assign n32423 = ~n29365 & ~n32422;
  assign n32424 = ~n29259 & n29382;
  assign n32425 = ~n32423 & ~n32424;
  assign n32426 = ~n32421 & ~n32425;
  assign n32427 = n32419 & ~n32426;
  assign n32428 = n29359 & n29364;
  assign n32429 = ~n29370 & ~n29382;
  assign n32430 = ~n32428 & n32429;
  assign n32431 = ~n29259 & ~n32430;
  assign n32432 = ~n29370 & ~n32428;
  assign n32433 = n29382 & ~n32432;
  assign n32434 = ~n32431 & ~n32433;
  assign n32435 = ~n32419 & ~n32434;
  assign n32436 = ~n32427 & ~n32435;
  assign n32437 = n29258 & ~n29418;
  assign n32438 = ~n29258 & n29418;
  assign n32439 = n29402 & ~n32438;
  assign n32440 = ~n32437 & ~n32439;
  assign n32441 = n32436 & ~n32440;
  assign n32442 = ~n29258 & ~n32249;
  assign n32443 = ~n32248 & ~n32442;
  assign n32444 = ~n32436 & ~n32443;
  assign n32445 = ~n32441 & ~n32444;
  assign n32446 = n32396 & n32445;
  assign n32447 = ~n32396 & ~n32445;
  assign n32448 = ~n32446 & ~n32447;
  assign n32449 = pi273 & pi275;
  assign n32450 = n10889 & n32449;
  assign n32451 = pi144 & pi273;
  assign n32452 = pi142 & pi275;
  assign n32453 = ~n32451 & ~n32452;
  assign n32454 = ~n32450 & ~n32453;
  assign n32455 = ~n32448 & ~n32454;
  assign n32456 = n32396 & ~n32445;
  assign n32457 = ~n32396 & n32445;
  assign n32458 = ~n32456 & ~n32457;
  assign n32459 = pi275 & ~n32451;
  assign n32460 = pi142 & n32459;
  assign n32461 = pi273 & ~n32452;
  assign n32462 = pi144 & n32461;
  assign n32463 = ~n32460 & ~n32462;
  assign n32464 = ~n32458 & ~n32463;
  assign n32465 = ~n32455 & ~n32464;
  assign n32466 = n32392 & ~n32465;
  assign n32467 = ~n32392 & n32465;
  assign n32468 = ~n32466 & ~n32467;
  assign n32469 = n29594 & ~n29605;
  assign n32470 = ~n29594 & n29605;
  assign n32471 = ~n29596 & ~n32470;
  assign n32472 = ~n32469 & ~n32471;
  assign n32473 = pi266 & ~n32472;
  assign n32474 = pi151 & n32473;
  assign n32475 = pi151 & pi266;
  assign n32476 = n32472 & ~n32475;
  assign n32477 = ~n32474 & ~n32476;
  assign n32478 = ~n32468 & ~n32477;
  assign n32479 = ~n32392 & ~n32465;
  assign n32480 = n32392 & n32465;
  assign n32481 = ~n32479 & ~n32480;
  assign n32482 = ~n32472 & ~n32475;
  assign n32483 = pi266 & n32472;
  assign n32484 = pi151 & n32483;
  assign n32485 = ~n32482 & ~n32484;
  assign n32486 = ~n32481 & ~n32485;
  assign n32487 = ~n32478 & ~n32486;
  assign n32488 = ~n32388 & n32487;
  assign n32489 = n32388 & ~n32487;
  assign n32490 = ~n32488 & ~n32489;
  assign n32491 = pi153 & pi155;
  assign n32492 = pi262 & pi264;
  assign n32493 = n32491 & n32492;
  assign n32494 = pi155 & pi262;
  assign n32495 = pi153 & pi264;
  assign n32496 = ~n32494 & ~n32495;
  assign n32497 = ~n32493 & ~n32496;
  assign n32498 = ~n32490 & ~n32497;
  assign n32499 = ~n32388 & ~n32487;
  assign n32500 = n32388 & n32487;
  assign n32501 = ~n32499 & ~n32500;
  assign n32502 = pi264 & ~n32494;
  assign n32503 = pi153 & n32502;
  assign n32504 = pi262 & ~n32495;
  assign n32505 = pi155 & n32504;
  assign n32506 = ~n32503 & ~n32505;
  assign n32507 = ~n32501 & ~n32506;
  assign n32508 = ~n32498 & ~n32507;
  assign n32509 = pi263 & ~n32508;
  assign n32510 = pi154 & n32509;
  assign n32511 = pi154 & pi263;
  assign n32512 = n32508 & ~n32511;
  assign n32513 = ~n32510 & ~n32512;
  assign n32514 = ~n32380 & ~n32513;
  assign n32515 = n32219 & ~n32377;
  assign n32516 = ~n32219 & n32377;
  assign n32517 = ~n32515 & ~n32516;
  assign n32518 = ~n32508 & ~n32511;
  assign n32519 = pi263 & n32508;
  assign n32520 = pi154 & n32519;
  assign n32521 = ~n32518 & ~n32520;
  assign n32522 = ~n32517 & ~n32521;
  assign n32523 = ~n32514 & ~n32522;
  assign n32524 = ~n32173 & ~n32174;
  assign n32525 = ~n29645 & ~n29646;
  assign n32526 = n29645 & n29646;
  assign n32527 = ~n29651 & ~n32526;
  assign n32528 = ~n32525 & ~n32527;
  assign n32529 = n28259 & n28264;
  assign n32530 = ~n28259 & ~n28264;
  assign n32531 = n28255 & ~n32530;
  assign n32532 = ~n32529 & ~n32531;
  assign n32533 = ~n29438 & n32532;
  assign n32534 = n29438 & ~n32532;
  assign n32535 = ~n29449 & ~n32534;
  assign n32536 = ~n32533 & ~n32535;
  assign n32537 = pi277 & ~n32536;
  assign n32538 = pi140 & n32537;
  assign n32539 = pi140 & pi277;
  assign n32540 = ~n29437 & ~n32539;
  assign n32541 = ~n32533 & n32540;
  assign n32542 = ~n32532 & ~n32539;
  assign n32543 = n29438 & n32542;
  assign n32544 = ~n32541 & ~n32543;
  assign n32545 = ~n32538 & n32544;
  assign n32546 = pi136 & pi281;
  assign n32547 = pi132 & pi285;
  assign n32548 = pi129 & pi288;
  assign n32549 = pi289 & ~n32548;
  assign n32550 = pi128 & n32549;
  assign n32551 = pi128 & pi289;
  assign n32552 = pi288 & ~n32551;
  assign n32553 = pi129 & n32552;
  assign n32554 = ~n32550 & ~n32553;
  assign n32555 = ~n32547 & ~n32554;
  assign n32556 = pi288 & pi289;
  assign n32557 = n1175 & n32556;
  assign n32558 = ~n32548 & ~n32551;
  assign n32559 = ~n32557 & ~n32558;
  assign n32560 = pi285 & ~n32559;
  assign n32561 = pi132 & n32560;
  assign n32562 = ~n32555 & ~n32561;
  assign n32563 = pi283 & n32562;
  assign n32564 = pi134 & n32563;
  assign n32565 = pi134 & pi283;
  assign n32566 = ~n32562 & ~n32565;
  assign n32567 = ~n32564 & ~n32566;
  assign n32568 = ~n32546 & ~n32567;
  assign n32569 = pi283 & ~n32562;
  assign n32570 = pi134 & n32569;
  assign n32571 = n32562 & ~n32565;
  assign n32572 = ~n32570 & ~n32571;
  assign n32573 = pi281 & ~n32572;
  assign n32574 = pi136 & n32573;
  assign n32575 = ~n32568 & ~n32574;
  assign n32576 = ~n32545 & ~n32575;
  assign n32577 = n32545 & n32575;
  assign n32578 = ~n32576 & ~n32577;
  assign n32579 = n28319 & n28324;
  assign n32580 = ~n28319 & ~n28324;
  assign n32581 = n28315 & ~n32580;
  assign n32582 = ~n32579 & ~n32581;
  assign n32583 = n29490 & ~n32582;
  assign n32584 = ~n29490 & n32582;
  assign n32585 = ~n29489 & ~n32584;
  assign n32586 = ~n32583 & ~n32585;
  assign n32587 = pi279 & n32586;
  assign n32588 = pi138 & n32587;
  assign n32589 = pi138 & pi279;
  assign n32590 = ~n32586 & ~n32589;
  assign n32591 = ~n32588 & ~n32590;
  assign n32592 = ~n32578 & ~n32591;
  assign n32593 = n32545 & ~n32575;
  assign n32594 = ~n32545 & n32575;
  assign n32595 = ~n32593 & ~n32594;
  assign n32596 = n32586 & ~n32589;
  assign n32597 = pi279 & ~n32586;
  assign n32598 = pi138 & n32597;
  assign n32599 = ~n32596 & ~n32598;
  assign n32600 = ~n32595 & ~n32599;
  assign n32601 = ~n32592 & ~n32600;
  assign n32602 = ~n28379 & n28384;
  assign n32603 = n28379 & ~n28384;
  assign n32604 = ~n28375 & ~n32603;
  assign n32605 = ~n32602 & ~n32604;
  assign n32606 = n29542 & ~n32605;
  assign n32607 = ~n29542 & n32605;
  assign n32608 = ~n29553 & ~n32607;
  assign n32609 = ~n32606 & ~n32608;
  assign n32610 = ~n32601 & ~n32609;
  assign n32611 = ~n29541 & ~n32606;
  assign n32612 = ~n32607 & ~n32611;
  assign n32613 = n32601 & ~n32612;
  assign n32614 = ~n32610 & ~n32613;
  assign n32615 = n32528 & n32614;
  assign n32616 = ~n32528 & ~n32614;
  assign n32617 = ~n32615 & ~n32616;
  assign n32618 = pi268 & pi270;
  assign n32619 = n16970 & n32618;
  assign n32620 = pi149 & pi268;
  assign n32621 = pi147 & pi270;
  assign n32622 = ~n32620 & ~n32621;
  assign n32623 = ~n32619 & ~n32622;
  assign n32624 = ~n32617 & ~n32623;
  assign n32625 = n32528 & ~n32614;
  assign n32626 = ~n32528 & n32614;
  assign n32627 = ~n32625 & ~n32626;
  assign n32628 = pi270 & ~n32620;
  assign n32629 = pi147 & n32628;
  assign n32630 = pi268 & ~n32621;
  assign n32631 = pi149 & n32630;
  assign n32632 = ~n32629 & ~n32631;
  assign n32633 = ~n32627 & ~n32632;
  assign n32634 = ~n32624 & ~n32633;
  assign n32635 = ~n29672 & n29694;
  assign n32636 = ~n32634 & ~n32635;
  assign n32637 = n29253 & n32636;
  assign n32638 = n29672 & ~n29694;
  assign n32639 = n32634 & ~n32638;
  assign n32640 = ~n29253 & n32639;
  assign n32641 = ~n32637 & ~n32640;
  assign n32642 = ~n32524 & ~n32641;
  assign n32643 = ~n29694 & ~n32634;
  assign n32644 = n29672 & n32643;
  assign n32645 = n29694 & n32634;
  assign n32646 = ~n29672 & n32645;
  assign n32647 = ~n32644 & ~n32646;
  assign n32648 = ~n29662 & ~n29678;
  assign n32649 = n29662 & n29678;
  assign n32650 = ~n32648 & ~n32649;
  assign n32651 = n29253 & n32639;
  assign n32652 = ~n29253 & n32636;
  assign n32653 = ~n32651 & ~n32652;
  assign n32654 = ~n32650 & ~n32653;
  assign n32655 = n32647 & ~n32654;
  assign n32656 = ~n32642 & n32655;
  assign n32657 = ~n32523 & ~n32656;
  assign n32658 = n32523 & n32656;
  assign n32659 = ~n32657 & ~n32658;
  assign n32660 = n29749 & n29754;
  assign n32661 = ~n29760 & ~n29763;
  assign n32662 = ~n32660 & ~n32661;
  assign n32663 = pi261 & n32662;
  assign n32664 = pi156 & n32663;
  assign n32665 = pi156 & pi261;
  assign n32666 = ~n32662 & ~n32665;
  assign n32667 = ~n32664 & ~n32666;
  assign n32668 = ~n32659 & ~n32667;
  assign n32669 = n32523 & ~n32656;
  assign n32670 = ~n32523 & n32656;
  assign n32671 = ~n32669 & ~n32670;
  assign n32672 = n32662 & ~n32665;
  assign n32673 = pi261 & ~n32662;
  assign n32674 = pi156 & n32673;
  assign n32675 = ~n32672 & ~n32674;
  assign n32676 = ~n32671 & ~n32675;
  assign n32677 = ~n32668 & ~n32676;
  assign n32678 = n32208 & ~n32677;
  assign n32679 = ~n32208 & n32677;
  assign n32680 = ~n32678 & ~n32679;
  assign n32681 = pi159 & pi258;
  assign n32682 = pi259 & ~n32681;
  assign n32683 = pi158 & n32682;
  assign n32684 = pi158 & pi259;
  assign n32685 = pi258 & ~n32684;
  assign n32686 = pi159 & n32685;
  assign n32687 = ~n32683 & ~n32686;
  assign n32688 = ~n29766 & n29785;
  assign n32689 = n29766 & ~n29785;
  assign n32690 = n29794 & ~n32689;
  assign n32691 = ~n32688 & ~n32690;
  assign n32692 = n32687 & ~n32691;
  assign n32693 = ~n29794 & ~n32688;
  assign n32694 = ~n32689 & ~n32693;
  assign n32695 = ~n32687 & ~n32694;
  assign n32696 = ~n32692 & ~n32695;
  assign n32697 = ~n32680 & ~n32696;
  assign n32698 = n32208 & n32677;
  assign n32699 = ~n32208 & ~n32677;
  assign n32700 = ~n32698 & ~n32699;
  assign n32701 = ~n32687 & ~n32691;
  assign n32702 = n32687 & ~n32694;
  assign n32703 = ~n32701 & ~n32702;
  assign n32704 = ~n32700 & ~n32703;
  assign n32705 = ~n32697 & ~n32704;
  assign n32706 = n29780 & n32705;
  assign n32707 = ~n29766 & ~n29794;
  assign n32708 = n29766 & n29794;
  assign n32709 = ~n32707 & ~n32708;
  assign n32710 = ~n29788 & ~n32709;
  assign n32711 = ~n29766 & n29794;
  assign n32712 = n29766 & ~n29794;
  assign n32713 = ~n32711 & ~n32712;
  assign n32714 = pi258 & ~n29785;
  assign n32715 = pi158 & n32714;
  assign n32716 = pi259 & ~n29784;
  assign n32717 = pi157 & n32716;
  assign n32718 = ~n32715 & ~n32717;
  assign n32719 = ~n32713 & ~n32718;
  assign n32720 = ~n32710 & ~n32719;
  assign n32721 = ~n29780 & ~n32705;
  assign n32722 = n32720 & n32721;
  assign n32723 = ~n32706 & ~n32722;
  assign n32724 = ~n29801 & ~n32723;
  assign n32725 = n29780 & n32720;
  assign n32726 = ~n29780 & ~n32720;
  assign n32727 = ~n32725 & ~n32726;
  assign n32728 = n32705 & ~n32727;
  assign n32729 = ~n29780 & n32705;
  assign n32730 = n29780 & ~n32705;
  assign n32731 = ~n32720 & n32730;
  assign n32732 = ~n32729 & ~n32731;
  assign n32733 = n29801 & ~n32732;
  assign n32734 = ~n32728 & ~n32733;
  assign n32735 = ~n32724 & n32734;
  assign n32736 = pi322 & ~n32735;
  assign n32737 = n32065 & n32736;
  assign n32738 = ~n32065 & ~n32736;
  assign n32739 = ~n32737 & ~n32738;
  assign n32740 = ~n29217 & n29854;
  assign n32741 = n29217 & ~n29854;
  assign n32742 = ~n32740 & ~n32741;
  assign n32743 = ~n29838 & n29859;
  assign n32744 = n29838 & ~n29859;
  assign n32745 = ~n32743 & ~n32744;
  assign n32746 = ~n32742 & ~n32745;
  assign n32747 = n29217 & n29854;
  assign n32748 = ~n29217 & ~n29854;
  assign n32749 = ~n32747 & ~n32748;
  assign n32750 = ~n29838 & ~n29859;
  assign n32751 = n29838 & n29859;
  assign n32752 = ~n32750 & ~n32751;
  assign n32753 = ~n32749 & ~n32752;
  assign n32754 = ~n32746 & ~n32753;
  assign n32755 = pi323 & n29822;
  assign n32756 = n26706 & ~n32755;
  assign n32757 = pi326 & n32756;
  assign n32758 = ~n32754 & n32757;
  assign n32759 = n29858 & ~n32754;
  assign n32760 = n29822 & ~n32759;
  assign n32761 = pi323 & n32760;
  assign n32762 = ~n32758 & ~n32761;
  assign n32763 = pi326 & n26175;
  assign n32764 = ~n32762 & ~n32763;
  assign n32765 = n32762 & n32763;
  assign n32766 = ~n32764 & ~n32765;
  assign n32767 = n28628 & ~n32766;
  assign n32768 = pi324 & n32767;
  assign n32769 = pi324 & n28628;
  assign n32770 = n32762 & ~n32763;
  assign n32771 = ~n32762 & n32763;
  assign n32772 = ~n32770 & ~n32771;
  assign n32773 = ~n32769 & ~n32772;
  assign n32774 = ~n32768 & ~n32773;
  assign n32775 = ~n32739 & ~n32774;
  assign n32776 = n32065 & ~n32736;
  assign n32777 = ~n32065 & n32736;
  assign n32778 = ~n32776 & ~n32777;
  assign n32779 = n28628 & ~n32772;
  assign n32780 = pi324 & n32779;
  assign n32781 = ~n32766 & ~n32769;
  assign n32782 = ~n32780 & ~n32781;
  assign n32783 = ~n32778 & ~n32782;
  assign n32784 = ~n32775 & ~n32783;
  assign n32785 = ~n32059 & ~n32784;
  assign n32786 = n32059 & n32784;
  assign n32787 = ~n32785 & ~n32786;
  assign n32788 = n19970 & n32754;
  assign n32789 = pi329 & n32788;
  assign n32790 = pi329 & n19970;
  assign n32791 = ~n29237 & ~n32790;
  assign n32792 = ~n32754 & n32791;
  assign n32793 = ~n32789 & ~n32792;
  assign n32794 = ~n29858 & ~n32793;
  assign n32795 = ~n29237 & ~n32759;
  assign n32796 = n19970 & ~n32795;
  assign n32797 = pi329 & n32796;
  assign n32798 = n26706 & ~n32790;
  assign n32799 = pi326 & n32798;
  assign n32800 = ~n29237 & n32799;
  assign n32801 = n32754 & n32800;
  assign n32802 = ~n32797 & ~n32801;
  assign n32803 = ~n32794 & n32802;
  assign n32804 = pi328 & n21479;
  assign n32805 = ~n32803 & ~n32804;
  assign n32806 = n21479 & n32803;
  assign n32807 = pi328 & n32806;
  assign n32808 = ~n32805 & ~n32807;
  assign n32809 = ~n32787 & ~n32808;
  assign n32810 = n32059 & ~n32784;
  assign n32811 = ~n32059 & n32784;
  assign n32812 = ~n32810 & ~n32811;
  assign n32813 = n32803 & ~n32804;
  assign n32814 = n21479 & ~n32803;
  assign n32815 = pi328 & n32814;
  assign n32816 = ~n32813 & ~n32815;
  assign n32817 = ~n32812 & ~n32816;
  assign n32818 = ~n32809 & ~n32817;
  assign n32819 = ~n32027 & ~n32818;
  assign n32820 = n32027 & n32818;
  assign n32821 = ~n32819 & ~n32820;
  assign n32822 = ~n31997 & ~n32821;
  assign n32823 = n32027 & ~n32818;
  assign n32824 = ~n32027 & n32818;
  assign n32825 = ~n32823 & ~n32824;
  assign n32826 = n31992 & ~n31993;
  assign n32827 = n19539 & ~n31992;
  assign n32828 = pi331 & n32827;
  assign n32829 = ~n32826 & ~n32828;
  assign n32830 = ~n32825 & ~n32829;
  assign n32831 = ~n32822 & ~n32830;
  assign n32832 = n31982 & n32831;
  assign n32833 = ~n31982 & ~n32831;
  assign n32834 = ~n32832 & ~n32833;
  assign n32835 = n29145 & ~n31714;
  assign n32836 = ~n29145 & ~n31704;
  assign n32837 = ~n32835 & ~n32836;
  assign n32838 = n27911 & ~n29134;
  assign n32839 = ~n27911 & ~n29124;
  assign n32840 = ~n32838 & ~n32839;
  assign n32841 = ~n29988 & ~n32840;
  assign n32842 = ~n29991 & ~n32841;
  assign n32843 = ~n29987 & n32842;
  assign n32844 = ~n32837 & ~n32843;
  assign n32845 = n29987 & ~n32842;
  assign n32846 = ~n32844 & ~n32845;
  assign n32847 = pi336 & n11384;
  assign n32848 = ~n32846 & ~n32847;
  assign n32849 = n32846 & n32847;
  assign n32850 = ~n32848 & ~n32849;
  assign n32851 = n11711 & ~n32850;
  assign n32852 = pi335 & n32851;
  assign n32853 = pi335 & n11711;
  assign n32854 = n32846 & ~n32847;
  assign n32855 = ~n32846 & n32847;
  assign n32856 = ~n32854 & ~n32855;
  assign n32857 = ~n32853 & ~n32856;
  assign n32858 = ~n32852 & ~n32857;
  assign n32859 = ~n32834 & ~n32858;
  assign n32860 = n31982 & ~n32831;
  assign n32861 = ~n31982 & n32831;
  assign n32862 = ~n32860 & ~n32861;
  assign n32863 = n11711 & ~n32856;
  assign n32864 = pi335 & n32863;
  assign n32865 = ~n32850 & ~n32853;
  assign n32866 = ~n32864 & ~n32865;
  assign n32867 = ~n32862 & ~n32866;
  assign n32868 = ~n32859 & ~n32867;
  assign n32869 = ~n31971 & ~n32868;
  assign n32870 = n31971 & n32868;
  assign n32871 = ~n32869 & ~n32870;
  assign n32872 = ~n31952 & ~n32871;
  assign n32873 = n31971 & ~n32868;
  assign n32874 = ~n31971 & n32868;
  assign n32875 = ~n32873 & ~n32874;
  assign n32876 = ~n31947 & ~n31948;
  assign n32877 = n9205 & n31947;
  assign n32878 = pi339 & n32877;
  assign n32879 = ~n32876 & ~n32878;
  assign n32880 = ~n32875 & ~n32879;
  assign n32881 = ~n32872 & ~n32880;
  assign n32882 = n31941 & ~n32881;
  assign n32883 = ~n31941 & n32881;
  assign n32884 = ~n32882 & ~n32883;
  assign n32885 = n2887 & ~n30139;
  assign n32886 = ~n30140 & ~n32885;
  assign n32887 = n4596 & ~n32886;
  assign n32888 = pi344 & n32887;
  assign n32889 = pi343 & n5714;
  assign n32890 = ~n4596 & ~n32885;
  assign n32891 = pi344 & ~n32890;
  assign n32892 = ~n30140 & ~n32891;
  assign n32893 = n30127 & ~n32892;
  assign n32894 = ~n32889 & ~n32893;
  assign n32895 = ~n32888 & n32894;
  assign n32896 = ~n32888 & ~n32893;
  assign n32897 = n32889 & ~n32896;
  assign n32898 = ~n32895 & ~n32897;
  assign n32899 = ~n32884 & ~n32898;
  assign n32900 = n31941 & n32881;
  assign n32901 = ~n31941 & ~n32881;
  assign n32902 = ~n32900 & ~n32901;
  assign n32903 = n32889 & ~n32893;
  assign n32904 = ~n32888 & n32903;
  assign n32905 = ~n32889 & ~n32896;
  assign n32906 = ~n32904 & ~n32905;
  assign n32907 = ~n32902 & ~n32906;
  assign n32908 = ~n32899 & ~n32907;
  assign n32909 = pi346 & n2887;
  assign n32910 = ~n32908 & ~n32909;
  assign n32911 = n2887 & n32908;
  assign n32912 = pi346 & n32911;
  assign n32913 = ~n32910 & ~n32912;
  assign n32914 = ~n31927 & ~n32913;
  assign n32915 = ~n29089 & ~n31643;
  assign n32916 = ~n31642 & ~n32915;
  assign n32917 = n32908 & ~n32909;
  assign n32918 = n2887 & ~n32908;
  assign n32919 = pi346 & n32918;
  assign n32920 = ~n32917 & ~n32919;
  assign n32921 = ~n32916 & ~n32920;
  assign n32922 = ~n32914 & ~n32921;
  assign n32923 = n31925 & ~n32922;
  assign n32924 = ~n31925 & n32922;
  assign n32925 = ~n32923 & ~n32924;
  assign n32926 = ~n31918 & ~n32925;
  assign n32927 = ~n31925 & ~n32922;
  assign n32928 = n31925 & n32922;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = ~n31651 & ~n31916;
  assign n32931 = n31651 & ~n31912;
  assign n32932 = ~n32930 & ~n32931;
  assign n32933 = ~n32929 & ~n32932;
  assign n32934 = ~n32926 & ~n32933;
  assign n32935 = n31631 & ~n32934;
  assign n32936 = ~n31631 & n32934;
  assign n32937 = ~n32935 & ~n32936;
  assign n32938 = pi350 & n1442;
  assign n32939 = pi289 & n32938;
  assign n32940 = ~pi289 & ~n32938;
  assign n32941 = ~n32939 & ~n32940;
  assign n32942 = ~n30232 & ~n30238;
  assign n32943 = ~n30237 & ~n32942;
  assign n32944 = n1729 & ~n32943;
  assign n32945 = pi349 & n32944;
  assign n32946 = pi349 & n1729;
  assign n32947 = ~n30251 & ~n32946;
  assign n32948 = ~n30237 & n32947;
  assign n32949 = n30236 & ~n32946;
  assign n32950 = n30235 & n32949;
  assign n32951 = ~n32948 & ~n32950;
  assign n32952 = ~n32945 & n32951;
  assign n32953 = n32941 & n32952;
  assign n32954 = ~n32941 & ~n32952;
  assign n32955 = ~n32953 & ~n32954;
  assign n32956 = ~n30239 & ~n30251;
  assign n32957 = ~n30232 & ~n30245;
  assign n32958 = ~n32956 & ~n32957;
  assign n32959 = n1156 & ~n32958;
  assign n32960 = pi352 & n32959;
  assign n32961 = pi294 & n1533;
  assign n32962 = ~n30953 & ~n30967;
  assign n32963 = ~n30954 & ~n32962;
  assign n32964 = pi293 & n1553;
  assign n32965 = n32963 & ~n32964;
  assign n32966 = n1553 & ~n32963;
  assign n32967 = pi293 & n32966;
  assign n32968 = ~n32965 & ~n32967;
  assign n32969 = ~n32961 & ~n32968;
  assign n32970 = ~n32963 & ~n32964;
  assign n32971 = n1553 & n32963;
  assign n32972 = pi293 & n32971;
  assign n32973 = ~n32970 & ~n32972;
  assign n32974 = n1533 & ~n32973;
  assign n32975 = pi294 & n32974;
  assign n32976 = ~n32969 & ~n32975;
  assign n32977 = n32960 & ~n32976;
  assign n32978 = ~n32960 & n32976;
  assign n32979 = ~n32977 & ~n32978;
  assign n32980 = ~n32955 & ~n32979;
  assign n32981 = ~n32941 & n32952;
  assign n32982 = n32941 & ~n32952;
  assign n32983 = ~n32981 & ~n32982;
  assign n32984 = ~n32960 & ~n32976;
  assign n32985 = n32960 & n32976;
  assign n32986 = ~n32984 & ~n32985;
  assign n32987 = ~n32983 & ~n32986;
  assign n32988 = ~n32980 & ~n32987;
  assign n32989 = ~n32937 & ~n32988;
  assign n32990 = n31631 & n32934;
  assign n32991 = ~n31631 & ~n32934;
  assign n32992 = ~n32990 & ~n32991;
  assign n32993 = ~n32979 & ~n32983;
  assign n32994 = ~n32955 & ~n32986;
  assign n32995 = ~n32993 & ~n32994;
  assign n32996 = ~n32992 & ~n32995;
  assign n32997 = ~n32989 & ~n32996;
  assign n32998 = ~n30261 & n30973;
  assign n32999 = n30261 & ~n30973;
  assign n33000 = ~n31606 & ~n31607;
  assign n33001 = pi288 & ~n33000;
  assign n33002 = n30257 & ~n30979;
  assign n33003 = ~n30257 & n30979;
  assign n33004 = ~n33002 & ~n33003;
  assign n33005 = ~pi288 & ~n33004;
  assign n33006 = ~n33001 & ~n33005;
  assign n33007 = ~n32999 & ~n33006;
  assign n33008 = ~n32998 & ~n33007;
  assign n33009 = ~n32997 & n33008;
  assign n33010 = n32997 & ~n33008;
  assign n33011 = ~n33009 & ~n33010;
  assign n33012 = ~n31617 & ~n33011;
  assign n33013 = ~n32997 & ~n33008;
  assign n33014 = n32997 & n33008;
  assign n33015 = ~n33013 & ~n33014;
  assign n33016 = n31617 & ~n33015;
  assign n33017 = ~n33012 & ~n33016;
  assign n33018 = n31048 & ~n33017;
  assign n33019 = ~n31048 & n33017;
  assign n33020 = ~n33018 & ~n33019;
  assign n33021 = ~n831 & n33020;
  assign n33022 = n31006 & ~n33021;
  assign n33023 = ~n31004 & ~n33022;
  assign po224 = ~pi160 & ~n33023;
  assign n33025 = pi063 & ~pi161;
  assign n33026 = pi319 & ~n1692;
  assign n33027 = ~pi319 & n1692;
  assign n33028 = pi321 & n1156;
  assign n33029 = n1699 & ~n33028;
  assign n33030 = pi320 & ~n33029;
  assign n33031 = pi321 & n1700;
  assign n33032 = ~n33030 & ~n33031;
  assign n33033 = ~n33027 & ~n33032;
  assign n33034 = ~n33026 & ~n33033;
  assign n33035 = ~n1679 & ~n33034;
  assign n33036 = n1679 & n33034;
  assign n33037 = pi318 & ~n33036;
  assign n33038 = ~n33035 & ~n33037;
  assign n33039 = ~n2070 & ~n33038;
  assign n33040 = n2070 & n33038;
  assign n33041 = pi317 & ~n33040;
  assign n33042 = ~n33039 & ~n33041;
  assign n33043 = ~n2432 & ~n33042;
  assign n33044 = n2432 & n33042;
  assign n33045 = pi316 & ~n33044;
  assign n33046 = ~n33043 & ~n33045;
  assign n33047 = ~n2852 & ~n33046;
  assign n33048 = n2852 & n33046;
  assign n33049 = pi315 & ~n33048;
  assign n33050 = ~n33047 & ~n33049;
  assign n33051 = ~n3331 & ~n33050;
  assign n33052 = n3331 & n33050;
  assign n33053 = pi314 & ~n33052;
  assign n33054 = ~n33051 & ~n33053;
  assign n33055 = ~n3319 & ~n33054;
  assign n33056 = n3319 & n33054;
  assign n33057 = pi313 & ~n33056;
  assign n33058 = ~n33055 & ~n33057;
  assign n33059 = ~n3909 & ~n33058;
  assign n33060 = n3909 & n33058;
  assign n33061 = pi312 & ~n33060;
  assign n33062 = ~n33059 & ~n33061;
  assign n33063 = ~n4558 & ~n33062;
  assign n33064 = n4558 & n33062;
  assign n33065 = pi311 & ~n33064;
  assign n33066 = ~n33063 & ~n33065;
  assign n33067 = ~n5723 & ~n33066;
  assign n33068 = n5723 & n33066;
  assign n33069 = pi310 & ~n33068;
  assign n33070 = ~n33067 & ~n33069;
  assign n33071 = ~n6523 & ~n33070;
  assign n33072 = n6523 & n33070;
  assign n33073 = pi309 & ~n33072;
  assign n33074 = ~n33071 & ~n33073;
  assign n33075 = ~n7364 & ~n33074;
  assign n33076 = n7364 & n33074;
  assign n33077 = pi308 & ~n33076;
  assign n33078 = ~n33075 & ~n33077;
  assign n33079 = ~n7601 & ~n33078;
  assign n33080 = n7601 & n33078;
  assign n33081 = pi307 & ~n33080;
  assign n33082 = ~n33079 & ~n33081;
  assign n33083 = ~n8513 & ~n33082;
  assign n33084 = n8513 & n33082;
  assign n33085 = pi306 & ~n33084;
  assign n33086 = ~n33083 & ~n33085;
  assign n33087 = ~n9167 & ~n33086;
  assign n33088 = n9167 & n33086;
  assign n33089 = pi305 & ~n33088;
  assign n33090 = ~n33087 & ~n33089;
  assign n33091 = ~n11375 & ~n33090;
  assign n33092 = n11375 & n33090;
  assign n33093 = pi304 & ~n33092;
  assign n33094 = ~n33091 & ~n33093;
  assign n33095 = ~n12895 & ~n33094;
  assign n33096 = n12895 & n33094;
  assign n33097 = pi303 & ~n33096;
  assign n33098 = ~n33095 & ~n33097;
  assign n33099 = ~n13729 & ~n33098;
  assign n33100 = n13729 & n33098;
  assign n33101 = pi302 & ~n33100;
  assign n33102 = ~n33099 & ~n33101;
  assign n33103 = ~n15166 & ~n33102;
  assign n33104 = n15166 & n33102;
  assign n33105 = pi301 & ~n33104;
  assign n33106 = ~n33103 & ~n33105;
  assign n33107 = ~n15616 & ~n33106;
  assign n33108 = n15616 & n33106;
  assign n33109 = pi300 & ~n33108;
  assign n33110 = ~n33107 & ~n33109;
  assign n33111 = ~n16527 & ~n33110;
  assign n33112 = n16527 & n33110;
  assign n33113 = pi299 & ~n33112;
  assign n33114 = ~n33111 & ~n33113;
  assign n33115 = ~n19548 & ~n33114;
  assign n33116 = n19548 & n33114;
  assign n33117 = pi298 & ~n33116;
  assign n33118 = ~n33115 & ~n33117;
  assign n33119 = ~n21446 & ~n33118;
  assign n33120 = n21446 & n33118;
  assign n33121 = pi297 & ~n33120;
  assign n33122 = ~n33119 & ~n33121;
  assign n33123 = ~n22557 & ~n33122;
  assign n33124 = n22557 & n33122;
  assign n33125 = pi296 & ~n33124;
  assign n33126 = ~n33123 & ~n33125;
  assign n33127 = ~n22545 & ~n33126;
  assign n33128 = n22545 & n33126;
  assign n33129 = pi295 & ~n33128;
  assign n33130 = ~n33127 & ~n33129;
  assign n33131 = ~n24906 & ~n33130;
  assign n33132 = n24906 & n33130;
  assign n33133 = pi294 & ~n33132;
  assign n33134 = ~n33131 & ~n33133;
  assign n33135 = ~n26683 & ~n33134;
  assign n33136 = n26683 & n33134;
  assign n33137 = pi293 & ~n33136;
  assign n33138 = ~n33135 & ~n33137;
  assign n33139 = ~n29801 & ~n33138;
  assign n33140 = n29801 & n33138;
  assign n33141 = pi292 & ~n33140;
  assign n33142 = ~n33139 & ~n33141;
  assign n33143 = ~n32720 & ~n33142;
  assign n33144 = n32720 & n33142;
  assign n33145 = pi291 & ~n33144;
  assign n33146 = ~n33143 & ~n33145;
  assign n33147 = n32705 & ~n33146;
  assign n33148 = ~pi291 & ~n33143;
  assign n33149 = ~n33144 & ~n33148;
  assign n33150 = ~n32705 & ~n33149;
  assign n33151 = ~n33147 & ~n33150;
  assign n33152 = ~n831 & n33151;
  assign n33153 = ~pi290 & n33152;
  assign n33154 = pi290 & ~n33152;
  assign n33155 = ~n33153 & ~n33154;
  assign n33156 = pi161 & ~n33155;
  assign n33157 = ~n33025 & ~n33156;
  assign po225 = ~pi160 & ~n33157;
  assign n33159 = n32720 & ~n33142;
  assign n33160 = ~n32720 & n33142;
  assign n33161 = ~n33159 & ~n33160;
  assign n33162 = ~n831 & ~n33161;
  assign n33163 = ~pi291 & n33162;
  assign n33164 = ~n33143 & ~n33144;
  assign n33165 = ~n831 & n33164;
  assign n33166 = pi291 & ~n33165;
  assign n33167 = ~n33163 & ~n33166;
  assign n33168 = pi161 & ~n33167;
  assign n33169 = pi062 & ~pi161;
  assign n33170 = ~n33168 & ~n33169;
  assign po226 = ~pi160 & ~n33170;
  assign n33172 = n29801 & ~n33138;
  assign n33173 = ~n29801 & n33138;
  assign n33174 = ~n33172 & ~n33173;
  assign n33175 = ~n831 & ~n33174;
  assign n33176 = ~pi292 & n33175;
  assign n33177 = ~n33139 & ~n33140;
  assign n33178 = ~n831 & n33177;
  assign n33179 = pi292 & ~n33178;
  assign n33180 = ~n33176 & ~n33179;
  assign n33181 = pi161 & ~n33180;
  assign n33182 = pi061 & ~pi161;
  assign n33183 = ~n33181 & ~n33182;
  assign po227 = ~pi160 & ~n33183;
  assign n33185 = ~pi060 & ~pi161;
  assign n33186 = ~n33135 & ~n33136;
  assign n33187 = ~n831 & n33186;
  assign n33188 = ~pi293 & ~n33187;
  assign n33189 = n26683 & ~n33134;
  assign n33190 = ~n26683 & n33134;
  assign n33191 = ~n33189 & ~n33190;
  assign n33192 = ~n831 & ~n33191;
  assign n33193 = pi293 & n33192;
  assign n33194 = ~n33188 & ~n33193;
  assign n33195 = pi161 & ~n33194;
  assign n33196 = ~n33185 & ~n33195;
  assign po228 = ~pi160 & n33196;
  assign n33198 = ~pi059 & ~pi161;
  assign n33199 = ~n33131 & ~n33132;
  assign n33200 = ~n831 & n33199;
  assign n33201 = ~pi294 & ~n33200;
  assign n33202 = n24906 & ~n33130;
  assign n33203 = ~n24906 & n33130;
  assign n33204 = ~n33202 & ~n33203;
  assign n33205 = ~n831 & ~n33204;
  assign n33206 = pi294 & n33205;
  assign n33207 = ~n33201 & ~n33206;
  assign n33208 = pi161 & ~n33207;
  assign n33209 = ~n33198 & ~n33208;
  assign po229 = ~pi160 & n33209;
  assign n33211 = n22545 & ~n33126;
  assign n33212 = ~n22545 & n33126;
  assign n33213 = ~n33211 & ~n33212;
  assign n33214 = ~n831 & ~n33213;
  assign n33215 = ~pi295 & n33214;
  assign n33216 = ~n33127 & ~n33128;
  assign n33217 = ~n831 & n33216;
  assign n33218 = pi295 & ~n33217;
  assign n33219 = ~n33215 & ~n33218;
  assign n33220 = pi161 & ~n33219;
  assign n33221 = pi058 & ~pi161;
  assign n33222 = ~n33220 & ~n33221;
  assign po230 = ~pi160 & ~n33222;
  assign n33224 = n22557 & ~n33122;
  assign n33225 = ~n22557 & n33122;
  assign n33226 = ~n33224 & ~n33225;
  assign n33227 = ~n831 & ~n33226;
  assign n33228 = ~pi296 & n33227;
  assign n33229 = ~n33123 & ~n33124;
  assign n33230 = ~n831 & n33229;
  assign n33231 = pi296 & ~n33230;
  assign n33232 = ~n33228 & ~n33231;
  assign n33233 = pi161 & ~n33232;
  assign n33234 = pi057 & ~pi161;
  assign n33235 = ~n33233 & ~n33234;
  assign po231 = ~pi160 & ~n33235;
  assign n33237 = n21446 & ~n33118;
  assign n33238 = ~n21446 & n33118;
  assign n33239 = ~n33237 & ~n33238;
  assign n33240 = ~n831 & ~n33239;
  assign n33241 = ~pi297 & n33240;
  assign n33242 = ~n33119 & ~n33120;
  assign n33243 = ~n831 & n33242;
  assign n33244 = pi297 & ~n33243;
  assign n33245 = ~n33241 & ~n33244;
  assign n33246 = pi161 & ~n33245;
  assign n33247 = pi056 & ~pi161;
  assign n33248 = ~n33246 & ~n33247;
  assign po232 = ~pi160 & ~n33248;
  assign n33250 = n19548 & ~n33114;
  assign n33251 = ~n19548 & n33114;
  assign n33252 = ~n33250 & ~n33251;
  assign n33253 = ~n831 & ~n33252;
  assign n33254 = ~pi298 & n33253;
  assign n33255 = ~n33115 & ~n33116;
  assign n33256 = ~n831 & n33255;
  assign n33257 = pi298 & ~n33256;
  assign n33258 = ~n33254 & ~n33257;
  assign n33259 = pi161 & ~n33258;
  assign n33260 = pi055 & ~pi161;
  assign n33261 = ~n33259 & ~n33260;
  assign po233 = ~pi160 & ~n33261;
  assign n33263 = n16527 & ~n33110;
  assign n33264 = ~n16527 & n33110;
  assign n33265 = ~n33263 & ~n33264;
  assign n33266 = ~n831 & ~n33265;
  assign n33267 = ~pi299 & n33266;
  assign n33268 = ~n33111 & ~n33112;
  assign n33269 = ~n831 & n33268;
  assign n33270 = pi299 & ~n33269;
  assign n33271 = ~n33267 & ~n33270;
  assign n33272 = pi161 & ~n33271;
  assign n33273 = pi054 & ~pi161;
  assign n33274 = ~n33272 & ~n33273;
  assign po234 = ~pi160 & ~n33274;
  assign n33276 = n15616 & ~n33106;
  assign n33277 = ~n15616 & n33106;
  assign n33278 = ~n33276 & ~n33277;
  assign n33279 = ~n831 & ~n33278;
  assign n33280 = ~pi300 & n33279;
  assign n33281 = ~n33107 & ~n33108;
  assign n33282 = ~n831 & n33281;
  assign n33283 = pi300 & ~n33282;
  assign n33284 = ~n33280 & ~n33283;
  assign n33285 = pi161 & ~n33284;
  assign n33286 = pi053 & ~pi161;
  assign n33287 = ~n33285 & ~n33286;
  assign po235 = ~pi160 & ~n33287;
  assign n33289 = n15166 & ~n33102;
  assign n33290 = ~n15166 & n33102;
  assign n33291 = ~n33289 & ~n33290;
  assign n33292 = ~n831 & ~n33291;
  assign n33293 = ~pi301 & n33292;
  assign n33294 = ~n33103 & ~n33104;
  assign n33295 = ~n831 & n33294;
  assign n33296 = pi301 & ~n33295;
  assign n33297 = ~n33293 & ~n33296;
  assign n33298 = pi161 & ~n33297;
  assign n33299 = pi052 & ~pi161;
  assign n33300 = ~n33298 & ~n33299;
  assign po236 = ~pi160 & ~n33300;
  assign n33302 = n13729 & ~n33098;
  assign n33303 = ~n13729 & n33098;
  assign n33304 = ~n33302 & ~n33303;
  assign n33305 = ~n831 & ~n33304;
  assign n33306 = ~pi302 & n33305;
  assign n33307 = ~n33099 & ~n33100;
  assign n33308 = ~n831 & n33307;
  assign n33309 = pi302 & ~n33308;
  assign n33310 = ~n33306 & ~n33309;
  assign n33311 = pi161 & ~n33310;
  assign n33312 = pi051 & ~pi161;
  assign n33313 = ~n33311 & ~n33312;
  assign po237 = ~pi160 & ~n33313;
  assign n33315 = n12895 & ~n33094;
  assign n33316 = ~n12895 & n33094;
  assign n33317 = ~n33315 & ~n33316;
  assign n33318 = ~n831 & ~n33317;
  assign n33319 = ~pi303 & n33318;
  assign n33320 = ~n33095 & ~n33096;
  assign n33321 = ~n831 & n33320;
  assign n33322 = pi303 & ~n33321;
  assign n33323 = ~n33319 & ~n33322;
  assign n33324 = pi161 & ~n33323;
  assign n33325 = pi050 & ~pi161;
  assign n33326 = ~n33324 & ~n33325;
  assign po238 = ~pi160 & ~n33326;
  assign n33328 = n11375 & ~n33090;
  assign n33329 = ~n11375 & n33090;
  assign n33330 = ~n33328 & ~n33329;
  assign n33331 = ~n831 & ~n33330;
  assign n33332 = ~pi304 & n33331;
  assign n33333 = ~n33091 & ~n33092;
  assign n33334 = ~n831 & n33333;
  assign n33335 = pi304 & ~n33334;
  assign n33336 = ~n33332 & ~n33335;
  assign n33337 = pi161 & ~n33336;
  assign n33338 = pi049 & ~pi161;
  assign n33339 = ~n33337 & ~n33338;
  assign po239 = ~pi160 & ~n33339;
  assign n33341 = n9167 & ~n33086;
  assign n33342 = ~n9167 & n33086;
  assign n33343 = ~n33341 & ~n33342;
  assign n33344 = ~n831 & ~n33343;
  assign n33345 = ~pi305 & n33344;
  assign n33346 = ~n33087 & ~n33088;
  assign n33347 = ~n831 & n33346;
  assign n33348 = pi305 & ~n33347;
  assign n33349 = ~n33345 & ~n33348;
  assign n33350 = pi161 & ~n33349;
  assign n33351 = pi048 & ~pi161;
  assign n33352 = ~n33350 & ~n33351;
  assign po240 = ~pi160 & ~n33352;
  assign n33354 = n8513 & ~n33082;
  assign n33355 = ~n8513 & n33082;
  assign n33356 = ~n33354 & ~n33355;
  assign n33357 = ~n831 & ~n33356;
  assign n33358 = ~pi306 & n33357;
  assign n33359 = ~n33083 & ~n33084;
  assign n33360 = ~n831 & n33359;
  assign n33361 = pi306 & ~n33360;
  assign n33362 = ~n33358 & ~n33361;
  assign n33363 = pi161 & ~n33362;
  assign n33364 = pi047 & ~pi161;
  assign n33365 = ~n33363 & ~n33364;
  assign po241 = ~pi160 & ~n33365;
  assign n33367 = n7601 & ~n33078;
  assign n33368 = ~n7601 & n33078;
  assign n33369 = ~n33367 & ~n33368;
  assign n33370 = ~n831 & ~n33369;
  assign n33371 = ~pi307 & n33370;
  assign n33372 = ~n33079 & ~n33080;
  assign n33373 = ~n831 & n33372;
  assign n33374 = pi307 & ~n33373;
  assign n33375 = ~n33371 & ~n33374;
  assign n33376 = pi161 & ~n33375;
  assign n33377 = pi046 & ~pi161;
  assign n33378 = ~n33376 & ~n33377;
  assign po242 = ~pi160 & ~n33378;
  assign n33380 = n7364 & ~n33074;
  assign n33381 = ~n7364 & n33074;
  assign n33382 = ~n33380 & ~n33381;
  assign n33383 = ~n831 & ~n33382;
  assign n33384 = ~pi308 & n33383;
  assign n33385 = ~n33075 & ~n33076;
  assign n33386 = ~n831 & n33385;
  assign n33387 = pi308 & ~n33386;
  assign n33388 = ~n33384 & ~n33387;
  assign n33389 = pi161 & ~n33388;
  assign n33390 = pi045 & ~pi161;
  assign n33391 = ~n33389 & ~n33390;
  assign po243 = ~pi160 & ~n33391;
  assign n33393 = n6523 & ~n33070;
  assign n33394 = ~n6523 & n33070;
  assign n33395 = ~n33393 & ~n33394;
  assign n33396 = ~n831 & ~n33395;
  assign n33397 = ~pi309 & n33396;
  assign n33398 = ~n33071 & ~n33072;
  assign n33399 = ~n831 & n33398;
  assign n33400 = pi309 & ~n33399;
  assign n33401 = ~n33397 & ~n33400;
  assign n33402 = pi161 & ~n33401;
  assign n33403 = pi044 & ~pi161;
  assign n33404 = ~n33402 & ~n33403;
  assign po244 = ~pi160 & ~n33404;
  assign n33406 = n5723 & ~n33066;
  assign n33407 = ~n5723 & n33066;
  assign n33408 = ~n33406 & ~n33407;
  assign n33409 = ~n831 & ~n33408;
  assign n33410 = ~pi310 & n33409;
  assign n33411 = ~n33067 & ~n33068;
  assign n33412 = ~n831 & n33411;
  assign n33413 = pi310 & ~n33412;
  assign n33414 = ~n33410 & ~n33413;
  assign n33415 = pi161 & ~n33414;
  assign n33416 = pi043 & ~pi161;
  assign n33417 = ~n33415 & ~n33416;
  assign po245 = ~pi160 & ~n33417;
  assign n33419 = n4558 & ~n33062;
  assign n33420 = ~n4558 & n33062;
  assign n33421 = ~n33419 & ~n33420;
  assign n33422 = ~n831 & ~n33421;
  assign n33423 = ~pi311 & n33422;
  assign n33424 = ~n33063 & ~n33064;
  assign n33425 = ~n831 & n33424;
  assign n33426 = pi311 & ~n33425;
  assign n33427 = ~n33423 & ~n33426;
  assign n33428 = pi161 & ~n33427;
  assign n33429 = pi042 & ~pi161;
  assign n33430 = ~n33428 & ~n33429;
  assign po246 = ~pi160 & ~n33430;
  assign n33432 = n3909 & ~n33058;
  assign n33433 = ~n3909 & n33058;
  assign n33434 = ~n33432 & ~n33433;
  assign n33435 = ~n831 & ~n33434;
  assign n33436 = ~pi312 & n33435;
  assign n33437 = ~n33059 & ~n33060;
  assign n33438 = ~n831 & n33437;
  assign n33439 = pi312 & ~n33438;
  assign n33440 = ~n33436 & ~n33439;
  assign n33441 = pi161 & ~n33440;
  assign n33442 = pi041 & ~pi161;
  assign n33443 = ~n33441 & ~n33442;
  assign po247 = ~pi160 & ~n33443;
  assign n33445 = ~pi040 & ~pi161;
  assign n33446 = ~n33055 & ~n33056;
  assign n33447 = ~n831 & n33446;
  assign n33448 = ~pi313 & ~n33447;
  assign n33449 = n3319 & ~n33054;
  assign n33450 = ~n3319 & n33054;
  assign n33451 = ~n33449 & ~n33450;
  assign n33452 = ~n831 & ~n33451;
  assign n33453 = pi313 & n33452;
  assign n33454 = ~n33448 & ~n33453;
  assign n33455 = pi161 & ~n33454;
  assign n33456 = ~n33445 & ~n33455;
  assign po248 = ~pi160 & n33456;
  assign n33458 = ~pi039 & ~pi161;
  assign n33459 = ~n33051 & ~n33052;
  assign n33460 = ~n831 & n33459;
  assign n33461 = ~pi314 & ~n33460;
  assign n33462 = n3331 & ~n33050;
  assign n33463 = ~n3331 & n33050;
  assign n33464 = ~n33462 & ~n33463;
  assign n33465 = ~n831 & ~n33464;
  assign n33466 = pi314 & n33465;
  assign n33467 = ~n33461 & ~n33466;
  assign n33468 = pi161 & ~n33467;
  assign n33469 = ~n33458 & ~n33468;
  assign po249 = ~pi160 & n33469;
  assign n33471 = ~pi038 & ~pi161;
  assign n33472 = ~n33047 & ~n33048;
  assign n33473 = ~n831 & n33472;
  assign n33474 = ~pi315 & ~n33473;
  assign n33475 = n2852 & ~n33046;
  assign n33476 = ~n2852 & n33046;
  assign n33477 = ~n33475 & ~n33476;
  assign n33478 = ~n831 & ~n33477;
  assign n33479 = pi315 & n33478;
  assign n33480 = ~n33474 & ~n33479;
  assign n33481 = pi161 & ~n33480;
  assign n33482 = ~n33471 & ~n33481;
  assign po250 = ~pi160 & n33482;
  assign n33484 = ~pi037 & ~pi161;
  assign n33485 = ~n33043 & ~n33044;
  assign n33486 = ~n831 & n33485;
  assign n33487 = ~pi316 & ~n33486;
  assign n33488 = n2432 & ~n33042;
  assign n33489 = ~n2432 & n33042;
  assign n33490 = ~n33488 & ~n33489;
  assign n33491 = ~n831 & ~n33490;
  assign n33492 = pi316 & n33491;
  assign n33493 = ~n33487 & ~n33492;
  assign n33494 = pi161 & ~n33493;
  assign n33495 = ~n33484 & ~n33494;
  assign po251 = ~pi160 & n33495;
  assign n33497 = ~pi036 & ~pi161;
  assign n33498 = ~n33039 & ~n33040;
  assign n33499 = ~n831 & n33498;
  assign n33500 = ~pi317 & ~n33499;
  assign n33501 = n2070 & ~n33038;
  assign n33502 = ~n2070 & n33038;
  assign n33503 = ~n33501 & ~n33502;
  assign n33504 = ~n831 & ~n33503;
  assign n33505 = pi317 & n33504;
  assign n33506 = ~n33500 & ~n33505;
  assign n33507 = pi161 & ~n33506;
  assign n33508 = ~n33497 & ~n33507;
  assign po252 = ~pi160 & n33508;
  assign n33510 = pi035 & ~pi161;
  assign n33511 = pi318 & n831;
  assign n33512 = ~n1679 & n33034;
  assign n33513 = n1679 & ~n33034;
  assign n33514 = ~n33512 & ~n33513;
  assign n33515 = pi318 & ~n33514;
  assign n33516 = ~n33035 & ~n33036;
  assign n33517 = ~pi318 & ~n33516;
  assign n33518 = ~n33515 & ~n33517;
  assign n33519 = ~n831 & n33518;
  assign n33520 = ~n33511 & ~n33519;
  assign n33521 = pi161 & ~n33520;
  assign n33522 = ~n33510 & ~n33521;
  assign po253 = ~pi160 & ~n33522;
  assign n33524 = pi034 & ~pi161;
  assign n33525 = pi319 & n831;
  assign n33526 = pi319 & n1692;
  assign n33527 = ~pi319 & ~n1692;
  assign n33528 = ~n33526 & ~n33527;
  assign n33529 = ~n33032 & ~n33528;
  assign n33530 = pi320 & ~n1699;
  assign n33531 = ~n33026 & ~n33027;
  assign n33532 = ~n33028 & ~n33531;
  assign n33533 = ~n33530 & n33532;
  assign n33534 = n1699 & ~n33531;
  assign n33535 = ~pi320 & n33534;
  assign n33536 = ~n33533 & ~n33535;
  assign n33537 = ~n33529 & n33536;
  assign n33538 = ~n831 & n33537;
  assign n33539 = ~n33525 & ~n33538;
  assign n33540 = pi161 & ~n33539;
  assign n33541 = ~n33524 & ~n33540;
  assign po254 = ~pi160 & ~n33541;
  assign n33543 = pi033 & ~pi161;
  assign n33544 = pi320 & n831;
  assign n33545 = pi320 & n1699;
  assign n33546 = ~pi320 & ~n1699;
  assign n33547 = ~n33545 & ~n33546;
  assign n33548 = pi258 & ~n33547;
  assign n33549 = pi128 & n33548;
  assign n33550 = pi321 & n33549;
  assign n33551 = ~pi320 & n1699;
  assign n33552 = ~n33530 & ~n33551;
  assign n33553 = ~n33028 & ~n33552;
  assign n33554 = ~n33550 & ~n33553;
  assign n33555 = ~n831 & n33554;
  assign n33556 = ~n33544 & ~n33555;
  assign n33557 = pi161 & ~n33556;
  assign n33558 = ~n33543 & ~n33557;
  assign po255 = ~pi160 & ~n33558;
  assign n33560 = pi032 & ~pi161;
  assign n33561 = ~n831 & n1156;
  assign n33562 = ~pi321 & n33561;
  assign n33563 = pi321 & ~n33561;
  assign n33564 = ~n33562 & ~n33563;
  assign n33565 = pi161 & ~n33564;
  assign n33566 = ~n33560 & ~n33565;
  assign po256 = ~pi160 & ~n33566;
  assign n33568 = pi000 & ~pi161;
  assign n33569 = ~pi322 & ~n831;
  assign n33570 = pi128 & n33569;
  assign n33571 = pi128 & ~n831;
  assign n33572 = pi322 & ~n33571;
  assign n33573 = ~n33570 & ~n33572;
  assign n33574 = pi161 & ~n33573;
  assign n33575 = ~n33568 & ~n33574;
  assign po257 = ~pi160 & ~n33575;
  assign n33577 = pi001 & ~pi161;
  assign n33578 = pi323 & n831;
  assign n33579 = ~pi129 & pi323;
  assign n33580 = pi129 & ~pi323;
  assign n33581 = ~n33579 & ~n33580;
  assign n33582 = pi322 & ~n33581;
  assign n33583 = pi128 & n33582;
  assign n33584 = pi129 & pi323;
  assign n33585 = ~pi129 & ~pi323;
  assign n33586 = ~n33584 & ~n33585;
  assign n33587 = pi128 & pi322;
  assign n33588 = ~n33586 & ~n33587;
  assign n33589 = ~n33583 & ~n33588;
  assign n33590 = ~n831 & n33589;
  assign n33591 = ~n33578 & ~n33590;
  assign n33592 = pi161 & ~n33591;
  assign n33593 = ~n33577 & ~n33592;
  assign po258 = ~pi160 & ~n33593;
  assign n33595 = pi002 & ~pi161;
  assign n33596 = pi324 & n831;
  assign n33597 = pi130 & ~pi324;
  assign n33598 = ~pi130 & pi324;
  assign n33599 = ~n33597 & ~n33598;
  assign n33600 = pi322 & ~n33585;
  assign n33601 = pi128 & n33600;
  assign n33602 = ~n33584 & ~n33601;
  assign n33603 = ~n33599 & ~n33602;
  assign n33604 = pi130 & pi324;
  assign n33605 = ~pi130 & ~pi324;
  assign n33606 = ~n33604 & ~n33605;
  assign n33607 = ~n33584 & ~n33587;
  assign n33608 = ~n33585 & ~n33607;
  assign n33609 = ~n33606 & ~n33608;
  assign n33610 = ~n33603 & ~n33609;
  assign n33611 = ~n831 & n33610;
  assign n33612 = ~n33596 & ~n33611;
  assign n33613 = pi161 & ~n33612;
  assign n33614 = ~n33595 & ~n33613;
  assign po259 = ~pi160 & ~n33614;
  assign n33616 = pi003 & ~pi161;
  assign n33617 = pi325 & n831;
  assign n33618 = ~n33602 & ~n33605;
  assign n33619 = ~n33604 & ~n33618;
  assign n33620 = pi325 & n33619;
  assign n33621 = ~pi325 & ~n33619;
  assign n33622 = ~n33620 & ~n33621;
  assign n33623 = pi131 & ~n33622;
  assign n33624 = pi325 & ~n33619;
  assign n33625 = ~pi325 & n33619;
  assign n33626 = ~n33624 & ~n33625;
  assign n33627 = ~pi131 & ~n33626;
  assign n33628 = ~n33623 & ~n33627;
  assign n33629 = ~n831 & n33628;
  assign n33630 = ~n33617 & ~n33629;
  assign n33631 = pi161 & ~n33630;
  assign n33632 = ~n33616 & ~n33631;
  assign po260 = ~pi160 & ~n33632;
  assign n33634 = pi004 & ~pi161;
  assign n33635 = pi326 & n831;
  assign n33636 = ~pi132 & pi326;
  assign n33637 = pi132 & ~pi326;
  assign n33638 = ~n33636 & ~n33637;
  assign n33639 = pi131 & ~n33625;
  assign n33640 = ~n33624 & ~n33639;
  assign n33641 = ~n33638 & ~n33640;
  assign n33642 = pi132 & pi326;
  assign n33643 = ~pi132 & ~pi326;
  assign n33644 = ~n33642 & ~n33643;
  assign n33645 = ~pi131 & ~n33624;
  assign n33646 = ~n33625 & ~n33645;
  assign n33647 = ~n33644 & ~n33646;
  assign n33648 = ~n33641 & ~n33647;
  assign n33649 = ~n831 & n33648;
  assign n33650 = ~n33635 & ~n33649;
  assign n33651 = pi161 & ~n33650;
  assign n33652 = ~n33634 & ~n33651;
  assign po261 = ~pi160 & ~n33652;
  assign n33654 = pi005 & ~pi161;
  assign n33655 = pi327 & n831;
  assign n33656 = ~n33640 & ~n33643;
  assign n33657 = ~n33642 & ~n33656;
  assign n33658 = pi327 & n33657;
  assign n33659 = ~pi327 & ~n33657;
  assign n33660 = ~n33658 & ~n33659;
  assign n33661 = pi133 & ~n33660;
  assign n33662 = pi327 & ~n33657;
  assign n33663 = ~pi327 & n33657;
  assign n33664 = ~n33662 & ~n33663;
  assign n33665 = ~pi133 & ~n33664;
  assign n33666 = ~n33661 & ~n33665;
  assign n33667 = ~n831 & n33666;
  assign n33668 = ~n33655 & ~n33667;
  assign n33669 = pi161 & ~n33668;
  assign n33670 = ~n33654 & ~n33669;
  assign po262 = ~pi160 & ~n33670;
  assign n33672 = ~pi006 & ~pi161;
  assign n33673 = pi133 & ~n33663;
  assign n33674 = ~n33662 & ~n33673;
  assign n33675 = ~pi328 & ~n33674;
  assign n33676 = ~n831 & n33674;
  assign n33677 = pi328 & n33676;
  assign n33678 = ~n33675 & ~n33677;
  assign n33679 = pi134 & ~n33678;
  assign n33680 = ~pi328 & n831;
  assign n33681 = ~pi328 & n33674;
  assign n33682 = ~n831 & ~n33674;
  assign n33683 = pi328 & n33682;
  assign n33684 = ~n33681 & ~n33683;
  assign n33685 = ~pi134 & ~n33684;
  assign n33686 = ~n33680 & ~n33685;
  assign n33687 = ~n33679 & n33686;
  assign n33688 = pi161 & ~n33687;
  assign n33689 = ~n33672 & ~n33688;
  assign po263 = ~pi160 & n33689;
  assign n33691 = pi007 & ~pi161;
  assign n33692 = pi329 & n831;
  assign n33693 = pi328 & ~n33674;
  assign n33694 = pi134 & ~n33681;
  assign n33695 = ~n33693 & ~n33694;
  assign n33696 = pi329 & n33695;
  assign n33697 = ~pi329 & ~n33695;
  assign n33698 = ~n33696 & ~n33697;
  assign n33699 = pi135 & ~n33698;
  assign n33700 = pi329 & ~n33695;
  assign n33701 = ~pi329 & n33695;
  assign n33702 = ~n33700 & ~n33701;
  assign n33703 = ~pi135 & ~n33702;
  assign n33704 = ~n33699 & ~n33703;
  assign n33705 = ~n831 & n33704;
  assign n33706 = ~n33692 & ~n33705;
  assign n33707 = pi161 & ~n33706;
  assign n33708 = ~n33691 & ~n33707;
  assign po264 = ~pi160 & ~n33708;
  assign n33710 = pi008 & ~pi161;
  assign n33711 = pi330 & n831;
  assign n33712 = pi135 & ~n33701;
  assign n33713 = ~n33700 & ~n33712;
  assign n33714 = pi330 & n33713;
  assign n33715 = ~pi330 & ~n33713;
  assign n33716 = ~n33714 & ~n33715;
  assign n33717 = pi136 & ~n33716;
  assign n33718 = pi330 & ~n33713;
  assign n33719 = ~pi330 & n33713;
  assign n33720 = ~n33718 & ~n33719;
  assign n33721 = ~pi136 & ~n33720;
  assign n33722 = ~n33717 & ~n33721;
  assign n33723 = ~n831 & n33722;
  assign n33724 = ~n33711 & ~n33723;
  assign n33725 = pi161 & ~n33724;
  assign n33726 = ~n33710 & ~n33725;
  assign po265 = ~pi160 & ~n33726;
  assign n33728 = ~pi009 & ~pi161;
  assign n33729 = pi136 & ~n33719;
  assign n33730 = ~n33718 & ~n33729;
  assign n33731 = ~pi331 & ~n33730;
  assign n33732 = ~n831 & n33730;
  assign n33733 = pi331 & n33732;
  assign n33734 = ~n33731 & ~n33733;
  assign n33735 = pi137 & ~n33734;
  assign n33736 = ~pi331 & n831;
  assign n33737 = ~pi331 & n33730;
  assign n33738 = ~n831 & ~n33730;
  assign n33739 = pi331 & n33738;
  assign n33740 = ~n33737 & ~n33739;
  assign n33741 = ~pi137 & ~n33740;
  assign n33742 = ~n33736 & ~n33741;
  assign n33743 = ~n33735 & n33742;
  assign n33744 = pi161 & ~n33743;
  assign n33745 = ~n33728 & ~n33744;
  assign po266 = ~pi160 & n33745;
  assign n33747 = ~pi010 & ~pi161;
  assign n33748 = pi331 & ~n33730;
  assign n33749 = pi137 & ~n33737;
  assign n33750 = ~n33748 & ~n33749;
  assign n33751 = ~pi332 & ~n33750;
  assign n33752 = ~n831 & n33750;
  assign n33753 = pi332 & n33752;
  assign n33754 = ~n33751 & ~n33753;
  assign n33755 = pi138 & ~n33754;
  assign n33756 = ~pi332 & n831;
  assign n33757 = ~pi332 & n33750;
  assign n33758 = ~n831 & ~n33750;
  assign n33759 = pi332 & n33758;
  assign n33760 = ~n33757 & ~n33759;
  assign n33761 = ~pi138 & ~n33760;
  assign n33762 = ~n33756 & ~n33761;
  assign n33763 = ~n33755 & n33762;
  assign n33764 = pi161 & ~n33763;
  assign n33765 = ~n33747 & ~n33764;
  assign po267 = ~pi160 & n33765;
  assign n33767 = ~pi011 & ~pi161;
  assign n33768 = pi332 & ~n33750;
  assign n33769 = pi138 & ~n33757;
  assign n33770 = ~n33768 & ~n33769;
  assign n33771 = ~pi333 & ~n33770;
  assign n33772 = ~n831 & n33770;
  assign n33773 = pi333 & n33772;
  assign n33774 = ~n33771 & ~n33773;
  assign n33775 = pi139 & ~n33774;
  assign n33776 = ~pi333 & n831;
  assign n33777 = ~pi333 & n33770;
  assign n33778 = ~n831 & ~n33770;
  assign n33779 = pi333 & n33778;
  assign n33780 = ~n33777 & ~n33779;
  assign n33781 = ~pi139 & ~n33780;
  assign n33782 = ~n33776 & ~n33781;
  assign n33783 = ~n33775 & n33782;
  assign n33784 = pi161 & ~n33783;
  assign n33785 = ~n33767 & ~n33784;
  assign po268 = ~pi160 & n33785;
  assign n33787 = ~pi012 & ~pi161;
  assign n33788 = pi333 & ~n33770;
  assign n33789 = pi139 & ~n33777;
  assign n33790 = ~n33788 & ~n33789;
  assign n33791 = ~pi334 & ~n33790;
  assign n33792 = ~n831 & n33790;
  assign n33793 = pi334 & n33792;
  assign n33794 = ~n33791 & ~n33793;
  assign n33795 = pi140 & ~n33794;
  assign n33796 = ~pi334 & n831;
  assign n33797 = ~pi334 & n33790;
  assign n33798 = ~n831 & ~n33790;
  assign n33799 = pi334 & n33798;
  assign n33800 = ~n33797 & ~n33799;
  assign n33801 = ~pi140 & ~n33800;
  assign n33802 = ~n33796 & ~n33801;
  assign n33803 = ~n33795 & n33802;
  assign n33804 = pi161 & ~n33803;
  assign n33805 = ~n33787 & ~n33804;
  assign po269 = ~pi160 & n33805;
  assign n33807 = ~pi013 & ~pi161;
  assign n33808 = pi334 & ~n33790;
  assign n33809 = pi140 & ~n33797;
  assign n33810 = ~n33808 & ~n33809;
  assign n33811 = ~pi335 & ~n33810;
  assign n33812 = ~n831 & n33810;
  assign n33813 = pi335 & n33812;
  assign n33814 = ~n33811 & ~n33813;
  assign n33815 = pi141 & ~n33814;
  assign n33816 = ~pi335 & n831;
  assign n33817 = ~pi335 & n33810;
  assign n33818 = ~n831 & ~n33810;
  assign n33819 = pi335 & n33818;
  assign n33820 = ~n33817 & ~n33819;
  assign n33821 = ~pi141 & ~n33820;
  assign n33822 = ~n33816 & ~n33821;
  assign n33823 = ~n33815 & n33822;
  assign n33824 = pi161 & ~n33823;
  assign n33825 = ~n33807 & ~n33824;
  assign po270 = ~pi160 & n33825;
  assign n33827 = ~pi014 & ~pi161;
  assign n33828 = pi335 & ~n33810;
  assign n33829 = pi141 & ~n33817;
  assign n33830 = ~n33828 & ~n33829;
  assign n33831 = ~pi336 & ~n33830;
  assign n33832 = ~n831 & n33830;
  assign n33833 = pi336 & n33832;
  assign n33834 = ~n33831 & ~n33833;
  assign n33835 = pi142 & ~n33834;
  assign n33836 = ~pi336 & n831;
  assign n33837 = ~pi336 & n33830;
  assign n33838 = ~n831 & ~n33830;
  assign n33839 = pi336 & n33838;
  assign n33840 = ~n33837 & ~n33839;
  assign n33841 = ~pi142 & ~n33840;
  assign n33842 = ~n33836 & ~n33841;
  assign n33843 = ~n33835 & n33842;
  assign n33844 = pi161 & ~n33843;
  assign n33845 = ~n33827 & ~n33844;
  assign po271 = ~pi160 & n33845;
  assign n33847 = ~pi015 & ~pi161;
  assign n33848 = pi336 & ~n33830;
  assign n33849 = pi142 & ~n33837;
  assign n33850 = ~n33848 & ~n33849;
  assign n33851 = ~pi337 & ~n33850;
  assign n33852 = ~n831 & n33850;
  assign n33853 = pi337 & n33852;
  assign n33854 = ~n33851 & ~n33853;
  assign n33855 = pi143 & ~n33854;
  assign n33856 = ~pi337 & n831;
  assign n33857 = ~pi337 & n33850;
  assign n33858 = ~n831 & ~n33850;
  assign n33859 = pi337 & n33858;
  assign n33860 = ~n33857 & ~n33859;
  assign n33861 = ~pi143 & ~n33860;
  assign n33862 = ~n33856 & ~n33861;
  assign n33863 = ~n33855 & n33862;
  assign n33864 = pi161 & ~n33863;
  assign n33865 = ~n33847 & ~n33864;
  assign po272 = ~pi160 & n33865;
  assign n33867 = ~pi016 & ~pi161;
  assign n33868 = pi337 & ~n33850;
  assign n33869 = pi143 & ~n33857;
  assign n33870 = ~n33868 & ~n33869;
  assign n33871 = ~pi338 & ~n33870;
  assign n33872 = ~n831 & n33870;
  assign n33873 = pi338 & n33872;
  assign n33874 = ~n33871 & ~n33873;
  assign n33875 = pi144 & ~n33874;
  assign n33876 = ~pi338 & n831;
  assign n33877 = ~pi338 & n33870;
  assign n33878 = ~n831 & ~n33870;
  assign n33879 = pi338 & n33878;
  assign n33880 = ~n33877 & ~n33879;
  assign n33881 = ~pi144 & ~n33880;
  assign n33882 = ~n33876 & ~n33881;
  assign n33883 = ~n33875 & n33882;
  assign n33884 = pi161 & ~n33883;
  assign n33885 = ~n33867 & ~n33884;
  assign po273 = ~pi160 & n33885;
  assign n33887 = ~pi017 & ~pi161;
  assign n33888 = pi338 & ~n33870;
  assign n33889 = pi144 & ~n33877;
  assign n33890 = ~n33888 & ~n33889;
  assign n33891 = ~pi339 & ~n33890;
  assign n33892 = ~n831 & n33890;
  assign n33893 = pi339 & n33892;
  assign n33894 = ~n33891 & ~n33893;
  assign n33895 = pi145 & ~n33894;
  assign n33896 = ~pi339 & n831;
  assign n33897 = ~pi339 & n33890;
  assign n33898 = ~n831 & ~n33890;
  assign n33899 = pi339 & n33898;
  assign n33900 = ~n33897 & ~n33899;
  assign n33901 = ~pi145 & ~n33900;
  assign n33902 = ~n33896 & ~n33901;
  assign n33903 = ~n33895 & n33902;
  assign n33904 = pi161 & ~n33903;
  assign n33905 = ~n33887 & ~n33904;
  assign po274 = ~pi160 & n33905;
  assign n33907 = ~pi018 & ~pi161;
  assign n33908 = pi339 & ~n33890;
  assign n33909 = pi145 & ~n33897;
  assign n33910 = ~n33908 & ~n33909;
  assign n33911 = ~pi340 & ~n33910;
  assign n33912 = ~n831 & n33910;
  assign n33913 = pi340 & n33912;
  assign n33914 = ~n33911 & ~n33913;
  assign n33915 = pi146 & ~n33914;
  assign n33916 = ~pi340 & n831;
  assign n33917 = ~pi340 & n33910;
  assign n33918 = ~n831 & ~n33910;
  assign n33919 = pi340 & n33918;
  assign n33920 = ~n33917 & ~n33919;
  assign n33921 = ~pi146 & ~n33920;
  assign n33922 = ~n33916 & ~n33921;
  assign n33923 = ~n33915 & n33922;
  assign n33924 = pi161 & ~n33923;
  assign n33925 = ~n33907 & ~n33924;
  assign po275 = ~pi160 & n33925;
  assign n33927 = ~pi019 & ~pi161;
  assign n33928 = pi340 & ~n33910;
  assign n33929 = pi146 & ~n33917;
  assign n33930 = ~n33928 & ~n33929;
  assign n33931 = ~pi341 & ~n33930;
  assign n33932 = ~n831 & n33930;
  assign n33933 = pi341 & n33932;
  assign n33934 = ~n33931 & ~n33933;
  assign n33935 = pi147 & ~n33934;
  assign n33936 = ~pi341 & n831;
  assign n33937 = ~pi341 & n33930;
  assign n33938 = ~n831 & ~n33930;
  assign n33939 = pi341 & n33938;
  assign n33940 = ~n33937 & ~n33939;
  assign n33941 = ~pi147 & ~n33940;
  assign n33942 = ~n33936 & ~n33941;
  assign n33943 = ~n33935 & n33942;
  assign n33944 = pi161 & ~n33943;
  assign n33945 = ~n33927 & ~n33944;
  assign po276 = ~pi160 & n33945;
  assign n33947 = ~pi020 & ~pi161;
  assign n33948 = pi341 & ~n33930;
  assign n33949 = pi147 & ~n33937;
  assign n33950 = ~n33948 & ~n33949;
  assign n33951 = ~pi342 & ~n33950;
  assign n33952 = ~n831 & n33950;
  assign n33953 = pi342 & n33952;
  assign n33954 = ~n33951 & ~n33953;
  assign n33955 = pi148 & ~n33954;
  assign n33956 = ~pi342 & n831;
  assign n33957 = ~pi342 & n33950;
  assign n33958 = ~n831 & ~n33950;
  assign n33959 = pi342 & n33958;
  assign n33960 = ~n33957 & ~n33959;
  assign n33961 = ~pi148 & ~n33960;
  assign n33962 = ~n33956 & ~n33961;
  assign n33963 = ~n33955 & n33962;
  assign n33964 = pi161 & ~n33963;
  assign n33965 = ~n33947 & ~n33964;
  assign po277 = ~pi160 & n33965;
  assign n33967 = ~pi021 & ~pi161;
  assign n33968 = pi342 & ~n33950;
  assign n33969 = pi148 & ~n33957;
  assign n33970 = ~n33968 & ~n33969;
  assign n33971 = ~pi343 & ~n33970;
  assign n33972 = ~n831 & n33970;
  assign n33973 = pi343 & n33972;
  assign n33974 = ~n33971 & ~n33973;
  assign n33975 = pi149 & ~n33974;
  assign n33976 = ~pi343 & n831;
  assign n33977 = ~pi343 & n33970;
  assign n33978 = ~n831 & ~n33970;
  assign n33979 = pi343 & n33978;
  assign n33980 = ~n33977 & ~n33979;
  assign n33981 = ~pi149 & ~n33980;
  assign n33982 = ~n33976 & ~n33981;
  assign n33983 = ~n33975 & n33982;
  assign n33984 = pi161 & ~n33983;
  assign n33985 = ~n33967 & ~n33984;
  assign po278 = ~pi160 & n33985;
  assign n33987 = ~pi022 & ~pi161;
  assign n33988 = pi343 & ~n33970;
  assign n33989 = pi149 & ~n33977;
  assign n33990 = ~n33988 & ~n33989;
  assign n33991 = ~pi344 & ~n33990;
  assign n33992 = ~n831 & n33990;
  assign n33993 = pi344 & n33992;
  assign n33994 = ~n33991 & ~n33993;
  assign n33995 = pi150 & ~n33994;
  assign n33996 = ~pi344 & n831;
  assign n33997 = ~pi344 & n33990;
  assign n33998 = ~n831 & ~n33990;
  assign n33999 = pi344 & n33998;
  assign n34000 = ~n33997 & ~n33999;
  assign n34001 = ~pi150 & ~n34000;
  assign n34002 = ~n33996 & ~n34001;
  assign n34003 = ~n33995 & n34002;
  assign n34004 = pi161 & ~n34003;
  assign n34005 = ~n33987 & ~n34004;
  assign po279 = ~pi160 & n34005;
  assign n34007 = ~pi023 & ~pi161;
  assign n34008 = pi344 & ~n33990;
  assign n34009 = pi150 & ~n33997;
  assign n34010 = ~n34008 & ~n34009;
  assign n34011 = ~pi345 & ~n34010;
  assign n34012 = ~n831 & n34010;
  assign n34013 = pi345 & n34012;
  assign n34014 = ~n34011 & ~n34013;
  assign n34015 = pi151 & ~n34014;
  assign n34016 = ~pi345 & n831;
  assign n34017 = ~pi345 & n34010;
  assign n34018 = ~n831 & ~n34010;
  assign n34019 = pi345 & n34018;
  assign n34020 = ~n34017 & ~n34019;
  assign n34021 = ~pi151 & ~n34020;
  assign n34022 = ~n34016 & ~n34021;
  assign n34023 = ~n34015 & n34022;
  assign n34024 = pi161 & ~n34023;
  assign n34025 = ~n34007 & ~n34024;
  assign po280 = ~pi160 & n34025;
  assign n34027 = ~pi024 & ~pi161;
  assign n34028 = pi345 & ~n34010;
  assign n34029 = pi151 & ~n34017;
  assign n34030 = ~n34028 & ~n34029;
  assign n34031 = ~pi346 & ~n34030;
  assign n34032 = ~n831 & n34030;
  assign n34033 = pi346 & n34032;
  assign n34034 = ~n34031 & ~n34033;
  assign n34035 = pi152 & ~n34034;
  assign n34036 = ~pi346 & n831;
  assign n34037 = ~pi346 & n34030;
  assign n34038 = ~n831 & ~n34030;
  assign n34039 = pi346 & n34038;
  assign n34040 = ~n34037 & ~n34039;
  assign n34041 = ~pi152 & ~n34040;
  assign n34042 = ~n34036 & ~n34041;
  assign n34043 = ~n34035 & n34042;
  assign n34044 = pi161 & ~n34043;
  assign n34045 = ~n34027 & ~n34044;
  assign po281 = ~pi160 & n34045;
  assign n34047 = ~pi025 & ~pi161;
  assign n34048 = pi346 & ~n34030;
  assign n34049 = pi152 & ~n34037;
  assign n34050 = ~n34048 & ~n34049;
  assign n34051 = ~pi347 & ~n34050;
  assign n34052 = ~n831 & n34050;
  assign n34053 = pi347 & n34052;
  assign n34054 = ~n34051 & ~n34053;
  assign n34055 = pi153 & ~n34054;
  assign n34056 = ~pi347 & n831;
  assign n34057 = ~pi347 & n34050;
  assign n34058 = ~n831 & ~n34050;
  assign n34059 = pi347 & n34058;
  assign n34060 = ~n34057 & ~n34059;
  assign n34061 = ~pi153 & ~n34060;
  assign n34062 = ~n34056 & ~n34061;
  assign n34063 = ~n34055 & n34062;
  assign n34064 = pi161 & ~n34063;
  assign n34065 = ~n34047 & ~n34064;
  assign po282 = ~pi160 & n34065;
  assign n34067 = ~pi026 & ~pi161;
  assign n34068 = pi347 & ~n34050;
  assign n34069 = pi153 & ~n34057;
  assign n34070 = ~n34068 & ~n34069;
  assign n34071 = ~pi348 & ~n34070;
  assign n34072 = ~n831 & n34070;
  assign n34073 = pi348 & n34072;
  assign n34074 = ~n34071 & ~n34073;
  assign n34075 = pi154 & ~n34074;
  assign n34076 = ~pi348 & n831;
  assign n34077 = ~pi348 & n34070;
  assign n34078 = ~n831 & ~n34070;
  assign n34079 = pi348 & n34078;
  assign n34080 = ~n34077 & ~n34079;
  assign n34081 = ~pi154 & ~n34080;
  assign n34082 = ~n34076 & ~n34081;
  assign n34083 = ~n34075 & n34082;
  assign n34084 = pi161 & ~n34083;
  assign n34085 = ~n34067 & ~n34084;
  assign po283 = ~pi160 & n34085;
  assign n34087 = ~pi027 & ~pi161;
  assign n34088 = pi348 & ~n34070;
  assign n34089 = pi154 & ~n34077;
  assign n34090 = ~n34088 & ~n34089;
  assign n34091 = ~pi349 & ~n34090;
  assign n34092 = ~n831 & n34090;
  assign n34093 = pi349 & n34092;
  assign n34094 = ~n34091 & ~n34093;
  assign n34095 = pi155 & ~n34094;
  assign n34096 = ~pi349 & n831;
  assign n34097 = ~pi349 & n34090;
  assign n34098 = ~n831 & ~n34090;
  assign n34099 = pi349 & n34098;
  assign n34100 = ~n34097 & ~n34099;
  assign n34101 = ~pi155 & ~n34100;
  assign n34102 = ~n34096 & ~n34101;
  assign n34103 = ~n34095 & n34102;
  assign n34104 = pi161 & ~n34103;
  assign n34105 = ~n34087 & ~n34104;
  assign po284 = ~pi160 & n34105;
  assign n34107 = ~pi028 & ~pi161;
  assign n34108 = pi349 & ~n34090;
  assign n34109 = pi155 & ~n34097;
  assign n34110 = ~n34108 & ~n34109;
  assign n34111 = ~pi350 & ~n34110;
  assign n34112 = ~n831 & n34110;
  assign n34113 = pi350 & n34112;
  assign n34114 = ~n34111 & ~n34113;
  assign n34115 = pi156 & ~n34114;
  assign n34116 = ~pi350 & n831;
  assign n34117 = ~pi350 & n34110;
  assign n34118 = ~n831 & ~n34110;
  assign n34119 = pi350 & n34118;
  assign n34120 = ~n34117 & ~n34119;
  assign n34121 = ~pi156 & ~n34120;
  assign n34122 = ~n34116 & ~n34121;
  assign n34123 = ~n34115 & n34122;
  assign n34124 = pi161 & ~n34123;
  assign n34125 = ~n34107 & ~n34124;
  assign po285 = ~pi160 & n34125;
  assign n34127 = ~pi029 & ~pi161;
  assign n34128 = pi350 & ~n34110;
  assign n34129 = pi156 & ~n34117;
  assign n34130 = ~n34128 & ~n34129;
  assign n34131 = ~pi351 & ~n34130;
  assign n34132 = ~n831 & n34130;
  assign n34133 = pi351 & n34132;
  assign n34134 = ~n34131 & ~n34133;
  assign n34135 = pi157 & ~n34134;
  assign n34136 = ~pi351 & n831;
  assign n34137 = ~pi351 & n34130;
  assign n34138 = ~n831 & ~n34130;
  assign n34139 = pi351 & n34138;
  assign n34140 = ~n34137 & ~n34139;
  assign n34141 = ~pi157 & ~n34140;
  assign n34142 = ~n34136 & ~n34141;
  assign n34143 = ~n34135 & n34142;
  assign n34144 = pi161 & ~n34143;
  assign n34145 = ~n34127 & ~n34144;
  assign po286 = ~pi160 & n34145;
  assign n34147 = pi030 & ~pi161;
  assign n34148 = pi351 & ~n34130;
  assign n34149 = pi157 & ~n34137;
  assign n34150 = ~n34148 & ~n34149;
  assign n34151 = pi352 & ~n34150;
  assign n34152 = ~pi352 & n34150;
  assign n34153 = ~n34151 & ~n34152;
  assign n34154 = pi158 & ~n34153;
  assign n34155 = ~pi352 & ~n34150;
  assign n34156 = pi352 & n34150;
  assign n34157 = ~n34155 & ~n34156;
  assign n34158 = ~pi158 & ~n34157;
  assign n34159 = ~n34154 & ~n34158;
  assign n34160 = ~n831 & ~n34159;
  assign n34161 = ~n1006 & ~n34160;
  assign n34162 = pi161 & ~n34161;
  assign n34163 = ~n34147 & ~n34162;
  assign po287 = ~pi160 & ~n34163;
  assign n34165 = pi031 & ~pi161;
  assign n34166 = pi158 & ~n34152;
  assign n34167 = ~n34151 & ~n34166;
  assign n34168 = ~pi159 & ~n34167;
  assign n34169 = ~pi158 & ~n34151;
  assign n34170 = ~n34152 & ~n34169;
  assign n34171 = pi159 & ~n34170;
  assign n34172 = ~n34168 & ~n34171;
  assign n34173 = ~n831 & ~n34172;
  assign n34174 = ~pi353 & n34173;
  assign n34175 = pi353 & ~n34173;
  assign n34176 = ~n34174 & ~n34175;
  assign n34177 = pi161 & ~n34176;
  assign n34178 = ~n34165 & ~n34177;
  assign po288 = ~pi160 & ~n34178;
  assign po000 = pi194;
  assign po001 = pi195;
  assign po002 = pi206;
  assign po003 = pi217;
  assign po004 = pi220;
  assign po005 = pi221;
  assign po006 = pi222;
  assign po007 = pi223;
  assign po008 = pi224;
  assign po009 = pi225;
  assign po010 = pi196;
  assign po011 = pi197;
  assign po012 = pi198;
  assign po013 = pi199;
  assign po014 = pi200;
  assign po015 = pi201;
  assign po016 = pi202;
  assign po017 = pi203;
  assign po018 = pi204;
  assign po019 = pi205;
  assign po020 = pi207;
  assign po021 = pi208;
  assign po022 = pi209;
  assign po023 = pi210;
  assign po024 = pi211;
  assign po025 = pi212;
  assign po026 = pi213;
  assign po027 = pi214;
  assign po028 = pi215;
  assign po029 = pi216;
  assign po030 = pi218;
  assign po031 = pi219;
  assign po032 = pi226;
  assign po033 = pi227;
  assign po034 = pi238;
  assign po035 = pi249;
  assign po036 = pi252;
  assign po037 = pi253;
  assign po038 = pi254;
  assign po039 = pi255;
  assign po040 = pi256;
  assign po041 = pi257;
  assign po042 = pi228;
  assign po043 = pi229;
  assign po044 = pi230;
  assign po045 = pi231;
  assign po046 = pi232;
  assign po047 = pi233;
  assign po048 = pi234;
  assign po049 = pi235;
  assign po050 = pi236;
  assign po051 = pi237;
  assign po052 = pi239;
  assign po053 = pi240;
  assign po054 = pi241;
  assign po055 = pi242;
  assign po056 = pi243;
  assign po057 = pi244;
  assign po058 = pi245;
  assign po059 = pi246;
  assign po060 = pi247;
  assign po061 = pi248;
  assign po062 = pi250;
  assign po063 = pi251;
  assign po064 = pi162;
  assign po065 = pi163;
  assign po066 = pi174;
  assign po067 = pi185;
  assign po068 = pi188;
  assign po069 = pi189;
  assign po070 = pi190;
  assign po071 = pi191;
  assign po072 = pi192;
  assign po073 = pi193;
  assign po074 = pi164;
  assign po075 = pi165;
  assign po076 = pi166;
  assign po077 = pi167;
  assign po078 = pi168;
  assign po079 = pi169;
  assign po080 = pi170;
  assign po081 = pi171;
  assign po082 = pi172;
  assign po083 = pi173;
  assign po084 = pi175;
  assign po085 = pi176;
  assign po086 = pi177;
  assign po087 = pi178;
  assign po088 = pi179;
  assign po089 = pi180;
  assign po090 = pi181;
  assign po091 = pi182;
  assign po092 = pi183;
  assign po093 = pi184;
  assign po094 = pi186;
  assign po095 = pi187;
endmodule


