//Written by the Majority Logic Package Thu Apr 30 23:14:44 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89, pi90, pi91, pi92, pi93, pi94, pi95;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, v802, v803, v804, v805, v806, v807, v808, v809, v810, v811, v812, v813, v814, v815, v816, v817, v818, v819, v820, v821, v822, v823, v824, v825, v826, v827, v828, v829, v830, v831, v832, v833, v834, v835, v836, v837, v838, v839, v840, v841, v842, v843, v844, v845, v846, v847, v848, v849, v850, v851, v852, v853, v854, v855, v856, v857, v858, v859, v860, v861, v862, v863, v864, v865, v866, v867, v868, v869, v870, v871, v872, v873, v874, v875, v876, v877, v878, v879, v880, v881, v882, v883, v884, v885, v886, v887, v888, v889, v890, v891, v892, v893, v894, v895, v896, v897, v898, v899, v900, v901, v902, v903, v904, v905, v906, v907, v908, v909, v910, v911, v912, v913, v914, v915, v916, v917, v918, v919, v920, v921, v922, v923, v924, v925, v926, v927, v928, v929, v930, v931, v932, v933, v934, v935, v936, v937, v938, v939, v940, v941, v942, v943, v944, v945, v946, v947, v948, v949, v950, v951, v952, v953, v954, v955, v956, v957, v958, v959, v960, v961, v962, v963, v964, v965, v966, v967, v968, v969, v970, v971, v972, v973, v974, v975, v976, v977, v978, v979, v980, v981, v982, v983, v984, v985, v986, v987, v988, v989, v990, v991, v992, v993, v994, v995, v996, v997, v998, v999, v1000, v1001, v1002, v1003, v1004, v1005, v1006, v1007, v1008, v1009, v1010, v1011, v1012, v1013, v1014, v1015, v1016, v1017, v1018, v1019, v1020, v1021, v1022, v1023, v1024, v1025, v1026, v1027, v1028, v1029, v1030, v1031, v1032, v1033, v1034, v1035, v1036, v1037, v1038, v1039, v1040, v1041, v1042, v1043, v1044, v1045, v1046, v1047, v1048, v1049, v1050, v1051, v1052, v1053, v1054, v1055, v1056, v1057, v1058, v1059, v1060, v1061, v1062, v1063, v1064, v1065, v1066, v1067, v1068, v1069, v1070, v1071, v1072, v1073, v1074, v1075, v1076, v1077, v1078, v1079, v1080, v1081, v1082, v1083, v1084, v1085, v1086, v1087, v1088, v1089, v1090, v1091, v1092, v1093, v1094, v1095, v1096, v1097, v1098, v1099, v1100, v1101, v1102, v1103, v1104, v1105, v1106, v1107, v1108, v1109, v1110, v1111, v1112, v1113, v1114, v1115, v1116, v1117, v1118, v1119, v1120, v1121, v1122, v1123, v1124, v1125, v1126, v1127, v1128, v1129, v1130, v1131, v1132, v1133, v1134, v1135, v1136, v1137, v1138, v1139, v1140, v1141, v1142, v1143, v1144, v1145, v1146, v1147, v1148, v1149, v1150, v1151, v1152, v1153, v1154, v1155, v1156, v1157, v1158, v1159, v1160, v1161, v1162, v1163, v1164, v1165, v1166, v1167, v1168, v1169, v1170, v1171, v1172, v1173, v1174, v1175, v1176, v1177, v1178, v1179, v1180, v1181, v1182, v1183, v1184, v1185, v1186, v1187, v1188, v1189, v1190, v1191, v1192, v1193, v1194, v1195, v1196, v1197, v1198, v1199, v1200, v1201, v1202, v1203, v1204, v1205, v1206, v1207, v1208, v1209, v1210, v1211, v1212, v1213, v1214, v1215, v1216, v1217, v1218, v1219, v1220, v1221, v1222, v1223, v1224, v1225, v1226, v1227, v1228, v1229, v1230, v1231, v1232, v1233, v1234, v1235, v1236, v1237, v1238, v1239, v1240, v1241, v1242, v1243, v1244, v1245, v1246, v1247, v1248, v1249, v1250, v1251, v1252, v1253, v1254, v1255, v1256, v1257, v1258, v1259, v1260, v1261, v1262, v1263, v1264, v1265, v1266, v1267, v1268, v1269, v1270, v1271, v1272, v1273, v1274, v1275, v1276, v1277, v1278, v1279, v1280, v1281, v1282, v1283, v1284, v1285, v1286, v1287, v1288, v1289, v1290, v1291, v1292, v1293, v1294, v1295, v1296, v1297, v1298, v1299, v1300, v1301, v1302, v1303, v1304, v1305, v1306, v1307, v1308, v1309, v1310, v1311, v1312, v1313, v1314, v1315, v1316, v1317, v1318, v1319, v1320, v1321, v1322, v1323, v1324, v1325, v1326, v1327, v1328, v1329, v1330, v1331, v1332, v1333, v1334, v1335, v1336, v1337, v1338, v1339, v1340, v1341, v1342, v1343, v1344, v1345, v1346, v1347, v1348, v1349, v1350, v1351, v1352, v1353, v1354, v1355, v1356, v1357, v1358, v1359, v1360, v1361, v1362, v1363, v1364, v1365, v1366, v1367, v1368, v1369, v1370, v1371, v1372, v1373, v1374, v1375, v1376, v1377, v1378, v1379, v1380, v1381, v1382, v1383, v1384, v1385, v1386, v1387, v1388, v1389, v1390, v1391, v1392, v1393, v1394, v1395, v1396, v1397, v1398, v1399, v1400, v1401, v1402, v1403, v1404, v1405, v1406, v1407, v1408, v1409, v1410, v1411, v1412, v1413, v1414, v1415, v1416, v1417, v1418, v1419, v1420, v1421, v1422, v1423, v1424, v1425, v1426, v1427, v1428, v1429, v1430, v1431, v1432, v1433, v1434, v1435, v1436, v1437, v1438, v1439, v1440, v1441, v1442, v1443, v1444, v1445, v1446, v1447, v1448, v1449, v1450, v1451, v1452, v1453, v1454, v1455, v1456, v1457, v1458, v1459, v1460, v1461, v1462, v1463, v1464, v1465, v1466, v1467, v1468, v1469, v1470, v1471, v1472, v1473, v1474, v1475, v1476, v1477, v1478, v1479, v1480, v1481, v1482, v1483, v1484, v1485, v1486, v1487, v1488, v1489, v1490, v1491, v1492, v1493, v1494, v1495, v1496, v1497, v1498, v1499, v1500, v1501, v1502, v1503, v1504, v1505, v1506, v1507, v1508, v1509, v1510, v1511, v1512, v1513, v1514, v1515, v1516, v1517, v1518, v1519, v1520, v1521, v1522, v1523, v1524, v1525, v1526, v1527, v1528, v1529, v1530, v1531, v1532, v1533, v1534, v1535, v1536, v1537, v1538, v1539, v1540, v1541, v1542, v1543, v1544, v1545, v1546, v1547, v1548, v1549, v1550, v1551, v1552, v1553, v1554, v1555, v1556, v1557, v1558, v1559, v1560, v1561, v1562, v1563, v1564, v1565, v1566, v1567, v1568, v1569, v1570, v1571, v1572, v1573, v1574, v1575, v1576, v1577, v1578, v1579, v1580, v1581, v1582, v1583, v1584, v1585, v1586, v1587, v1588, v1589, v1590, v1591, v1592, v1593, v1594, v1595, v1596, v1597, v1598, v1599, v1600, v1601, v1602, v1603, v1604, v1605, v1606, v1607, v1608, v1609, v1610, v1611, v1612, v1613, v1614, v1615, v1616, v1617, v1618, v1619, v1620, v1621, v1622, v1623, v1624, v1625, v1626, v1627, v1628, v1629, v1630, v1631, v1632, v1633, v1634, v1635, v1636, v1637, v1638, v1639, v1640, v1641, v1642, v1643, v1644, v1645, v1646, v1647, v1648, v1649, v1650, v1651, v1652, v1653, v1654, v1655, v1656, v1657, v1658, v1659, v1660, v1661, v1662, v1663, v1664, v1665, v1666, v1667, v1668, v1669, v1670, v1671, v1672, v1673, v1674, v1675, v1676, v1677, v1678, v1679, v1680, v1681, v1682, v1683, v1684, v1685, v1686, v1687, v1688, v1689, v1690, v1691, v1692, v1693, v1694, v1695, v1696, v1697, v1698, v1699, v1700, v1701, v1702, v1703, v1704, v1705, v1706, v1707, v1708, v1709, v1710, v1711, v1712, v1713, v1714, v1715, v1716, v1717, v1718, v1719, v1720, v1721, v1722, v1723, v1724, v1725, v1726, v1727, v1728, v1729, v1730, v1731, v1732, v1733, v1734, v1735, v1736, v1737, v1738, v1739, v1740, v1741, v1742, v1743, v1744, v1745, v1746, v1747, v1748, v1749, v1750, v1751, v1752, v1753, v1754, v1755, v1756, v1757, v1758, v1759, v1760, v1761, v1762, v1763, v1764, v1765, v1766, v1767, v1768, v1769, v1770, v1771, v1772, v1773, v1774, v1775, v1776, v1777, v1778, v1779, v1780, v1781, v1782, v1783, v1784, v1785, v1786, v1787, v1788, v1789, v1790, v1791, v1792, v1793, v1794, v1795, v1796, v1797, v1798, v1799, v1800, v1801, v1802, v1803, v1804, v1805, v1806, v1807, v1808, v1809, v1810, v1811, v1812, v1813, v1814, v1815, v1816, v1817, v1818, v1819, v1820, v1821, v1822, v1823, v1824, v1825, v1826, v1827, v1828, v1829, v1830, v1831, v1832, v1833, v1834, v1835, v1836, v1837, v1838, v1839, v1840, v1841, v1842, v1843, v1844, v1845, v1846, v1847, v1848, v1849, v1850, v1851, v1852, v1853, v1854, v1855, v1856, v1857, v1858, v1859, v1860, v1861, v1862, v1863, v1864, v1865, v1866, v1867, v1868, v1869, v1870, v1871, v1872, v1873, v1874, v1875, v1876, v1877, v1878, v1879, v1880, v1881, v1882, v1883, v1884, v1885, v1886, v1887, v1888, v1889, v1890, v1891, v1892, v1893, v1894, v1895, v1896, v1897, v1898, v1899, v1900, v1901, v1902, v1903, v1904, v1905, v1906, v1907, v1908, v1909, v1910, v1911, v1912, v1913, v1914, v1915, v1916, v1917, v1918, v1919, v1920, v1921, v1922, v1923, v1924, v1925, v1926, v1927, v1928, v1929, v1930, v1931, v1932, v1933, v1934, v1935, v1936, v1937, v1938, v1939, v1940, v1941, v1942, v1943, v1944, v1945, v1946, v1947, v1948, v1949, v1950, v1951, v1952, v1953, v1954, v1955, v1956, v1957, v1958, v1959, v1960, v1961, v1962, v1963, v1964, v1965, v1966, v1967, v1968, v1969, v1970, v1971, v1972, v1973, v1974, v1975, v1976, v1977, v1978, v1979, v1980, v1981, v1982, v1983, v1984, v1985, v1986, v1987, v1988, v1989, v1990, v1991, v1992, v1993, v1994, v1995, v1996, v1997, v1998, v1999, v2000, v2001, v2002, v2003, v2004, v2005, v2006, v2007, v2008, v2009, v2010, v2011, v2012, v2013, v2014, v2015, v2016, v2017, v2018, v2019, v2020, v2021, v2022, v2023, v2024, v2025, v2026, v2027, v2028, v2029, v2030, v2031, v2032, v2033, v2034, v2035, v2036, v2037, v2038, v2039, v2040, v2041, v2042, v2043, v2044, v2045, v2046, v2047, v2048, v2049, v2050, v2051, v2052, v2053, v2054, v2055, v2056, v2057, v2058, v2059, v2060, v2061, v2062, v2063, v2064, v2065, v2066, v2067, v2068, v2069, v2070, v2071, v2072, v2073, v2074, v2075, v2076, v2077, v2078, v2079, v2080, v2081, v2082, v2083, v2084, v2085, v2086, v2087, v2088, v2089, v2090, v2091, v2092, v2093, v2094, v2095, v2096, v2097, v2098, v2099, v2100, v2101, v2102, v2103, v2104, v2105, v2106, v2107, v2108, v2109, v2110, v2111, v2112, v2113, v2114, v2115, v2116, v2117, v2118, v2119, v2120, v2121, v2122, v2123, v2124, v2125, v2126, v2127, v2128, v2129, v2130, v2131, v2132, v2133, v2134, v2135, v2136, v2137, v2138, v2139, v2140, v2141, v2142, v2143, v2144, v2145, v2146, v2147, v2148, v2149, v2150, v2151, v2152, v2153, v2154, v2155, v2156, v2157, v2158, v2159, v2160, v2161, v2162, v2163, v2164, v2165, v2166, v2167, v2168, v2169, v2170, v2171, v2172, v2173, v2174, v2175, v2176, v2177, v2178, v2179, v2180, v2181, v2182, v2183, v2184, v2185, v2186, v2187, v2188, v2189, v2190, v2191, v2192, v2193, v2194, v2195, v2196, v2197, v2198, v2199, v2200, v2201, v2202, v2203, v2204, v2205, v2206, v2207, v2208, v2209, v2210, v2211, v2212, v2213, v2214, v2215, v2216, v2217, v2218, v2219, v2220, v2221, v2222, v2223, v2224, v2225, v2226, v2227, v2228, v2229, v2230, v2231, v2232, v2233, v2234, v2235, v2236, v2237, v2238, v2239, v2240, v2241, v2242, v2243, v2244, v2245, v2246, v2247, v2248, v2249, v2250, v2251, v2252, v2253, v2254, v2255, v2256, v2257, v2258, v2259, v2260, v2261, v2262, v2263, v2264, v2265, v2266, v2267, v2268, v2269, v2270, v2271, v2272, v2273, v2274, v2275, v2276, v2277, v2278, v2279, v2280, v2281, v2282, v2283, v2284, v2285, v2286, v2287, v2288, v2289, v2290, v2291, v2292, v2293, v2294, v2295, v2296, v2297, v2298, v2299, v2300, v2301, v2302, v2303, v2304, v2305, v2306, v2307, v2308, v2309, v2310, v2311, v2312, v2313, v2314, v2315, v2316, v2317, v2318, v2319, v2320, v2321, v2322, v2323, v2324, v2325, v2326, v2327, v2328, v2329, v2330, v2331, v2332, v2333, v2334, v2335, v2336, v2337, v2338, v2339, v2340, v2341, v2342, v2343, v2344, v2345, v2346, v2347, v2348, v2349, v2350, v2351, v2352, v2353, v2354, v2355, v2356, v2357, v2358, v2359, v2360, v2361, v2362, v2363, v2364, v2365, v2366, v2367, v2368, v2369, v2370, v2371, v2372, v2373, v2374, v2375, v2376, v2377, v2378, v2379, v2380, v2381, v2382, v2383, v2384, v2385, v2386, v2387, v2388, v2389, v2390, v2391, v2392, v2393, v2394, v2395, v2396, v2397, v2398, v2399, v2400, v2401, v2402, v2403, v2404, v2405, v2406, v2407, v2408, v2409, v2410, v2411, v2412, v2413, v2414, v2415, v2416, v2417, v2418, v2419, v2420, v2421, v2422, v2423, v2424, v2425, v2426, v2427, v2428, v2429, v2430, v2431, v2432, v2433, v2434, v2435, v2436, v2437, v2438, v2439, v2440, v2441, v2442, v2443, v2444, v2445, v2446, v2447, v2448, v2449, v2450, v2451, v2452, v2453, v2454, v2455, v2456, v2457, v2458, v2459, v2460, v2461, v2462, v2463, v2464, v2465, v2466, v2467, v2468, v2469, v2470, v2471, v2472, v2473, v2474, v2475, v2476, v2477, v2478, v2479, v2480, v2481, v2482, v2483, v2484, v2485, v2486, v2487, v2488, v2489, v2490, v2491, v2492, v2493, v2494, v2495, v2496, v2497, v2498, v2499, v2500, v2501, v2502, v2503, v2504, v2505, v2506, v2507, v2508, v2509, v2510, v2511, v2512, v2513, v2514, v2515, v2516, v2517, v2518, v2519, v2520, v2521, v2522, v2523, v2524, v2525, v2526, v2527, v2528, v2529, v2530, v2531, v2532, v2533, v2534, v2535, v2536, v2537, v2538, v2539, v2540, v2541, v2542, v2543, v2544, v2545, v2546, v2547, v2548, v2549, v2550, v2551, v2552, v2553, v2554, v2555, v2556, v2557, v2558, v2559, v2560, v2561, v2562, v2563, v2564, v2565, v2566, v2567, v2568, v2569, v2570, v2571, v2572, v2573, v2574, v2575, v2576, v2577, v2578, v2579, v2580, v2581, v2582, v2583, v2584, v2585, v2586, v2587, v2588, v2589, v2590, v2591, v2592, v2593, v2594, v2595, v2596, v2597, v2598, v2599, v2600, v2601, v2602, v2603, v2604, v2605, v2606, v2607, v2608, v2609, v2610, v2611, v2612, v2613, v2614, v2615, v2616, v2617, v2618, v2619, v2620, v2621, v2622, v2623, v2624, v2625, v2626, v2627, v2628, v2629, v2630, v2631, v2632, v2633, v2634, v2635, v2636, v2637, v2638, v2639, v2640, v2641, v2642, v2643, v2644, v2645, v2646, v2647, v2648, v2649, v2650, v2651, v2652, v2653, v2654, v2655, v2656, v2657, v2658, v2659, v2660, v2661, v2662, v2663, v2664, v2665, v2666, v2667, v2668, v2669, v2670, v2671, v2672, v2673, v2674, v2675, v2676, v2677, v2678, v2679, v2680, v2681, v2682, v2683, v2684, v2685, v2686, v2687, v2688, v2689, v2690, v2691, v2692, v2693, v2694, v2695, v2696, v2697, v2698, v2699, v2700, v2701, v2702, v2703, v2704, v2705, v2706, v2707, v2708, v2709, v2710, v2711, v2712, v2713, v2714, v2715, v2716, v2717, v2718, v2719, v2720, v2721, v2722, v2723, v2724, v2725, v2726, v2727, v2728, v2729, v2730, v2731, v2732, v2733, v2734, v2735, v2736, v2737, v2738, v2739, v2740, v2741, v2742, v2743, v2744, v2745, v2746, v2747, v2748, v2749, v2750, v2751, v2752, v2753, v2754, v2755, v2756, v2757, v2758, v2759, v2760, v2761, v2762, v2763, v2764, v2765, v2766, v2767, v2768, v2769, v2770, v2771, v2772, v2773, v2774, v2775, v2776, v2777, v2778, v2779, v2780, v2781, v2782, v2783, v2784, v2785, v2786, v2787, v2788, v2789, v2790, v2791, v2792, v2793, v2794, v2795, v2796, v2797, v2798, v2799, v2800, v2801, v2802, v2803, v2804, v2805, v2806, v2807, v2808, v2809, v2810, v2811, v2812, v2813, v2814, v2815, v2816, v2817, v2818, v2819, v2820, v2821, v2822, v2823, v2824, v2825, v2826, v2827, v2828, v2829, v2830, v2831, v2832, v2833, v2834, v2835, v2836, v2837, v2838, v2839, v2840, v2841, v2842, v2843, v2844, v2845, v2846, v2847, v2848, v2849, v2850, v2851, v2852, v2853, v2854, v2855, v2856, v2857, v2858, v2859, v2860, v2861, v2862, v2863, v2864, v2865, v2866, v2867, v2868, v2869, v2870, v2871, v2872, v2873, v2874, v2875, v2876, v2877, v2878, v2879, v2880, v2881, v2882, v2883, v2884, v2885, v2886, v2887, v2888, v2889, v2890, v2891, v2892, v2893, v2894, v2895, v2896, v2897, v2898, v2899, v2900, v2901, v2902, v2903, v2904, v2905, v2906, v2907, v2908, v2909, v2910, v2911, v2912, v2913, v2914, v2915, v2916, v2917, v2918, v2919, v2920, v2921, v2922, v2923, v2924, v2925, v2926, v2927, v2928, v2929, v2930, v2931, v2932, v2933, v2934, v2935, v2936, v2937, v2938, v2939, v2940, v2941, v2942, v2943, v2944, v2945, v2946, v2947, v2948, v2949, v2950, v2951, v2952, v2953, v2954, v2955, v2956, v2957, v2958, v2959, v2960, v2961, v2962, v2963, v2964, v2965, v2966, v2967, v2968, v2969, v2970, v2971, v2972, v2973, v2974, v2975, v2976, v2977, v2978, v2979, v2980, v2981, v2982, v2983, v2984, v2985, v2986, v2987, v2988, v2989, v2990, v2991, v2992, v2993, v2994, v2995, v2996, v2997, v2998, v2999, v3000, v3001, v3002, v3003, v3004, v3005, v3006, v3007, v3008, v3009, v3010, v3011, v3012, v3013, v3014, v3015, v3016, v3017, v3018, v3019, v3020, v3021, v3022, v3023, v3024, v3025, v3026, v3027, v3028, v3029, v3030, v3031, v3032, v3033, v3034, v3035, v3036, v3037, v3038, v3039, v3040, v3041, v3042, v3043, v3044, v3045, v3046, v3047, v3048, v3049, v3050, v3051, v3052, v3053, v3054, v3055, v3056, v3057, v3058, v3059, v3060, v3061, v3062, v3063, v3064, v3065, v3066, v3067, v3068, v3069, v3070, v3071, v3072, v3073, v3074, v3075, v3076, v3077, v3078, v3079, v3080, v3081, v3082, v3083, v3084, v3085, v3086, v3087, v3088, v3089, v3090, v3091, v3092, v3093, v3094, v3095, v3096, v3097, v3098, v3099, v3100, v3101, v3102, v3103, v3104, v3105, v3106, v3107, v3108, v3109, v3110, v3111, v3112, v3113, v3114, v3115, v3116, v3117, v3118, v3119, v3120, v3121, v3122, v3123, v3124, v3125, v3126, v3127, v3128, v3129, v3130, v3131, v3132, v3133, v3134, v3135, v3136, v3137, v3138, v3139, v3140, v3141, v3142, v3143, v3144, v3145, v3146, v3147, v3148, v3149, v3150, v3151, v3152, v3153, v3154, v3155, v3156, v3157, v3158, v3159, v3160, v3161, v3162, v3163, v3164, v3165, v3166, v3167, v3168, v3169, v3170, v3171, v3172, v3173, v3174, v3175, v3176, v3177, v3178, v3179, v3180, v3181, v3182, v3183, v3184, v3185, v3186, v3187, v3188, v3189, v3190, v3191, v3192, v3193, v3194, v3195, v3196, v3197, v3198, v3199, v3200, v3201, v3202, v3203, v3204, v3205, v3206, v3207, v3208, v3209, v3210, v3211, v3212, v3213, v3214, v3215, v3216, v3217, v3218, v3219, v3220, v3221, v3222, v3223, v3224, v3225, v3226, v3227, v3228, v3229, v3230, v3231, v3232, v3233, v3234, v3235, v3236, v3237, v3238, v3239, v3240, v3241, v3242, v3243, v3244, v3245, v3246, v3247, v3248, v3249, v3250, v3251, v3252, v3253, v3254, v3255, v3256, v3257, v3258, v3259, v3260, v3261, v3262, v3263, v3264, v3265, v3266, v3267, v3268, v3269, v3270, v3271, v3272, v3273, v3274, v3275, v3276, v3277, v3278, v3279, v3280, v3281, v3282, v3283, v3284, v3285, v3286, v3287, v3288, v3289, v3290, v3291, v3292, v3293, v3294, v3295, v3296, v3297, v3298, v3299, v3300, v3301, v3302, v3303, v3304, v3305, v3306, v3307, v3308, v3309, v3310, v3311, v3312, v3313, v3314, v3315, v3316, v3317, v3318, v3319, v3320, v3321, v3322, v3323, v3324, v3325, v3326, v3327, v3328, v3329, v3330, v3331, v3332, v3333, v3334, v3335, v3336, v3337, v3338, v3339, v3340, v3341, v3342, v3343, v3344, v3345, v3346, v3347, v3348, v3349, v3350, v3351, v3352, v3353, v3354, v3355, v3356, v3357, v3358, v3359, v3360, v3361, v3362, v3363, v3364, v3365, v3366, v3367, v3368, v3369, v3370, v3371, v3372, v3373, v3374, v3375, v3376, v3377, v3378, v3379, v3380, v3381, v3382, v3383, v3384, v3385, v3386, v3387, v3388, v3389, v3390, v3391, v3392, v3393, v3394, v3395, v3396, v3397, v3398, v3399, v3400, v3401, v3402, v3403, v3404, v3405, v3406, v3407, v3408, v3409, v3410, v3411, v3412, v3413, v3414, v3415, v3416, v3417, v3418, v3419, v3420, v3421, v3422, v3423, v3424, v3425, v3426, v3427, v3428, v3429, v3430, v3431, v3432, v3433, v3434, v3435, v3436, v3437, v3438, v3439, v3440, v3441, v3442, v3443, v3444, v3445, v3446, v3447, v3448, v3449, v3450, v3451, v3452, v3453, v3454, v3455, v3456, v3457, v3458, v3459, v3460, v3461, v3462, v3463, v3464, v3465, v3466, v3467, v3468, v3469, v3470, v3471, v3472, v3473, v3474, v3475, v3476, v3477, v3478, v3479, v3480, v3481, v3482, v3483, v3484, v3485, v3486, v3487, v3488, v3489, v3490, v3491, v3492, v3493, v3494, v3495, v3496, v3497, v3498, v3499, v3500, v3501, v3502, v3503, v3504, v3505, v3506, v3507, v3508, v3509, v3510, v3511, v3512, v3513, v3514, v3515, v3516, v3517, v3518, v3519, v3520, v3521, v3522, v3523, v3524, v3525, v3526, v3527, v3528, v3529, v3530, v3531, v3532, v3533, v3534, v3535, v3536, v3537, v3538, v3539, v3540, v3541, v3542, v3543, v3544, v3545, v3546, v3547, v3548, v3549, v3550, v3551, v3552, v3553, v3554, v3555, v3556, v3557, v3558, v3559, v3560, v3561, v3562, v3563, v3564, v3565, v3566, v3567, v3568, v3569, v3570, v3571, v3572, v3573, v3574, v3575, v3576, v3577, v3578, v3579, v3580, v3581, v3582, v3583, v3584, v3585, v3586, v3587, v3588, v3589, v3590, v3591, v3592, v3593, v3594, v3595, v3596, v3597, v3598, v3599, v3600, v3601, v3602, v3603, v3604, v3605, v3606, v3607, v3608, v3609, v3610, v3611, v3612, v3613, v3614, v3615, v3616, v3617, v3618, v3619, v3620, v3621, v3622, v3623, v3624, v3625, v3626, v3627, v3628, v3629, v3630, v3631, v3632, v3633, v3634, v3635, v3636, v3637, v3638, v3639, v3640, v3641, v3642, v3643, v3644, v3645, v3646, v3647, v3648, v3649, v3650, v3651, v3652, v3653, v3654, v3655, v3656, v3657, v3658, v3659, v3660, v3661, v3662, v3663, v3664, v3665, v3666, v3667, v3668, v3669, v3670, v3671, v3672, v3673, v3674, v3675, v3676, v3677, v3678, v3679, v3680, v3681, v3682, v3683, v3684, v3685, v3686, v3687, v3688, v3689, v3690, v3691, v3692, v3693, v3694, v3695, v3696, v3697, v3698, v3699, v3700, v3701, v3702, v3703, v3704, v3705, v3706, v3707, v3708, v3709, v3710, v3711, v3712, v3713, v3714, v3715, v3716, v3717, v3718, v3719, v3720, v3721, v3722, v3723, v3724, v3725, v3726, v3727, v3728, v3729, v3730, v3731, v3732, v3733, v3734, v3735, v3736, v3737, v3738, v3739, v3740, v3741, v3742, v3743, v3744, v3745, v3746, v3747, v3748, v3749, v3750, v3751, v3752, v3753, v3754, v3755, v3756, v3757, v3758, v3759, v3760, v3761, v3762, v3763, v3764, v3765, v3766, v3767, v3768, v3769, v3770, v3771, v3772, v3773, v3774, v3775, v3776, v3777, v3778, v3779, v3780, v3781, v3782, v3783, v3784, v3785, v3786, v3787, v3788, v3789, v3790, v3791, v3792, v3793, v3794, v3795, v3796, v3797, v3798, v3799, v3800, v3801, v3802, v3803, v3804, v3805, v3806, v3807, v3808, v3809, v3810, v3811, v3812, v3813, v3814, v3815, v3816, v3817, v3818, v3819, v3820, v3821, v3822, v3823, v3824, v3825, v3826, v3827, v3828, v3829, v3830, v3831, v3832, v3833, v3834, v3835, v3836, v3837, v3838, v3839, v3840, v3841, v3842, v3843, v3844, v3845, v3846, v3847, v3848, v3849, v3850, v3851, v3852, v3853, v3854, v3855, v3856, v3857, v3858, v3859, v3860, v3861, v3862, v3863, v3864, v3865, v3866, v3867, v3868, v3869, v3870, v3871, v3872, v3873, v3874, v3875, v3876, v3877, v3878, v3879, v3880, v3881, v3882, v3883, v3884, v3885, v3886, v3887, v3888, v3889, v3890, v3891, v3892, v3893, v3894, v3895, v3896, v3897, v3898, v3899, v3900, v3901, v3902, v3903, v3904, v3905, v3906, v3907, v3908, v3909, v3910, v3911, v3912, v3913, v3914, v3915, v3916, v3917, v3918, v3919, v3920, v3921, v3922, v3923, v3924, v3925, v3926, v3927, v3928, v3929, v3930, v3931, v3932, v3933, v3934, v3935, v3936, v3937, v3938, v3939, v3940, v3941, v3942, v3943, v3944, v3945, v3946, v3947, v3948, v3949, v3950, v3951, v3952, v3953, v3954, v3955, v3956, v3957, v3958, v3959, v3960, v3961, v3962, v3963, v3964, v3965, v3966, v3967, v3968, v3969, v3970, v3971, v3972, v3973, v3974, v3975, v3976, v3977, v3978, v3979, v3980, v3981, v3982, v3983, v3984, v3985, v3986, v3987, v3988, v3989, v3990, v3991, v3992, v3993, v3994, v3995, v3996, v3997, v3998, v3999, v4000, v4001, v4002, v4003, v4004, v4005, v4006, v4007, v4008, v4009, v4010, v4011, v4012, v4013, v4014, v4015, v4016, v4017, v4018, v4019, v4020, v4021, v4022, v4023, v4024, v4025, v4026, v4027, v4028, v4029, 
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325;
assign w0 = pi00 & pi32;
assign w1 = pi64 & w0;
assign v0 = ~(pi64 | w0);
assign w2 = v0;
assign v1 = ~(w1 | w2);
assign w3 = v1;
assign w4 = pi00 & pi33;
assign w5 = pi01 & pi32;
assign w6 = pi65 & w5;
assign v2 = ~(pi65 | w5);
assign w7 = v2;
assign v3 = ~(w6 | w7);
assign w8 = v3;
assign w9 = w4 & w8;
assign v4 = ~(w4 | w8);
assign w10 = v4;
assign v5 = ~(w9 | w10);
assign w11 = v5;
assign w12 = w1 & w11;
assign v6 = ~(w1 | w11);
assign w13 = v6;
assign v7 = ~(w12 | w13);
assign w14 = v7;
assign w15 = (~w9 & ~w11) | (~w9 & w8577) | (~w11 & w8577);
assign w16 = pi01 & pi33;
assign w17 = pi00 & pi34;
assign v8 = ~(w16 | w17);
assign w18 = v8;
assign w19 = pi01 & pi34;
assign w20 = w4 & w19;
assign v9 = ~(w18 | w20);
assign w21 = v9;
assign w22 = pi02 & pi32;
assign w23 = pi66 & w22;
assign v10 = ~(pi66 | w22);
assign w24 = v10;
assign v11 = ~(w23 | w24);
assign w25 = v11;
assign w26 = w21 & w25;
assign v12 = ~(w21 | w25);
assign w27 = v12;
assign v13 = ~(w26 | w27);
assign w28 = v13;
assign w29 = w6 & w28;
assign v14 = ~(w6 | w28);
assign w30 = v14;
assign v15 = ~(w29 | w30);
assign w31 = v15;
assign w32 = ~w15 & w31;
assign w33 = w15 & ~w31;
assign v16 = ~(w32 | w33);
assign w34 = v16;
assign w35 = (~w29 & ~w31) | (~w29 & w8578) | (~w31 & w8578);
assign v17 = ~(w20 | w26);
assign w36 = v17;
assign w37 = pi00 & pi35;
assign w38 = w23 & w37;
assign v18 = ~(w23 | w37);
assign w39 = v18;
assign v19 = ~(w38 | w39);
assign w40 = v19;
assign w41 = pi03 & pi32;
assign w42 = pi67 & w41;
assign v20 = ~(pi67 | w41);
assign w43 = v20;
assign v21 = ~(w42 | w43);
assign w44 = v21;
assign w45 = pi02 & pi33;
assign v22 = ~(w19 | w45);
assign w46 = v22;
assign w47 = pi02 & pi34;
assign w48 = w16 & w47;
assign v23 = ~(w46 | w48);
assign w49 = v23;
assign w50 = w44 & ~w49;
assign w51 = ~w44 & w49;
assign v24 = ~(w50 | w51);
assign w52 = v24;
assign w53 = w40 & ~w52;
assign w54 = ~w40 & w52;
assign v25 = ~(w53 | w54);
assign w55 = v25;
assign w56 = ~w36 & w55;
assign w57 = w36 & ~w55;
assign v26 = ~(w56 | w57);
assign w58 = v26;
assign w59 = w35 & ~w58;
assign w60 = ~w35 & w58;
assign v27 = ~(w59 | w60);
assign w61 = v27;
assign v28 = ~(w38 | w53);
assign w62 = v28;
assign w63 = pi00 & pi36;
assign w64 = w44 & ~w46;
assign w65 = w42 & ~w48;
assign w66 = w43 & w48;
assign v29 = ~(w65 | w66);
assign w67 = v29;
assign w68 = ~w64 & w67;
assign w69 = w63 & ~w68;
assign w70 = ~w63 & w68;
assign v30 = ~(w69 | w70);
assign w71 = v30;
assign w72 = pi01 & pi35;
assign v31 = ~(w47 | w72);
assign w73 = v31;
assign w74 = pi02 & pi35;
assign w75 = w19 & w74;
assign v32 = ~(w73 | w75);
assign w76 = v32;
assign w77 = pi03 & pi33;
assign w78 = pi04 & pi32;
assign w79 = pi68 & w78;
assign v33 = ~(pi68 | w78);
assign w80 = v33;
assign v34 = ~(w79 | w80);
assign w81 = v34;
assign w82 = w77 & ~w81;
assign w83 = ~w77 & w81;
assign v35 = ~(w82 | w83);
assign w84 = v35;
assign w85 = w76 & ~w84;
assign w86 = ~w76 & w84;
assign v36 = ~(w85 | w86);
assign w87 = v36;
assign w88 = w71 & w87;
assign v37 = ~(w71 | w87);
assign w89 = v37;
assign v38 = ~(w88 | w89);
assign w90 = v38;
assign w91 = w62 & ~w90;
assign w92 = ~w62 & w90;
assign v39 = ~(w91 | w92);
assign w93 = v39;
assign w94 = (~w56 & ~w58) | (~w56 & w8579) | (~w58 & w8579);
assign w95 = ~w93 & w94;
assign w96 = w93 & ~w94;
assign v40 = ~(w95 | w96);
assign w97 = v40;
assign v41 = ~(w69 | w88);
assign w98 = v41;
assign w99 = w42 & w48;
assign w100 = pi05 & pi32;
assign w101 = pi69 & w100;
assign v42 = ~(pi69 | w100);
assign w102 = v42;
assign v43 = ~(w101 | w102);
assign w103 = v43;
assign w104 = pi04 & pi33;
assign w105 = pi00 & pi37;
assign v44 = ~(w104 | w105);
assign w106 = v44;
assign w107 = ~w103 & w106;
assign w108 = ~w102 & w104;
assign v45 = ~(w101 | w105);
assign w109 = v45;
assign w110 = w108 & w109;
assign v46 = ~(w107 | w110);
assign w111 = v46;
assign w112 = ~w104 & w105;
assign w113 = w103 & ~w112;
assign w114 = pi04 & pi37;
assign w115 = w4 & w114;
assign v47 = ~(w103 | w115);
assign w116 = v47;
assign v48 = ~(w113 | w116);
assign w117 = v48;
assign w118 = w111 & ~w117;
assign w119 = pi01 & pi36;
assign w120 = pi03 & pi34;
assign v49 = ~(w74 | w120);
assign w121 = v49;
assign w122 = pi03 & pi35;
assign w123 = w47 & w122;
assign v50 = ~(w121 | w123);
assign w124 = v50;
assign w125 = w119 & ~w124;
assign w126 = ~w119 & w124;
assign v51 = ~(w125 | w126);
assign w127 = v51;
assign w128 = ~w118 & w127;
assign w129 = w118 & ~w127;
assign v52 = ~(w128 | w129);
assign w130 = v52;
assign w131 = w99 & w130;
assign v53 = ~(w99 | w130);
assign w132 = v53;
assign v54 = ~(w131 | w132);
assign w133 = v54;
assign v55 = ~(w75 | w85);
assign w134 = v55;
assign v56 = ~(w77 | w79);
assign w135 = v56;
assign v57 = ~(w80 | w135);
assign w136 = v57;
assign w137 = ~w134 & w136;
assign w138 = w134 & ~w136;
assign v58 = ~(w137 | w138);
assign w139 = v58;
assign w140 = w133 & w139;
assign v59 = ~(w133 | w139);
assign w141 = v59;
assign v60 = ~(w140 | w141);
assign w142 = v60;
assign w143 = w98 & ~w142;
assign w144 = ~w98 & w142;
assign v61 = ~(w143 | w144);
assign w145 = v61;
assign w146 = ~w92 & w94;
assign v62 = ~(w91 | w146);
assign w147 = v62;
assign w148 = w145 & ~w147;
assign w149 = ~w145 & w147;
assign v63 = ~(w148 | w149);
assign w150 = v63;
assign w151 = w111 & ~w127;
assign v64 = ~(w117 | w151);
assign w152 = v64;
assign v65 = ~(w101 | w108);
assign w153 = v65;
assign w154 = w119 & ~w121;
assign v66 = ~(w123 | w154);
assign w155 = v66;
assign v67 = ~(w153 | w155);
assign w156 = v67;
assign w157 = w153 & w155;
assign v68 = ~(w156 | w157);
assign w158 = v68;
assign w159 = ~w152 & w158;
assign w160 = w152 & ~w158;
assign v69 = ~(w159 | w160);
assign w161 = v69;
assign w162 = w137 & w161;
assign v70 = ~(w137 | w161);
assign w163 = v70;
assign v71 = ~(w162 | w163);
assign w164 = v71;
assign w165 = pi06 & pi32;
assign w166 = pi70 & w165;
assign v72 = ~(pi70 | w165);
assign w167 = v72;
assign v73 = ~(w166 | w167);
assign w168 = v73;
assign w169 = pi05 & pi33;
assign w170 = pi04 & pi34;
assign v74 = ~(w169 | w170);
assign w171 = v74;
assign w172 = pi05 & pi34;
assign w173 = w104 & w172;
assign v75 = ~(w171 | w173);
assign w174 = v75;
assign w175 = w122 & ~w174;
assign w176 = ~w122 & w174;
assign v76 = ~(w175 | w176);
assign w177 = v76;
assign w178 = ~w168 & w177;
assign w179 = w168 & ~w177;
assign v77 = ~(w178 | w179);
assign w180 = v77;
assign w181 = pi00 & pi38;
assign w182 = pi01 & pi37;
assign w183 = pi02 & pi36;
assign v78 = ~(w182 | w183);
assign w184 = v78;
assign w185 = pi02 & pi37;
assign w186 = w119 & w185;
assign v79 = ~(w184 | w186);
assign w187 = v79;
assign w188 = w181 & ~w187;
assign w189 = ~w181 & w187;
assign v80 = ~(w188 | w189);
assign w190 = v80;
assign w191 = w180 & w190;
assign v81 = ~(w180 | w190);
assign w192 = v81;
assign v82 = ~(w191 | w192);
assign w193 = v82;
assign w194 = w164 & ~w193;
assign w195 = ~w164 & w193;
assign v83 = ~(w194 | w195);
assign w196 = v83;
assign v84 = ~(w131 | w140);
assign w197 = v84;
assign w198 = ~w196 & w197;
assign w199 = w196 & ~w197;
assign v85 = ~(w198 | w199);
assign w200 = v85;
assign v86 = ~(w144 | w147);
assign w201 = v86;
assign v87 = ~(w143 | w201);
assign w202 = v87;
assign w203 = ~w200 & w202;
assign w204 = w200 & ~w202;
assign v88 = ~(w203 | w204);
assign w205 = v88;
assign v89 = ~(w198 | w204);
assign w206 = v89;
assign w207 = (~w162 & ~w164) | (~w162 & w8665) | (~w164 & w8665);
assign w208 = w181 & ~w184;
assign v90 = ~(w186 | w208);
assign w209 = v90;
assign w210 = w122 & ~w171;
assign v91 = ~(w173 | w210);
assign w211 = v91;
assign v92 = ~(w209 | w211);
assign w212 = v92;
assign w213 = w209 & w211;
assign v93 = ~(w212 | w213);
assign w214 = v93;
assign w215 = (~w178 & ~w180) | (~w178 & w8666) | (~w180 & w8666);
assign w216 = w214 & w215;
assign v94 = ~(w214 | w215);
assign w217 = v94;
assign v95 = ~(w216 | w217);
assign w218 = v95;
assign w219 = (~w156 & w152) | (~w156 & w8667) | (w152 & w8667);
assign w220 = pi07 & pi32;
assign w221 = pi71 & w220;
assign v96 = ~(pi71 | w220);
assign w222 = v96;
assign v97 = ~(w221 | w222);
assign w223 = v97;
assign w224 = pi06 & pi33;
assign v98 = ~(w172 | w224);
assign w225 = v98;
assign w226 = pi06 & pi34;
assign w227 = w169 & w226;
assign v99 = ~(w225 | w227);
assign w228 = v99;
assign w229 = w223 & ~w228;
assign w230 = ~w223 & w228;
assign v100 = ~(w229 | w230);
assign w231 = v100;
assign w232 = pi00 & pi39;
assign w233 = pi01 & pi38;
assign v101 = ~(w232 | w233);
assign w234 = v101;
assign w235 = pi01 & pi39;
assign w236 = w181 & w235;
assign v102 = ~(w234 | w236);
assign w237 = v102;
assign w238 = w166 & ~w237;
assign w239 = ~w166 & w237;
assign v103 = ~(w238 | w239);
assign w240 = v103;
assign w241 = w231 & w240;
assign v104 = ~(w231 | w240);
assign w242 = v104;
assign v105 = ~(w241 | w242);
assign w243 = v105;
assign w244 = pi03 & pi36;
assign w245 = pi04 & pi35;
assign v106 = ~(w244 | w245);
assign w246 = v106;
assign w247 = pi04 & pi36;
assign w248 = w122 & w247;
assign v107 = ~(w246 | w248);
assign w249 = v107;
assign w250 = w185 & ~w249;
assign w251 = ~w185 & w249;
assign v108 = ~(w250 | w251);
assign w252 = v108;
assign w253 = w243 & ~w252;
assign w254 = ~w243 & w252;
assign v109 = ~(w253 | w254);
assign w255 = v109;
assign w256 = ~w219 & w255;
assign w257 = w219 & ~w255;
assign v110 = ~(w256 | w257);
assign w258 = v110;
assign w259 = w218 & ~w258;
assign w260 = ~w218 & w258;
assign v111 = ~(w259 | w260);
assign w261 = v111;
assign v112 = ~(w207 | w261);
assign w262 = v112;
assign w263 = w207 & w261;
assign v113 = ~(w262 | w263);
assign w264 = v113;
assign w265 = w206 & w264;
assign v114 = ~(w206 | w264);
assign w266 = v114;
assign v115 = ~(w265 | w266);
assign w267 = v115;
assign v116 = ~(w198 | w263);
assign w268 = v116;
assign w269 = (~w262 & w204) | (~w262 & w8580) | (w204 & w8580);
assign v117 = ~(w212 | w216);
assign w270 = v117;
assign w271 = pi05 & pi35;
assign v118 = ~(w226 | w271);
assign w272 = v118;
assign w273 = pi06 & pi35;
assign w274 = w172 & w273;
assign v119 = ~(w272 | w274);
assign w275 = v119;
assign w276 = pi07 & pi33;
assign w277 = pi08 & pi32;
assign w278 = pi72 & w277;
assign v120 = ~(pi72 | w277);
assign w279 = v120;
assign v121 = ~(w278 | w279);
assign w280 = v121;
assign w281 = w276 & w280;
assign v122 = ~(w276 | w280);
assign w282 = v122;
assign v123 = ~(w281 | w282);
assign w283 = v123;
assign w284 = w275 & w283;
assign v124 = ~(w275 | w283);
assign w285 = v124;
assign v125 = ~(w284 | w285);
assign w286 = v125;
assign w287 = pi02 & pi38;
assign w288 = pi03 & pi37;
assign v126 = ~(w247 | w288);
assign w289 = v126;
assign w290 = w114 & w244;
assign v127 = ~(w289 | w290);
assign w291 = v127;
assign w292 = w287 & ~w291;
assign w293 = ~w287 & w291;
assign v128 = ~(w292 | w293);
assign w294 = v128;
assign w295 = ~w286 & w294;
assign w296 = w286 & ~w294;
assign v129 = ~(w295 | w296);
assign w297 = v129;
assign w298 = pi00 & pi40;
assign v130 = ~(w235 | w298);
assign w299 = v130;
assign w300 = pi01 & pi40;
assign w301 = w232 & w300;
assign v131 = ~(w299 | w301);
assign w302 = v131;
assign w303 = w221 & w227;
assign v132 = ~(w221 | w227);
assign w304 = v132;
assign v133 = ~(w303 | w304);
assign w305 = v133;
assign w306 = w223 & ~w225;
assign v134 = ~(w305 | w306);
assign w307 = v134;
assign w308 = w302 & ~w307;
assign w309 = ~w302 & w307;
assign v135 = ~(w308 | w309);
assign w310 = v135;
assign w311 = w297 & ~w310;
assign w312 = ~w297 & w310;
assign v136 = ~(w311 | w312);
assign w313 = v136;
assign w314 = (~w242 & ~w243) | (~w242 & w8668) | (~w243 & w8668);
assign w315 = w166 & ~w234;
assign v137 = ~(w236 | w315);
assign w316 = v137;
assign w317 = w185 & ~w246;
assign v138 = ~(w248 | w317);
assign w318 = v138;
assign v139 = ~(w316 | w318);
assign w319 = v139;
assign w320 = w316 & w318;
assign v140 = ~(w319 | w320);
assign w321 = v140;
assign w322 = ~w314 & w321;
assign w323 = w314 & ~w321;
assign v141 = ~(w322 | w323);
assign w324 = v141;
assign w325 = w313 & ~w324;
assign w326 = ~w313 & w324;
assign v142 = ~(w325 | w326);
assign w327 = v142;
assign w328 = w270 & ~w327;
assign w329 = ~w270 & w327;
assign v143 = ~(w328 | w329);
assign w330 = v143;
assign v144 = ~(w257 | w260);
assign w331 = v144;
assign w332 = w330 & w331;
assign v145 = ~(w330 | w331);
assign w333 = v145;
assign v146 = ~(w332 | w333);
assign w334 = v146;
assign w335 = ~w269 & w334;
assign w336 = w269 & ~w334;
assign v147 = ~(w335 | w336);
assign w337 = v147;
assign w338 = pi00 & pi41;
assign w339 = w303 & w338;
assign v148 = ~(w303 | w338);
assign w340 = v148;
assign v149 = ~(w339 | w340);
assign w341 = v149;
assign v150 = ~(w278 | w281);
assign w342 = v150;
assign w343 = (~w274 & ~w283) | (~w274 & w8581) | (~w283 & w8581);
assign v151 = ~(w342 | w343);
assign w344 = v151;
assign w345 = w342 & w343;
assign v152 = ~(w344 | w345);
assign w346 = v152;
assign w347 = w341 & w346;
assign v153 = ~(w341 | w346);
assign w348 = v153;
assign v154 = ~(w347 | w348);
assign w349 = v154;
assign w350 = pi03 & pi38;
assign w351 = pi02 & pi39;
assign v155 = ~(w350 | w351);
assign w352 = v155;
assign w353 = pi03 & pi39;
assign w354 = w287 & w353;
assign v156 = ~(w352 | w354);
assign w355 = v156;
assign w356 = w300 & ~w355;
assign w357 = ~w300 & w355;
assign v157 = ~(w356 | w357);
assign w358 = v157;
assign w359 = pi08 & pi33;
assign w360 = pi09 & pi32;
assign w361 = pi73 & w360;
assign v158 = ~(pi73 | w360);
assign w362 = v158;
assign v159 = ~(w361 | w362);
assign w363 = v159;
assign w364 = w359 & w363;
assign v160 = ~(w359 | w363);
assign w365 = v160;
assign v161 = ~(w364 | w365);
assign w366 = v161;
assign v162 = ~(w114 | w366);
assign w367 = v162;
assign w368 = w114 & w366;
assign v163 = ~(w367 | w368);
assign w369 = v163;
assign w370 = pi05 & pi36;
assign w371 = pi07 & pi34;
assign v164 = ~(w273 | w371);
assign w372 = v164;
assign w373 = pi07 & pi35;
assign w374 = w226 & w373;
assign v165 = ~(w372 | w374);
assign w375 = v165;
assign w376 = w370 & ~w375;
assign w377 = ~w370 & w375;
assign v166 = ~(w376 | w377);
assign w378 = v166;
assign w379 = w369 & ~w378;
assign w380 = ~w369 & w378;
assign v167 = ~(w379 | w380);
assign w381 = v167;
assign w382 = ~w358 & w381;
assign w383 = w358 & ~w381;
assign v168 = ~(w382 | w383);
assign w384 = v168;
assign w385 = w349 & w384;
assign v169 = ~(w349 | w384);
assign w386 = v169;
assign v170 = ~(w385 | w386);
assign w387 = v170;
assign v171 = ~(w319 | w322);
assign w388 = v171;
assign w389 = (~w295 & ~w297) | (~w295 & w8582) | (~w297 & w8582);
assign v172 = ~(w301 | w308);
assign w390 = v172;
assign w391 = w287 & ~w289;
assign v173 = ~(w290 | w391);
assign w392 = v173;
assign v174 = ~(w390 | w392);
assign w393 = v174;
assign w394 = w390 & w392;
assign v175 = ~(w393 | w394);
assign w395 = v175;
assign w396 = w389 & w395;
assign v176 = ~(w389 | w395);
assign w397 = v176;
assign v177 = ~(w396 | w397);
assign w398 = v177;
assign w399 = ~w388 & w398;
assign w400 = w388 & ~w398;
assign v178 = ~(w399 | w400);
assign w401 = v178;
assign w402 = w387 & w401;
assign v179 = ~(w387 | w401);
assign w403 = v179;
assign v180 = ~(w402 | w403);
assign w404 = v180;
assign v181 = ~(w326 | w329);
assign w405 = v181;
assign w406 = ~w404 & w405;
assign w407 = w404 & ~w405;
assign v182 = ~(w406 | w407);
assign w408 = v182;
assign v183 = ~(w332 | w335);
assign w409 = v183;
assign w410 = w408 & w409;
assign v184 = ~(w408 | w409);
assign w411 = v184;
assign v185 = ~(w410 | w411);
assign w412 = v185;
assign v186 = ~(w332 | w407);
assign w413 = v186;
assign w414 = ~w335 & w413;
assign v187 = ~(w406 | w414);
assign w415 = v187;
assign v188 = ~(w399 | w402);
assign w416 = v188;
assign v189 = ~(w393 | w396);
assign w417 = v189;
assign w418 = (~w382 & ~w384) | (~w382 & w8583) | (~w384 & w8583);
assign w419 = (~w339 & ~w346) | (~w339 & w8669) | (~w346 & w8669);
assign w420 = w300 & ~w352;
assign v190 = ~(w354 | w420);
assign w421 = v190;
assign v191 = ~(w419 | w421);
assign w422 = v191;
assign w423 = w419 & w421;
assign v192 = ~(w422 | w423);
assign w424 = v192;
assign w425 = ~w418 & w424;
assign w426 = w418 & ~w424;
assign v193 = ~(w425 | w426);
assign w427 = v193;
assign w428 = ~w417 & w427;
assign w429 = w417 & ~w427;
assign v194 = ~(w428 | w429);
assign w430 = v194;
assign w431 = pi04 & pi38;
assign v195 = ~(w353 | w431);
assign w432 = v195;
assign w433 = pi04 & pi39;
assign w434 = w350 & w433;
assign v196 = ~(w432 | w434);
assign w435 = v196;
assign w436 = pi00 & pi42;
assign w437 = pi01 & pi41;
assign w438 = pi02 & pi40;
assign v197 = ~(w437 | w438);
assign w439 = v197;
assign w440 = pi02 & pi41;
assign w441 = w300 & w440;
assign v198 = ~(w439 | w441);
assign w442 = v198;
assign w443 = w436 & ~w442;
assign w444 = ~w436 & w442;
assign v199 = ~(w443 | w444);
assign w445 = v199;
assign w446 = w435 & ~w445;
assign w447 = ~w435 & w445;
assign v200 = ~(w446 | w447);
assign w448 = v200;
assign w449 = pi05 & pi37;
assign w450 = pi09 & pi33;
assign w451 = pi10 & pi32;
assign w452 = pi74 & w451;
assign v201 = ~(pi74 | w451);
assign w453 = v201;
assign v202 = ~(w452 | w453);
assign w454 = v202;
assign w455 = w450 & w454;
assign v203 = ~(w450 | w454);
assign w456 = v203;
assign v204 = ~(w455 | w456);
assign w457 = v204;
assign w458 = w449 & w457;
assign v205 = ~(w449 | w457);
assign w459 = v205;
assign v206 = ~(w458 | w459);
assign w460 = v206;
assign w461 = pi06 & pi36;
assign w462 = pi08 & pi34;
assign v207 = ~(w373 | w462);
assign w463 = v207;
assign w464 = pi08 & pi35;
assign w465 = w371 & w464;
assign v208 = ~(w463 | w465);
assign w466 = v208;
assign w467 = w461 & ~w466;
assign w468 = ~w461 & w466;
assign v209 = ~(w467 | w468);
assign w469 = v209;
assign w470 = w460 & ~w469;
assign w471 = ~w460 & w469;
assign v210 = ~(w470 | w471);
assign w472 = v210;
assign w473 = (~w361 & ~w363) | (~w361 & w8670) | (~w363 & w8670);
assign w474 = w370 & ~w372;
assign v211 = ~(w374 | w474);
assign w475 = v211;
assign v212 = ~(w473 | w475);
assign w476 = v212;
assign w477 = w473 & w475;
assign v213 = ~(w476 | w477);
assign w478 = v213;
assign w479 = ~w368 & w378;
assign v214 = ~(w367 | w479);
assign w480 = v214;
assign w481 = ~w479 & w8671;
assign w482 = (~w478 & w479) | (~w478 & w8672) | (w479 & w8672);
assign v215 = ~(w481 | w482);
assign w483 = v215;
assign w484 = w344 & w483;
assign v216 = ~(w344 | w483);
assign w485 = v216;
assign v217 = ~(w484 | w485);
assign w486 = v217;
assign w487 = w472 & w486;
assign v218 = ~(w472 | w486);
assign w488 = v218;
assign v219 = ~(w487 | w488);
assign w489 = v219;
assign w490 = w448 & w489;
assign v220 = ~(w448 | w489);
assign w491 = v220;
assign v221 = ~(w490 | w491);
assign w492 = v221;
assign w493 = w430 & w492;
assign v222 = ~(w430 | w492);
assign w494 = v222;
assign v223 = ~(w493 | w494);
assign w495 = v223;
assign w496 = ~w416 & w495;
assign w497 = w416 & ~w495;
assign v224 = ~(w496 | w497);
assign w498 = v224;
assign v225 = ~(w415 | w498);
assign w499 = v225;
assign w500 = w415 & w498;
assign v226 = ~(w499 | w500);
assign w501 = v226;
assign v227 = ~(w496 | w500);
assign w502 = v227;
assign v228 = ~(w428 | w493);
assign w503 = v228;
assign v229 = ~(w422 | w425);
assign w504 = v229;
assign w505 = pi06 & pi37;
assign w506 = pi10 & pi33;
assign w507 = pi11 & pi32;
assign w508 = pi75 & w507;
assign v230 = ~(pi75 | w507);
assign w509 = v230;
assign v231 = ~(w508 | w509);
assign w510 = v231;
assign w511 = w506 & w510;
assign v232 = ~(w506 | w510);
assign w512 = v232;
assign v233 = ~(w511 | w512);
assign w513 = v233;
assign w514 = w505 & w513;
assign v234 = ~(w505 | w513);
assign w515 = v234;
assign v235 = ~(w514 | w515);
assign w516 = v235;
assign w517 = pi07 & pi36;
assign w518 = pi09 & pi34;
assign v236 = ~(w464 | w518);
assign w519 = v236;
assign w520 = pi09 & pi35;
assign w521 = w462 & w520;
assign v237 = ~(w519 | w521);
assign w522 = v237;
assign w523 = w517 & ~w522;
assign w524 = ~w517 & w522;
assign v238 = ~(w523 | w524);
assign w525 = v238;
assign w526 = w516 & ~w525;
assign w527 = ~w516 & w525;
assign v239 = ~(w526 | w527);
assign w528 = v239;
assign w529 = (~w458 & ~w460) | (~w458 & w8673) | (~w460 & w8673);
assign w530 = (~w452 & ~w454) | (~w452 & w8674) | (~w454 & w8674);
assign w531 = w461 & ~w463;
assign v240 = ~(w465 | w531);
assign w532 = v240;
assign v241 = ~(w530 | w532);
assign w533 = v241;
assign w534 = w530 & w532;
assign v242 = ~(w533 | w534);
assign w535 = v242;
assign w536 = ~w434 & w535;
assign w537 = w434 & ~w535;
assign v243 = ~(w536 | w537);
assign w538 = v243;
assign w539 = w529 & ~w538;
assign w540 = ~w529 & w538;
assign v244 = ~(w539 | w540);
assign w541 = v244;
assign w542 = w528 & ~w541;
assign w543 = ~w528 & w541;
assign v245 = ~(w542 | w543);
assign w544 = v245;
assign w545 = pi00 & pi43;
assign w546 = pi01 & pi42;
assign v246 = ~(w545 | w546);
assign w547 = v246;
assign w548 = pi01 & pi43;
assign w549 = w436 & w548;
assign v247 = ~(w547 | w549);
assign w550 = v247;
assign w551 = (w480 & w8675) | (w480 & w8676) | (w8675 & w8676);
assign w552 = ~w550 & w9294;
assign v248 = ~(w551 | w552);
assign w553 = v248;
assign w554 = pi03 & pi40;
assign w555 = pi05 & pi38;
assign v249 = ~(w433 | w555);
assign w556 = v249;
assign w557 = pi05 & pi39;
assign w558 = w431 & w557;
assign v250 = ~(w556 | w558);
assign w559 = v250;
assign w560 = w554 & w559;
assign v251 = ~(w554 | w559);
assign w561 = v251;
assign v252 = ~(w560 | w561);
assign w562 = v252;
assign w563 = w440 & w562;
assign v253 = ~(w440 | w562);
assign w564 = v253;
assign v254 = ~(w563 | w564);
assign w565 = v254;
assign w566 = w553 & w565;
assign v255 = ~(w553 | w565);
assign w567 = v255;
assign v256 = ~(w566 | w567);
assign w568 = v256;
assign w569 = w544 & w568;
assign v257 = ~(w544 | w568);
assign w570 = v257;
assign v258 = ~(w569 | w570);
assign w571 = v258;
assign w572 = w504 & ~w571;
assign w573 = ~w504 & w571;
assign v259 = ~(w572 | w573);
assign w574 = v259;
assign w575 = (~w446 & ~w489) | (~w446 & w8585) | (~w489 & w8585);
assign w576 = (~w484 & ~w486) | (~w484 & w8586) | (~w486 & w8586);
assign w577 = w436 & ~w439;
assign v260 = ~(w441 | w577);
assign w578 = v260;
assign v261 = ~(w576 | w578);
assign w579 = v261;
assign w580 = w576 & w578;
assign v262 = ~(w579 | w580);
assign w581 = v262;
assign w582 = ~w575 & w581;
assign w583 = w575 & ~w581;
assign v263 = ~(w582 | w583);
assign w584 = v263;
assign w585 = w574 & ~w584;
assign w586 = ~w574 & w584;
assign v264 = ~(w585 | w586);
assign w587 = v264;
assign v265 = ~(w503 | w587);
assign w588 = v265;
assign w589 = w503 & w587;
assign v266 = ~(w588 | w589);
assign w590 = v266;
assign w591 = w502 & w590;
assign v267 = ~(w502 | w590);
assign w592 = v267;
assign v268 = ~(w591 | w592);
assign w593 = v268;
assign v269 = ~(w496 | w588);
assign w594 = v269;
assign w595 = (~w589 & w500) | (~w589 & w8677) | (w500 & w8677);
assign v270 = ~(w579 | w582);
assign w596 = v270;
assign w597 = pi07 & pi37;
assign w598 = pi11 & pi33;
assign w599 = pi12 & pi32;
assign w600 = pi76 & w599;
assign v271 = ~(pi76 | w599);
assign w601 = v271;
assign v272 = ~(w600 | w601);
assign w602 = v272;
assign w603 = w598 & w602;
assign v273 = ~(w598 | w602);
assign w604 = v273;
assign v274 = ~(w603 | w604);
assign w605 = v274;
assign w606 = w597 & w605;
assign v275 = ~(w597 | w605);
assign w607 = v275;
assign v276 = ~(w606 | w607);
assign w608 = v276;
assign w609 = pi08 & pi36;
assign w610 = pi10 & pi34;
assign v277 = ~(w520 | w610);
assign w611 = v277;
assign w612 = pi10 & pi35;
assign w613 = w518 & w612;
assign v278 = ~(w611 | w613);
assign w614 = v278;
assign w615 = w609 & ~w614;
assign w616 = ~w609 & w614;
assign v279 = ~(w615 | w616);
assign w617 = v279;
assign w618 = w608 & ~w617;
assign w619 = ~w608 & w617;
assign v280 = ~(w618 | w619);
assign w620 = v280;
assign w621 = (~w514 & ~w516) | (~w514 & w8678) | (~w516 & w8678);
assign w622 = w562 & w8587;
assign w623 = w440 & w554;
assign w624 = w558 & ~w623;
assign v281 = ~(w560 | w624);
assign w625 = v281;
assign w626 = ~w622 & w625;
assign w627 = (~w508 & ~w510) | (~w508 & w8679) | (~w510 & w8679);
assign w628 = w517 & ~w519;
assign v282 = ~(w521 | w628);
assign w629 = v282;
assign v283 = ~(w627 | w629);
assign w630 = v283;
assign w631 = w627 & w629;
assign v284 = ~(w630 | w631);
assign w632 = v284;
assign w633 = w626 & ~w632;
assign w634 = ~w626 & w632;
assign v285 = ~(w633 | w634);
assign w635 = v285;
assign w636 = w621 & ~w635;
assign w637 = ~w621 & w635;
assign v286 = ~(w636 | w637);
assign w638 = v286;
assign w639 = w620 & w638;
assign v287 = ~(w620 | w638);
assign w640 = v287;
assign v288 = ~(w639 | w640);
assign w641 = v288;
assign v289 = ~(w529 | w534);
assign w642 = v289;
assign v290 = ~(w533 | w642);
assign w643 = v290;
assign w644 = pi00 & pi44;
assign v291 = ~(w548 | w644);
assign w645 = v291;
assign w646 = pi01 & pi44;
assign w647 = w545 & w646;
assign v292 = ~(w645 | w647);
assign w648 = v292;
assign w649 = pi03 & pi41;
assign w650 = pi02 & pi42;
assign v293 = ~(w649 | w650);
assign w651 = v293;
assign w652 = pi03 & pi42;
assign w653 = w440 & w652;
assign v294 = ~(w651 | w653);
assign w654 = v294;
assign w655 = pi04 & pi40;
assign w656 = pi06 & pi38;
assign v295 = ~(w557 | w656);
assign w657 = v295;
assign w658 = pi06 & pi39;
assign w659 = w555 & w658;
assign v296 = ~(w657 | w659);
assign w660 = v296;
assign w661 = w655 & ~w660;
assign w662 = ~w655 & w660;
assign v297 = ~(w661 | w662);
assign w663 = v297;
assign w664 = w654 & ~w663;
assign w665 = ~w654 & w663;
assign v298 = ~(w664 | w665);
assign w666 = v298;
assign w667 = w648 & ~w666;
assign w668 = ~w648 & w666;
assign v299 = ~(w667 | w668);
assign w669 = v299;
assign w670 = w643 & w669;
assign v300 = ~(w643 | w669);
assign w671 = v300;
assign v301 = ~(w670 | w671);
assign w672 = v301;
assign w673 = w641 & w672;
assign v302 = ~(w641 | w672);
assign w674 = v302;
assign v303 = ~(w673 | w674);
assign w675 = v303;
assign w676 = ~w596 & w675;
assign w677 = w596 & ~w675;
assign v304 = ~(w676 | w677);
assign w678 = v304;
assign v305 = ~(w566 | w569);
assign w679 = v305;
assign v306 = ~(w549 | w551);
assign w680 = v306;
assign w681 = w434 & w541;
assign v307 = ~(w542 | w681);
assign w682 = v307;
assign v308 = ~(w680 | w682);
assign w683 = v308;
assign w684 = w680 & w682;
assign v309 = ~(w683 | w684);
assign w685 = v309;
assign w686 = w679 & ~w685;
assign w687 = ~w679 & w685;
assign v310 = ~(w686 | w687);
assign w688 = v310;
assign w689 = w678 & ~w688;
assign w690 = ~w678 & w688;
assign v311 = ~(w689 | w690);
assign w691 = v311;
assign v312 = ~(w572 | w585);
assign w692 = v312;
assign w693 = w691 & ~w692;
assign w694 = ~w691 & w692;
assign v313 = ~(w693 | w694);
assign w695 = v313;
assign w696 = w595 & ~w695;
assign w697 = ~w595 & w695;
assign v314 = ~(w696 | w697);
assign w698 = v314;
assign v315 = ~(w595 | w694);
assign w699 = v315;
assign v316 = ~(w693 | w699);
assign w700 = v316;
assign v317 = ~(w677 | w689);
assign w701 = v317;
assign w702 = pi05 & pi40;
assign w703 = pi07 & pi38;
assign v318 = ~(w658 | w703);
assign w704 = v318;
assign w705 = pi07 & pi39;
assign w706 = w656 & w705;
assign v319 = ~(w704 | w706);
assign w707 = v319;
assign w708 = w702 & ~w707;
assign w709 = ~w702 & w707;
assign v320 = ~(w708 | w709);
assign w710 = v320;
assign w711 = w646 & ~w710;
assign w712 = ~w646 & w710;
assign v321 = ~(w711 | w712);
assign w713 = v321;
assign w714 = pi02 & pi43;
assign w715 = pi04 & pi41;
assign v322 = ~(w652 | w715);
assign w716 = v322;
assign w717 = pi04 & pi42;
assign w718 = w649 & w717;
assign v323 = ~(w716 | w718);
assign w719 = v323;
assign w720 = w714 & ~w719;
assign w721 = ~w714 & w719;
assign v324 = ~(w720 | w721);
assign w722 = v324;
assign w723 = w713 & ~w722;
assign w724 = ~w713 & w722;
assign v325 = ~(w723 | w724);
assign w725 = v325;
assign w726 = pi00 & pi45;
assign w727 = w558 & w623;
assign w728 = w726 & w727;
assign v326 = ~(w726 | w727);
assign w729 = v326;
assign v327 = ~(w728 | w729);
assign w730 = v327;
assign w731 = (~w630 & w621) | (~w630 & w9234) | (w621 & w9234);
assign w732 = ~w730 & w731;
assign w733 = w730 & ~w731;
assign v328 = ~(w732 | w733);
assign w734 = v328;
assign w735 = w725 & w734;
assign v329 = ~(w725 | w734);
assign w736 = v329;
assign v330 = ~(w735 | w736);
assign w737 = v330;
assign w738 = (~w606 & ~w608) | (~w606 & w8680) | (~w608 & w8680);
assign v331 = ~(w600 | w603);
assign w739 = v331;
assign w740 = w609 & ~w611;
assign v332 = ~(w613 | w740);
assign w741 = v332;
assign v333 = ~(w739 | w741);
assign w742 = v333;
assign w743 = w739 & w741;
assign v334 = ~(w742 | w743);
assign w744 = v334;
assign w745 = ~w738 & w744;
assign w746 = w738 & ~w744;
assign v335 = ~(w745 | w746);
assign w747 = v335;
assign w748 = pi08 & pi37;
assign w749 = pi12 & pi33;
assign w750 = pi13 & pi32;
assign w751 = pi77 & w750;
assign v336 = ~(pi77 | w750);
assign w752 = v336;
assign v337 = ~(w751 | w752);
assign w753 = v337;
assign w754 = w749 & w753;
assign v338 = ~(w749 | w753);
assign w755 = v338;
assign v339 = ~(w754 | w755);
assign w756 = v339;
assign w757 = w748 & w756;
assign v340 = ~(w748 | w756);
assign w758 = v340;
assign v341 = ~(w757 | w758);
assign w759 = v341;
assign w760 = pi09 & pi36;
assign w761 = pi11 & pi34;
assign v342 = ~(w612 | w761);
assign w762 = v342;
assign w763 = pi11 & pi35;
assign w764 = w610 & w763;
assign v343 = ~(w762 | w764);
assign w765 = v343;
assign w766 = w760 & ~w765;
assign w767 = ~w760 & w765;
assign v344 = ~(w766 | w767);
assign w768 = v344;
assign w769 = w759 & ~w768;
assign w770 = ~w759 & w768;
assign v345 = ~(w769 | w770);
assign w771 = v345;
assign w772 = (~w653 & w663) | (~w653 & w9235) | (w663 & w9235);
assign w773 = w655 & ~w657;
assign v346 = ~(w659 | w773);
assign w774 = v346;
assign v347 = ~(w772 | w774);
assign w775 = v347;
assign w776 = w772 & w774;
assign v348 = ~(w775 | w776);
assign w777 = v348;
assign v349 = ~(w771 | w777);
assign w778 = v349;
assign w779 = w771 & w777;
assign v350 = ~(w778 | w779);
assign w780 = v350;
assign w781 = w747 & ~w780;
assign w782 = ~w747 & w780;
assign v351 = ~(w781 | w782);
assign w783 = v351;
assign w784 = w737 & ~w783;
assign w785 = ~w737 & w783;
assign v352 = ~(w784 | w785);
assign w786 = v352;
assign w787 = w666 & ~w672;
assign v353 = ~(w673 | w787);
assign w788 = v353;
assign v354 = ~(w626 | w638);
assign w789 = v354;
assign v355 = ~(w639 | w789);
assign w790 = v355;
assign v356 = ~(w643 | w645);
assign w791 = v356;
assign v357 = ~(w647 | w791);
assign w792 = v357;
assign v358 = ~(w790 | w792);
assign w793 = v358;
assign w794 = w790 & w792;
assign v359 = ~(w793 | w794);
assign w795 = v359;
assign w796 = ~w788 & w795;
assign w797 = w788 & ~w795;
assign v360 = ~(w796 | w797);
assign w798 = v360;
assign v361 = ~(w683 | w687);
assign w799 = v361;
assign w800 = ~w798 & w799;
assign w801 = w798 & ~w799;
assign v362 = ~(w800 | w801);
assign w802 = v362;
assign w803 = w786 & ~w802;
assign w804 = ~w786 & w802;
assign v363 = ~(w803 | w804);
assign w805 = v363;
assign w806 = w701 & ~w805;
assign w807 = ~w701 & w805;
assign v364 = ~(w806 | w807);
assign w808 = v364;
assign v365 = ~(w700 | w808);
assign w809 = v365;
assign w810 = ~w693 & w808;
assign w811 = ~w699 & w810;
assign v366 = ~(w809 | w811);
assign w812 = v366;
assign v367 = ~(w806 | w811);
assign w813 = v367;
assign w814 = pi08 & pi38;
assign w815 = pi09 & pi37;
assign w816 = pi10 & pi36;
assign v368 = ~(w815 | w816);
assign w817 = v368;
assign w818 = pi10 & pi37;
assign w819 = w760 & w818;
assign v369 = ~(w817 | w819);
assign w820 = v369;
assign w821 = w814 & ~w820;
assign w822 = ~w814 & w820;
assign v370 = ~(w821 | w822);
assign w823 = v370;
assign w824 = pi12 & pi34;
assign w825 = pi13 & pi33;
assign v371 = ~(w824 | w825);
assign w826 = v371;
assign w827 = pi13 & pi34;
assign w828 = w749 & w827;
assign v372 = ~(w826 | w828);
assign w829 = v372;
assign w830 = ~w705 & w763;
assign w831 = w705 & ~w763;
assign v373 = ~(w830 | w831);
assign w832 = v373;
assign w833 = w829 & w832;
assign v374 = ~(w829 | w832);
assign w834 = v374;
assign v375 = ~(w833 | w834);
assign w835 = v375;
assign v376 = ~(w823 | w835);
assign w836 = v376;
assign w837 = w823 & w835;
assign v377 = ~(w836 | w837);
assign w838 = v377;
assign w839 = (~w757 & ~w759) | (~w757 & w8588) | (~w759 & w8588);
assign w840 = (~w751 & ~w753) | (~w751 & w9236) | (~w753 & w9236);
assign w841 = w760 & ~w762;
assign v378 = ~(w764 | w841);
assign w842 = v378;
assign v379 = ~(w840 | w842);
assign w843 = v379;
assign w844 = w840 & w842;
assign v380 = ~(w843 | w844);
assign w845 = v380;
assign w846 = ~w839 & w845;
assign w847 = w839 & ~w845;
assign v381 = ~(w846 | w847);
assign w848 = v381;
assign w849 = (~w711 & ~w713) | (~w711 & w8681) | (~w713 & w8681);
assign w850 = w714 & ~w716;
assign v382 = ~(w718 | w850);
assign w851 = v382;
assign w852 = w702 & ~w704;
assign v383 = ~(w706 | w852);
assign w853 = v383;
assign v384 = ~(w851 | w853);
assign w854 = v384;
assign w855 = w851 & w853;
assign v385 = ~(w854 | w855);
assign w856 = v385;
assign w857 = w849 & ~w856;
assign w858 = ~w849 & w856;
assign v386 = ~(w857 | w858);
assign w859 = v386;
assign w860 = w848 & w859;
assign v387 = ~(w848 | w859);
assign w861 = v387;
assign v388 = ~(w860 | w861);
assign w862 = v388;
assign w863 = w838 & w862;
assign v389 = ~(w838 | w862);
assign w864 = v389;
assign v390 = ~(w863 | w864);
assign w865 = v390;
assign w866 = pi00 & pi46;
assign w867 = pi05 & pi41;
assign w868 = pi06 & pi40;
assign v391 = ~(w867 | w868);
assign w869 = v391;
assign w870 = pi06 & pi41;
assign w871 = w702 & w870;
assign v392 = ~(w869 | w871);
assign w872 = v392;
assign w873 = w717 & ~w872;
assign w874 = ~w717 & w872;
assign v393 = ~(w873 | w874);
assign w875 = v393;
assign w876 = w866 & ~w875;
assign w877 = ~w866 & w875;
assign v394 = ~(w876 | w877);
assign w878 = v394;
assign w879 = pi01 & pi45;
assign w880 = pi02 & pi44;
assign w881 = pi03 & pi43;
assign v395 = ~(w880 | w881);
assign w882 = v395;
assign w883 = pi03 & pi44;
assign w884 = w714 & w883;
assign v396 = ~(w882 | w884);
assign w885 = v396;
assign w886 = w879 & ~w885;
assign w887 = ~w879 & w885;
assign v397 = ~(w886 | w887);
assign w888 = v397;
assign w889 = w878 & ~w888;
assign w890 = ~w878 & w888;
assign v398 = ~(w889 | w890);
assign w891 = v398;
assign w892 = (~w742 & w738) | (~w742 & w9237) | (w738 & w9237);
assign w893 = pi14 & pi32;
assign w894 = pi78 & w893;
assign v399 = ~(pi78 | w893);
assign w895 = v399;
assign v400 = ~(w894 | w895);
assign w896 = v400;
assign v401 = ~(w775 | w896);
assign w897 = v401;
assign w898 = w775 & w896;
assign v402 = ~(w897 | w898);
assign w899 = v402;
assign w900 = w892 & ~w899;
assign w901 = ~w892 & w899;
assign v403 = ~(w900 | w901);
assign w902 = v403;
assign w903 = w891 & w902;
assign v404 = ~(w891 | w902);
assign w904 = v404;
assign v405 = ~(w903 | w904);
assign w905 = v405;
assign w906 = w865 & w905;
assign v406 = ~(w865 | w905);
assign w907 = v406;
assign v407 = ~(w906 | w907);
assign w908 = v407;
assign v408 = ~(w793 | w796);
assign w909 = v408;
assign v409 = ~(w735 | w784);
assign w910 = v409;
assign v410 = ~(w778 | w782);
assign w911 = v410;
assign v411 = ~(w728 | w733);
assign w912 = v411;
assign w913 = w911 & ~w912;
assign w914 = ~w911 & w912;
assign v412 = ~(w913 | w914);
assign w915 = v412;
assign w916 = ~w910 & w915;
assign w917 = w910 & ~w915;
assign v413 = ~(w916 | w917);
assign w918 = v413;
assign w919 = ~w909 & w918;
assign w920 = w909 & ~w918;
assign v414 = ~(w919 | w920);
assign w921 = v414;
assign w922 = w908 & w921;
assign v415 = ~(w908 | w921);
assign w923 = v415;
assign v416 = ~(w922 | w923);
assign w924 = v416;
assign v417 = ~(w800 | w804);
assign w925 = v417;
assign w926 = w924 & w925;
assign v418 = ~(w924 | w925);
assign w927 = v418;
assign v419 = ~(w926 | w927);
assign w928 = v419;
assign w929 = w813 & ~w928;
assign w930 = ~w813 & w928;
assign v420 = ~(w929 | w930);
assign w931 = v420;
assign v421 = ~(w806 | w926);
assign w932 = v421;
assign w933 = (~w927 & w811) | (~w927 & w8682) | (w811 & w8682);
assign v422 = ~(w919 | w922);
assign w934 = v422;
assign v423 = ~(w913 | w916);
assign w935 = v423;
assign w936 = (~w903 & ~w865) | (~w903 & w9238) | (~w865 & w9238);
assign w937 = (~w860 & ~w862) | (~w860 & w9239) | (~w862 & w9239);
assign v424 = ~(w898 | w901);
assign w938 = v424;
assign v425 = ~(w937 | w938);
assign w939 = v425;
assign w940 = w937 & w938;
assign v426 = ~(w939 | w940);
assign w941 = v426;
assign w942 = ~w936 & w941;
assign w943 = w936 & ~w941;
assign v427 = ~(w942 | w943);
assign w944 = v427;
assign w945 = w935 & ~w944;
assign w946 = ~w935 & w944;
assign v428 = ~(w945 | w946);
assign w947 = v428;
assign w948 = pi04 & pi43;
assign w949 = pi05 & pi42;
assign v429 = ~(w948 | w949);
assign w950 = v429;
assign w951 = pi05 & pi43;
assign w952 = w717 & w951;
assign v430 = ~(w950 | w952);
assign w953 = v430;
assign w954 = w883 & ~w953;
assign w955 = ~w883 & w953;
assign v431 = ~(w954 | w955);
assign w956 = v431;
assign w957 = w894 & ~w956;
assign w958 = ~w894 & w956;
assign v432 = ~(w957 | w958);
assign w959 = v432;
assign w960 = pi00 & pi47;
assign w961 = pi01 & pi46;
assign w962 = pi02 & pi45;
assign v433 = ~(w961 | w962);
assign w963 = v433;
assign w964 = pi02 & pi46;
assign w965 = w879 & w964;
assign v434 = ~(w963 | w965);
assign w966 = v434;
assign w967 = w960 & ~w966;
assign w968 = ~w960 & w966;
assign v435 = ~(w967 | w968);
assign w969 = v435;
assign w970 = w959 & ~w969;
assign w971 = ~w959 & w969;
assign v436 = ~(w970 | w971);
assign w972 = v436;
assign w973 = pi15 & pi32;
assign v437 = ~(pi79 | w973);
assign w974 = v437;
assign w975 = pi79 & w973;
assign v438 = ~(w974 | w975);
assign w976 = v438;
assign w977 = pi14 & pi33;
assign v439 = ~(w827 | w977);
assign w978 = v439;
assign w979 = w827 & w977;
assign v440 = ~(w978 | w979);
assign w980 = v440;
assign w981 = w976 & ~w980;
assign w982 = ~w976 & w980;
assign v441 = ~(w981 | w982);
assign w983 = v441;
assign w984 = ~w844 & w983;
assign w985 = (w984 & ~w839) | (w984 & w8683) | (~w839 & w8683);
assign v442 = ~(w843 | w983);
assign w986 = v442;
assign w987 = (w986 & w839) | (w986 & w8684) | (w839 & w8684);
assign v443 = ~(w985 | w987);
assign w988 = v443;
assign w989 = (~w854 & w849) | (~w854 & w9240) | (w849 & w9240);
assign w990 = ~w988 & w989;
assign w991 = w988 & ~w989;
assign v444 = ~(w990 | w991);
assign w992 = v444;
assign w993 = w972 & ~w992;
assign w994 = ~w972 & w992;
assign v445 = ~(w993 | w994);
assign w995 = v445;
assign w996 = pi11 & pi36;
assign w997 = pi12 & pi35;
assign v446 = ~(w996 | w997);
assign w998 = v446;
assign w999 = pi12 & pi36;
assign w1000 = w763 & w999;
assign v447 = ~(w998 | w1000);
assign w1001 = v447;
assign w1002 = w818 & ~w1001;
assign w1003 = ~w818 & w1001;
assign v448 = ~(w1002 | w1003);
assign w1004 = v448;
assign w1005 = w870 & ~w1004;
assign w1006 = ~w870 & w1004;
assign v449 = ~(w1005 | w1006);
assign w1007 = v449;
assign w1008 = pi07 & pi40;
assign w1009 = pi08 & pi39;
assign w1010 = pi09 & pi38;
assign v450 = ~(w1009 | w1010);
assign w1011 = v450;
assign w1012 = pi09 & pi39;
assign w1013 = w814 & w1012;
assign v451 = ~(w1011 | w1013);
assign w1014 = v451;
assign w1015 = w1008 & ~w1014;
assign w1016 = ~w1008 & w1014;
assign v452 = ~(w1015 | w1016);
assign w1017 = v452;
assign w1018 = w1007 & ~w1017;
assign w1019 = ~w1007 & w1017;
assign v453 = ~(w1018 | w1019);
assign w1020 = v453;
assign w1021 = (~w876 & ~w878) | (~w876 & w8685) | (~w878 & w8685);
assign w1022 = w879 & ~w882;
assign v454 = ~(w884 | w1022);
assign w1023 = v454;
assign w1024 = w717 & ~w869;
assign v455 = ~(w871 | w1024);
assign w1025 = v455;
assign v456 = ~(w1023 | w1025);
assign w1026 = v456;
assign w1027 = w1023 & w1025;
assign v457 = ~(w1026 | w1027);
assign w1028 = v457;
assign w1029 = ~w1021 & w1028;
assign w1030 = w1021 & ~w1028;
assign v458 = ~(w1029 | w1030);
assign w1031 = v458;
assign w1032 = w763 & ~w826;
assign v459 = ~(w828 | w1032);
assign w1033 = v459;
assign w1034 = w814 & ~w817;
assign v460 = ~(w819 | w1034);
assign w1035 = v460;
assign v461 = ~(w1033 | w1035);
assign w1036 = v461;
assign w1037 = w1033 & w1035;
assign v462 = ~(w1036 | w1037);
assign w1038 = v462;
assign w1039 = w705 & w835;
assign v463 = ~(w836 | w1039);
assign w1040 = v463;
assign w1041 = w1038 & ~w1040;
assign w1042 = ~w1038 & w1040;
assign v464 = ~(w1041 | w1042);
assign w1043 = v464;
assign w1044 = w1031 & w1043;
assign v465 = ~(w1031 | w1043);
assign w1045 = v465;
assign v466 = ~(w1044 | w1045);
assign w1046 = v466;
assign w1047 = w1020 & ~w1046;
assign w1048 = ~w1020 & w1046;
assign v467 = ~(w1047 | w1048);
assign w1049 = v467;
assign w1050 = ~w995 & w1049;
assign w1051 = w995 & ~w1049;
assign v468 = ~(w1050 | w1051);
assign w1052 = v468;
assign w1053 = w947 & ~w1052;
assign w1054 = ~w947 & w1052;
assign v469 = ~(w1053 | w1054);
assign w1055 = v469;
assign v470 = ~(w934 | w1055);
assign w1056 = v470;
assign w1057 = w934 & w1055;
assign v471 = ~(w1056 | w1057);
assign w1058 = v471;
assign w1059 = w933 & ~w1058;
assign w1060 = ~w933 & w1058;
assign v472 = ~(w1059 | w1060);
assign w1061 = v472;
assign w1062 = (~w1026 & w1021) | (~w1026 & w9241) | (w1021 & w9241);
assign w1063 = pi14 & pi34;
assign w1064 = pi13 & pi35;
assign v473 = ~(w1063 | w1064);
assign w1065 = v473;
assign w1066 = pi14 & pi35;
assign w1067 = w827 & w1066;
assign v474 = ~(w1065 | w1067);
assign w1068 = v474;
assign w1069 = pi15 & pi33;
assign w1070 = pi16 & pi32;
assign w1071 = pi80 & w1070;
assign v475 = ~(pi80 | w1070);
assign w1072 = v475;
assign v476 = ~(w1071 | w1072);
assign w1073 = v476;
assign w1074 = w1069 & ~w1073;
assign w1075 = ~w1069 & w1073;
assign v477 = ~(w1074 | w1075);
assign w1076 = v477;
assign w1077 = w1068 & ~w1076;
assign w1078 = ~w1068 & w1076;
assign v478 = ~(w1077 | w1078);
assign w1079 = v478;
assign w1080 = (~w1036 & w1040) | (~w1036 & w8686) | (w1040 & w8686);
assign w1081 = w1079 & ~w1080;
assign w1082 = ~w1079 & w1080;
assign v479 = ~(w1081 | w1082);
assign w1083 = v479;
assign w1084 = ~w1062 & w1083;
assign w1085 = w1062 & ~w1083;
assign v480 = ~(w1084 | w1085);
assign w1086 = v480;
assign w1087 = pi03 & pi45;
assign w1088 = pi04 & pi44;
assign v481 = ~(w951 | w1088);
assign w1089 = v481;
assign w1090 = pi05 & pi44;
assign w1091 = w948 & w1090;
assign v482 = ~(w1089 | w1091);
assign w1092 = v482;
assign w1093 = w1087 & ~w1092;
assign w1094 = ~w1087 & w1092;
assign v483 = ~(w1093 | w1094);
assign w1095 = v483;
assign w1096 = w976 & ~w978;
assign w1097 = w975 & ~w979;
assign w1098 = w974 & w979;
assign v484 = ~(w1097 | w1098);
assign w1099 = v484;
assign w1100 = ~w1096 & w1099;
assign v485 = ~(w1095 | w1100);
assign w1101 = v485;
assign w1102 = w1095 & w1100;
assign v486 = ~(w1101 | w1102);
assign w1103 = v486;
assign w1104 = pi00 & pi48;
assign w1105 = pi01 & pi47;
assign v487 = ~(w964 | w1105);
assign w1106 = v487;
assign w1107 = pi02 & pi47;
assign w1108 = w961 & w1107;
assign v488 = ~(w1106 | w1108);
assign w1109 = v488;
assign w1110 = w1104 & ~w1109;
assign w1111 = ~w1104 & w1109;
assign v489 = ~(w1110 | w1111);
assign w1112 = v489;
assign w1113 = w1103 & w1112;
assign v490 = ~(w1103 | w1112);
assign w1114 = v490;
assign v491 = ~(w1113 | w1114);
assign w1115 = v491;
assign w1116 = w1086 & ~w1115;
assign w1117 = ~w1086 & w1115;
assign v492 = ~(w1116 | w1117);
assign w1118 = v492;
assign w1119 = pi06 & pi42;
assign w1120 = pi11 & pi37;
assign v493 = ~(w999 | w1120);
assign w1121 = v493;
assign w1122 = pi12 & pi37;
assign w1123 = w996 & w1122;
assign v494 = ~(w1121 | w1123);
assign w1124 = v494;
assign w1125 = pi10 & pi38;
assign w1126 = ~w1124 & w1125;
assign w1127 = w1124 & ~w1125;
assign v495 = ~(w1126 | w1127);
assign w1128 = v495;
assign w1129 = w1119 & ~w1128;
assign w1130 = ~w1119 & w1128;
assign v496 = ~(w1129 | w1130);
assign w1131 = v496;
assign w1132 = pi07 & pi41;
assign w1133 = pi08 & pi40;
assign v497 = ~(w1012 | w1133);
assign w1134 = v497;
assign w1135 = pi09 & pi40;
assign w1136 = w1009 & w1135;
assign v498 = ~(w1134 | w1136);
assign w1137 = v498;
assign w1138 = w1132 & ~w1137;
assign w1139 = ~w1132 & w1137;
assign v499 = ~(w1138 | w1139);
assign w1140 = v499;
assign w1141 = w1131 & ~w1140;
assign w1142 = ~w1131 & w1140;
assign v500 = ~(w1141 | w1142);
assign w1143 = v500;
assign w1144 = (~w957 & ~w959) | (~w957 & w8687) | (~w959 & w8687);
assign w1145 = w960 & ~w963;
assign v501 = ~(w965 | w1145);
assign w1146 = v501;
assign w1147 = w883 & ~w950;
assign v502 = ~(w952 | w1147);
assign w1148 = v502;
assign v503 = ~(w1146 | w1148);
assign w1149 = v503;
assign w1150 = w1146 & w1148;
assign v504 = ~(w1149 | w1150);
assign w1151 = v504;
assign w1152 = ~w1144 & w1151;
assign w1153 = w1144 & ~w1151;
assign v505 = ~(w1152 | w1153);
assign w1154 = v505;
assign w1155 = w818 & ~w998;
assign v506 = ~(w1000 | w1155);
assign w1156 = v506;
assign w1157 = w1008 & ~w1011;
assign v507 = ~(w1013 | w1157);
assign w1158 = v507;
assign v508 = ~(w1156 | w1158);
assign w1159 = v508;
assign w1160 = w1156 & w1158;
assign v509 = ~(w1159 | w1160);
assign w1161 = v509;
assign w1162 = (~w1005 & ~w1007) | (~w1005 & w8688) | (~w1007 & w8688);
assign w1163 = w1161 & ~w1162;
assign w1164 = ~w1161 & w1162;
assign v510 = ~(w1163 | w1164);
assign w1165 = v510;
assign v511 = ~(w1154 | w1165);
assign w1166 = v511;
assign w1167 = w1154 & w1165;
assign v512 = ~(w1166 | w1167);
assign w1168 = v512;
assign w1169 = w1143 & ~w1168;
assign w1170 = ~w1143 & w1168;
assign v513 = ~(w1169 | w1170);
assign w1171 = v513;
assign w1172 = w1118 & ~w1171;
assign w1173 = ~w1118 & w1171;
assign v514 = ~(w1172 | w1173);
assign w1174 = v514;
assign v515 = ~(w939 | w942);
assign w1175 = v515;
assign v516 = ~(w993 | w1051);
assign w1176 = v516;
assign w1177 = w983 & ~w985;
assign v517 = ~(w990 | w1177);
assign w1178 = v517;
assign w1179 = (~w1045 & ~w1046) | (~w1045 & w9242) | (~w1046 & w9242);
assign w1180 = w1178 & w1179;
assign v518 = ~(w1178 | w1179);
assign w1181 = v518;
assign v519 = ~(w1180 | w1181);
assign w1182 = v519;
assign w1183 = w1176 & ~w1182;
assign w1184 = ~w1176 & w1182;
assign v520 = ~(w1183 | w1184);
assign w1185 = v520;
assign w1186 = w1175 & ~w1185;
assign w1187 = ~w1175 & w1185;
assign v521 = ~(w1186 | w1187);
assign w1188 = v521;
assign w1189 = w1174 & ~w1188;
assign w1190 = ~w1174 & w1188;
assign v522 = ~(w1189 | w1190);
assign w1191 = v522;
assign v523 = ~(w945 | w1053);
assign w1192 = v523;
assign w1193 = ~w1191 & w1192;
assign w1194 = w1191 & ~w1192;
assign v524 = ~(w1193 | w1194);
assign w1195 = v524;
assign v525 = ~(w1056 | w933);
assign w1196 = v525;
assign v526 = ~(w1057 | w1196);
assign w1197 = v526;
assign v527 = ~(w1195 | w1197);
assign w1198 = v527;
assign w1199 = w1195 & w1197;
assign v528 = ~(w1198 | w1199);
assign w1200 = v528;
assign v529 = ~(w1193 | w1199);
assign w1201 = v529;
assign w1202 = pi11 & pi38;
assign w1203 = pi10 & pi39;
assign v530 = ~(w1202 | w1203);
assign w1204 = v530;
assign w1205 = pi11 & pi39;
assign w1206 = w1125 & w1205;
assign v531 = ~(w1204 | w1206);
assign w1207 = v531;
assign w1208 = w1135 & ~w1207;
assign w1209 = ~w1135 & w1207;
assign v532 = ~(w1208 | w1209);
assign w1210 = v532;
assign w1211 = w1090 & ~w1210;
assign w1212 = ~w1090 & w1210;
assign v533 = ~(w1211 | w1212);
assign w1213 = v533;
assign w1214 = pi06 & pi43;
assign w1215 = pi07 & pi42;
assign w1216 = pi08 & pi41;
assign v534 = ~(w1215 | w1216);
assign w1217 = v534;
assign w1218 = pi08 & pi42;
assign w1219 = w1132 & w1218;
assign v535 = ~(w1217 | w1219);
assign w1220 = v535;
assign w1221 = w1214 & ~w1220;
assign w1222 = ~w1214 & w1220;
assign v536 = ~(w1221 | w1222);
assign w1223 = v536;
assign w1224 = w1213 & ~w1223;
assign w1225 = ~w1213 & w1223;
assign v537 = ~(w1224 | w1225);
assign w1226 = v537;
assign w1227 = ~w1121 & w1125;
assign v538 = ~(w1123 | w1227);
assign w1228 = v538;
assign w1229 = w1132 & ~w1134;
assign v539 = ~(w1136 | w1229);
assign w1230 = v539;
assign v540 = ~(w1228 | w1230);
assign w1231 = v540;
assign w1232 = w1228 & w1230;
assign v541 = ~(w1231 | w1232);
assign w1233 = v541;
assign w1234 = (~w1129 & ~w1131) | (~w1129 & w8689) | (~w1131 & w8689);
assign w1235 = w1233 & ~w1234;
assign w1236 = ~w1233 & w1234;
assign v542 = ~(w1235 | w1236);
assign w1237 = v542;
assign w1238 = w1104 & ~w1106;
assign v543 = ~(w1108 | w1238);
assign w1239 = v543;
assign w1240 = w1087 & ~w1089;
assign v544 = ~(w1091 | w1240);
assign w1241 = v544;
assign v545 = ~(w1239 | w1241);
assign w1242 = v545;
assign w1243 = w1239 & w1241;
assign v546 = ~(w1242 | w1243);
assign w1244 = v546;
assign v547 = ~(w1102 | w1113);
assign w1245 = v547;
assign w1246 = w1244 & w1245;
assign v548 = ~(w1244 | w1245);
assign w1247 = v548;
assign v549 = ~(w1246 | w1247);
assign w1248 = v549;
assign w1249 = w1237 & w1248;
assign v550 = ~(w1237 | w1248);
assign w1250 = v550;
assign v551 = ~(w1249 | w1250);
assign w1251 = v551;
assign w1252 = w1226 & w1251;
assign v552 = ~(w1226 | w1251);
assign w1253 = v552;
assign v553 = ~(w1252 | w1253);
assign w1254 = v553;
assign v554 = ~(w1149 | w1152);
assign w1255 = v554;
assign w1256 = pi13 & pi36;
assign w1257 = pi15 & pi34;
assign v555 = ~(w1066 | w1257);
assign w1258 = v555;
assign w1259 = pi15 & pi35;
assign w1260 = w1063 & w1259;
assign v556 = ~(w1258 | w1260);
assign w1261 = v556;
assign w1262 = w1256 & ~w1261;
assign w1263 = ~w1256 & w1261;
assign v557 = ~(w1262 | w1263);
assign w1264 = v557;
assign w1265 = pi17 & pi32;
assign w1266 = pi81 & w1265;
assign v558 = ~(pi81 | w1265);
assign w1267 = v558;
assign v559 = ~(w1266 | w1267);
assign w1268 = v559;
assign w1269 = pi16 & pi33;
assign w1270 = ~w1122 & w1269;
assign w1271 = w1122 & ~w1269;
assign v560 = ~(w1270 | w1271);
assign w1272 = v560;
assign w1273 = w1268 & w1272;
assign v561 = ~(w1268 | w1272);
assign w1274 = v561;
assign v562 = ~(w1273 | w1274);
assign w1275 = v562;
assign v563 = ~(w1264 | w1275);
assign w1276 = v563;
assign w1277 = w1264 & w1275;
assign v564 = ~(w1276 | w1277);
assign w1278 = v564;
assign w1279 = (~w1159 & w1162) | (~w1159 & w9243) | (w1162 & w9243);
assign w1280 = ~w1278 & w1279;
assign w1281 = w1278 & ~w1279;
assign v565 = ~(w1280 | w1281);
assign w1282 = v565;
assign w1283 = w1255 & w1282;
assign v566 = ~(w1255 | w1282);
assign w1284 = v566;
assign v567 = ~(w1283 | w1284);
assign w1285 = v567;
assign v568 = ~(w1069 | w1071);
assign w1286 = v568;
assign v569 = ~(w1072 | w1286);
assign w1287 = v569;
assign w1288 = (w1076 & w8690) | (w1076 & w8691) | (w8690 & w8691);
assign w1289 = (~w1076 & w8692) | (~w1076 & w8693) | (w8692 & w8693);
assign v570 = ~(w1288 | w1289);
assign w1290 = v570;
assign w1291 = pi03 & pi46;
assign w1292 = pi04 & pi45;
assign v571 = ~(w1291 | w1292);
assign w1293 = v571;
assign w1294 = pi04 & pi46;
assign w1295 = w1087 & w1294;
assign v572 = ~(w1293 | w1295);
assign w1296 = v572;
assign w1297 = w1107 & ~w1296;
assign w1298 = ~w1107 & w1296;
assign v573 = ~(w1297 | w1298);
assign w1299 = v573;
assign w1300 = w1290 & ~w1299;
assign w1301 = ~w1290 & w1299;
assign v574 = ~(w1300 | w1301);
assign w1302 = v574;
assign w1303 = pi00 & pi49;
assign w1304 = pi01 & pi48;
assign v575 = ~(w1303 | w1304);
assign w1305 = v575;
assign w1306 = pi01 & pi49;
assign w1307 = w1104 & w1306;
assign v576 = ~(w1305 | w1307);
assign w1308 = v576;
assign w1309 = w975 & w979;
assign w1310 = ~w1308 & w1309;
assign w1311 = w1308 & ~w1309;
assign v577 = ~(w1310 | w1311);
assign w1312 = v577;
assign w1313 = w1302 & w1312;
assign v578 = ~(w1302 | w1312);
assign w1314 = v578;
assign v579 = ~(w1313 | w1314);
assign w1315 = v579;
assign v580 = ~(w1285 | w1315);
assign w1316 = v580;
assign w1317 = w1285 & w1315;
assign v581 = ~(w1316 | w1317);
assign w1318 = v581;
assign w1319 = w1254 & w1318;
assign v582 = ~(w1254 | w1318);
assign w1320 = v582;
assign v583 = ~(w1319 | w1320);
assign w1321 = v583;
assign w1322 = (~w1180 & w1176) | (~w1180 & w9244) | (w1176 & w9244);
assign w1323 = w1321 & ~w1322;
assign w1324 = ~w1321 & w1322;
assign v584 = ~(w1323 | w1324);
assign w1325 = v584;
assign v585 = ~(w1116 | w1172);
assign w1326 = v585;
assign v586 = ~(w1081 | w1084);
assign w1327 = v586;
assign w1328 = (~w1166 & ~w1168) | (~w1166 & w9245) | (~w1168 & w9245);
assign w1329 = ~w1327 & w1328;
assign w1330 = w1327 & ~w1328;
assign v587 = ~(w1329 | w1330);
assign w1331 = v587;
assign w1332 = w1326 & w1331;
assign v588 = ~(w1326 | w1331);
assign w1333 = v588;
assign v589 = ~(w1332 | w1333);
assign w1334 = v589;
assign w1335 = w1325 & ~w1334;
assign w1336 = ~w1325 & w1334;
assign v590 = ~(w1335 | w1336);
assign w1337 = v590;
assign w1338 = (~w1186 & ~w1188) | (~w1186 & w9246) | (~w1188 & w9246);
assign v591 = ~(w1337 | w1338);
assign w1339 = v591;
assign w1340 = w1337 & w1338;
assign v592 = ~(w1339 | w1340);
assign w1341 = v592;
assign w1342 = w1201 & w1341;
assign v593 = ~(w1201 | w1341);
assign w1343 = v593;
assign v594 = ~(w1342 | w1343);
assign w1344 = v594;
assign v595 = ~(w1323 | w1335);
assign w1345 = v595;
assign v596 = ~(w1316 | w1319);
assign w1346 = v596;
assign v597 = ~(w1280 | w1283);
assign w1347 = v597;
assign v598 = ~(w1249 | w1252);
assign w1348 = v598;
assign w1349 = w1347 & ~w1348;
assign w1350 = ~w1347 & w1348;
assign v599 = ~(w1349 | w1350);
assign w1351 = v599;
assign w1352 = ~w1346 & w1351;
assign w1353 = w1346 & ~w1351;
assign v600 = ~(w1352 | w1353);
assign w1354 = v600;
assign v601 = ~(w1242 | w1246);
assign w1355 = v601;
assign w1356 = pi12 & pi38;
assign v602 = ~(w1205 | w1356);
assign w1357 = v602;
assign w1358 = pi12 & pi39;
assign w1359 = w1202 & w1358;
assign v603 = ~(w1357 | w1359);
assign w1360 = v603;
assign w1361 = (~w1231 & w1234) | (~w1231 & w9247) | (w1234 & w9247);
assign w1362 = ~w1360 & w1361;
assign w1363 = w1360 & ~w1361;
assign v604 = ~(w1362 | w1363);
assign w1364 = v604;
assign w1365 = w1355 & w1364;
assign v605 = ~(w1355 | w1364);
assign w1366 = v605;
assign v606 = ~(w1365 | w1366);
assign w1367 = v606;
assign w1368 = pi14 & pi36;
assign w1369 = pi16 & pi34;
assign v607 = ~(w1259 | w1369);
assign w1370 = v607;
assign w1371 = pi16 & pi35;
assign w1372 = w1257 & w1371;
assign v608 = ~(w1370 | w1372);
assign w1373 = v608;
assign w1374 = w1368 & ~w1373;
assign w1375 = ~w1368 & w1373;
assign v609 = ~(w1374 | w1375);
assign w1376 = v609;
assign w1377 = pi18 & pi32;
assign w1378 = pi82 & w1377;
assign v610 = ~(pi82 | w1377);
assign w1379 = v610;
assign v611 = ~(w1378 | w1379);
assign w1380 = v611;
assign w1381 = pi13 & pi37;
assign w1382 = pi17 & pi33;
assign w1383 = ~w1381 & w1382;
assign w1384 = w1381 & ~w1382;
assign v612 = ~(w1383 | w1384);
assign w1385 = v612;
assign w1386 = w1380 & w1385;
assign v613 = ~(w1380 | w1385);
assign w1387 = v613;
assign v614 = ~(w1386 | w1387);
assign w1388 = v614;
assign w1389 = w1376 & w1388;
assign v615 = ~(w1376 | w1388);
assign w1390 = v615;
assign v616 = ~(w1389 | w1390);
assign w1391 = v616;
assign w1392 = pi02 & pi48;
assign w1393 = pi03 & pi47;
assign v617 = ~(w1392 | w1393);
assign w1394 = v617;
assign w1395 = pi03 & pi48;
assign w1396 = w1107 & w1395;
assign v618 = ~(w1394 | w1396);
assign w1397 = v618;
assign w1398 = w1306 & ~w1397;
assign w1399 = ~w1306 & w1397;
assign v619 = ~(w1398 | w1399);
assign w1400 = v619;
assign w1401 = w1391 & ~w1400;
assign w1402 = ~w1391 & w1400;
assign v620 = ~(w1401 | w1402);
assign w1403 = v620;
assign w1404 = w1256 & ~w1258;
assign v621 = ~(w1260 | w1404);
assign w1405 = v621;
assign v622 = ~(w1266 | w1269);
assign w1406 = v622;
assign v623 = ~(w1267 | w1406);
assign w1407 = v623;
assign w1408 = ~w1405 & w1407;
assign w1409 = w1405 & ~w1407;
assign v624 = ~(w1408 | w1409);
assign w1410 = v624;
assign w1411 = w1122 & w1275;
assign v625 = ~(w1276 | w1411);
assign w1412 = v625;
assign w1413 = w1410 & ~w1412;
assign w1414 = ~w1410 & w1412;
assign v626 = ~(w1413 | w1414);
assign w1415 = v626;
assign w1416 = pi00 & pi50;
assign v627 = ~(w1289 | w1416);
assign w1417 = v627;
assign w1418 = w1289 & w1416;
assign v628 = ~(w1417 | w1418);
assign w1419 = v628;
assign w1420 = ~w1415 & w1419;
assign w1421 = w1415 & ~w1419;
assign v629 = ~(w1420 | w1421);
assign w1422 = v629;
assign w1423 = w1403 & ~w1422;
assign w1424 = ~w1403 & w1422;
assign v630 = ~(w1423 | w1424);
assign w1425 = v630;
assign w1426 = w1367 & ~w1425;
assign w1427 = ~w1367 & w1425;
assign v631 = ~(w1426 | w1427);
assign w1428 = v631;
assign w1429 = (~w1211 & ~w1213) | (~w1211 & w9248) | (~w1213 & w9248);
assign w1430 = w1214 & ~w1217;
assign v632 = ~(w1219 | w1430);
assign w1431 = v632;
assign w1432 = w1135 & ~w1204;
assign v633 = ~(w1206 | w1432);
assign w1433 = v633;
assign v634 = ~(w1431 | w1433);
assign w1434 = v634;
assign w1435 = w1431 & w1433;
assign v635 = ~(w1434 | w1435);
assign w1436 = v635;
assign w1437 = ~w1429 & w1436;
assign w1438 = w1429 & ~w1436;
assign v636 = ~(w1437 | w1438);
assign w1439 = v636;
assign w1440 = pi09 & pi41;
assign w1441 = pi10 & pi40;
assign v637 = ~(w1440 | w1441);
assign w1442 = v637;
assign w1443 = pi10 & pi41;
assign w1444 = w1135 & w1443;
assign v638 = ~(w1442 | w1444);
assign w1445 = v638;
assign w1446 = w1218 & ~w1445;
assign w1447 = ~w1218 & w1445;
assign v639 = ~(w1446 | w1447);
assign w1448 = v639;
assign w1449 = w1294 & ~w1448;
assign w1450 = ~w1294 & w1448;
assign v640 = ~(w1449 | w1450);
assign w1451 = v640;
assign w1452 = pi05 & pi45;
assign w1453 = pi06 & pi44;
assign w1454 = pi07 & pi43;
assign v641 = ~(w1453 | w1454);
assign w1455 = v641;
assign w1456 = pi07 & pi44;
assign w1457 = w1214 & w1456;
assign v642 = ~(w1455 | w1457);
assign w1458 = v642;
assign w1459 = w1452 & ~w1458;
assign w1460 = ~w1452 & w1458;
assign v643 = ~(w1459 | w1460);
assign w1461 = v643;
assign w1462 = w1451 & ~w1461;
assign w1463 = ~w1451 & w1461;
assign v644 = ~(w1462 | w1463);
assign w1464 = v644;
assign w1465 = w1439 & w1464;
assign v645 = ~(w1439 | w1464);
assign w1466 = v645;
assign v646 = ~(w1465 | w1466);
assign w1467 = v646;
assign w1468 = w1107 & ~w1293;
assign v647 = ~(w1295 | w1468);
assign w1469 = v647;
assign w1470 = ~w1305 & w1309;
assign v648 = ~(w1307 | w1470);
assign w1471 = v648;
assign v649 = ~(w1469 | w1471);
assign w1472 = v649;
assign w1473 = w1469 & w1471;
assign v650 = ~(w1472 | w1473);
assign w1474 = v650;
assign w1475 = (~w1301 & ~w1302) | (~w1301 & w9249) | (~w1302 & w9249);
assign w1476 = w1474 & w1475;
assign v651 = ~(w1474 | w1475);
assign w1477 = v651;
assign v652 = ~(w1476 | w1477);
assign w1478 = v652;
assign w1479 = w1467 & ~w1478;
assign w1480 = ~w1467 & w1478;
assign v653 = ~(w1479 | w1480);
assign w1481 = v653;
assign w1482 = w1428 & w1481;
assign v654 = ~(w1428 | w1481);
assign w1483 = v654;
assign v655 = ~(w1482 | w1483);
assign w1484 = v655;
assign w1485 = (~w1330 & ~w1326) | (~w1330 & w9250) | (~w1326 & w9250);
assign w1486 = ~w1484 & w1485;
assign w1487 = w1484 & ~w1485;
assign v656 = ~(w1486 | w1487);
assign w1488 = v656;
assign w1489 = w1354 & ~w1488;
assign w1490 = ~w1354 & w1488;
assign v657 = ~(w1489 | w1490);
assign w1491 = v657;
assign v658 = ~(w1345 | w1491);
assign w1492 = v658;
assign w1493 = w1345 & w1491;
assign v659 = ~(w1492 | w1493);
assign w1494 = v659;
assign v660 = ~(w1339 | w1342);
assign w1495 = v660;
assign w1496 = w1494 & w1495;
assign v661 = ~(w1494 | w1495);
assign w1497 = v661;
assign v662 = ~(w1496 | w1497);
assign w1498 = v662;
assign v663 = ~(w1492 | w1496);
assign w1499 = v663;
assign w1500 = pi14 & pi37;
assign w1501 = pi18 & pi33;
assign w1502 = pi19 & pi32;
assign w1503 = pi83 & w1502;
assign v664 = ~(pi83 | w1502);
assign w1504 = v664;
assign v665 = ~(w1503 | w1504);
assign w1505 = v665;
assign w1506 = w1501 & w1505;
assign v666 = ~(w1501 | w1505);
assign w1507 = v666;
assign v667 = ~(w1506 | w1507);
assign w1508 = v667;
assign w1509 = w1500 & w1508;
assign v668 = ~(w1500 | w1508);
assign w1510 = v668;
assign v669 = ~(w1509 | w1510);
assign w1511 = v669;
assign w1512 = pi15 & pi36;
assign w1513 = pi17 & pi34;
assign v670 = ~(w1371 | w1513);
assign w1514 = v670;
assign w1515 = pi17 & pi35;
assign w1516 = w1369 & w1515;
assign v671 = ~(w1514 | w1516);
assign w1517 = v671;
assign w1518 = w1512 & ~w1517;
assign w1519 = ~w1512 & w1517;
assign v672 = ~(w1518 | w1519);
assign w1520 = v672;
assign w1521 = w1511 & ~w1520;
assign w1522 = ~w1511 & w1520;
assign v673 = ~(w1521 | w1522);
assign w1523 = v673;
assign w1524 = pi00 & pi51;
assign w1525 = pi01 & pi50;
assign w1526 = pi02 & pi49;
assign v674 = ~(w1525 | w1526);
assign w1527 = v674;
assign w1528 = pi02 & pi50;
assign w1529 = w1306 & w1528;
assign v675 = ~(w1527 | w1529);
assign w1530 = v675;
assign w1531 = w1524 & ~w1530;
assign w1532 = ~w1524 & w1530;
assign v676 = ~(w1531 | w1532);
assign w1533 = v676;
assign w1534 = w1523 & ~w1533;
assign w1535 = ~w1523 & w1533;
assign v677 = ~(w1534 | w1535);
assign w1536 = v677;
assign w1537 = w1368 & ~w1370;
assign v678 = ~(w1372 | w1537);
assign w1538 = v678;
assign v679 = ~(w1378 | w1382);
assign w1539 = v679;
assign v680 = ~(w1379 | w1539);
assign w1540 = v680;
assign w1541 = ~w1538 & w1540;
assign w1542 = w1538 & ~w1540;
assign v681 = ~(w1541 | w1542);
assign w1543 = v681;
assign w1544 = w1381 & w1388;
assign v682 = ~(w1390 | w1544);
assign w1545 = v682;
assign w1546 = w1543 & ~w1545;
assign w1547 = ~w1543 & w1545;
assign v683 = ~(w1546 | w1547);
assign w1548 = v683;
assign w1549 = (~w1408 & w1412) | (~w1408 & w8590) | (w1412 & w8590);
assign w1550 = w1359 & ~w1549;
assign w1551 = ~w1359 & w1549;
assign v684 = ~(w1550 | w1551);
assign w1552 = v684;
assign w1553 = w1548 & w1552;
assign v685 = ~(w1548 | w1552);
assign w1554 = v685;
assign v686 = ~(w1553 | w1554);
assign w1555 = v686;
assign w1556 = w1536 & w1555;
assign v687 = ~(w1536 | w1555);
assign w1557 = v687;
assign v688 = ~(w1556 | w1557);
assign w1558 = v688;
assign v689 = ~(w1434 | w1437);
assign w1559 = v689;
assign w1560 = pi11 & pi40;
assign w1561 = pi13 & pi38;
assign v690 = ~(w1358 | w1561);
assign w1562 = v690;
assign w1563 = pi13 & pi39;
assign w1564 = w1356 & w1563;
assign v691 = ~(w1562 | w1564);
assign w1565 = v691;
assign w1566 = w1560 & w1565;
assign v692 = ~(w1560 | w1565);
assign w1567 = v692;
assign v693 = ~(w1566 | w1567);
assign w1568 = v693;
assign w1569 = w1443 & w1568;
assign v694 = ~(w1443 | w1568);
assign w1570 = v694;
assign v695 = ~(w1569 | w1570);
assign w1571 = v695;
assign w1572 = ~w1559 & w1571;
assign w1573 = w1559 & ~w1571;
assign v696 = ~(w1572 | w1573);
assign w1574 = v696;
assign v697 = ~(w1472 | w1476);
assign w1575 = v697;
assign w1576 = w1574 & ~w1575;
assign w1577 = ~w1574 & w1575;
assign v698 = ~(w1576 | w1577);
assign w1578 = v698;
assign w1579 = w1558 & w1578;
assign v699 = ~(w1558 | w1578);
assign w1580 = v699;
assign v700 = ~(w1579 | w1580);
assign w1581 = v700;
assign v701 = ~(w1449 | w1462);
assign w1582 = v701;
assign w1583 = w1452 & ~w1455;
assign v702 = ~(w1457 | w1583);
assign w1584 = v702;
assign w1585 = w1218 & ~w1442;
assign v703 = ~(w1444 | w1585);
assign w1586 = v703;
assign v704 = ~(w1584 | w1586);
assign w1587 = v704;
assign w1588 = w1584 & w1586;
assign v705 = ~(w1587 | w1588);
assign w1589 = v705;
assign w1590 = ~w1582 & w1589;
assign w1591 = w1582 & ~w1589;
assign v706 = ~(w1590 | w1591);
assign w1592 = v706;
assign w1593 = pi08 & pi43;
assign w1594 = pi09 & pi42;
assign v707 = ~(w1593 | w1594);
assign w1595 = v707;
assign w1596 = pi09 & pi43;
assign w1597 = w1218 & w1596;
assign v708 = ~(w1595 | w1597);
assign w1598 = v708;
assign w1599 = w1456 & ~w1598;
assign w1600 = ~w1456 & w1598;
assign v709 = ~(w1599 | w1600);
assign w1601 = v709;
assign w1602 = w1395 & ~w1601;
assign w1603 = ~w1395 & w1601;
assign v710 = ~(w1602 | w1603);
assign w1604 = v710;
assign w1605 = pi04 & pi47;
assign w1606 = pi05 & pi46;
assign w1607 = pi06 & pi45;
assign v711 = ~(w1606 | w1607);
assign w1608 = v711;
assign w1609 = pi06 & pi46;
assign w1610 = w1452 & w1609;
assign v712 = ~(w1608 | w1610);
assign w1611 = v712;
assign w1612 = w1605 & ~w1611;
assign w1613 = ~w1605 & w1611;
assign v713 = ~(w1612 | w1613);
assign w1614 = v713;
assign w1615 = w1604 & ~w1614;
assign w1616 = ~w1604 & w1614;
assign v714 = ~(w1615 | w1616);
assign w1617 = v714;
assign w1618 = w1592 & w1617;
assign v715 = ~(w1592 | w1617);
assign w1619 = v715;
assign v716 = ~(w1618 | w1619);
assign w1620 = v716;
assign w1621 = (~w1401 & w1422) | (~w1401 & w8694) | (w1422 & w8694);
assign w1622 = w1306 & ~w1394;
assign v717 = ~(w1396 | w1622);
assign w1623 = v717;
assign w1624 = (~w1623 & w1289) | (~w1623 & w9251) | (w1289 & w9251);
assign w1625 = (w1624 & w1415) | (w1624 & w8695) | (w1415 & w8695);
assign w1626 = ~w1418 & w1623;
assign v718 = ~(w1625 | w1626);
assign w1627 = v718;
assign w1628 = w1415 & w9252;
assign v719 = ~(w1627 | w1628);
assign w1629 = v719;
assign v720 = ~(w1621 | w1629);
assign w1630 = v720;
assign w1631 = w1621 & w1629;
assign v721 = ~(w1630 | w1631);
assign w1632 = v721;
assign w1633 = w1620 & ~w1632;
assign w1634 = ~w1620 & w1632;
assign v722 = ~(w1633 | w1634);
assign w1635 = v722;
assign w1636 = w1581 & ~w1635;
assign w1637 = ~w1581 & w1635;
assign v723 = ~(w1636 | w1637);
assign w1638 = v723;
assign v724 = ~(w1349 | w1352);
assign w1639 = v724;
assign v725 = ~(w1426 | w1482);
assign w1640 = v725;
assign v726 = ~(w1362 | w1365);
assign w1641 = v726;
assign v727 = ~(w1466 | w1479);
assign w1642 = v727;
assign w1643 = w1641 & w1642;
assign v728 = ~(w1641 | w1642);
assign w1644 = v728;
assign v729 = ~(w1643 | w1644);
assign w1645 = v729;
assign w1646 = w1640 & w1645;
assign v730 = ~(w1640 | w1645);
assign w1647 = v730;
assign v731 = ~(w1646 | w1647);
assign w1648 = v731;
assign w1649 = ~w1639 & w1648;
assign w1650 = w1639 & ~w1648;
assign v732 = ~(w1649 | w1650);
assign w1651 = v732;
assign w1652 = w1638 & w1651;
assign v733 = ~(w1638 | w1651);
assign w1653 = v733;
assign v734 = ~(w1652 | w1653);
assign w1654 = v734;
assign v735 = ~(w1487 | w1490);
assign w1655 = v735;
assign v736 = ~(w1654 | w1655);
assign w1656 = v736;
assign w1657 = w1654 & w1655;
assign v737 = ~(w1656 | w1657);
assign w1658 = v737;
assign w1659 = w1499 & ~w1658;
assign w1660 = ~w1499 & w1658;
assign v738 = ~(w1659 | w1660);
assign w1661 = v738;
assign w1662 = ~w1057 & w1195;
assign w1663 = w1341 & w1494;
assign w1664 = w1662 & w1663;
assign w1665 = w1658 & w1664;
assign w1666 = ~w1196 & w1665;
assign v739 = ~(w1193 | w1340);
assign w1667 = v739;
assign v740 = ~(w1339 | w1493);
assign w1668 = v740;
assign w1669 = ~w1667 & w1668;
assign v741 = ~(w1492 | w1657);
assign w1670 = v741;
assign w1671 = ~w1669 & w1670;
assign v742 = ~(w1656 | w1671);
assign w1672 = v742;
assign v743 = ~(w1666 | w1672);
assign w1673 = v743;
assign v744 = ~(w1649 | w1652);
assign w1674 = v744;
assign v745 = ~(w1643 | w1646);
assign w1675 = v745;
assign v746 = ~(w1579 | w1636);
assign w1676 = v746;
assign v747 = ~(w1572 | w1576);
assign w1677 = v747;
assign v748 = ~(w1619 | w1633);
assign w1678 = v748;
assign w1679 = ~w1677 & w1678;
assign w1680 = w1677 & ~w1678;
assign v749 = ~(w1679 | w1680);
assign w1681 = v749;
assign w1682 = ~w1676 & w1681;
assign w1683 = w1676 & ~w1681;
assign v750 = ~(w1682 | w1683);
assign w1684 = v750;
assign w1685 = ~w1675 & w1684;
assign w1686 = w1675 & ~w1684;
assign v751 = ~(w1685 | w1686);
assign w1687 = v751;
assign v752 = ~(w1587 | w1590);
assign w1688 = v752;
assign w1689 = pi11 & pi41;
assign w1690 = pi10 & pi42;
assign v753 = ~(w1689 | w1690);
assign w1691 = v753;
assign w1692 = pi11 & pi42;
assign w1693 = w1443 & w1692;
assign v754 = ~(w1691 | w1693);
assign w1694 = v754;
assign w1695 = pi12 & pi40;
assign w1696 = pi14 & pi38;
assign v755 = ~(w1563 | w1696);
assign w1697 = v755;
assign w1698 = pi14 & pi39;
assign w1699 = w1561 & w1698;
assign v756 = ~(w1697 | w1699);
assign w1700 = v756;
assign w1701 = w1695 & ~w1700;
assign w1702 = ~w1695 & w1700;
assign v757 = ~(w1701 | w1702);
assign w1703 = v757;
assign w1704 = w1694 & ~w1703;
assign w1705 = ~w1694 & w1703;
assign v758 = ~(w1704 | w1705);
assign w1706 = v758;
assign w1707 = ~w1688 & w1706;
assign w1708 = w1688 & ~w1706;
assign v759 = ~(w1707 | w1708);
assign w1709 = v759;
assign v760 = ~(w1625 | w1630);
assign w1710 = v760;
assign w1711 = w1709 & ~w1710;
assign w1712 = ~w1709 & w1710;
assign v761 = ~(w1711 | w1712);
assign w1713 = v761;
assign w1714 = pi15 & pi37;
assign w1715 = pi19 & pi33;
assign w1716 = pi20 & pi32;
assign w1717 = pi84 & w1716;
assign v762 = ~(pi84 | w1716);
assign w1718 = v762;
assign v763 = ~(w1717 | w1718);
assign w1719 = v763;
assign w1720 = w1715 & w1719;
assign v764 = ~(w1715 | w1719);
assign w1721 = v764;
assign v765 = ~(w1720 | w1721);
assign w1722 = v765;
assign w1723 = w1714 & w1722;
assign v766 = ~(w1714 | w1722);
assign w1724 = v766;
assign v767 = ~(w1723 | w1724);
assign w1725 = v767;
assign w1726 = pi16 & pi36;
assign w1727 = pi18 & pi34;
assign v768 = ~(w1515 | w1727);
assign w1728 = v768;
assign w1729 = pi18 & pi35;
assign w1730 = w1513 & w1729;
assign v769 = ~(w1728 | w1730);
assign w1731 = v769;
assign w1732 = w1726 & ~w1731;
assign w1733 = ~w1726 & w1731;
assign v770 = ~(w1732 | w1733);
assign w1734 = v770;
assign w1735 = w1725 & ~w1734;
assign w1736 = ~w1725 & w1734;
assign v771 = ~(w1735 | w1736);
assign w1737 = v771;
assign w1738 = pi00 & pi52;
assign w1739 = pi01 & pi51;
assign v772 = ~(w1528 | w1739);
assign w1740 = v772;
assign w1741 = pi02 & pi51;
assign w1742 = w1525 & w1741;
assign v773 = ~(w1740 | w1742);
assign w1743 = v773;
assign w1744 = w1738 & ~w1743;
assign w1745 = ~w1738 & w1743;
assign v774 = ~(w1744 | w1745);
assign w1746 = v774;
assign w1747 = w1737 & ~w1746;
assign w1748 = ~w1737 & w1746;
assign v775 = ~(w1747 | w1748);
assign w1749 = v775;
assign w1750 = (~w1509 & ~w1511) | (~w1509 & w8591) | (~w1511 & w8591);
assign w1751 = (~w1503 & ~w1505) | (~w1503 & w9253) | (~w1505 & w9253);
assign w1752 = w1512 & ~w1514;
assign v776 = ~(w1516 | w1752);
assign w1753 = v776;
assign v777 = ~(w1751 | w1753);
assign w1754 = v777;
assign w1755 = w1751 & w1753;
assign v778 = ~(w1754 | w1755);
assign w1756 = v778;
assign w1757 = ~w1750 & w1756;
assign w1758 = w1750 & ~w1756;
assign v779 = ~(w1757 | w1758);
assign w1759 = v779;
assign w1760 = (~w1541 & w1545) | (~w1541 & w8592) | (w1545 & w8592);
assign w1761 = (~w1564 & ~w1568) | (~w1564 & w8593) | (~w1568 & w8593);
assign w1762 = w1568 & w8594;
assign v780 = ~(w1761 | w1762);
assign w1763 = v780;
assign v781 = ~(w1566 | w1763);
assign w1764 = v781;
assign w1765 = w1760 & w1764;
assign v782 = ~(w1760 | w1764);
assign w1766 = v782;
assign v783 = ~(w1765 | w1766);
assign w1767 = v783;
assign w1768 = w1759 & ~w1767;
assign w1769 = ~w1759 & w1767;
assign v784 = ~(w1768 | w1769);
assign w1770 = v784;
assign w1771 = w1749 & ~w1770;
assign w1772 = ~w1749 & w1770;
assign v785 = ~(w1771 | w1772);
assign w1773 = v785;
assign w1774 = w1713 & w1773;
assign v786 = ~(w1713 | w1773);
assign w1775 = v786;
assign v787 = ~(w1774 | w1775);
assign w1776 = v787;
assign w1777 = (~w1534 & ~w1555) | (~w1534 & w8696) | (~w1555 & w8696);
assign w1778 = (~w1550 & ~w1552) | (~w1550 & w8697) | (~w1552 & w8697);
assign w1779 = w1524 & ~w1527;
assign v788 = ~(w1529 | w1779);
assign w1780 = v788;
assign v789 = ~(w1778 | w1780);
assign w1781 = v789;
assign w1782 = w1778 & w1780;
assign v790 = ~(w1781 | w1782);
assign w1783 = v790;
assign w1784 = ~w1777 & w1783;
assign w1785 = w1777 & ~w1783;
assign v791 = ~(w1784 | w1785);
assign w1786 = v791;
assign w1787 = pi03 & pi49;
assign w1788 = pi07 & pi45;
assign w1789 = pi08 & pi44;
assign v792 = ~(w1596 | w1789);
assign w1790 = v792;
assign w1791 = pi09 & pi44;
assign w1792 = w1593 & w1791;
assign v793 = ~(w1790 | w1792);
assign w1793 = v793;
assign w1794 = w1788 & ~w1793;
assign w1795 = ~w1788 & w1793;
assign v794 = ~(w1794 | w1795);
assign w1796 = v794;
assign w1797 = w1787 & ~w1796;
assign w1798 = ~w1787 & w1796;
assign v795 = ~(w1797 | w1798);
assign w1799 = v795;
assign w1800 = pi04 & pi48;
assign w1801 = pi05 & pi47;
assign v796 = ~(w1609 | w1801);
assign w1802 = v796;
assign w1803 = pi06 & pi47;
assign w1804 = w1606 & w1803;
assign v797 = ~(w1802 | w1804);
assign w1805 = v797;
assign w1806 = w1800 & ~w1805;
assign w1807 = ~w1800 & w1805;
assign v798 = ~(w1806 | w1807);
assign w1808 = v798;
assign w1809 = w1799 & ~w1808;
assign w1810 = ~w1799 & w1808;
assign v799 = ~(w1809 | w1810);
assign w1811 = v799;
assign v800 = ~(w1602 | w1615);
assign w1812 = v800;
assign w1813 = w1605 & ~w1608;
assign v801 = ~(w1610 | w1813);
assign w1814 = v801;
assign w1815 = w1456 & ~w1595;
assign v802 = ~(w1597 | w1815);
assign w1816 = v802;
assign v803 = ~(w1814 | w1816);
assign w1817 = v803;
assign w1818 = w1814 & w1816;
assign v804 = ~(w1817 | w1818);
assign w1819 = v804;
assign w1820 = ~w1812 & w1819;
assign w1821 = w1812 & ~w1819;
assign v805 = ~(w1820 | w1821);
assign w1822 = v805;
assign w1823 = w1811 & w1822;
assign v806 = ~(w1811 | w1822);
assign w1824 = v806;
assign v807 = ~(w1823 | w1824);
assign w1825 = v807;
assign v808 = ~(w1786 | w1825);
assign w1826 = v808;
assign w1827 = w1786 & w1825;
assign v809 = ~(w1826 | w1827);
assign w1828 = v809;
assign w1829 = w1776 & w1828;
assign v810 = ~(w1776 | w1828);
assign w1830 = v810;
assign v811 = ~(w1829 | w1830);
assign w1831 = v811;
assign w1832 = w1687 & w1831;
assign v812 = ~(w1687 | w1831);
assign w1833 = v812;
assign v813 = ~(w1832 | w1833);
assign w1834 = v813;
assign w1835 = ~w1674 & w1834;
assign w1836 = w1674 & ~w1834;
assign v814 = ~(w1835 | w1836);
assign w1837 = v814;
assign w1838 = ~w1673 & w1837;
assign w1839 = w1673 & ~w1837;
assign v815 = ~(w1838 | w1839);
assign w1840 = v815;
assign v816 = ~(w1685 | w1832);
assign w1841 = v816;
assign w1842 = pi16 & pi37;
assign w1843 = pi20 & pi33;
assign w1844 = pi21 & pi32;
assign w1845 = pi85 & w1844;
assign v817 = ~(pi85 | w1844);
assign w1846 = v817;
assign v818 = ~(w1845 | w1846);
assign w1847 = v818;
assign w1848 = w1843 & w1847;
assign v819 = ~(w1843 | w1847);
assign w1849 = v819;
assign v820 = ~(w1848 | w1849);
assign w1850 = v820;
assign w1851 = w1842 & w1850;
assign v821 = ~(w1842 | w1850);
assign w1852 = v821;
assign v822 = ~(w1851 | w1852);
assign w1853 = v822;
assign w1854 = pi17 & pi36;
assign w1855 = pi19 & pi34;
assign v823 = ~(w1729 | w1855);
assign w1856 = v823;
assign w1857 = pi19 & pi35;
assign w1858 = w1727 & w1857;
assign v824 = ~(w1856 | w1858);
assign w1859 = v824;
assign w1860 = w1854 & ~w1859;
assign w1861 = ~w1854 & w1859;
assign v825 = ~(w1860 | w1861);
assign w1862 = v825;
assign w1863 = w1853 & ~w1862;
assign w1864 = ~w1853 & w1862;
assign v826 = ~(w1863 | w1864);
assign w1865 = v826;
assign w1866 = pi00 & pi53;
assign w1867 = pi01 & pi52;
assign v827 = ~(w1866 | w1867);
assign w1868 = v827;
assign w1869 = pi01 & pi53;
assign w1870 = w1738 & w1869;
assign v828 = ~(w1868 | w1870);
assign w1871 = v828;
assign w1872 = w1871 & w9295;
assign w1873 = (w1750 & w9254) | (w1750 & w9255) | (w9254 & w9255);
assign v829 = ~(w1872 | w1873);
assign w1874 = v829;
assign w1875 = w1865 & w1874;
assign v830 = ~(w1865 | w1874);
assign w1876 = v830;
assign v831 = ~(w1875 | w1876);
assign w1877 = v831;
assign w1878 = (~w1693 & w1703) | (~w1693 & w8699) | (w1703 & w8699);
assign w1879 = w1695 & ~w1697;
assign v832 = ~(w1699 | w1879);
assign w1880 = v832;
assign v833 = ~(w1878 | w1880);
assign w1881 = v833;
assign w1882 = w1878 & w1880;
assign v834 = ~(w1881 | w1882);
assign w1883 = v834;
assign w1884 = (~w1723 & ~w1725) | (~w1723 & w8595) | (~w1725 & w8595);
assign w1885 = (~w1717 & ~w1719) | (~w1717 & w8596) | (~w1719 & w8596);
assign w1886 = w1726 & ~w1728;
assign v835 = ~(w1730 | w1886);
assign w1887 = v835;
assign v836 = ~(w1885 | w1887);
assign w1888 = v836;
assign w1889 = w1885 & w1887;
assign v837 = ~(w1888 | w1889);
assign w1890 = v837;
assign w1891 = w1884 & ~w1890;
assign w1892 = ~w1884 & w1890;
assign v838 = ~(w1891 | w1892);
assign w1893 = v838;
assign w1894 = w1762 & w1893;
assign v839 = ~(w1762 | w1893);
assign w1895 = v839;
assign v840 = ~(w1894 | w1895);
assign w1896 = v840;
assign w1897 = w1883 & ~w1896;
assign w1898 = ~w1883 & w1896;
assign v841 = ~(w1897 | w1898);
assign w1899 = v841;
assign w1900 = w1877 & ~w1899;
assign w1901 = ~w1877 & w1899;
assign v842 = ~(w1900 | w1901);
assign w1902 = v842;
assign v843 = ~(w1817 | w1820);
assign w1903 = v843;
assign w1904 = pi13 & pi40;
assign w1905 = pi15 & pi38;
assign v844 = ~(w1698 | w1905);
assign w1906 = v844;
assign w1907 = pi15 & pi39;
assign w1908 = w1696 & w1907;
assign v845 = ~(w1906 | w1908);
assign w1909 = v845;
assign w1910 = w1904 & ~w1909;
assign w1911 = ~w1904 & w1909;
assign v846 = ~(w1910 | w1911);
assign w1912 = v846;
assign w1913 = w1791 & ~w1912;
assign w1914 = ~w1791 & w1912;
assign v847 = ~(w1913 | w1914);
assign w1915 = v847;
assign w1916 = pi10 & pi43;
assign w1917 = pi12 & pi41;
assign v848 = ~(w1692 | w1917);
assign w1918 = v848;
assign w1919 = pi12 & pi42;
assign w1920 = w1689 & w1919;
assign v849 = ~(w1918 | w1920);
assign w1921 = v849;
assign w1922 = w1916 & ~w1921;
assign w1923 = ~w1916 & w1921;
assign v850 = ~(w1922 | w1923);
assign w1924 = v850;
assign w1925 = w1915 & ~w1924;
assign w1926 = ~w1915 & w1924;
assign v851 = ~(w1925 | w1926);
assign w1927 = v851;
assign w1928 = ~w1903 & w1927;
assign w1929 = w1903 & ~w1927;
assign v852 = ~(w1928 | w1929);
assign w1930 = v852;
assign w1931 = (w1930 & w1784) | (w1930 & w9256) | (w1784 & w9256);
assign w1932 = ~w1784 & w9257;
assign v853 = ~(w1931 | w1932);
assign w1933 = v853;
assign w1934 = w1902 & w1933;
assign v854 = ~(w1902 | w1933);
assign w1935 = v854;
assign v855 = ~(w1934 | w1935);
assign w1936 = v855;
assign w1937 = pi08 & pi45;
assign w1938 = pi07 & pi46;
assign v856 = ~(w1937 | w1938);
assign w1939 = v856;
assign w1940 = pi08 & pi46;
assign w1941 = w1788 & w1940;
assign v857 = ~(w1939 | w1941);
assign w1942 = v857;
assign w1943 = w1803 & ~w1942;
assign w1944 = ~w1803 & w1942;
assign v858 = ~(w1943 | w1944);
assign w1945 = v858;
assign w1946 = w1741 & ~w1945;
assign w1947 = ~w1741 & w1945;
assign v859 = ~(w1946 | w1947);
assign w1948 = v859;
assign w1949 = pi03 & pi50;
assign w1950 = pi04 & pi49;
assign w1951 = pi05 & pi48;
assign v860 = ~(w1950 | w1951);
assign w1952 = v860;
assign w1953 = pi05 & pi49;
assign w1954 = w1800 & w1953;
assign v861 = ~(w1952 | w1954);
assign w1955 = v861;
assign w1956 = w1949 & ~w1955;
assign w1957 = ~w1949 & w1955;
assign v862 = ~(w1956 | w1957);
assign w1958 = v862;
assign w1959 = w1948 & ~w1958;
assign w1960 = ~w1948 & w1958;
assign v863 = ~(w1959 | w1960);
assign w1961 = v863;
assign v864 = ~(w1797 | w1809);
assign w1962 = v864;
assign w1963 = w1800 & ~w1802;
assign v865 = ~(w1804 | w1963);
assign w1964 = v865;
assign w1965 = w1788 & ~w1790;
assign v866 = ~(w1792 | w1965);
assign w1966 = v866;
assign v867 = ~(w1964 | w1966);
assign w1967 = v867;
assign w1968 = w1964 & w1966;
assign v868 = ~(w1967 | w1968);
assign w1969 = v868;
assign w1970 = ~w1962 & w1969;
assign w1971 = w1962 & ~w1969;
assign v869 = ~(w1970 | w1971);
assign w1972 = v869;
assign w1973 = (~w1747 & w1770) | (~w1747 & w8700) | (w1770 & w8700);
assign w1974 = w1738 & ~w1740;
assign v870 = ~(w1742 | w1974);
assign w1975 = v870;
assign w1976 = ~w1769 & w8701;
assign w1977 = (w1975 & w1769) | (w1975 & w8702) | (w1769 & w8702);
assign v871 = ~(w1976 | w1977);
assign w1978 = v871;
assign w1979 = ~w1973 & w1978;
assign w1980 = w1973 & ~w1978;
assign v872 = ~(w1979 | w1980);
assign w1981 = v872;
assign w1982 = w1972 & w1981;
assign v873 = ~(w1972 | w1981);
assign w1983 = v873;
assign v874 = ~(w1982 | w1983);
assign w1984 = v874;
assign w1985 = w1961 & ~w1984;
assign w1986 = ~w1961 & w1984;
assign v875 = ~(w1985 | w1986);
assign w1987 = v875;
assign w1988 = w1936 & ~w1987;
assign w1989 = ~w1936 & w1987;
assign v876 = ~(w1988 | w1989);
assign w1990 = v876;
assign v877 = ~(w1679 | w1682);
assign w1991 = v877;
assign v878 = ~(w1707 | w1711);
assign w1992 = v878;
assign w1993 = (~w1823 & ~w1786) | (~w1823 & w9258) | (~w1786 & w9258);
assign v879 = ~(w1992 | w1993);
assign w1994 = v879;
assign w1995 = w1992 & w1993;
assign v880 = ~(w1994 | w1995);
assign w1996 = v880;
assign v881 = ~(w1774 | w1828);
assign w1997 = v881;
assign v882 = ~(w1775 | w1997);
assign w1998 = v882;
assign w1999 = w1996 & w1998;
assign v883 = ~(w1996 | w1998);
assign w2000 = v883;
assign v884 = ~(w1999 | w2000);
assign w2001 = v884;
assign w2002 = ~w1991 & w2001;
assign w2003 = w1991 & ~w2001;
assign v885 = ~(w2002 | w2003);
assign w2004 = v885;
assign w2005 = w1990 & w2004;
assign v886 = ~(w1990 | w2004);
assign w2006 = v886;
assign v887 = ~(w2005 | w2006);
assign w2007 = v887;
assign w2008 = w1841 & ~w2007;
assign w2009 = ~w1841 & w2007;
assign v888 = ~(w2008 | w2009);
assign w2010 = v888;
assign v889 = ~(w1835 | w1838);
assign w2011 = v889;
assign w2012 = w2010 & w2011;
assign v890 = ~(w2010 | w2011);
assign w2013 = v890;
assign v891 = ~(w2012 | w2013);
assign w2014 = v891;
assign w2015 = (~w2002 & ~w2004) | (~w2002 & w9259) | (~w2004 & w9259);
assign w2016 = (~w1934 & w1987) | (~w1934 & w9260) | (w1987 & w9260);
assign v892 = ~(w1928 | w1931);
assign w2017 = v892;
assign w2018 = (~w1983 & ~w1984) | (~w1983 & w9261) | (~w1984 & w9261);
assign w2019 = ~w2017 & w2018;
assign w2020 = w2017 & ~w2018;
assign v893 = ~(w2019 | w2020);
assign w2021 = v893;
assign w2022 = ~w2016 & w2021;
assign w2023 = w2016 & ~w2021;
assign v894 = ~(w2022 | w2023);
assign w2024 = v894;
assign w2025 = (~w1994 & ~w1998) | (~w1994 & w9262) | (~w1998 & w9262);
assign w2026 = pi00 & pi54;
assign w2027 = (~w1889 & w1735) | (~w1889 & w8597) | (w1735 & w8597);
assign w2028 = (w1735 & w8703) | (w1735 & w8704) | (w8703 & w8704);
assign w2029 = ~w1723 & w8598;
assign w2030 = w1889 & w2026;
assign w2031 = (~w2030 & w1735) | (~w2030 & w8599) | (w1735 & w8599);
assign w2032 = w1881 & w2031;
assign w2033 = ~w2028 & w2032;
assign v895 = ~(w1881 | w2031);
assign w2034 = v895;
assign v896 = ~(w1881 | w2026);
assign w2035 = v896;
assign w2036 = w2027 & w2035;
assign v897 = ~(w2034 | w2036);
assign w2037 = v897;
assign w2038 = ~w2033 & w2037;
assign w2039 = pi10 & pi44;
assign w2040 = pi14 & pi40;
assign w2041 = pi16 & pi38;
assign v898 = ~(w1907 | w2041);
assign w2042 = v898;
assign w2043 = pi16 & pi39;
assign w2044 = w1905 & w2043;
assign v899 = ~(w2042 | w2044);
assign w2045 = v899;
assign w2046 = w2040 & ~w2045;
assign w2047 = ~w2040 & w2045;
assign v900 = ~(w2046 | w2047);
assign w2048 = v900;
assign w2049 = w2039 & ~w2048;
assign w2050 = ~w2039 & w2048;
assign v901 = ~(w2049 | w2050);
assign w2051 = v901;
assign w2052 = pi11 & pi43;
assign w2053 = pi13 & pi41;
assign v902 = ~(w1919 | w2053);
assign w2054 = v902;
assign w2055 = pi13 & pi42;
assign w2056 = w1917 & w2055;
assign v903 = ~(w2054 | w2056);
assign w2057 = v903;
assign w2058 = w2052 & ~w2057;
assign w2059 = ~w2052 & w2057;
assign v904 = ~(w2058 | w2059);
assign w2060 = v904;
assign w2061 = w2051 & ~w2060;
assign w2062 = ~w2051 & w2060;
assign v905 = ~(w2061 | w2062);
assign w2063 = v905;
assign w2064 = ~w2038 & w2063;
assign w2065 = w2038 & ~w2063;
assign v906 = ~(w2064 | w2065);
assign w2066 = v906;
assign w2067 = pi17 & pi37;
assign w2068 = pi21 & pi33;
assign w2069 = pi22 & pi32;
assign w2070 = pi86 & w2069;
assign v907 = ~(pi86 | w2069);
assign w2071 = v907;
assign v908 = ~(w2070 | w2071);
assign w2072 = v908;
assign w2073 = w2068 & w2072;
assign v909 = ~(w2068 | w2072);
assign w2074 = v909;
assign v910 = ~(w2073 | w2074);
assign w2075 = v910;
assign w2076 = w2067 & w2075;
assign v911 = ~(w2067 | w2075);
assign w2077 = v911;
assign v912 = ~(w2076 | w2077);
assign w2078 = v912;
assign w2079 = pi18 & pi36;
assign w2080 = pi20 & pi34;
assign v913 = ~(w1857 | w2080);
assign w2081 = v913;
assign w2082 = pi20 & pi35;
assign w2083 = w1855 & w2082;
assign v914 = ~(w2081 | w2083);
assign w2084 = v914;
assign w2085 = w2079 & ~w2084;
assign w2086 = ~w2079 & w2084;
assign v915 = ~(w2085 | w2086);
assign w2087 = v915;
assign w2088 = w2078 & ~w2087;
assign w2089 = ~w2078 & w2087;
assign v916 = ~(w2088 | w2089);
assign w2090 = v916;
assign w2091 = (~w1913 & ~w1915) | (~w1913 & w8600) | (~w1915 & w8600);
assign w2092 = w1916 & ~w1918;
assign v917 = ~(w1920 | w2092);
assign w2093 = v917;
assign w2094 = w1904 & ~w1906;
assign v918 = ~(w1908 | w2094);
assign w2095 = v918;
assign w2096 = w2093 & w2095;
assign v919 = ~(w2093 | w2095);
assign w2097 = v919;
assign v920 = ~(w2096 | w2097);
assign w2098 = v920;
assign w2099 = w2091 & ~w2098;
assign w2100 = ~w2091 & w2098;
assign v921 = ~(w2099 | w2100);
assign w2101 = v921;
assign w2102 = (~w1851 & ~w1853) | (~w1851 & w8601) | (~w1853 & w8601);
assign v922 = ~(w1845 | w1848);
assign w2103 = v922;
assign w2104 = w1854 & ~w1856;
assign v923 = ~(w1858 | w2104);
assign w2105 = v923;
assign v924 = ~(w2103 | w2105);
assign w2106 = v924;
assign w2107 = w2103 & w2105;
assign v925 = ~(w2106 | w2107);
assign w2108 = v925;
assign w2109 = w2102 & ~w2108;
assign w2110 = ~w2102 & w2108;
assign v926 = ~(w2109 | w2110);
assign w2111 = v926;
assign v927 = ~(w2101 | w2111);
assign w2112 = v927;
assign w2113 = w2101 & w2111;
assign v928 = ~(w2112 | w2113);
assign w2114 = v928;
assign w2115 = w2090 & ~w2114;
assign w2116 = ~w2090 & w2114;
assign v929 = ~(w2115 | w2116);
assign w2117 = v929;
assign w2118 = w2066 & ~w2117;
assign w2119 = ~w2066 & w2117;
assign v930 = ~(w2118 | w2119);
assign w2120 = v930;
assign w2121 = pi09 & pi45;
assign v931 = ~(w1940 | w2121);
assign w2122 = v931;
assign w2123 = pi09 & pi46;
assign w2124 = w1937 & w2123;
assign v932 = ~(w2122 | w2124);
assign w2125 = v932;
assign v933 = ~(w1967 | w1970);
assign w2126 = v933;
assign w2127 = w2125 & ~w2126;
assign w2128 = ~w2125 & w2126;
assign v934 = ~(w2127 | w2128);
assign w2129 = v934;
assign w2130 = (w2129 & w1979) | (w2129 & w9263) | (w1979 & w9263);
assign w2131 = ~w1979 & w9264;
assign v935 = ~(w2130 | w2131);
assign w2132 = v935;
assign w2133 = w2120 & w2132;
assign v936 = ~(w2120 | w2132);
assign w2134 = v936;
assign v937 = ~(w2133 | w2134);
assign w2135 = v937;
assign w2136 = (~w1875 & w1899) | (~w1875 & w8705) | (w1899 & w8705);
assign v938 = ~(w1870 | w1872);
assign w2137 = v938;
assign w2138 = ~w2137 & w9296;
assign w2139 = (w1896 & w9265) | (w1896 & w9266) | (w9265 & w9266);
assign v939 = ~(w2138 | w2139);
assign w2140 = v939;
assign w2141 = ~w2136 & w2140;
assign w2142 = w2136 & ~w2140;
assign v940 = ~(w2141 | w2142);
assign w2143 = v940;
assign v941 = ~(w1946 | w1959);
assign w2144 = v941;
assign w2145 = w1949 & ~w1952;
assign v942 = ~(w1954 | w2145);
assign w2146 = v942;
assign w2147 = w1803 & ~w1939;
assign v943 = ~(w1941 | w2147);
assign w2148 = v943;
assign v944 = ~(w2146 | w2148);
assign w2149 = v944;
assign w2150 = w2146 & w2148;
assign v945 = ~(w2149 | w2150);
assign w2151 = v945;
assign w2152 = ~w2144 & w2151;
assign w2153 = w2144 & ~w2151;
assign v946 = ~(w2152 | w2153);
assign w2154 = v946;
assign w2155 = pi06 & pi48;
assign w2156 = pi07 & pi47;
assign v947 = ~(w2155 | w2156);
assign w2157 = v947;
assign w2158 = pi07 & pi48;
assign w2159 = w1803 & w2158;
assign v948 = ~(w2157 | w2159);
assign w2160 = v948;
assign w2161 = w1953 & ~w2160;
assign w2162 = ~w1953 & w2160;
assign v949 = ~(w2161 | w2162);
assign w2163 = v949;
assign w2164 = w1869 & ~w2163;
assign w2165 = ~w1869 & w2163;
assign v950 = ~(w2164 | w2165);
assign w2166 = v950;
assign w2167 = pi02 & pi52;
assign w2168 = pi03 & pi51;
assign w2169 = pi04 & pi50;
assign v951 = ~(w2168 | w2169);
assign w2170 = v951;
assign w2171 = pi04 & pi51;
assign w2172 = w1949 & w2171;
assign v952 = ~(w2170 | w2172);
assign w2173 = v952;
assign w2174 = w2167 & ~w2173;
assign w2175 = ~w2167 & w2173;
assign v953 = ~(w2174 | w2175);
assign w2176 = v953;
assign w2177 = w2166 & ~w2176;
assign w2178 = ~w2166 & w2176;
assign v954 = ~(w2177 | w2178);
assign w2179 = v954;
assign w2180 = w2154 & w2179;
assign v955 = ~(w2154 | w2179);
assign w2181 = v955;
assign v956 = ~(w2180 | w2181);
assign w2182 = v956;
assign w2183 = w2143 & ~w2182;
assign w2184 = ~w2143 & w2182;
assign v957 = ~(w2183 | w2184);
assign w2185 = v957;
assign w2186 = w2135 & ~w2185;
assign w2187 = ~w2135 & w2185;
assign v958 = ~(w2186 | w2187);
assign w2188 = v958;
assign w2189 = ~w2025 & w2188;
assign w2190 = w2025 & ~w2188;
assign v959 = ~(w2189 | w2190);
assign w2191 = v959;
assign w2192 = w2024 & w2191;
assign v960 = ~(w2024 | w2191);
assign w2193 = v960;
assign v961 = ~(w2192 | w2193);
assign w2194 = v961;
assign w2195 = ~w2015 & w2194;
assign w2196 = w2015 & ~w2194;
assign v962 = ~(w2195 | w2196);
assign w2197 = v962;
assign v963 = ~(w2008 | w2012);
assign w2198 = v963;
assign v964 = ~(w2197 | w2198);
assign w2199 = v964;
assign w2200 = ~w2008 & w2197;
assign v965 = ~(w1835 | w2009);
assign w2201 = v965;
assign w2202 = w2200 & ~w2201;
assign w2203 = w2197 & w9267;
assign w2204 = ~w1673 & w2203;
assign v966 = ~(w2202 | w2204);
assign w2205 = v966;
assign w2206 = ~w2199 & w2205;
assign w2207 = ~w2195 & w2205;
assign v967 = ~(w2149 | w2152);
assign w2208 = v967;
assign w2209 = pi08 & pi47;
assign w2210 = pi10 & pi45;
assign v968 = ~(w2123 | w2210);
assign w2211 = v968;
assign w2212 = pi10 & pi46;
assign w2213 = w2121 & w2212;
assign v969 = ~(w2211 | w2213);
assign w2214 = v969;
assign w2215 = w2209 & w2214;
assign v970 = ~(w2209 | w2214);
assign w2216 = v970;
assign v971 = ~(w2215 | w2216);
assign w2217 = v971;
assign w2218 = w2158 & w2217;
assign v972 = ~(w2158 | w2217);
assign w2219 = v972;
assign v973 = ~(w2218 | w2219);
assign w2220 = v973;
assign w2221 = ~w2208 & w2220;
assign w2222 = w2208 & ~w2220;
assign v974 = ~(w2221 | w2222);
assign w2223 = v974;
assign w2224 = ~w2138 & w2223;
assign w2225 = ~w2141 & w2224;
assign w2226 = w2136 & ~w2138;
assign v975 = ~(w2139 | w2223);
assign w2227 = v975;
assign w2228 = ~w2226 & w2227;
assign v976 = ~(w2225 | w2228);
assign w2229 = v976;
assign w2230 = pi18 & pi37;
assign w2231 = pi22 & pi33;
assign w2232 = pi23 & pi32;
assign w2233 = pi87 & w2232;
assign v977 = ~(pi87 | w2232);
assign w2234 = v977;
assign v978 = ~(w2233 | w2234);
assign w2235 = v978;
assign w2236 = w2231 & w2235;
assign v979 = ~(w2231 | w2235);
assign w2237 = v979;
assign v980 = ~(w2236 | w2237);
assign w2238 = v980;
assign w2239 = w2230 & w2238;
assign v981 = ~(w2230 | w2238);
assign w2240 = v981;
assign v982 = ~(w2239 | w2240);
assign w2241 = v982;
assign w2242 = pi19 & pi36;
assign w2243 = pi21 & pi34;
assign v983 = ~(w2082 | w2243);
assign w2244 = v983;
assign w2245 = pi21 & pi35;
assign w2246 = w2080 & w2245;
assign v984 = ~(w2244 | w2246);
assign w2247 = v984;
assign w2248 = w2242 & ~w2247;
assign w2249 = ~w2242 & w2247;
assign v985 = ~(w2248 | w2249);
assign w2250 = v985;
assign w2251 = w2241 & ~w2250;
assign w2252 = ~w2241 & w2250;
assign v986 = ~(w2251 | w2252);
assign w2253 = v986;
assign w2254 = (~w2049 & ~w2051) | (~w2049 & w8602) | (~w2051 & w8602);
assign w2255 = w2052 & ~w2054;
assign v987 = ~(w2056 | w2255);
assign w2256 = v987;
assign w2257 = w2040 & ~w2042;
assign v988 = ~(w2044 | w2257);
assign w2258 = v988;
assign v989 = ~(w2256 | w2258);
assign w2259 = v989;
assign w2260 = w2256 & w2258;
assign v990 = ~(w2259 | w2260);
assign w2261 = v990;
assign w2262 = w2254 & ~w2261;
assign w2263 = ~w2254 & w2261;
assign v991 = ~(w2262 | w2263);
assign w2264 = v991;
assign w2265 = w2124 & w2264;
assign v992 = ~(w2124 | w2264);
assign w2266 = v992;
assign v993 = ~(w2265 | w2266);
assign w2267 = v993;
assign w2268 = w2253 & w2267;
assign v994 = ~(w2253 | w2267);
assign w2269 = v994;
assign v995 = ~(w2268 | w2269);
assign w2270 = v995;
assign w2271 = pi11 & pi44;
assign w2272 = pi15 & pi40;
assign w2273 = pi17 & pi38;
assign v996 = ~(w2043 | w2273);
assign w2274 = v996;
assign w2275 = pi17 & pi39;
assign w2276 = w2041 & w2275;
assign v997 = ~(w2274 | w2276);
assign w2277 = v997;
assign w2278 = w2272 & ~w2277;
assign w2279 = ~w2272 & w2277;
assign v998 = ~(w2278 | w2279);
assign w2280 = v998;
assign w2281 = w2271 & ~w2280;
assign w2282 = ~w2271 & w2280;
assign v999 = ~(w2281 | w2282);
assign w2283 = v999;
assign w2284 = pi12 & pi43;
assign w2285 = pi14 & pi41;
assign v1000 = ~(w2055 | w2285);
assign w2286 = v1000;
assign w2287 = pi14 & pi42;
assign w2288 = w2053 & w2287;
assign v1001 = ~(w2286 | w2288);
assign w2289 = v1001;
assign w2290 = w2284 & ~w2289;
assign w2291 = ~w2284 & w2289;
assign v1002 = ~(w2290 | w2291);
assign w2292 = v1002;
assign w2293 = w2283 & ~w2292;
assign w2294 = ~w2283 & w2292;
assign v1003 = ~(w2293 | w2294);
assign w2295 = v1003;
assign w2296 = (~w2097 & w2091) | (~w2097 & w8707) | (w2091 & w8707);
assign w2297 = (~w2106 & w2102) | (~w2106 & w8708) | (w2102 & w8708);
assign v1004 = ~(w2296 | w2297);
assign w2298 = v1004;
assign w2299 = w2296 & w2297;
assign v1005 = ~(w2298 | w2299);
assign w2300 = v1005;
assign w2301 = (~w2076 & ~w2078) | (~w2076 & w8603) | (~w2078 & w8603);
assign v1006 = ~(w2070 | w2073);
assign w2302 = v1006;
assign w2303 = w2079 & ~w2081;
assign v1007 = ~(w2083 | w2303);
assign w2304 = v1007;
assign v1008 = ~(w2302 | w2304);
assign w2305 = v1008;
assign w2306 = w2302 & w2304;
assign v1009 = ~(w2305 | w2306);
assign w2307 = v1009;
assign w2308 = w2301 & ~w2307;
assign w2309 = ~w2301 & w2307;
assign v1010 = ~(w2308 | w2309);
assign w2310 = v1010;
assign w2311 = w2300 & w2310;
assign v1011 = ~(w2300 | w2310);
assign w2312 = v1011;
assign v1012 = ~(w2311 | w2312);
assign w2313 = v1012;
assign v1013 = ~(w2295 | w2313);
assign w2314 = v1013;
assign w2315 = w2295 & w2313;
assign v1014 = ~(w2314 | w2315);
assign w2316 = v1014;
assign w2317 = w2270 & ~w2316;
assign w2318 = ~w2270 & w2316;
assign v1015 = ~(w2317 | w2318);
assign w2319 = v1015;
assign v1016 = ~(w2229 | w2319);
assign w2320 = v1016;
assign w2321 = w2229 & w2319;
assign v1017 = ~(w2320 | w2321);
assign w2322 = v1017;
assign v1018 = ~(w2064 | w2118);
assign w2323 = v1018;
assign w2324 = (~w2112 & ~w2114) | (~w2112 & w8709) | (~w2114 & w8709);
assign w2325 = w1881 & ~w2031;
assign w2326 = w2027 & ~w2035;
assign v1019 = ~(w2325 | w2326);
assign w2327 = v1019;
assign w2328 = w2324 & ~w2327;
assign w2329 = ~w2324 & w2327;
assign v1020 = ~(w2328 | w2329);
assign w2330 = v1020;
assign w2331 = ~w2323 & w2330;
assign w2332 = w2323 & ~w2330;
assign v1021 = ~(w2331 | w2332);
assign w2333 = v1021;
assign w2334 = pi00 & pi55;
assign w2335 = pi05 & pi50;
assign w2336 = pi06 & pi49;
assign v1022 = ~(w2335 | w2336);
assign w2337 = v1022;
assign w2338 = pi06 & pi50;
assign w2339 = w1953 & w2338;
assign v1023 = ~(w2337 | w2339);
assign w2340 = v1023;
assign w2341 = w2171 & ~w2340;
assign w2342 = ~w2171 & w2340;
assign v1024 = ~(w2341 | w2342);
assign w2343 = v1024;
assign w2344 = w2334 & ~w2343;
assign w2345 = ~w2334 & w2343;
assign v1025 = ~(w2344 | w2345);
assign w2346 = v1025;
assign w2347 = pi01 & pi54;
assign w2348 = pi02 & pi53;
assign w2349 = pi03 & pi52;
assign v1026 = ~(w2348 | w2349);
assign w2350 = v1026;
assign w2351 = pi03 & pi53;
assign w2352 = w2167 & w2351;
assign v1027 = ~(w2350 | w2352);
assign w2353 = v1027;
assign w2354 = w2347 & ~w2353;
assign w2355 = ~w2347 & w2353;
assign v1028 = ~(w2354 | w2355);
assign w2356 = v1028;
assign w2357 = w2346 & ~w2356;
assign w2358 = ~w2346 & w2356;
assign v1029 = ~(w2357 | w2358);
assign w2359 = v1029;
assign v1030 = ~(w2164 | w2177);
assign w2360 = v1030;
assign w2361 = w2167 & ~w2170;
assign v1031 = ~(w2172 | w2361);
assign w2362 = v1031;
assign w2363 = w1953 & ~w2157;
assign v1032 = ~(w2159 | w2363);
assign w2364 = v1032;
assign v1033 = ~(w2362 | w2364);
assign w2365 = v1033;
assign w2366 = w2362 & w2364;
assign v1034 = ~(w2365 | w2366);
assign w2367 = v1034;
assign w2368 = ~w2360 & w2367;
assign w2369 = w2360 & ~w2367;
assign v1035 = ~(w2368 | w2369);
assign w2370 = v1035;
assign w2371 = w2359 & w2370;
assign v1036 = ~(w2359 | w2370);
assign w2372 = v1036;
assign v1037 = ~(w2371 | w2372);
assign w2373 = v1037;
assign w2374 = w2333 & ~w2373;
assign w2375 = ~w2333 & w2373;
assign v1038 = ~(w2374 | w2375);
assign w2376 = v1038;
assign w2377 = w2322 & ~w2376;
assign w2378 = ~w2322 & w2376;
assign v1039 = ~(w2377 | w2378);
assign w2379 = v1039;
assign v1040 = ~(w2019 | w2022);
assign w2380 = v1040;
assign v1041 = ~(w2133 | w2186);
assign w2381 = v1041;
assign v1042 = ~(w2127 | w2130);
assign w2382 = v1042;
assign v1043 = ~(w2181 | w2184);
assign w2383 = v1043;
assign w2384 = ~w2382 & w2383;
assign w2385 = w2382 & ~w2383;
assign v1044 = ~(w2384 | w2385);
assign w2386 = v1044;
assign w2387 = w2381 & ~w2386;
assign w2388 = ~w2381 & w2386;
assign v1045 = ~(w2387 | w2388);
assign w2389 = v1045;
assign w2390 = ~w2380 & w2389;
assign w2391 = w2380 & ~w2389;
assign v1046 = ~(w2390 | w2391);
assign w2392 = v1046;
assign w2393 = w2379 & w2392;
assign v1047 = ~(w2379 | w2392);
assign w2394 = v1047;
assign v1048 = ~(w2393 | w2394);
assign w2395 = v1048;
assign v1049 = ~(w2189 | w2192);
assign w2396 = v1049;
assign w2397 = w2395 & ~w2396;
assign w2398 = ~w2395 & w2396;
assign v1050 = ~(w2397 | w2398);
assign w2399 = v1050;
assign w2400 = w2207 & w2399;
assign v1051 = ~(w2207 | w2399);
assign w2401 = v1051;
assign v1052 = ~(w2400 | w2401);
assign w2402 = v1052;
assign v1053 = ~(w2195 | w2397);
assign w2403 = v1053;
assign w2404 = ~w2204 & w9268;
assign v1054 = ~(w2398 | w2404);
assign w2405 = v1054;
assign v1055 = ~(w2390 | w2393);
assign w2406 = v1055;
assign v1056 = ~(w2365 | w2368);
assign w2407 = v1056;
assign w2408 = pi08 & pi48;
assign w2409 = pi07 & pi49;
assign v1057 = ~(w2408 | w2409);
assign w2410 = v1057;
assign w2411 = pi08 & pi49;
assign w2412 = w2158 & w2411;
assign v1058 = ~(w2410 | w2412);
assign w2413 = v1058;
assign w2414 = pi09 & pi47;
assign w2415 = pi11 & pi45;
assign v1059 = ~(w2212 | w2415);
assign w2416 = v1059;
assign w2417 = pi11 & pi46;
assign w2418 = w2210 & w2417;
assign v1060 = ~(w2416 | w2418);
assign w2419 = v1060;
assign w2420 = w2414 & ~w2419;
assign w2421 = ~w2414 & w2419;
assign v1061 = ~(w2420 | w2421);
assign w2422 = v1061;
assign w2423 = w2413 & ~w2422;
assign w2424 = ~w2413 & w2422;
assign v1062 = ~(w2423 | w2424);
assign w2425 = v1062;
assign w2426 = ~w2407 & w2425;
assign w2427 = w2407 & ~w2425;
assign v1063 = ~(w2426 | w2427);
assign w2428 = v1063;
assign w2429 = ~w2328 & w2428;
assign w2430 = (w2429 & w2323) | (w2429 & w8710) | (w2323 & w8710);
assign w2431 = ~w2118 & w8711;
assign v1064 = ~(w2329 | w2428);
assign w2432 = v1064;
assign w2433 = ~w2431 & w2432;
assign v1065 = ~(w2430 | w2433);
assign w2434 = v1065;
assign w2435 = pi19 & pi37;
assign w2436 = pi23 & pi33;
assign w2437 = pi24 & pi32;
assign w2438 = pi88 & w2437;
assign v1066 = ~(pi88 | w2437);
assign w2439 = v1066;
assign v1067 = ~(w2438 | w2439);
assign w2440 = v1067;
assign w2441 = w2436 & w2440;
assign v1068 = ~(w2436 | w2440);
assign w2442 = v1068;
assign v1069 = ~(w2441 | w2442);
assign w2443 = v1069;
assign w2444 = w2435 & w2443;
assign v1070 = ~(w2435 | w2443);
assign w2445 = v1070;
assign v1071 = ~(w2444 | w2445);
assign w2446 = v1071;
assign w2447 = pi20 & pi36;
assign w2448 = pi22 & pi34;
assign v1072 = ~(w2245 | w2448);
assign w2449 = v1072;
assign w2450 = pi22 & pi35;
assign w2451 = w2243 & w2450;
assign v1073 = ~(w2449 | w2451);
assign w2452 = v1073;
assign w2453 = w2447 & ~w2452;
assign w2454 = ~w2447 & w2452;
assign v1074 = ~(w2453 | w2454);
assign w2455 = v1074;
assign w2456 = w2446 & ~w2455;
assign w2457 = ~w2446 & w2455;
assign v1075 = ~(w2456 | w2457);
assign w2458 = v1075;
assign w2459 = (~w2281 & ~w2283) | (~w2281 & w8604) | (~w2283 & w8604);
assign w2460 = w2284 & ~w2286;
assign v1076 = ~(w2288 | w2460);
assign w2461 = v1076;
assign w2462 = w2272 & ~w2274;
assign v1077 = ~(w2276 | w2462);
assign w2463 = v1077;
assign v1078 = ~(w2461 | w2463);
assign w2464 = v1078;
assign w2465 = w2461 & w2463;
assign v1079 = ~(w2464 | w2465);
assign w2466 = v1079;
assign w2467 = ~w2459 & w2466;
assign w2468 = w2459 & ~w2466;
assign v1080 = ~(w2467 | w2468);
assign w2469 = v1080;
assign v1081 = ~(w2213 | w2218);
assign w2470 = v1081;
assign w2471 = w2213 & w2218;
assign v1082 = ~(w2470 | w2471);
assign w2472 = v1082;
assign v1083 = ~(w2215 | w2472);
assign w2473 = v1083;
assign w2474 = w2469 & ~w2473;
assign w2475 = ~w2469 & w2473;
assign v1084 = ~(w2474 | w2475);
assign w2476 = v1084;
assign w2477 = w2458 & w2476;
assign v1085 = ~(w2458 | w2476);
assign w2478 = v1085;
assign v1086 = ~(w2477 | w2478);
assign w2479 = v1086;
assign w2480 = pi12 & pi44;
assign w2481 = pi16 & pi40;
assign w2482 = pi18 & pi38;
assign v1087 = ~(w2275 | w2482);
assign w2483 = v1087;
assign w2484 = pi18 & pi39;
assign w2485 = w2273 & w2484;
assign v1088 = ~(w2483 | w2485);
assign w2486 = v1088;
assign w2487 = w2481 & ~w2486;
assign w2488 = ~w2481 & w2486;
assign v1089 = ~(w2487 | w2488);
assign w2489 = v1089;
assign w2490 = w2480 & ~w2489;
assign w2491 = ~w2480 & w2489;
assign v1090 = ~(w2490 | w2491);
assign w2492 = v1090;
assign w2493 = pi13 & pi43;
assign w2494 = pi15 & pi41;
assign v1091 = ~(w2287 | w2494);
assign w2495 = v1091;
assign w2496 = pi15 & pi42;
assign w2497 = w2285 & w2496;
assign v1092 = ~(w2495 | w2497);
assign w2498 = v1092;
assign w2499 = w2493 & ~w2498;
assign w2500 = ~w2493 & w2498;
assign v1093 = ~(w2499 | w2500);
assign w2501 = v1093;
assign w2502 = w2492 & ~w2501;
assign w2503 = ~w2492 & w2501;
assign v1094 = ~(w2502 | w2503);
assign w2504 = v1094;
assign w2505 = (~w2239 & ~w2241) | (~w2239 & w8605) | (~w2241 & w8605);
assign v1095 = ~(w2233 | w2236);
assign w2506 = v1095;
assign w2507 = w2242 & ~w2244;
assign v1096 = ~(w2246 | w2507);
assign w2508 = v1096;
assign v1097 = ~(w2506 | w2508);
assign w2509 = v1097;
assign w2510 = w2506 & w2508;
assign v1098 = ~(w2509 | w2510);
assign w2511 = v1098;
assign w2512 = ~w2505 & w2511;
assign w2513 = w2505 & ~w2511;
assign v1099 = ~(w2512 | w2513);
assign w2514 = v1099;
assign w2515 = (~w2259 & w2254) | (~w2259 & w8712) | (w2254 & w8712);
assign w2516 = (~w2305 & w2301) | (~w2305 & w8713) | (w2301 & w8713);
assign v1100 = ~(w2515 | w2516);
assign w2517 = v1100;
assign w2518 = w2515 & w2516;
assign v1101 = ~(w2517 | w2518);
assign w2519 = v1101;
assign w2520 = w2514 & w2519;
assign v1102 = ~(w2514 | w2519);
assign w2521 = v1102;
assign v1103 = ~(w2520 | w2521);
assign w2522 = v1103;
assign v1104 = ~(w2504 | w2522);
assign w2523 = v1104;
assign w2524 = w2504 & w2522;
assign v1105 = ~(w2523 | w2524);
assign w2525 = v1105;
assign w2526 = w2479 & ~w2525;
assign w2527 = ~w2479 & w2525;
assign v1106 = ~(w2526 | w2527);
assign w2528 = v1106;
assign v1107 = ~(w2434 | w2528);
assign w2529 = v1107;
assign w2530 = w2434 & w2528;
assign v1108 = ~(w2529 | w2530);
assign w2531 = v1108;
assign v1109 = ~(w2265 | w2268);
assign w2532 = v1109;
assign v1110 = ~(w2298 | w2311);
assign w2533 = v1110;
assign v1111 = ~(w2532 | w2533);
assign w2534 = v1111;
assign w2535 = w2532 & w2533;
assign v1112 = ~(w2534 | w2535);
assign w2536 = v1112;
assign w2537 = w2270 & ~w2314;
assign v1113 = ~(w2315 | w2537);
assign w2538 = v1113;
assign w2539 = w2536 & ~w2538;
assign w2540 = ~w2536 & w2538;
assign v1114 = ~(w2539 | w2540);
assign w2541 = v1114;
assign v1115 = ~(w2344 | w2357);
assign w2542 = v1115;
assign w2543 = w2347 & ~w2350;
assign v1116 = ~(w2352 | w2543);
assign w2544 = v1116;
assign w2545 = w2171 & ~w2337;
assign v1117 = ~(w2339 | w2545);
assign w2546 = v1117;
assign v1118 = ~(w2544 | w2546);
assign w2547 = v1118;
assign w2548 = w2544 & w2546;
assign v1119 = ~(w2547 | w2548);
assign w2549 = v1119;
assign w2550 = ~w2542 & w2549;
assign w2551 = w2542 & ~w2549;
assign v1120 = ~(w2550 | w2551);
assign w2552 = v1120;
assign w2553 = pi00 & pi56;
assign w2554 = pi04 & pi52;
assign w2555 = pi05 & pi51;
assign v1121 = ~(w2338 | w2555);
assign w2556 = v1121;
assign w2557 = pi06 & pi51;
assign w2558 = w2335 & w2557;
assign v1122 = ~(w2556 | w2558);
assign w2559 = v1122;
assign w2560 = w2554 & ~w2559;
assign w2561 = ~w2554 & w2559;
assign v1123 = ~(w2560 | w2561);
assign w2562 = v1123;
assign w2563 = w2553 & ~w2562;
assign w2564 = ~w2553 & w2562;
assign v1124 = ~(w2563 | w2564);
assign w2565 = v1124;
assign w2566 = pi01 & pi55;
assign w2567 = pi02 & pi54;
assign v1125 = ~(w2351 | w2567);
assign w2568 = v1125;
assign w2569 = pi03 & pi54;
assign w2570 = w2348 & w2569;
assign v1126 = ~(w2568 | w2570);
assign w2571 = v1126;
assign w2572 = w2566 & ~w2571;
assign w2573 = ~w2566 & w2571;
assign v1127 = ~(w2572 | w2573);
assign w2574 = v1127;
assign w2575 = w2565 & ~w2574;
assign w2576 = ~w2565 & w2574;
assign v1128 = ~(w2575 | w2576);
assign w2577 = v1128;
assign w2578 = w2552 & w2577;
assign v1129 = ~(w2552 | w2577);
assign w2579 = v1129;
assign v1130 = ~(w2578 | w2579);
assign w2580 = v1130;
assign w2581 = w2541 & w2580;
assign v1131 = ~(w2541 | w2580);
assign w2582 = v1131;
assign v1132 = ~(w2581 | w2582);
assign w2583 = v1132;
assign w2584 = w2531 & w2583;
assign v1133 = ~(w2531 | w2583);
assign w2585 = v1133;
assign v1134 = ~(w2584 | w2585);
assign w2586 = v1134;
assign v1135 = ~(w2320 | w2377);
assign w2587 = v1135;
assign v1136 = ~(w2372 | w2375);
assign w2588 = v1136;
assign v1137 = ~(w2222 | w2225);
assign w2589 = v1137;
assign w2590 = w2588 & w2589;
assign v1138 = ~(w2588 | w2589);
assign w2591 = v1138;
assign v1139 = ~(w2590 | w2591);
assign w2592 = v1139;
assign w2593 = ~w2587 & w2592;
assign w2594 = w2587 & ~w2592;
assign v1140 = ~(w2593 | w2594);
assign w2595 = v1140;
assign v1141 = ~(w2384 | w2388);
assign w2596 = v1141;
assign w2597 = w2595 & ~w2596;
assign w2598 = ~w2595 & w2596;
assign v1142 = ~(w2597 | w2598);
assign w2599 = v1142;
assign w2600 = w2586 & w2599;
assign v1143 = ~(w2586 | w2599);
assign w2601 = v1143;
assign v1144 = ~(w2600 | w2601);
assign w2602 = v1144;
assign w2603 = ~w2406 & w2602;
assign w2604 = w2406 & ~w2602;
assign v1145 = ~(w2603 | w2604);
assign w2605 = v1145;
assign w2606 = w2405 & w2605;
assign v1146 = ~(w2405 | w2605);
assign w2607 = v1146;
assign v1147 = ~(w2606 | w2607);
assign w2608 = v1147;
assign v1148 = ~(w2597 | w2600);
assign w2609 = v1148;
assign v1149 = ~(w2474 | w2477);
assign w2610 = v1149;
assign v1150 = ~(w2517 | w2520);
assign w2611 = v1150;
assign v1151 = ~(w2610 | w2611);
assign w2612 = v1151;
assign w2613 = w2610 & w2611;
assign v1152 = ~(w2612 | w2613);
assign w2614 = v1152;
assign w2615 = w2479 & ~w2523;
assign v1153 = ~(w2524 | w2615);
assign w2616 = v1153;
assign w2617 = w2614 & ~w2616;
assign w2618 = ~w2614 & w2616;
assign v1154 = ~(w2617 | w2618);
assign w2619 = v1154;
assign w2620 = (~w2509 & w2505) | (~w2509 & w8714) | (w2505 & w8714);
assign w2621 = pi05 & pi52;
assign w2622 = pi04 & pi53;
assign v1155 = ~(w2621 | w2622);
assign w2623 = v1155;
assign w2624 = pi05 & pi53;
assign w2625 = w2554 & w2624;
assign v1156 = ~(w2623 | w2625);
assign w2626 = v1156;
assign w2627 = w2569 & ~w2626;
assign w2628 = ~w2569 & w2626;
assign v1157 = ~(w2627 | w2628);
assign w2629 = v1157;
assign v1158 = ~(w2620 | w2629);
assign w2630 = v1158;
assign w2631 = w2620 & w2629;
assign v1159 = ~(w2630 | w2631);
assign w2632 = v1159;
assign w2633 = pi00 & pi57;
assign w2634 = pi01 & pi56;
assign w2635 = pi02 & pi55;
assign v1160 = ~(w2634 | w2635);
assign w2636 = v1160;
assign w2637 = pi02 & pi56;
assign w2638 = w2566 & w2637;
assign v1161 = ~(w2636 | w2638);
assign w2639 = v1161;
assign w2640 = w2633 & ~w2639;
assign w2641 = ~w2633 & w2639;
assign v1162 = ~(w2640 | w2641);
assign w2642 = v1162;
assign w2643 = w2632 & ~w2642;
assign w2644 = ~w2632 & w2642;
assign v1163 = ~(w2643 | w2644);
assign w2645 = v1163;
assign v1164 = ~(w2563 | w2575);
assign w2646 = v1164;
assign w2647 = w2566 & ~w2568;
assign v1165 = ~(w2570 | w2647);
assign w2648 = v1165;
assign w2649 = w2554 & ~w2556;
assign v1166 = ~(w2558 | w2649);
assign w2650 = v1166;
assign v1167 = ~(w2648 | w2650);
assign w2651 = v1167;
assign w2652 = w2648 & w2650;
assign v1168 = ~(w2651 | w2652);
assign w2653 = v1168;
assign w2654 = ~w2646 & w2653;
assign w2655 = w2646 & ~w2653;
assign v1169 = ~(w2654 | w2655);
assign w2656 = v1169;
assign w2657 = w2645 & w2656;
assign v1170 = ~(w2645 | w2656);
assign w2658 = v1170;
assign v1171 = ~(w2657 | w2658);
assign w2659 = v1171;
assign w2660 = w2619 & ~w2659;
assign w2661 = ~w2619 & w2659;
assign v1172 = ~(w2660 | w2661);
assign w2662 = v1172;
assign v1173 = ~(w2534 | w2539);
assign w2663 = v1173;
assign v1174 = ~(w2547 | w2550);
assign w2664 = v1174;
assign w2665 = pi10 & pi47;
assign w2666 = pi12 & pi45;
assign v1175 = ~(w2417 | w2666);
assign w2667 = v1175;
assign w2668 = pi12 & pi46;
assign w2669 = w2415 & w2668;
assign v1176 = ~(w2667 | w2669);
assign w2670 = v1176;
assign w2671 = w2665 & ~w2670;
assign w2672 = ~w2665 & w2670;
assign v1177 = ~(w2671 | w2672);
assign w2673 = v1177;
assign w2674 = w2557 & ~w2673;
assign w2675 = ~w2557 & w2673;
assign v1178 = ~(w2674 | w2675);
assign w2676 = v1178;
assign w2677 = pi07 & pi50;
assign w2678 = pi09 & pi48;
assign v1179 = ~(w2411 | w2678);
assign w2679 = v1179;
assign w2680 = pi09 & pi49;
assign w2681 = w2408 & w2680;
assign v1180 = ~(w2679 | w2681);
assign w2682 = v1180;
assign w2683 = w2677 & ~w2682;
assign w2684 = ~w2677 & w2682;
assign v1181 = ~(w2683 | w2684);
assign w2685 = v1181;
assign w2686 = w2676 & ~w2685;
assign w2687 = ~w2676 & w2685;
assign v1182 = ~(w2686 | w2687);
assign w2688 = v1182;
assign w2689 = ~w2664 & w2688;
assign w2690 = w2664 & ~w2688;
assign v1183 = ~(w2689 | w2690);
assign w2691 = v1183;
assign w2692 = pi13 & pi44;
assign w2693 = pi17 & pi40;
assign w2694 = pi19 & pi38;
assign v1184 = ~(w2484 | w2694);
assign w2695 = v1184;
assign w2696 = pi19 & pi39;
assign w2697 = w2482 & w2696;
assign v1185 = ~(w2695 | w2697);
assign w2698 = v1185;
assign w2699 = w2693 & ~w2698;
assign w2700 = ~w2693 & w2698;
assign v1186 = ~(w2699 | w2700);
assign w2701 = v1186;
assign w2702 = w2692 & ~w2701;
assign w2703 = ~w2692 & w2701;
assign v1187 = ~(w2702 | w2703);
assign w2704 = v1187;
assign w2705 = pi14 & pi43;
assign w2706 = pi16 & pi41;
assign v1188 = ~(w2496 | w2706);
assign w2707 = v1188;
assign w2708 = pi16 & pi42;
assign w2709 = w2494 & w2708;
assign v1189 = ~(w2707 | w2709);
assign w2710 = v1189;
assign w2711 = w2705 & ~w2710;
assign w2712 = ~w2705 & w2710;
assign v1190 = ~(w2711 | w2712);
assign w2713 = v1190;
assign w2714 = w2704 & ~w2713;
assign w2715 = ~w2704 & w2713;
assign v1191 = ~(w2714 | w2715);
assign w2716 = v1191;
assign w2717 = ~w2464 & w2471;
assign w2718 = ~w2467 & w2717;
assign w2719 = (~w2465 & w2293) | (~w2465 & w8606) | (w2293 & w8606);
assign w2720 = (w2293 & w8715) | (w2293 & w8716) | (w8715 & w8716);
assign v1192 = ~(w2718 | w2720);
assign w2721 = v1192;
assign w2722 = (~w2444 & ~w2446) | (~w2444 & w8717) | (~w2446 & w8717);
assign v1193 = ~(w2438 | w2441);
assign w2723 = v1193;
assign w2724 = w2447 & ~w2449;
assign v1194 = ~(w2451 | w2724);
assign w2725 = v1194;
assign v1195 = ~(w2723 | w2725);
assign w2726 = v1195;
assign w2727 = w2723 & w2725;
assign v1196 = ~(w2726 | w2727);
assign w2728 = v1196;
assign w2729 = ~w2722 & w2728;
assign w2730 = w2722 & ~w2728;
assign v1197 = ~(w2729 | w2730);
assign w2731 = v1197;
assign w2732 = ~w2721 & w2731;
assign w2733 = w2721 & ~w2731;
assign v1198 = ~(w2732 | w2733);
assign w2734 = v1198;
assign w2735 = w2716 & w2734;
assign v1199 = ~(w2716 | w2734);
assign w2736 = v1199;
assign v1200 = ~(w2735 | w2736);
assign w2737 = v1200;
assign w2738 = pi20 & pi37;
assign w2739 = pi24 & pi33;
assign w2740 = pi25 & pi32;
assign w2741 = pi89 & w2740;
assign v1201 = ~(pi89 | w2740);
assign w2742 = v1201;
assign v1202 = ~(w2741 | w2742);
assign w2743 = v1202;
assign w2744 = w2739 & w2743;
assign v1203 = ~(w2739 | w2743);
assign w2745 = v1203;
assign v1204 = ~(w2744 | w2745);
assign w2746 = v1204;
assign w2747 = w2738 & w2746;
assign v1205 = ~(w2738 | w2746);
assign w2748 = v1205;
assign v1206 = ~(w2747 | w2748);
assign w2749 = v1206;
assign w2750 = pi21 & pi36;
assign w2751 = pi23 & pi34;
assign v1207 = ~(w2450 | w2751);
assign w2752 = v1207;
assign w2753 = pi23 & pi35;
assign w2754 = w2448 & w2753;
assign v1208 = ~(w2752 | w2754);
assign w2755 = v1208;
assign w2756 = w2750 & ~w2755;
assign w2757 = ~w2750 & w2755;
assign v1209 = ~(w2756 | w2757);
assign w2758 = v1209;
assign w2759 = w2749 & ~w2758;
assign w2760 = ~w2749 & w2758;
assign v1210 = ~(w2759 | w2760);
assign w2761 = v1210;
assign w2762 = (~w2412 & w2422) | (~w2412 & w8607) | (w2422 & w8607);
assign w2763 = w2414 & ~w2416;
assign v1211 = ~(w2418 | w2763);
assign w2764 = v1211;
assign v1212 = ~(w2764 | w2762);
assign w2765 = v1212;
assign w2766 = w2762 & w2764;
assign v1213 = ~(w2765 | w2766);
assign w2767 = v1213;
assign w2768 = w2761 & w2767;
assign v1214 = ~(w2761 | w2767);
assign w2769 = v1214;
assign v1215 = ~(w2768 | w2769);
assign w2770 = v1215;
assign w2771 = (~w2490 & ~w2492) | (~w2490 & w9125) | (~w2492 & w9125);
assign w2772 = w2493 & ~w2495;
assign v1216 = ~(w2497 | w2772);
assign w2773 = v1216;
assign w2774 = w2481 & ~w2483;
assign v1217 = ~(w2485 | w2774);
assign w2775 = v1217;
assign v1218 = ~(w2773 | w2775);
assign w2776 = v1218;
assign w2777 = w2773 & w2775;
assign v1219 = ~(w2776 | w2777);
assign w2778 = v1219;
assign w2779 = ~w2771 & w2778;
assign w2780 = w2771 & ~w2778;
assign v1220 = ~(w2779 | w2780);
assign w2781 = v1220;
assign w2782 = w2770 & ~w2781;
assign w2783 = ~w2770 & w2781;
assign v1221 = ~(w2782 | w2783);
assign w2784 = v1221;
assign w2785 = w2737 & w2784;
assign v1222 = ~(w2737 | w2784);
assign w2786 = v1222;
assign v1223 = ~(w2785 | w2786);
assign w2787 = v1223;
assign w2788 = w2691 & ~w2787;
assign w2789 = ~w2691 & w2787;
assign v1224 = ~(w2788 | w2789);
assign w2790 = v1224;
assign w2791 = w2663 & w2790;
assign v1225 = ~(w2663 | w2790);
assign w2792 = v1225;
assign v1226 = ~(w2791 | w2792);
assign w2793 = v1226;
assign v1227 = ~(w2662 | w2793);
assign w2794 = v1227;
assign w2795 = w2662 & w2793;
assign v1228 = ~(w2794 | w2795);
assign w2796 = v1228;
assign v1229 = ~(w2590 | w2593);
assign w2797 = v1229;
assign v1230 = ~(w2529 | w2584);
assign w2798 = v1230;
assign v1231 = ~(w2427 | w2430);
assign w2799 = v1231;
assign v1232 = ~(w2578 | w2581);
assign w2800 = v1232;
assign w2801 = w2799 & ~w2800;
assign w2802 = ~w2799 & w2800;
assign v1233 = ~(w2801 | w2802);
assign w2803 = v1233;
assign w2804 = ~w2798 & w2803;
assign w2805 = w2798 & ~w2803;
assign v1234 = ~(w2804 | w2805);
assign w2806 = v1234;
assign w2807 = ~w2797 & w2806;
assign w2808 = w2797 & ~w2806;
assign v1235 = ~(w2807 | w2808);
assign w2809 = v1235;
assign w2810 = w2796 & w2809;
assign v1236 = ~(w2796 | w2809);
assign w2811 = v1236;
assign v1237 = ~(w2810 | w2811);
assign w2812 = v1237;
assign w2813 = w2609 & ~w2812;
assign w2814 = ~w2609 & w2812;
assign v1238 = ~(w2813 | w2814);
assign w2815 = v1238;
assign v1239 = ~(w2603 | w2606);
assign w2816 = v1239;
assign w2817 = w2815 & ~w2816;
assign w2818 = ~w2815 & w2816;
assign v1240 = ~(w2817 | w2818);
assign w2819 = v1240;
assign v1241 = ~(w2807 | w2810);
assign w2820 = v1241;
assign w2821 = w2471 & w2719;
assign v1242 = ~(w2732 | w2821);
assign w2822 = v1242;
assign v1243 = ~(w2769 | w2782);
assign w2823 = v1243;
assign w2824 = ~w2822 & w2823;
assign w2825 = w2822 & ~w2823;
assign v1244 = ~(w2824 | w2825);
assign w2826 = v1244;
assign v1245 = ~(w2736 | w2784);
assign w2827 = v1245;
assign v1246 = ~(w2735 | w2827);
assign w2828 = v1246;
assign w2829 = w2826 & ~w2828;
assign w2830 = ~w2826 & w2828;
assign v1247 = ~(w2829 | w2830);
assign w2831 = v1247;
assign v1248 = ~(w2630 | w2643);
assign w2832 = v1248;
assign w2833 = w2633 & ~w2636;
assign v1249 = ~(w2638 | w2833);
assign w2834 = v1249;
assign w2835 = w2569 & ~w2623;
assign v1250 = ~(w2625 | w2835);
assign w2836 = v1250;
assign v1251 = ~(w2834 | w2836);
assign w2837 = v1251;
assign w2838 = w2834 & w2836;
assign v1252 = ~(w2837 | w2838);
assign w2839 = v1252;
assign w2840 = ~w2832 & w2839;
assign w2841 = w2832 & ~w2839;
assign v1253 = ~(w2840 | w2841);
assign w2842 = v1253;
assign v1254 = ~(w2776 | w2779);
assign w2843 = v1254;
assign w2844 = pi03 & pi55;
assign w2845 = pi04 & pi54;
assign v1255 = ~(w2844 | w2845);
assign w2846 = v1255;
assign w2847 = pi04 & pi55;
assign w2848 = w2569 & w2847;
assign v1256 = ~(w2846 | w2848);
assign w2849 = v1256;
assign w2850 = w2637 & ~w2849;
assign w2851 = ~w2637 & w2849;
assign v1257 = ~(w2850 | w2851);
assign w2852 = v1257;
assign v1258 = ~(w2843 | w2852);
assign w2853 = v1258;
assign w2854 = w2843 & w2852;
assign v1259 = ~(w2853 | w2854);
assign w2855 = v1259;
assign w2856 = pi00 & pi58;
assign w2857 = pi01 & pi57;
assign v1260 = ~(w2856 | w2857);
assign w2858 = v1260;
assign w2859 = pi01 & pi58;
assign w2860 = w2633 & w2859;
assign v1261 = ~(w2858 | w2860);
assign w2861 = v1261;
assign v1262 = ~(w2726 | w2729);
assign w2862 = v1262;
assign w2863 = w2861 & ~w2862;
assign w2864 = ~w2861 & w2862;
assign v1263 = ~(w2863 | w2864);
assign w2865 = v1263;
assign w2866 = w2855 & w2865;
assign v1264 = ~(w2855 | w2865);
assign w2867 = v1264;
assign v1265 = ~(w2866 | w2867);
assign w2868 = v1265;
assign w2869 = w2842 & w2868;
assign v1266 = ~(w2842 | w2868);
assign w2870 = v1266;
assign v1267 = ~(w2869 | w2870);
assign w2871 = v1267;
assign w2872 = w2831 & w2871;
assign v1268 = ~(w2831 | w2871);
assign w2873 = v1268;
assign v1269 = ~(w2872 | w2873);
assign w2874 = v1269;
assign v1270 = ~(w2612 | w2617);
assign w2875 = v1270;
assign w2876 = pi06 & pi52;
assign v1271 = ~(w2624 | w2876);
assign w2877 = v1271;
assign w2878 = pi06 & pi53;
assign w2879 = w2621 & w2878;
assign v1272 = ~(w2877 | w2879);
assign w2880 = v1272;
assign v1273 = ~(w2651 | w2654);
assign w2881 = v1273;
assign w2882 = w2880 & ~w2881;
assign w2883 = ~w2880 & w2881;
assign v1274 = ~(w2882 | w2883);
assign w2884 = v1274;
assign w2885 = pi07 & pi51;
assign w2886 = pi11 & pi47;
assign w2887 = pi13 & pi45;
assign v1275 = ~(w2668 | w2887);
assign w2888 = v1275;
assign w2889 = pi13 & pi46;
assign w2890 = w2666 & w2889;
assign v1276 = ~(w2888 | w2890);
assign w2891 = v1276;
assign w2892 = w2886 & ~w2891;
assign w2893 = ~w2886 & w2891;
assign v1277 = ~(w2892 | w2893);
assign w2894 = v1277;
assign w2895 = w2885 & ~w2894;
assign w2896 = ~w2885 & w2894;
assign v1278 = ~(w2895 | w2896);
assign w2897 = v1278;
assign w2898 = pi08 & pi50;
assign w2899 = pi10 & pi48;
assign v1279 = ~(w2680 | w2899);
assign w2900 = v1279;
assign w2901 = pi10 & pi49;
assign w2902 = w2678 & w2901;
assign v1280 = ~(w2900 | w2902);
assign w2903 = v1280;
assign w2904 = w2898 & ~w2903;
assign w2905 = ~w2898 & w2903;
assign v1281 = ~(w2904 | w2905);
assign w2906 = v1281;
assign w2907 = w2897 & ~w2906;
assign w2908 = ~w2897 & w2906;
assign v1282 = ~(w2907 | w2908);
assign w2909 = v1282;
assign w2910 = (~w2702 & ~w2704) | (~w2702 & w8718) | (~w2704 & w8718);
assign w2911 = w2705 & ~w2707;
assign v1283 = ~(w2709 | w2911);
assign w2912 = v1283;
assign w2913 = w2693 & ~w2695;
assign v1284 = ~(w2697 | w2913);
assign w2914 = v1284;
assign v1285 = ~(w2912 | w2914);
assign w2915 = v1285;
assign w2916 = w2912 & w2914;
assign v1286 = ~(w2915 | w2916);
assign w2917 = v1286;
assign w2918 = ~w2910 & w2917;
assign w2919 = w2910 & ~w2917;
assign v1287 = ~(w2918 | w2919);
assign w2920 = v1287;
assign w2921 = (~w2747 & ~w2749) | (~w2747 & w8608) | (~w2749 & w8608);
assign w2922 = (~w2741 & ~w2743) | (~w2741 & w8719) | (~w2743 & w8719);
assign w2923 = w2750 & ~w2752;
assign v1288 = ~(w2754 | w2923);
assign w2924 = v1288;
assign v1289 = ~(w2922 | w2924);
assign w2925 = v1289;
assign w2926 = w2922 & w2924;
assign v1290 = ~(w2925 | w2926);
assign w2927 = v1290;
assign w2928 = w2765 & ~w2927;
assign w2929 = ~w2765 & w2927;
assign v1291 = ~(w2928 | w2929);
assign w2930 = v1291;
assign w2931 = w2921 & ~w2930;
assign w2932 = ~w2921 & w2930;
assign v1292 = ~(w2931 | w2932);
assign w2933 = v1292;
assign w2934 = w2920 & ~w2933;
assign w2935 = ~w2920 & w2933;
assign v1293 = ~(w2934 | w2935);
assign w2936 = v1293;
assign v1294 = ~(w2909 | w2936);
assign w2937 = v1294;
assign w2938 = w2909 & w2936;
assign v1295 = ~(w2937 | w2938);
assign w2939 = v1295;
assign w2940 = pi14 & pi44;
assign w2941 = pi18 & pi40;
assign w2942 = pi20 & pi38;
assign v1296 = ~(w2696 | w2942);
assign w2943 = v1296;
assign w2944 = pi20 & pi39;
assign w2945 = w2694 & w2944;
assign v1297 = ~(w2943 | w2945);
assign w2946 = v1297;
assign w2947 = w2941 & ~w2946;
assign w2948 = ~w2941 & w2946;
assign v1298 = ~(w2947 | w2948);
assign w2949 = v1298;
assign w2950 = w2940 & ~w2949;
assign w2951 = ~w2940 & w2949;
assign v1299 = ~(w2950 | w2951);
assign w2952 = v1299;
assign w2953 = pi15 & pi43;
assign w2954 = pi17 & pi41;
assign v1300 = ~(w2708 | w2954);
assign w2955 = v1300;
assign w2956 = pi17 & pi42;
assign w2957 = w2706 & w2956;
assign v1301 = ~(w2955 | w2957);
assign w2958 = v1301;
assign w2959 = w2953 & ~w2958;
assign w2960 = ~w2953 & w2958;
assign v1302 = ~(w2959 | w2960);
assign w2961 = v1302;
assign w2962 = w2952 & ~w2961;
assign w2963 = ~w2952 & w2961;
assign v1303 = ~(w2962 | w2963);
assign w2964 = v1303;
assign w2965 = pi21 & pi37;
assign w2966 = pi25 & pi33;
assign w2967 = pi26 & pi32;
assign w2968 = pi90 & w2967;
assign v1304 = ~(pi90 | w2967);
assign w2969 = v1304;
assign v1305 = ~(w2968 | w2969);
assign w2970 = v1305;
assign w2971 = w2966 & w2970;
assign v1306 = ~(w2966 | w2970);
assign w2972 = v1306;
assign v1307 = ~(w2971 | w2972);
assign w2973 = v1307;
assign w2974 = w2965 & w2973;
assign v1308 = ~(w2965 | w2973);
assign w2975 = v1308;
assign v1309 = ~(w2974 | w2975);
assign w2976 = v1309;
assign w2977 = pi22 & pi36;
assign w2978 = pi24 & pi34;
assign v1310 = ~(w2753 | w2978);
assign w2979 = v1310;
assign w2980 = pi24 & pi35;
assign w2981 = w2751 & w2980;
assign v1311 = ~(w2979 | w2981);
assign w2982 = v1311;
assign w2983 = w2977 & ~w2982;
assign w2984 = ~w2977 & w2982;
assign v1312 = ~(w2983 | w2984);
assign w2985 = v1312;
assign w2986 = w2976 & ~w2985;
assign w2987 = ~w2976 & w2985;
assign v1313 = ~(w2986 | w2987);
assign w2988 = v1313;
assign w2989 = (~w2674 & ~w2676) | (~w2674 & w8720) | (~w2676 & w8720);
assign w2990 = w2677 & ~w2679;
assign v1314 = ~(w2681 | w2990);
assign w2991 = v1314;
assign w2992 = w2665 & ~w2667;
assign v1315 = ~(w2669 | w2992);
assign w2993 = v1315;
assign v1316 = ~(w2991 | w2993);
assign w2994 = v1316;
assign w2995 = w2991 & w2993;
assign v1317 = ~(w2994 | w2995);
assign w2996 = v1317;
assign w2997 = ~w2989 & w2996;
assign w2998 = w2989 & ~w2996;
assign v1318 = ~(w2997 | w2998);
assign w2999 = v1318;
assign w3000 = w2988 & w2999;
assign v1319 = ~(w2988 | w2999);
assign w3001 = v1319;
assign v1320 = ~(w3000 | w3001);
assign w3002 = v1320;
assign w3003 = w2964 & w3002;
assign v1321 = ~(w2964 | w3002);
assign w3004 = v1321;
assign v1322 = ~(w3003 | w3004);
assign w3005 = v1322;
assign w3006 = w2939 & ~w3005;
assign w3007 = ~w2939 & w3005;
assign v1323 = ~(w3006 | w3007);
assign w3008 = v1323;
assign w3009 = w2884 & ~w3008;
assign w3010 = ~w2884 & w3008;
assign v1324 = ~(w3009 | w3010);
assign w3011 = v1324;
assign w3012 = w2875 & w3011;
assign v1325 = ~(w2875 | w3011);
assign w3013 = v1325;
assign v1326 = ~(w3012 | w3013);
assign w3014 = v1326;
assign w3015 = w2874 & ~w3014;
assign w3016 = ~w2874 & w3014;
assign v1327 = ~(w3015 | w3016);
assign w3017 = v1327;
assign v1328 = ~(w2801 | w2804);
assign w3018 = v1328;
assign w3019 = ~w2787 & w2793;
assign v1329 = ~(w2794 | w3019);
assign w3020 = v1329;
assign v1330 = ~(w2658 | w2661);
assign w3021 = v1330;
assign v1331 = ~(w2663 | w2690);
assign w3022 = v1331;
assign v1332 = ~(w2689 | w3022);
assign w3023 = v1332;
assign w3024 = w3021 & ~w3023;
assign w3025 = ~w3021 & w3023;
assign v1333 = ~(w3024 | w3025);
assign w3026 = v1333;
assign w3027 = ~w3020 & w3026;
assign w3028 = w3020 & ~w3026;
assign v1334 = ~(w3027 | w3028);
assign w3029 = v1334;
assign w3030 = ~w3018 & w3029;
assign w3031 = w3018 & ~w3029;
assign v1335 = ~(w3030 | w3031);
assign w3032 = v1335;
assign w3033 = w3017 & w3032;
assign v1336 = ~(w3017 | w3032);
assign w3034 = v1336;
assign v1337 = ~(w3033 | w3034);
assign w3035 = v1337;
assign w3036 = ~w2820 & w3035;
assign w3037 = w2820 & ~w3035;
assign v1338 = ~(w3036 | w3037);
assign w3038 = v1338;
assign v1339 = ~(w2814 | w2817);
assign w3039 = v1339;
assign w3040 = w3038 & ~w3039;
assign w3041 = ~w3038 & w3039;
assign v1340 = ~(w3040 | w3041);
assign w3042 = v1340;
assign v1341 = ~(w3036 | w3040);
assign w3043 = v1341;
assign w3044 = (~w3030 & ~w3032) | (~w3030 & w8721) | (~w3032 & w8721);
assign w3045 = pi22 & pi37;
assign w3046 = pi26 & pi33;
assign w3047 = pi27 & pi32;
assign w3048 = pi91 & w3047;
assign v1342 = ~(pi91 | w3047);
assign w3049 = v1342;
assign v1343 = ~(w3048 | w3049);
assign w3050 = v1343;
assign w3051 = w3046 & w3050;
assign v1344 = ~(w3046 | w3050);
assign w3052 = v1344;
assign v1345 = ~(w3051 | w3052);
assign w3053 = v1345;
assign w3054 = w3045 & w3053;
assign v1346 = ~(w3045 | w3053);
assign w3055 = v1346;
assign v1347 = ~(w3054 | w3055);
assign w3056 = v1347;
assign w3057 = pi23 & pi36;
assign w3058 = pi25 & pi34;
assign v1348 = ~(w2980 | w3058);
assign w3059 = v1348;
assign w3060 = pi25 & pi35;
assign w3061 = w2978 & w3060;
assign v1349 = ~(w3059 | w3061);
assign w3062 = v1349;
assign w3063 = w3057 & ~w3062;
assign w3064 = ~w3057 & w3062;
assign v1350 = ~(w3063 | w3064);
assign w3065 = v1350;
assign w3066 = w3056 & ~w3065;
assign w3067 = ~w3056 & w3065;
assign v1351 = ~(w3066 | w3067);
assign w3068 = v1351;
assign w3069 = w2879 & w3068;
assign v1352 = ~(w2879 | w3068);
assign w3070 = v1352;
assign v1353 = ~(w3069 | w3070);
assign w3071 = v1353;
assign w3072 = pi15 & pi44;
assign w3073 = pi19 & pi40;
assign w3074 = pi21 & pi38;
assign v1354 = ~(w2944 | w3074);
assign w3075 = v1354;
assign w3076 = pi21 & pi39;
assign w3077 = w2942 & w3076;
assign v1355 = ~(w3075 | w3077);
assign w3078 = v1355;
assign w3079 = w3073 & ~w3078;
assign w3080 = ~w3073 & w3078;
assign v1356 = ~(w3079 | w3080);
assign w3081 = v1356;
assign w3082 = w3072 & ~w3081;
assign w3083 = ~w3072 & w3081;
assign v1357 = ~(w3082 | w3083);
assign w3084 = v1357;
assign w3085 = pi16 & pi43;
assign w3086 = pi18 & pi41;
assign v1358 = ~(w2956 | w3086);
assign w3087 = v1358;
assign w3088 = pi18 & pi42;
assign w3089 = w2954 & w3088;
assign v1359 = ~(w3087 | w3089);
assign w3090 = v1359;
assign w3091 = w3085 & ~w3090;
assign w3092 = ~w3085 & w3090;
assign v1360 = ~(w3091 | w3092);
assign w3093 = v1360;
assign w3094 = w3084 & ~w3093;
assign w3095 = ~w3084 & w3093;
assign v1361 = ~(w3094 | w3095);
assign w3096 = v1361;
assign w3097 = w3071 & w3096;
assign v1362 = ~(w3071 | w3096);
assign w3098 = v1362;
assign v1363 = ~(w3097 | w3098);
assign w3099 = v1363;
assign w3100 = (~w2895 & ~w2897) | (~w2895 & w8918) | (~w2897 & w8918);
assign w3101 = w2898 & ~w2900;
assign v1364 = ~(w2902 | w3101);
assign w3102 = v1364;
assign w3103 = w2886 & ~w2888;
assign v1365 = ~(w2890 | w3103);
assign w3104 = v1365;
assign v1366 = ~(w3102 | w3104);
assign w3105 = v1366;
assign w3106 = w3102 & w3104;
assign v1367 = ~(w3105 | w3106);
assign w3107 = v1367;
assign w3108 = ~w3100 & w3107;
assign w3109 = w3100 & ~w3107;
assign v1368 = ~(w3108 | w3109);
assign w3110 = v1368;
assign w3111 = (~w2950 & ~w2952) | (~w2950 & w8609) | (~w2952 & w8609);
assign w3112 = w2953 & ~w2955;
assign v1369 = ~(w2957 | w3112);
assign w3113 = v1369;
assign w3114 = w2941 & ~w2943;
assign v1370 = ~(w2945 | w3114);
assign w3115 = v1370;
assign v1371 = ~(w3113 | w3115);
assign w3116 = v1371;
assign w3117 = w3113 & w3115;
assign v1372 = ~(w3116 | w3117);
assign w3118 = v1372;
assign w3119 = ~w3111 & w3118;
assign w3120 = w3111 & ~w3118;
assign v1373 = ~(w3119 | w3120);
assign w3121 = v1373;
assign w3122 = (~w2974 & ~w2976) | (~w2974 & w8610) | (~w2976 & w8610);
assign w3123 = (~w2968 & ~w2970) | (~w2968 & w8919) | (~w2970 & w8919);
assign w3124 = w2977 & ~w2979;
assign v1374 = ~(w2981 | w3124);
assign w3125 = v1374;
assign v1375 = ~(w3123 | w3125);
assign w3126 = v1375;
assign w3127 = w3123 & w3125;
assign v1376 = ~(w3126 | w3127);
assign w3128 = v1376;
assign w3129 = ~w3122 & w3128;
assign w3130 = w3122 & ~w3128;
assign v1377 = ~(w3129 | w3130);
assign w3131 = v1377;
assign w3132 = w3121 & w3131;
assign v1378 = ~(w3121 | w3131);
assign w3133 = v1378;
assign v1379 = ~(w3132 | w3133);
assign w3134 = v1379;
assign w3135 = w3110 & w3134;
assign v1380 = ~(w3110 | w3134);
assign w3136 = v1380;
assign v1381 = ~(w3135 | w3136);
assign w3137 = v1381;
assign w3138 = pi08 & pi51;
assign w3139 = pi12 & pi47;
assign w3140 = pi14 & pi45;
assign v1382 = ~(w2889 | w3140);
assign w3141 = v1382;
assign w3142 = pi14 & pi46;
assign w3143 = w2887 & w3142;
assign v1383 = ~(w3141 | w3143);
assign w3144 = v1383;
assign w3145 = w3139 & ~w3144;
assign w3146 = ~w3139 & w3144;
assign v1384 = ~(w3145 | w3146);
assign w3147 = v1384;
assign w3148 = w3138 & ~w3147;
assign w3149 = ~w3138 & w3147;
assign v1385 = ~(w3148 | w3149);
assign w3150 = v1385;
assign w3151 = pi09 & pi50;
assign w3152 = pi11 & pi48;
assign v1386 = ~(w2901 | w3152);
assign w3153 = v1386;
assign w3154 = pi11 & pi49;
assign w3155 = w2899 & w3154;
assign v1387 = ~(w3153 | w3155);
assign w3156 = v1387;
assign w3157 = w3151 & ~w3156;
assign w3158 = ~w3151 & w3156;
assign v1388 = ~(w3157 | w3158);
assign w3159 = v1388;
assign w3160 = w3150 & ~w3159;
assign w3161 = ~w3150 & w3159;
assign v1389 = ~(w3160 | w3161);
assign w3162 = v1389;
assign w3163 = w3137 & w3162;
assign v1390 = ~(w3137 | w3162);
assign w3164 = v1390;
assign v1391 = ~(w3163 | w3164);
assign w3165 = v1391;
assign w3166 = w3099 & w3165;
assign v1392 = ~(w3099 | w3165);
assign w3167 = v1392;
assign v1393 = ~(w3166 | w3167);
assign w3168 = v1393;
assign w3169 = (~w2824 & w2828) | (~w2824 & w8722) | (w2828 & w8722);
assign v1394 = ~(w2837 | w2840);
assign w3170 = v1394;
assign w3171 = pi05 & pi54;
assign w3172 = pi07 & pi52;
assign v1395 = ~(w2878 | w3172);
assign w3173 = v1395;
assign w3174 = pi07 & pi53;
assign w3175 = w2876 & w3174;
assign v1396 = ~(w3173 | w3175);
assign w3176 = v1396;
assign w3177 = w3171 & w3176;
assign v1397 = ~(w3171 | w3176);
assign w3178 = v1397;
assign v1398 = ~(w3177 | w3178);
assign w3179 = v1398;
assign w3180 = w2847 & w3179;
assign v1399 = ~(w2847 | w3179);
assign w3181 = v1399;
assign v1400 = ~(w3180 | w3181);
assign w3182 = v1400;
assign w3183 = ~w3170 & w3182;
assign w3184 = w3170 & ~w3182;
assign v1401 = ~(w3183 | w3184);
assign w3185 = v1401;
assign w3186 = ~w3169 & w3185;
assign w3187 = w3169 & ~w3185;
assign v1402 = ~(w3186 | w3187);
assign w3188 = v1402;
assign w3189 = w3168 & w3188;
assign v1403 = ~(w3168 | w3188);
assign w3190 = v1403;
assign v1404 = ~(w3189 | w3190);
assign w3191 = v1404;
assign v1405 = ~(w2853 | w2866);
assign w3192 = v1405;
assign v1406 = ~(w2860 | w2863);
assign w3193 = v1406;
assign w3194 = w2637 & ~w2846;
assign v1407 = ~(w2848 | w3194);
assign w3195 = v1407;
assign v1408 = ~(w3193 | w3195);
assign w3196 = v1408;
assign w3197 = w3193 & w3195;
assign v1409 = ~(w3196 | w3197);
assign w3198 = v1409;
assign w3199 = ~w3192 & w3198;
assign w3200 = w3192 & ~w3198;
assign v1410 = ~(w3199 | w3200);
assign w3201 = v1410;
assign w3202 = (~w2994 & w2989) | (~w2994 & w9126) | (w2989 & w9126);
assign w3203 = pi02 & pi57;
assign w3204 = pi03 & pi56;
assign v1411 = ~(w3203 | w3204);
assign w3205 = v1411;
assign w3206 = pi03 & pi57;
assign w3207 = w2637 & w3206;
assign v1412 = ~(w3205 | w3207);
assign w3208 = v1412;
assign w3209 = w2859 & ~w3208;
assign w3210 = ~w2859 & w3208;
assign v1413 = ~(w3209 | w3210);
assign w3211 = v1413;
assign w3212 = w3202 & w3211;
assign v1414 = ~(w3202 | w3211);
assign w3213 = v1414;
assign v1415 = ~(w3212 | w3213);
assign w3214 = v1415;
assign w3215 = (~w2915 & w2910) | (~w2915 & w9127) | (w2910 & w9127);
assign w3216 = pi00 & pi59;
assign w3217 = w3216 & w9297;
assign w3218 = (w2921 & w8920) | (w2921 & w8921) | (w8920 & w8921);
assign v1416 = ~(w3217 | w3218);
assign w3219 = v1416;
assign w3220 = ~w3215 & w3219;
assign w3221 = w3215 & ~w3219;
assign v1417 = ~(w3220 | w3221);
assign w3222 = v1417;
assign w3223 = w3214 & ~w3222;
assign w3224 = ~w3214 & w3222;
assign v1418 = ~(w3223 | w3224);
assign w3225 = v1418;
assign w3226 = w3201 & ~w3225;
assign w3227 = ~w3201 & w3225;
assign v1419 = ~(w3226 | w3227);
assign w3228 = v1419;
assign v1420 = ~(w2937 | w3006);
assign w3229 = v1420;
assign w3230 = w2765 & w2933;
assign v1421 = ~(w2934 | w3230);
assign w3231 = v1421;
assign v1422 = ~(w3000 | w3003);
assign w3232 = v1422;
assign v1423 = ~(w3231 | w3232);
assign w3233 = v1423;
assign w3234 = w3231 & w3232;
assign v1424 = ~(w3233 | w3234);
assign w3235 = v1424;
assign w3236 = w3229 & w3235;
assign v1425 = ~(w3229 | w3235);
assign w3237 = v1425;
assign v1426 = ~(w3236 | w3237);
assign w3238 = v1426;
assign w3239 = w3228 & ~w3238;
assign w3240 = ~w3228 & w3238;
assign v1427 = ~(w3239 | w3240);
assign w3241 = v1427;
assign w3242 = w3191 & ~w3241;
assign w3243 = ~w3191 & w3241;
assign v1428 = ~(w3242 | w3243);
assign w3244 = v1428;
assign w3245 = (~w3024 & w3020) | (~w3024 & w8724) | (w3020 & w8724);
assign w3246 = ~w3008 & w3014;
assign v1429 = ~(w3015 | w3246);
assign w3247 = v1429;
assign v1430 = ~(w2869 | w2872);
assign w3248 = v1430;
assign w3249 = w2875 & ~w2882;
assign v1431 = ~(w2883 | w3249);
assign w3250 = v1431;
assign w3251 = ~w3248 & w3250;
assign w3252 = w3248 & ~w3250;
assign v1432 = ~(w3251 | w3252);
assign w3253 = v1432;
assign w3254 = ~w3247 & w3253;
assign w3255 = w3247 & ~w3253;
assign v1433 = ~(w3254 | w3255);
assign w3256 = v1433;
assign w3257 = ~w3245 & w3256;
assign w3258 = w3245 & ~w3256;
assign v1434 = ~(w3257 | w3258);
assign w3259 = v1434;
assign w3260 = w3244 & w3259;
assign v1435 = ~(w3244 | w3259);
assign w3261 = v1435;
assign v1436 = ~(w3260 | w3261);
assign w3262 = v1436;
assign w3263 = ~w3044 & w3262;
assign w3264 = w3044 & ~w3262;
assign v1437 = ~(w3263 | w3264);
assign w3265 = v1437;
assign w3266 = w3043 & w3265;
assign v1438 = ~(w3043 | w3265);
assign w3267 = v1438;
assign v1439 = ~(w3266 | w3267);
assign w3268 = v1439;
assign v1440 = ~(w2603 | w2814);
assign w3269 = v1440;
assign v1441 = ~(w2813 | w3037);
assign w3270 = v1441;
assign w3271 = ~w3269 & w3270;
assign w3272 = (~w3264 & w3271) | (~w3264 & w8725) | (w3271 & w8725);
assign w3273 = w2605 & w2815;
assign w3274 = w3038 & w3265;
assign w3275 = w3273 & w3274;
assign w3276 = w2405 & w3275;
assign v1442 = ~(w3272 | w3276);
assign w3277 = v1442;
assign v1443 = ~(w3257 | w3260);
assign w3278 = v1443;
assign w3279 = (~w3105 & w3100) | (~w3105 & w9128) | (w3100 & w9128);
assign w3280 = pi01 & pi59;
assign w3281 = pi02 & pi58;
assign v1444 = ~(w3206 | w3281);
assign w3282 = v1444;
assign w3283 = pi03 & pi58;
assign w3284 = w3203 & w3283;
assign v1445 = ~(w3282 | w3284);
assign w3285 = v1445;
assign w3286 = w3280 & ~w3285;
assign w3287 = ~w3280 & w3285;
assign v1446 = ~(w3286 | w3287);
assign w3288 = v1446;
assign w3289 = w3279 & w3288;
assign v1447 = ~(w3279 | w3288);
assign w3290 = v1447;
assign v1448 = ~(w3289 | w3290);
assign w3291 = v1448;
assign w3292 = (~w3116 & w3111) | (~w3116 & w9129) | (w3111 & w9129);
assign w3293 = pi00 & pi60;
assign w3294 = (~w3122 & w8922) | (~w3122 & w8923) | (w8922 & w8923);
assign w3295 = (w3122 & w8924) | (w3122 & w8925) | (w8924 & w8925);
assign v1449 = ~(w3294 | w3295);
assign w3296 = v1449;
assign w3297 = ~w3292 & w3296;
assign w3298 = w3292 & ~w3296;
assign v1450 = ~(w3297 | w3298);
assign w3299 = v1450;
assign w3300 = w3291 & ~w3299;
assign w3301 = ~w3291 & w3299;
assign v1451 = ~(w3300 | w3301);
assign w3302 = v1451;
assign w3303 = (~w3212 & w3222) | (~w3212 & w9130) | (w3222 & w9130);
assign w3304 = (~w3217 & ~w3219) | (~w3217 & w9131) | (~w3219 & w9131);
assign w3305 = w2859 & ~w3205;
assign v1452 = ~(w3207 | w3305);
assign w3306 = v1452;
assign v1453 = ~(w3304 | w3306);
assign w3307 = v1453;
assign w3308 = w3304 & w3306;
assign v1454 = ~(w3307 | w3308);
assign w3309 = v1454;
assign w3310 = w3303 & w3309;
assign v1455 = ~(w3303 | w3309);
assign w3311 = v1455;
assign v1456 = ~(w3310 | w3311);
assign w3312 = v1456;
assign w3313 = (~w3163 & ~w3165) | (~w3163 & w8726) | (~w3165 & w8726);
assign v1457 = ~(w3069 | w3097);
assign w3314 = v1457;
assign w3315 = (~w3132 & ~w3134) | (~w3132 & w9132) | (~w3134 & w9132);
assign v1458 = ~(w3314 | w3315);
assign w3316 = v1458;
assign w3317 = w3314 & w3315;
assign v1459 = ~(w3316 | w3317);
assign w3318 = v1459;
assign w3319 = (w3165 & w9133) | (w3165 & w9134) | (w9133 & w9134);
assign w3320 = ~w3318 & w3313;
assign v1460 = ~(w3319 | w3320);
assign w3321 = v1460;
assign w3322 = w3312 & w3321;
assign v1461 = ~(w3312 | w3321);
assign w3323 = v1461;
assign v1462 = ~(w3322 | w3323);
assign w3324 = v1462;
assign w3325 = ~w3302 & w3324;
assign w3326 = w3302 & ~w3324;
assign v1463 = ~(w3325 | w3326);
assign w3327 = v1463;
assign w3328 = pi16 & pi44;
assign w3329 = pi20 & pi40;
assign w3330 = pi22 & pi38;
assign v1464 = ~(w3076 | w3330);
assign w3331 = v1464;
assign w3332 = pi22 & pi39;
assign w3333 = w3074 & w3332;
assign v1465 = ~(w3331 | w3333);
assign w3334 = v1465;
assign w3335 = w3329 & ~w3334;
assign w3336 = ~w3329 & w3334;
assign v1466 = ~(w3335 | w3336);
assign w3337 = v1466;
assign w3338 = w3328 & ~w3337;
assign w3339 = ~w3328 & w3337;
assign v1467 = ~(w3338 | w3339);
assign w3340 = v1467;
assign w3341 = pi17 & pi43;
assign w3342 = pi19 & pi41;
assign v1468 = ~(w3088 | w3342);
assign w3343 = v1468;
assign w3344 = pi19 & pi42;
assign w3345 = w3086 & w3344;
assign v1469 = ~(w3343 | w3345);
assign w3346 = v1469;
assign w3347 = w3341 & ~w3346;
assign w3348 = ~w3341 & w3346;
assign v1470 = ~(w3347 | w3348);
assign w3349 = v1470;
assign w3350 = w3340 & ~w3349;
assign w3351 = ~w3340 & w3349;
assign v1471 = ~(w3350 | w3351);
assign w3352 = v1471;
assign w3353 = pi23 & pi37;
assign w3354 = pi27 & pi33;
assign w3355 = pi28 & pi32;
assign w3356 = pi92 & w3355;
assign v1472 = ~(pi92 | w3355);
assign w3357 = v1472;
assign v1473 = ~(w3356 | w3357);
assign w3358 = v1473;
assign w3359 = w3354 & w3358;
assign v1474 = ~(w3354 | w3358);
assign w3360 = v1474;
assign v1475 = ~(w3359 | w3360);
assign w3361 = v1475;
assign w3362 = w3353 & w3361;
assign v1476 = ~(w3353 | w3361);
assign w3363 = v1476;
assign v1477 = ~(w3362 | w3363);
assign w3364 = v1477;
assign w3365 = pi24 & pi36;
assign w3366 = pi26 & pi34;
assign v1478 = ~(w3060 | w3366);
assign w3367 = v1478;
assign w3368 = pi26 & pi35;
assign w3369 = w3058 & w3368;
assign v1479 = ~(w3367 | w3369);
assign w3370 = v1479;
assign w3371 = w3365 & ~w3370;
assign w3372 = ~w3365 & w3370;
assign v1480 = ~(w3371 | w3372);
assign w3373 = v1480;
assign w3374 = w3364 & ~w3373;
assign w3375 = ~w3364 & w3373;
assign v1481 = ~(w3374 | w3375);
assign w3376 = v1481;
assign v1482 = ~(w3175 | w3180);
assign w3377 = v1482;
assign w3378 = w3175 & w3180;
assign v1483 = ~(w3377 | w3378);
assign w3379 = v1483;
assign v1484 = ~(w3177 | w3379);
assign w3380 = v1484;
assign w3381 = w3376 & ~w3380;
assign w3382 = ~w3376 & w3380;
assign v1485 = ~(w3381 | w3382);
assign w3383 = v1485;
assign w3384 = w3352 & w3383;
assign v1486 = ~(w3352 | w3383);
assign w3385 = v1486;
assign v1487 = ~(w3384 | w3385);
assign w3386 = v1487;
assign w3387 = (~w3148 & ~w3150) | (~w3148 & w8926) | (~w3150 & w8926);
assign w3388 = w3151 & ~w3153;
assign v1488 = ~(w3155 | w3388);
assign w3389 = v1488;
assign w3390 = w3139 & ~w3141;
assign v1489 = ~(w3143 | w3390);
assign w3391 = v1489;
assign v1490 = ~(w3389 | w3391);
assign w3392 = v1490;
assign w3393 = w3389 & w3391;
assign v1491 = ~(w3392 | w3393);
assign w3394 = v1491;
assign w3395 = ~w3387 & w3394;
assign w3396 = w3387 & ~w3394;
assign v1492 = ~(w3395 | w3396);
assign w3397 = v1492;
assign w3398 = (~w3082 & ~w3084) | (~w3082 & w8611) | (~w3084 & w8611);
assign w3399 = w3085 & ~w3087;
assign v1493 = ~(w3089 | w3399);
assign w3400 = v1493;
assign w3401 = w3073 & ~w3075;
assign v1494 = ~(w3077 | w3401);
assign w3402 = v1494;
assign v1495 = ~(w3400 | w3402);
assign w3403 = v1495;
assign w3404 = w3400 & w3402;
assign v1496 = ~(w3403 | w3404);
assign w3405 = v1496;
assign w3406 = ~w3398 & w3405;
assign w3407 = w3398 & ~w3405;
assign v1497 = ~(w3406 | w3407);
assign w3408 = v1497;
assign w3409 = (~w3054 & ~w3056) | (~w3054 & w8612) | (~w3056 & w8612);
assign w3410 = (~w3048 & ~w3050) | (~w3048 & w8927) | (~w3050 & w8927);
assign w3411 = w3057 & ~w3059;
assign v1498 = ~(w3061 | w3411);
assign w3412 = v1498;
assign v1499 = ~(w3410 | w3412);
assign w3413 = v1499;
assign w3414 = w3410 & w3412;
assign v1500 = ~(w3413 | w3414);
assign w3415 = v1500;
assign w3416 = ~w3409 & w3415;
assign w3417 = w3409 & ~w3415;
assign v1501 = ~(w3416 | w3417);
assign w3418 = v1501;
assign w3419 = w3408 & w3418;
assign v1502 = ~(w3408 | w3418);
assign w3420 = v1502;
assign v1503 = ~(w3419 | w3420);
assign w3421 = v1503;
assign w3422 = w3397 & w3421;
assign v1504 = ~(w3397 | w3421);
assign w3423 = v1504;
assign v1505 = ~(w3422 | w3423);
assign w3424 = v1505;
assign w3425 = pi09 & pi51;
assign w3426 = pi13 & pi47;
assign w3427 = pi15 & pi45;
assign v1506 = ~(w3142 | w3427);
assign w3428 = v1506;
assign w3429 = pi15 & pi46;
assign w3430 = w3140 & w3429;
assign v1507 = ~(w3428 | w3430);
assign w3431 = v1507;
assign w3432 = w3426 & ~w3431;
assign w3433 = ~w3426 & w3431;
assign v1508 = ~(w3432 | w3433);
assign w3434 = v1508;
assign w3435 = w3425 & ~w3434;
assign w3436 = ~w3425 & w3434;
assign v1509 = ~(w3435 | w3436);
assign w3437 = v1509;
assign w3438 = pi10 & pi50;
assign w3439 = pi12 & pi48;
assign v1510 = ~(w3154 | w3439);
assign w3440 = v1510;
assign w3441 = pi12 & pi49;
assign w3442 = w3152 & w3441;
assign v1511 = ~(w3440 | w3442);
assign w3443 = v1511;
assign w3444 = w3438 & ~w3443;
assign w3445 = ~w3438 & w3443;
assign v1512 = ~(w3444 | w3445);
assign w3446 = v1512;
assign w3447 = w3437 & ~w3446;
assign w3448 = ~w3437 & w3446;
assign v1513 = ~(w3447 | w3448);
assign w3449 = v1513;
assign w3450 = w3424 & w3449;
assign v1514 = ~(w3424 | w3449);
assign w3451 = v1514;
assign v1515 = ~(w3450 | w3451);
assign w3452 = v1515;
assign w3453 = w3386 & w3452;
assign v1516 = ~(w3386 | w3452);
assign w3454 = v1516;
assign v1517 = ~(w3453 | w3454);
assign w3455 = v1517;
assign v1518 = ~(w3196 | w3199);
assign w3456 = v1518;
assign w3457 = pi05 & pi55;
assign w3458 = pi04 & pi56;
assign v1519 = ~(w3457 | w3458);
assign w3459 = v1519;
assign w3460 = pi05 & pi56;
assign w3461 = w2847 & w3460;
assign v1520 = ~(w3459 | w3461);
assign w3462 = v1520;
assign w3463 = pi06 & pi54;
assign w3464 = pi08 & pi52;
assign v1521 = ~(w3174 | w3464);
assign w3465 = v1521;
assign w3466 = pi08 & pi53;
assign w3467 = w3172 & w3466;
assign v1522 = ~(w3465 | w3467);
assign w3468 = v1522;
assign w3469 = w3463 & ~w3468;
assign w3470 = ~w3463 & w3468;
assign v1523 = ~(w3469 | w3470);
assign w3471 = v1523;
assign w3472 = w3462 & ~w3471;
assign w3473 = ~w3462 & w3471;
assign v1524 = ~(w3472 | w3473);
assign w3474 = v1524;
assign w3475 = ~w3456 & w3474;
assign w3476 = w3456 & ~w3474;
assign v1525 = ~(w3475 | w3476);
assign w3477 = v1525;
assign v1526 = ~(w3233 | w3236);
assign w3478 = v1526;
assign w3479 = w3477 & ~w3478;
assign w3480 = ~w3477 & w3478;
assign v1527 = ~(w3479 | w3480);
assign w3481 = v1527;
assign w3482 = w3455 & w3481;
assign v1528 = ~(w3455 | w3481);
assign w3483 = v1528;
assign v1529 = ~(w3482 | w3483);
assign w3484 = v1529;
assign w3485 = w3327 & w3484;
assign v1530 = ~(w3327 | w3484);
assign w3486 = v1530;
assign v1531 = ~(w3485 | w3486);
assign w3487 = v1531;
assign v1532 = ~(w3251 | w3254);
assign w3488 = v1532;
assign v1533 = ~(w3183 | w3186);
assign w3489 = v1533;
assign v1534 = ~(w3227 | w3239);
assign w3490 = v1534;
assign w3491 = ~w3489 & w3490;
assign w3492 = w3489 & ~w3490;
assign v1535 = ~(w3491 | w3492);
assign w3493 = v1535;
assign v1536 = ~(w3189 | w3242);
assign w3494 = v1536;
assign w3495 = w3493 & ~w3494;
assign w3496 = ~w3493 & w3494;
assign v1537 = ~(w3495 | w3496);
assign w3497 = v1537;
assign w3498 = ~w3488 & w3497;
assign w3499 = w3488 & ~w3497;
assign v1538 = ~(w3498 | w3499);
assign w3500 = v1538;
assign w3501 = w3487 & w3500;
assign v1539 = ~(w3487 | w3500);
assign w3502 = v1539;
assign v1540 = ~(w3501 | w3502);
assign w3503 = v1540;
assign w3504 = ~w3278 & w3503;
assign w3505 = w3278 & ~w3503;
assign v1541 = ~(w3504 | w3505);
assign w3506 = v1541;
assign w3507 = ~w3277 & w3506;
assign w3508 = w3277 & ~w3506;
assign v1542 = ~(w3507 | w3508);
assign w3509 = v1542;
assign v1543 = ~(w3498 | w3501);
assign w3510 = v1543;
assign v1544 = ~(w3482 | w3485);
assign w3511 = v1544;
assign v1545 = ~(w3475 | w3479);
assign w3512 = v1545;
assign v1546 = ~(w3322 | w3325);
assign w3513 = v1546;
assign v1547 = ~(w3512 | w3513);
assign w3514 = v1547;
assign w3515 = w3512 & w3513;
assign v1548 = ~(w3514 | w3515);
assign w3516 = v1548;
assign w3517 = ~w3511 & w3516;
assign w3518 = w3511 & ~w3516;
assign v1549 = ~(w3517 | w3518);
assign w3519 = v1549;
assign v1550 = ~(w3491 | w3495);
assign w3520 = v1550;
assign w3521 = (~w3289 & w3299) | (~w3289 & w9135) | (w3299 & w9135);
assign w3522 = (~w3294 & ~w3296) | (~w3294 & w9136) | (~w3296 & w9136);
assign w3523 = w3280 & ~w3282;
assign v1551 = ~(w3284 | w3523);
assign w3524 = v1551;
assign v1552 = ~(w3522 | w3524);
assign w3525 = v1552;
assign w3526 = w3522 & w3524;
assign v1553 = ~(w3525 | w3526);
assign w3527 = v1553;
assign w3528 = w3521 & w3527;
assign v1554 = ~(w3521 | w3527);
assign w3529 = v1554;
assign v1555 = ~(w3528 | w3529);
assign w3530 = v1555;
assign w3531 = (~w3450 & ~w3452) | (~w3450 & w8727) | (~w3452 & w8727);
assign v1556 = ~(w3381 | w3384);
assign w3532 = v1556;
assign w3533 = (~w3419 & ~w3421) | (~w3419 & w9137) | (~w3421 & w9137);
assign v1557 = ~(w3532 | w3533);
assign w3534 = v1557;
assign w3535 = w3532 & w3533;
assign v1558 = ~(w3534 | w3535);
assign w3536 = v1558;
assign w3537 = (w3452 & w9138) | (w3452 & w9139) | (w9138 & w9139);
assign w3538 = ~w3536 & w3531;
assign v1559 = ~(w3537 | w3538);
assign w3539 = v1559;
assign w3540 = w3530 & w3539;
assign v1560 = ~(w3530 | w3539);
assign w3541 = v1560;
assign v1561 = ~(w3540 | w3541);
assign w3542 = v1561;
assign w3543 = pi00 & pi61;
assign w3544 = pi02 & pi59;
assign w3545 = pi01 & pi60;
assign v1562 = ~(w3544 | w3545);
assign w3546 = v1562;
assign w3547 = pi02 & pi60;
assign w3548 = w3280 & w3547;
assign v1563 = ~(w3546 | w3548);
assign w3549 = v1563;
assign w3550 = w3543 & ~w3549;
assign w3551 = ~w3543 & w3549;
assign v1564 = ~(w3550 | w3551);
assign w3552 = v1564;
assign w3553 = w3378 & ~w3552;
assign w3554 = ~w3378 & w3552;
assign v1565 = ~(w3553 | w3554);
assign w3555 = v1565;
assign w3556 = (~w3392 & w3387) | (~w3392 & w9140) | (w3387 & w9140);
assign w3557 = (~w3413 & w3409) | (~w3413 & w8728) | (w3409 & w8728);
assign w3558 = (~w3403 & w3398) | (~w3403 & w8729) | (w3398 & w8729);
assign v1566 = ~(w3557 | w3558);
assign w3559 = v1566;
assign w3560 = w3557 & w3558;
assign v1567 = ~(w3559 | w3560);
assign w3561 = v1567;
assign w3562 = ~w3556 & w3561;
assign w3563 = w3556 & ~w3561;
assign v1568 = ~(w3562 | w3563);
assign w3564 = v1568;
assign w3565 = w3555 & w3564;
assign v1569 = ~(w3555 | w3564);
assign w3566 = v1569;
assign v1570 = ~(w3565 | w3566);
assign w3567 = v1570;
assign w3568 = w3542 & w3567;
assign v1571 = ~(w3542 | w3567);
assign w3569 = v1571;
assign v1572 = ~(w3568 | w3569);
assign w3570 = v1572;
assign w3571 = pi17 & pi44;
assign w3572 = pi21 & pi40;
assign w3573 = pi23 & pi38;
assign v1573 = ~(w3332 | w3573);
assign w3574 = v1573;
assign w3575 = pi23 & pi39;
assign w3576 = w3330 & w3575;
assign v1574 = ~(w3574 | w3576);
assign w3577 = v1574;
assign w3578 = w3572 & ~w3577;
assign w3579 = ~w3572 & w3577;
assign v1575 = ~(w3578 | w3579);
assign w3580 = v1575;
assign w3581 = w3571 & ~w3580;
assign w3582 = ~w3571 & w3580;
assign v1576 = ~(w3581 | w3582);
assign w3583 = v1576;
assign w3584 = pi18 & pi43;
assign w3585 = pi20 & pi41;
assign v1577 = ~(w3344 | w3585);
assign w3586 = v1577;
assign w3587 = pi20 & pi42;
assign w3588 = w3342 & w3587;
assign v1578 = ~(w3586 | w3588);
assign w3589 = v1578;
assign w3590 = w3584 & ~w3589;
assign w3591 = ~w3584 & w3589;
assign v1579 = ~(w3590 | w3591);
assign w3592 = v1579;
assign w3593 = w3583 & ~w3592;
assign w3594 = ~w3583 & w3592;
assign v1580 = ~(w3593 | w3594);
assign w3595 = v1580;
assign w3596 = pi24 & pi37;
assign w3597 = pi28 & pi33;
assign w3598 = pi29 & pi32;
assign w3599 = pi93 & w3598;
assign v1581 = ~(pi93 | w3598);
assign w3600 = v1581;
assign v1582 = ~(w3599 | w3600);
assign w3601 = v1582;
assign w3602 = w3597 & w3601;
assign v1583 = ~(w3597 | w3601);
assign w3603 = v1583;
assign v1584 = ~(w3602 | w3603);
assign w3604 = v1584;
assign w3605 = w3596 & w3604;
assign v1585 = ~(w3596 | w3604);
assign w3606 = v1585;
assign v1586 = ~(w3605 | w3606);
assign w3607 = v1586;
assign w3608 = pi25 & pi36;
assign w3609 = pi27 & pi34;
assign v1587 = ~(w3368 | w3609);
assign w3610 = v1587;
assign w3611 = pi27 & pi35;
assign w3612 = w3366 & w3611;
assign v1588 = ~(w3610 | w3612);
assign w3613 = v1588;
assign w3614 = w3608 & ~w3613;
assign w3615 = ~w3608 & w3613;
assign v1589 = ~(w3614 | w3615);
assign w3616 = v1589;
assign w3617 = w3607 & ~w3616;
assign w3618 = ~w3607 & w3616;
assign v1590 = ~(w3617 | w3618);
assign w3619 = v1590;
assign v1591 = ~(w3461 | w3472);
assign w3620 = v1591;
assign w3621 = w3463 & ~w3465;
assign v1592 = ~(w3467 | w3621);
assign w3622 = v1592;
assign v1593 = ~(w3620 | w3622);
assign w3623 = v1593;
assign w3624 = w3620 & w3622;
assign v1594 = ~(w3623 | w3624);
assign w3625 = v1594;
assign v1595 = ~(w3619 | w3625);
assign w3626 = v1595;
assign w3627 = w3619 & w3625;
assign v1596 = ~(w3626 | w3627);
assign w3628 = v1596;
assign w3629 = ~w3595 & w3628;
assign w3630 = w3595 & ~w3628;
assign v1597 = ~(w3629 | w3630);
assign w3631 = v1597;
assign w3632 = (~w3435 & ~w3437) | (~w3435 & w8928) | (~w3437 & w8928);
assign w3633 = w3438 & ~w3440;
assign v1598 = ~(w3442 | w3633);
assign w3634 = v1598;
assign w3635 = w3426 & ~w3428;
assign v1599 = ~(w3430 | w3635);
assign w3636 = v1599;
assign v1600 = ~(w3634 | w3636);
assign w3637 = v1600;
assign w3638 = w3634 & w3636;
assign v1601 = ~(w3637 | w3638);
assign w3639 = v1601;
assign w3640 = ~w3632 & w3639;
assign w3641 = w3632 & ~w3639;
assign v1602 = ~(w3640 | w3641);
assign w3642 = v1602;
assign w3643 = (~w3338 & ~w3340) | (~w3338 & w8613) | (~w3340 & w8613);
assign w3644 = w3341 & ~w3343;
assign v1603 = ~(w3345 | w3644);
assign w3645 = v1603;
assign w3646 = w3329 & ~w3331;
assign v1604 = ~(w3333 | w3646);
assign w3647 = v1604;
assign v1605 = ~(w3645 | w3647);
assign w3648 = v1605;
assign w3649 = w3645 & w3647;
assign v1606 = ~(w3648 | w3649);
assign w3650 = v1606;
assign w3651 = ~w3643 & w3650;
assign w3652 = w3643 & ~w3650;
assign v1607 = ~(w3651 | w3652);
assign w3653 = v1607;
assign w3654 = (~w3362 & ~w3364) | (~w3362 & w8614) | (~w3364 & w8614);
assign w3655 = (~w3356 & ~w3358) | (~w3356 & w8929) | (~w3358 & w8929);
assign w3656 = w3365 & ~w3367;
assign v1608 = ~(w3369 | w3656);
assign w3657 = v1608;
assign v1609 = ~(w3655 | w3657);
assign w3658 = v1609;
assign w3659 = w3655 & w3657;
assign v1610 = ~(w3658 | w3659);
assign w3660 = v1610;
assign w3661 = ~w3654 & w3660;
assign w3662 = w3654 & ~w3660;
assign v1611 = ~(w3661 | w3662);
assign w3663 = v1611;
assign w3664 = w3653 & w3663;
assign v1612 = ~(w3653 | w3663);
assign w3665 = v1612;
assign v1613 = ~(w3664 | w3665);
assign w3666 = v1613;
assign w3667 = w3642 & w3666;
assign v1614 = ~(w3642 | w3666);
assign w3668 = v1614;
assign v1615 = ~(w3667 | w3668);
assign w3669 = v1615;
assign w3670 = pi10 & pi51;
assign w3671 = pi14 & pi47;
assign w3672 = pi16 & pi45;
assign v1616 = ~(w3429 | w3672);
assign w3673 = v1616;
assign w3674 = pi16 & pi46;
assign w3675 = w3427 & w3674;
assign v1617 = ~(w3673 | w3675);
assign w3676 = v1617;
assign w3677 = w3671 & ~w3676;
assign w3678 = ~w3671 & w3676;
assign v1618 = ~(w3677 | w3678);
assign w3679 = v1618;
assign w3680 = w3670 & ~w3679;
assign w3681 = ~w3670 & w3679;
assign v1619 = ~(w3680 | w3681);
assign w3682 = v1619;
assign w3683 = pi11 & pi50;
assign w3684 = pi13 & pi48;
assign v1620 = ~(w3441 | w3684);
assign w3685 = v1620;
assign w3686 = pi13 & pi49;
assign w3687 = w3439 & w3686;
assign v1621 = ~(w3685 | w3687);
assign w3688 = v1621;
assign w3689 = w3683 & ~w3688;
assign w3690 = ~w3683 & w3688;
assign v1622 = ~(w3689 | w3690);
assign w3691 = v1622;
assign w3692 = w3682 & ~w3691;
assign w3693 = ~w3682 & w3691;
assign v1623 = ~(w3692 | w3693);
assign w3694 = v1623;
assign w3695 = w3669 & w3694;
assign v1624 = ~(w3669 | w3694);
assign w3696 = v1624;
assign v1625 = ~(w3695 | w3696);
assign w3697 = v1625;
assign w3698 = ~w3631 & w3697;
assign w3699 = w3631 & ~w3697;
assign v1626 = ~(w3698 | w3699);
assign w3700 = v1626;
assign w3701 = (~w3316 & w3313) | (~w3316 & w8930) | (w3313 & w8930);
assign v1627 = ~(w3307 | w3310);
assign w3702 = v1627;
assign w3703 = pi07 & pi54;
assign w3704 = pi09 & pi52;
assign v1628 = ~(w3466 | w3704);
assign w3705 = v1628;
assign w3706 = pi09 & pi53;
assign w3707 = w3464 & w3706;
assign v1629 = ~(w3705 | w3707);
assign w3708 = v1629;
assign w3709 = w3703 & ~w3708;
assign w3710 = ~w3703 & w3708;
assign v1630 = ~(w3709 | w3710);
assign w3711 = v1630;
assign w3712 = w3283 & ~w3711;
assign w3713 = ~w3283 & w3711;
assign v1631 = ~(w3712 | w3713);
assign w3714 = v1631;
assign w3715 = pi04 & pi57;
assign w3716 = pi06 & pi55;
assign v1632 = ~(w3460 | w3716);
assign w3717 = v1632;
assign w3718 = pi06 & pi56;
assign w3719 = w3457 & w3718;
assign v1633 = ~(w3717 | w3719);
assign w3720 = v1633;
assign w3721 = w3715 & ~w3720;
assign w3722 = ~w3715 & w3720;
assign v1634 = ~(w3721 | w3722);
assign w3723 = v1634;
assign w3724 = w3714 & ~w3723;
assign w3725 = ~w3714 & w3723;
assign v1635 = ~(w3724 | w3725);
assign w3726 = v1635;
assign w3727 = w3702 & ~w3726;
assign w3728 = ~w3702 & w3726;
assign v1636 = ~(w3727 | w3728);
assign w3729 = v1636;
assign w3730 = w3701 & w3729;
assign v1637 = ~(w3701 | w3729);
assign w3731 = v1637;
assign v1638 = ~(w3730 | w3731);
assign w3732 = v1638;
assign w3733 = w3700 & ~w3732;
assign w3734 = ~w3700 & w3732;
assign v1639 = ~(w3733 | w3734);
assign w3735 = v1639;
assign w3736 = w3570 & w3735;
assign v1640 = ~(w3570 | w3735);
assign w3737 = v1640;
assign v1641 = ~(w3736 | w3737);
assign w3738 = v1641;
assign w3739 = ~w3520 & w3738;
assign w3740 = w3520 & ~w3738;
assign v1642 = ~(w3739 | w3740);
assign w3741 = v1642;
assign w3742 = w3519 & w3741;
assign v1643 = ~(w3519 | w3741);
assign w3743 = v1643;
assign v1644 = ~(w3742 | w3743);
assign w3744 = v1644;
assign w3745 = w3510 & ~w3744;
assign w3746 = ~w3510 & w3744;
assign v1645 = ~(w3745 | w3746);
assign w3747 = v1645;
assign v1646 = ~(w3504 | w3507);
assign w3748 = v1646;
assign w3749 = ~w3747 & w3748;
assign w3750 = w3747 & ~w3748;
assign v1647 = ~(w3749 | w3750);
assign w3751 = v1647;
assign w3752 = w3506 & w3747;
assign w3753 = w3272 & w3752;
assign w3754 = w3275 & w9269;
assign v1648 = ~(w3753 | w3754);
assign w3755 = v1648;
assign v1649 = ~(w3504 | w3746);
assign w3756 = v1649;
assign v1650 = ~(w3745 | w3756);
assign w3757 = v1650;
assign w3758 = w3755 & ~w3757;
assign w3759 = pi11 & pi51;
assign w3760 = pi15 & pi47;
assign w3761 = pi17 & pi45;
assign v1651 = ~(w3674 | w3761);
assign w3762 = v1651;
assign w3763 = pi17 & pi46;
assign w3764 = w3672 & w3763;
assign v1652 = ~(w3762 | w3764);
assign w3765 = v1652;
assign w3766 = w3760 & ~w3765;
assign w3767 = ~w3760 & w3765;
assign v1653 = ~(w3766 | w3767);
assign w3768 = v1653;
assign w3769 = w3759 & ~w3768;
assign w3770 = ~w3759 & w3768;
assign v1654 = ~(w3769 | w3770);
assign w3771 = v1654;
assign w3772 = pi12 & pi50;
assign w3773 = pi14 & pi48;
assign v1655 = ~(w3686 | w3773);
assign w3774 = v1655;
assign w3775 = pi14 & pi49;
assign w3776 = w3684 & w3775;
assign v1656 = ~(w3774 | w3776);
assign w3777 = v1656;
assign w3778 = w3772 & ~w3777;
assign w3779 = ~w3772 & w3777;
assign v1657 = ~(w3778 | w3779);
assign w3780 = v1657;
assign w3781 = w3771 & ~w3780;
assign w3782 = ~w3771 & w3780;
assign v1658 = ~(w3781 | w3782);
assign w3783 = v1658;
assign w3784 = pi18 & pi44;
assign w3785 = pi22 & pi40;
assign w3786 = pi24 & pi38;
assign v1659 = ~(w3575 | w3786);
assign w3787 = v1659;
assign w3788 = pi24 & pi39;
assign w3789 = w3573 & w3788;
assign v1660 = ~(w3787 | w3789);
assign w3790 = v1660;
assign w3791 = w3785 & ~w3790;
assign w3792 = ~w3785 & w3790;
assign v1661 = ~(w3791 | w3792);
assign w3793 = v1661;
assign w3794 = w3784 & ~w3793;
assign w3795 = ~w3784 & w3793;
assign v1662 = ~(w3794 | w3795);
assign w3796 = v1662;
assign w3797 = pi19 & pi43;
assign w3798 = pi21 & pi41;
assign v1663 = ~(w3587 | w3798);
assign w3799 = v1663;
assign w3800 = pi21 & pi42;
assign w3801 = w3585 & w3800;
assign v1664 = ~(w3799 | w3801);
assign w3802 = v1664;
assign w3803 = w3797 & ~w3802;
assign w3804 = ~w3797 & w3802;
assign v1665 = ~(w3803 | w3804);
assign w3805 = v1665;
assign w3806 = w3796 & ~w3805;
assign w3807 = ~w3796 & w3805;
assign v1666 = ~(w3806 | w3807);
assign w3808 = v1666;
assign w3809 = pi25 & pi37;
assign w3810 = pi29 & pi33;
assign w3811 = pi30 & pi32;
assign w3812 = pi94 & w3811;
assign v1667 = ~(pi94 | w3811);
assign w3813 = v1667;
assign v1668 = ~(w3812 | w3813);
assign w3814 = v1668;
assign w3815 = w3810 & w3814;
assign v1669 = ~(w3810 | w3814);
assign w3816 = v1669;
assign v1670 = ~(w3815 | w3816);
assign w3817 = v1670;
assign w3818 = w3809 & w3817;
assign v1671 = ~(w3809 | w3817);
assign w3819 = v1671;
assign v1672 = ~(w3818 | w3819);
assign w3820 = v1672;
assign w3821 = pi26 & pi36;
assign w3822 = pi28 & pi34;
assign v1673 = ~(w3611 | w3822);
assign w3823 = v1673;
assign w3824 = pi28 & pi35;
assign w3825 = w3609 & w3824;
assign v1674 = ~(w3823 | w3825);
assign w3826 = v1674;
assign w3827 = w3821 & ~w3826;
assign w3828 = ~w3821 & w3826;
assign v1675 = ~(w3827 | w3828);
assign w3829 = v1675;
assign w3830 = w3820 & ~w3829;
assign w3831 = ~w3820 & w3829;
assign v1676 = ~(w3830 | w3831);
assign w3832 = v1676;
assign w3833 = w3808 & w3832;
assign v1677 = ~(w3808 | w3832);
assign w3834 = v1677;
assign v1678 = ~(w3833 | w3834);
assign w3835 = v1678;
assign w3836 = w3783 & w3835;
assign v1679 = ~(w3783 | w3835);
assign w3837 = v1679;
assign v1680 = ~(w3836 | w3837);
assign w3838 = v1680;
assign w3839 = (~w3712 & ~w3714) | (~w3712 & w8615) | (~w3714 & w8615);
assign w3840 = w3715 & ~w3717;
assign v1681 = ~(w3719 | w3840);
assign w3841 = v1681;
assign w3842 = w3703 & ~w3705;
assign v1682 = ~(w3707 | w3842);
assign w3843 = v1682;
assign v1683 = ~(w3841 | w3843);
assign w3844 = v1683;
assign w3845 = w3841 & w3843;
assign v1684 = ~(w3844 | w3845);
assign w3846 = v1684;
assign w3847 = ~w3839 & w3846;
assign w3848 = w3839 & ~w3846;
assign v1685 = ~(w3847 | w3848);
assign w3849 = v1685;
assign w3850 = (~w3680 & ~w3682) | (~w3680 & w8616) | (~w3682 & w8616);
assign w3851 = w3683 & ~w3685;
assign v1686 = ~(w3687 | w3851);
assign w3852 = v1686;
assign w3853 = w3671 & ~w3673;
assign v1687 = ~(w3675 | w3853);
assign w3854 = v1687;
assign v1688 = ~(w3852 | w3854);
assign w3855 = v1688;
assign w3856 = w3852 & w3854;
assign v1689 = ~(w3855 | w3856);
assign w3857 = v1689;
assign w3858 = ~w3850 & w3857;
assign w3859 = w3850 & ~w3857;
assign v1690 = ~(w3858 | w3859);
assign w3860 = v1690;
assign w3861 = (~w3581 & ~w3583) | (~w3581 & w8617) | (~w3583 & w8617);
assign w3862 = w3584 & ~w3586;
assign v1691 = ~(w3588 | w3862);
assign w3863 = v1691;
assign w3864 = w3572 & ~w3574;
assign v1692 = ~(w3576 | w3864);
assign w3865 = v1692;
assign v1693 = ~(w3863 | w3865);
assign w3866 = v1693;
assign w3867 = w3863 & w3865;
assign v1694 = ~(w3866 | w3867);
assign w3868 = v1694;
assign w3869 = ~w3861 & w3868;
assign w3870 = w3861 & ~w3868;
assign v1695 = ~(w3869 | w3870);
assign w3871 = v1695;
assign w3872 = w3860 & w3871;
assign v1696 = ~(w3860 | w3871);
assign w3873 = v1696;
assign v1697 = ~(w3872 | w3873);
assign w3874 = v1697;
assign w3875 = w3849 & w3874;
assign v1698 = ~(w3849 | w3874);
assign w3876 = v1698;
assign v1699 = ~(w3875 | w3876);
assign w3877 = v1699;
assign w3878 = pi04 & pi58;
assign w3879 = pi08 & pi54;
assign w3880 = pi10 & pi52;
assign v1700 = ~(w3706 | w3880);
assign w3881 = v1700;
assign w3882 = pi10 & pi53;
assign w3883 = w3704 & w3882;
assign v1701 = ~(w3881 | w3883);
assign w3884 = v1701;
assign w3885 = w3879 & ~w3884;
assign w3886 = ~w3879 & w3884;
assign v1702 = ~(w3885 | w3886);
assign w3887 = v1702;
assign w3888 = w3878 & ~w3887;
assign w3889 = ~w3878 & w3887;
assign v1703 = ~(w3888 | w3889);
assign w3890 = v1703;
assign w3891 = pi05 & pi57;
assign w3892 = pi07 & pi55;
assign v1704 = ~(w3718 | w3892);
assign w3893 = v1704;
assign w3894 = pi07 & pi56;
assign w3895 = w3716 & w3894;
assign v1705 = ~(w3893 | w3895);
assign w3896 = v1705;
assign w3897 = w3891 & ~w3896;
assign w3898 = ~w3891 & w3896;
assign v1706 = ~(w3897 | w3898);
assign w3899 = v1706;
assign w3900 = w3890 & ~w3899;
assign w3901 = ~w3890 & w3899;
assign v1707 = ~(w3900 | w3901);
assign w3902 = v1707;
assign w3903 = w3877 & w3902;
assign v1708 = ~(w3877 | w3902);
assign w3904 = v1708;
assign v1709 = ~(w3903 | w3904);
assign w3905 = v1709;
assign w3906 = w3838 & w3905;
assign v1710 = ~(w3838 | w3905);
assign w3907 = v1710;
assign v1711 = ~(w3906 | w3907);
assign w3908 = v1711;
assign w3909 = (~w3534 & w3531) | (~w3534 & w8931) | (w3531 & w8931);
assign w3910 = pi03 & pi59;
assign v1712 = ~(w3547 | w3910);
assign w3911 = v1712;
assign w3912 = pi03 & pi60;
assign w3913 = w3544 & w3912;
assign v1713 = ~(w3911 | w3913);
assign w3914 = v1713;
assign v1714 = ~(w3525 | w3528);
assign w3915 = v1714;
assign w3916 = w3914 & ~w3915;
assign w3917 = ~w3914 & w3915;
assign v1715 = ~(w3916 | w3917);
assign w3918 = v1715;
assign w3919 = w3909 & w3918;
assign v1716 = ~(w3909 | w3918);
assign w3920 = v1716;
assign v1717 = ~(w3919 | w3920);
assign w3921 = v1717;
assign w3922 = w3908 & ~w3921;
assign w3923 = ~w3908 & w3921;
assign v1718 = ~(w3922 | w3923);
assign w3924 = v1718;
assign w3925 = (~w3605 & ~w3607) | (~w3605 & w8618) | (~w3607 & w8618);
assign w3926 = (~w3599 & ~w3601) | (~w3599 & w8932) | (~w3601 & w8932);
assign w3927 = w3608 & ~w3610;
assign v1719 = ~(w3612 | w3927);
assign w3928 = v1719;
assign v1720 = ~(w3926 | w3928);
assign w3929 = v1720;
assign w3930 = w3926 & w3928;
assign v1721 = ~(w3929 | w3930);
assign w3931 = v1721;
assign w3932 = ~w3925 & w3931;
assign w3933 = w3925 & ~w3931;
assign v1722 = ~(w3932 | w3933);
assign w3934 = v1722;
assign w3935 = pi01 & pi61;
assign w3936 = pi00 & pi62;
assign v1723 = ~(w3935 | w3936);
assign w3937 = v1723;
assign w3938 = pi01 & pi62;
assign w3939 = w3543 & w3938;
assign v1724 = ~(w3937 | w3939);
assign w3940 = v1724;
assign w3941 = (~w3654 & w8933) | (~w3654 & w8934) | (w8933 & w8934);
assign w3942 = (w3654 & w8935) | (w3654 & w8936) | (w8935 & w8936);
assign v1725 = ~(w3941 | w3942);
assign w3943 = v1725;
assign w3944 = w3934 & w3943;
assign v1726 = ~(w3934 | w3943);
assign w3945 = v1726;
assign v1727 = ~(w3944 | w3945);
assign w3946 = v1727;
assign w3947 = (~w3637 & w3632) | (~w3637 & w9141) | (w3632 & w9141);
assign w3948 = (~w3648 & w3643) | (~w3648 & w8730) | (w3643 & w8730);
assign w3949 = w3623 & ~w3948;
assign w3950 = ~w3623 & w3948;
assign v1728 = ~(w3949 | w3950);
assign w3951 = v1728;
assign v1729 = ~(w3947 | w3951);
assign w3952 = v1729;
assign w3953 = w3947 & w3951;
assign v1730 = ~(w3952 | w3953);
assign w3954 = v1730;
assign w3955 = w3946 & ~w3954;
assign w3956 = ~w3946 & w3954;
assign v1731 = ~(w3955 | w3956);
assign w3957 = v1731;
assign w3958 = (~w3553 & ~w3564) | (~w3553 & w8937) | (~w3564 & w8937);
assign w3959 = (~w3559 & ~w3561) | (~w3559 & w8938) | (~w3561 & w8938);
assign w3960 = w3543 & ~w3546;
assign v1732 = ~(w3548 | w3960);
assign w3961 = v1732;
assign v1733 = ~(w3959 | w3961);
assign w3962 = v1733;
assign w3963 = w3959 & w3961;
assign v1734 = ~(w3962 | w3963);
assign w3964 = v1734;
assign w3965 = ~w3958 & w3964;
assign w3966 = w3958 & ~w3964;
assign v1735 = ~(w3965 | w3966);
assign w3967 = v1735;
assign w3968 = (~w3695 & ~w3697) | (~w3695 & w8731) | (~w3697 & w8731);
assign v1736 = ~(w3626 | w3629);
assign w3969 = v1736;
assign w3970 = (~w3664 & ~w3666) | (~w3664 & w9142) | (~w3666 & w9142);
assign w3971 = w3969 & ~w3970;
assign w3972 = ~w3969 & w3970;
assign v1737 = ~(w3971 | w3972);
assign w3973 = v1737;
assign w3974 = w3973 & w3968;
assign w3975 = (w3697 & w9143) | (w3697 & w9144) | (w9143 & w9144);
assign v1738 = ~(w3974 | w3975);
assign w3976 = v1738;
assign w3977 = w3967 & ~w3976;
assign w3978 = ~w3967 & w3976;
assign v1739 = ~(w3977 | w3978);
assign w3979 = v1739;
assign w3980 = w3957 & ~w3979;
assign w3981 = ~w3957 & w3979;
assign v1740 = ~(w3980 | w3981);
assign w3982 = v1740;
assign w3983 = w3924 & ~w3982;
assign w3984 = ~w3924 & w3982;
assign v1741 = ~(w3983 | w3984);
assign w3985 = v1741;
assign v1742 = ~(w3514 | w3517);
assign w3986 = v1742;
assign w3987 = (~w3733 & ~w3570) | (~w3733 & w8939) | (~w3570 & w8939);
assign v1743 = ~(w3727 | w3730);
assign w3988 = v1743;
assign w3989 = (~w3540 & ~w3542) | (~w3540 & w8940) | (~w3542 & w8940);
assign w3990 = w3988 & ~w3989;
assign w3991 = ~w3988 & w3989;
assign v1744 = ~(w3990 | w3991);
assign w3992 = v1744;
assign w3993 = ~w3987 & w3992;
assign w3994 = w3987 & ~w3992;
assign v1745 = ~(w3993 | w3994);
assign w3995 = v1745;
assign w3996 = ~w3986 & w3995;
assign w3997 = w3986 & ~w3995;
assign v1746 = ~(w3996 | w3997);
assign w3998 = v1746;
assign w3999 = w3985 & w3998;
assign v1747 = ~(w3985 | w3998);
assign w4000 = v1747;
assign v1748 = ~(w3999 | w4000);
assign w4001 = v1748;
assign v1749 = ~(w3739 | w3742);
assign w4002 = v1749;
assign w4003 = w4001 & ~w4002;
assign w4004 = ~w4001 & w4002;
assign v1750 = ~(w4003 | w4004);
assign w4005 = v1750;
assign w4006 = ~w3758 & w4005;
assign w4007 = w3758 & ~w4005;
assign v1751 = ~(w4006 | w4007);
assign w4008 = v1751;
assign v1752 = ~(w3757 | w4003);
assign w4009 = v1752;
assign w4010 = ~w3754 & w8732;
assign v1753 = ~(w4004 | w4010);
assign w4011 = v1753;
assign v1754 = ~(w3996 | w3999);
assign w4012 = v1754;
assign w4013 = pi12 & pi51;
assign w4014 = pi16 & pi47;
assign w4015 = pi18 & pi45;
assign v1755 = ~(w3763 | w4015);
assign w4016 = v1755;
assign w4017 = pi18 & pi46;
assign w4018 = w3761 & w4017;
assign v1756 = ~(w4016 | w4018);
assign w4019 = v1756;
assign w4020 = w4014 & ~w4019;
assign w4021 = ~w4014 & w4019;
assign v1757 = ~(w4020 | w4021);
assign w4022 = v1757;
assign w4023 = w4013 & ~w4022;
assign w4024 = ~w4013 & w4022;
assign v1758 = ~(w4023 | w4024);
assign w4025 = v1758;
assign w4026 = pi13 & pi50;
assign w4027 = pi15 & pi48;
assign v1759 = ~(w3775 | w4027);
assign w4028 = v1759;
assign w4029 = pi15 & pi49;
assign w4030 = w3773 & w4029;
assign v1760 = ~(w4028 | w4030);
assign w4031 = v1760;
assign w4032 = w4026 & ~w4031;
assign w4033 = ~w4026 & w4031;
assign v1761 = ~(w4032 | w4033);
assign w4034 = v1761;
assign w4035 = w4025 & ~w4034;
assign w4036 = ~w4025 & w4034;
assign v1762 = ~(w4035 | w4036);
assign w4037 = v1762;
assign w4038 = pi19 & pi44;
assign w4039 = pi23 & pi40;
assign w4040 = pi25 & pi38;
assign v1763 = ~(w3788 | w4040);
assign w4041 = v1763;
assign w4042 = pi25 & pi39;
assign w4043 = w3786 & w4042;
assign v1764 = ~(w4041 | w4043);
assign w4044 = v1764;
assign w4045 = w4039 & ~w4044;
assign w4046 = ~w4039 & w4044;
assign v1765 = ~(w4045 | w4046);
assign w4047 = v1765;
assign w4048 = w4038 & ~w4047;
assign w4049 = ~w4038 & w4047;
assign v1766 = ~(w4048 | w4049);
assign w4050 = v1766;
assign w4051 = pi20 & pi43;
assign w4052 = pi22 & pi41;
assign v1767 = ~(w3800 | w4052);
assign w4053 = v1767;
assign w4054 = pi22 & pi42;
assign w4055 = w3798 & w4054;
assign v1768 = ~(w4053 | w4055);
assign w4056 = v1768;
assign w4057 = w4051 & ~w4056;
assign w4058 = ~w4051 & w4056;
assign v1769 = ~(w4057 | w4058);
assign w4059 = v1769;
assign w4060 = w4050 & ~w4059;
assign w4061 = ~w4050 & w4059;
assign v1770 = ~(w4060 | w4061);
assign w4062 = v1770;
assign w4063 = pi26 & pi37;
assign w4064 = pi30 & pi33;
assign w4065 = pi31 & pi32;
assign v1771 = ~(pi95 | w4065);
assign w4066 = v1771;
assign w4067 = pi95 & w4065;
assign v1772 = ~(w4066 | w4067);
assign w4068 = v1772;
assign w4069 = w4064 & w4068;
assign v1773 = ~(w4064 | w4068);
assign w4070 = v1773;
assign v1774 = ~(w4069 | w4070);
assign w4071 = v1774;
assign w4072 = w4063 & w4071;
assign v1775 = ~(w4063 | w4071);
assign w4073 = v1775;
assign v1776 = ~(w4072 | w4073);
assign w4074 = v1776;
assign w4075 = pi27 & pi36;
assign w4076 = pi29 & pi34;
assign v1777 = ~(w3824 | w4076);
assign w4077 = v1777;
assign w4078 = pi29 & pi35;
assign w4079 = w3822 & w4078;
assign v1778 = ~(w4077 | w4079);
assign w4080 = v1778;
assign w4081 = w4075 & ~w4080;
assign w4082 = ~w4075 & w4080;
assign v1779 = ~(w4081 | w4082);
assign w4083 = v1779;
assign w4084 = w4074 & ~w4083;
assign w4085 = ~w4074 & w4083;
assign v1780 = ~(w4084 | w4085);
assign w4086 = v1780;
assign w4087 = w4062 & w4086;
assign v1781 = ~(w4062 | w4086);
assign w4088 = v1781;
assign v1782 = ~(w4087 | w4088);
assign w4089 = v1782;
assign w4090 = w4037 & w4089;
assign v1783 = ~(w4037 | w4089);
assign w4091 = v1783;
assign v1784 = ~(w4090 | w4091);
assign w4092 = v1784;
assign w4093 = pi05 & pi58;
assign w4094 = pi09 & pi54;
assign w4095 = pi11 & pi52;
assign v1785 = ~(w3882 | w4095);
assign w4096 = v1785;
assign w4097 = pi11 & pi53;
assign w4098 = w3880 & w4097;
assign v1786 = ~(w4096 | w4098);
assign w4099 = v1786;
assign w4100 = w4094 & ~w4099;
assign w4101 = ~w4094 & w4099;
assign v1787 = ~(w4100 | w4101);
assign w4102 = v1787;
assign w4103 = w4093 & ~w4102;
assign w4104 = ~w4093 & w4102;
assign v1788 = ~(w4103 | w4104);
assign w4105 = v1788;
assign w4106 = pi06 & pi57;
assign w4107 = pi08 & pi55;
assign v1789 = ~(w3894 | w4107);
assign w4108 = v1789;
assign w4109 = pi08 & pi56;
assign w4110 = w3892 & w4109;
assign v1790 = ~(w4108 | w4110);
assign w4111 = v1790;
assign w4112 = w4106 & ~w4111;
assign w4113 = ~w4106 & w4111;
assign v1791 = ~(w4112 | w4113);
assign w4114 = v1791;
assign w4115 = w4105 & ~w4114;
assign w4116 = ~w4105 & w4114;
assign v1792 = ~(w4115 | w4116);
assign w4117 = v1792;
assign w4118 = (~w3888 & ~w3890) | (~w3888 & w8619) | (~w3890 & w8619);
assign w4119 = w3891 & ~w3893;
assign v1793 = ~(w3895 | w4119);
assign w4120 = v1793;
assign w4121 = w3879 & ~w3881;
assign v1794 = ~(w3883 | w4121);
assign w4122 = v1794;
assign v1795 = ~(w4120 | w4122);
assign w4123 = v1795;
assign w4124 = w4120 & w4122;
assign v1796 = ~(w4123 | w4124);
assign w4125 = v1796;
assign w4126 = ~w4118 & w4125;
assign w4127 = w4118 & ~w4125;
assign v1797 = ~(w4126 | w4127);
assign w4128 = v1797;
assign w4129 = (~w3769 & ~w3771) | (~w3769 & w8620) | (~w3771 & w8620);
assign w4130 = w3772 & ~w3774;
assign v1798 = ~(w3776 | w4130);
assign w4131 = v1798;
assign w4132 = w3760 & ~w3762;
assign v1799 = ~(w3764 | w4132);
assign w4133 = v1799;
assign v1800 = ~(w4131 | w4133);
assign w4134 = v1800;
assign w4135 = w4131 & w4133;
assign v1801 = ~(w4134 | w4135);
assign w4136 = v1801;
assign w4137 = ~w4129 & w4136;
assign w4138 = w4129 & ~w4136;
assign v1802 = ~(w4137 | w4138);
assign w4139 = v1802;
assign w4140 = w4128 & w4139;
assign v1803 = ~(w4128 | w4139);
assign w4141 = v1803;
assign v1804 = ~(w4140 | w4141);
assign w4142 = v1804;
assign w4143 = w3913 & ~w4142;
assign w4144 = ~w3913 & w4142;
assign v1805 = ~(w4143 | w4144);
assign w4145 = v1805;
assign w4146 = ~w4117 & w4145;
assign w4147 = w4117 & ~w4145;
assign v1806 = ~(w4146 | w4147);
assign w4148 = v1806;
assign w4149 = ~w4092 & w4148;
assign w4150 = w4092 & ~w4148;
assign v1807 = ~(w4149 | w4150);
assign w4151 = v1807;
assign w4152 = pi00 & pi63;
assign w4153 = w3938 & ~w4152;
assign w4154 = ~w3938 & w4152;
assign v1808 = ~(w4153 | w4154);
assign w4155 = v1808;
assign w4156 = pi02 & pi61;
assign w4157 = pi04 & pi59;
assign v1809 = ~(w3912 | w4157);
assign w4158 = v1809;
assign w4159 = pi04 & pi60;
assign w4160 = w3910 & w4159;
assign v1810 = ~(w4158 | w4160);
assign w4161 = v1810;
assign w4162 = w4156 & ~w4161;
assign w4163 = ~w4156 & w4161;
assign v1811 = ~(w4162 | w4163);
assign w4164 = v1811;
assign w4165 = w4155 & ~w4164;
assign w4166 = ~w4155 & w4164;
assign v1812 = ~(w4165 | w4166);
assign w4167 = v1812;
assign w4168 = (w4167 & w3965) | (w4167 & w9145) | (w3965 & w9145);
assign w4169 = ~w3965 & w9146;
assign v1813 = ~(w4168 | w4169);
assign w4170 = v1813;
assign w4171 = (~w3972 & ~w3968) | (~w3972 & w8941) | (~w3968 & w8941);
assign w4172 = w4170 & w4171;
assign v1814 = ~(w4170 | w4171);
assign w4173 = v1814;
assign v1815 = ~(w4172 | w4173);
assign w4174 = v1815;
assign w4175 = w4151 & ~w4174;
assign w4176 = ~w4151 & w4174;
assign v1816 = ~(w4175 | w4176);
assign w4177 = v1816;
assign w4178 = (~w3818 & ~w3820) | (~w3818 & w8733) | (~w3820 & w8733);
assign v1817 = ~(w3812 | w3815);
assign w4179 = v1817;
assign w4180 = w3821 & ~w3823;
assign v1818 = ~(w3825 | w4180);
assign w4181 = v1818;
assign v1819 = ~(w4179 | w4181);
assign w4182 = v1819;
assign w4183 = w4179 & w4181;
assign v1820 = ~(w4182 | w4183);
assign w4184 = v1820;
assign w4185 = ~w4178 & w4184;
assign w4186 = w4178 & ~w4184;
assign v1821 = ~(w4185 | w4186);
assign w4187 = v1821;
assign w4188 = (~w3855 & w3850) | (~w3855 & w8734) | (w3850 & w8734);
assign w4189 = (~w3844 & w3839) | (~w3844 & w8735) | (w3839 & w8735);
assign v1822 = ~(w4188 | w4189);
assign w4190 = v1822;
assign w4191 = w4188 & w4189;
assign v1823 = ~(w4190 | w4191);
assign w4192 = v1823;
assign w4193 = w4187 & w4192;
assign v1824 = ~(w4187 | w4192);
assign w4194 = v1824;
assign v1825 = ~(w4193 | w4194);
assign w4195 = v1825;
assign w4196 = (~w3794 & ~w3796) | (~w3794 & w8736) | (~w3796 & w8736);
assign w4197 = w3797 & ~w3799;
assign v1826 = ~(w3801 | w4197);
assign w4198 = v1826;
assign w4199 = w3785 & ~w3787;
assign v1827 = ~(w3789 | w4199);
assign w4200 = v1827;
assign v1828 = ~(w4198 | w4200);
assign w4201 = v1828;
assign w4202 = w4198 & w4200;
assign v1829 = ~(w4201 | w4202);
assign w4203 = v1829;
assign w4204 = ~w4196 & w4203;
assign w4205 = w4196 & ~w4203;
assign v1830 = ~(w4204 | w4205);
assign w4206 = v1830;
assign w4207 = (~w3866 & w3861) | (~w3866 & w8737) | (w3861 & w8737);
assign w4208 = (~w3929 & w3925) | (~w3929 & w8738) | (w3925 & w8738);
assign w4209 = w4207 & w4208;
assign v1831 = ~(w4207 | w4208);
assign w4210 = v1831;
assign v1832 = ~(w4209 | w4210);
assign w4211 = v1832;
assign w4212 = w4206 & ~w4211;
assign w4213 = ~w4206 & w4211;
assign v1833 = ~(w4212 | w4213);
assign w4214 = v1833;
assign w4215 = w4195 & w4214;
assign v1834 = ~(w4195 | w4214);
assign w4216 = v1834;
assign v1835 = ~(w4215 | w4216);
assign w4217 = v1835;
assign w4218 = (~w3944 & w3954) | (~w3944 & w8942) | (w3954 & w8942);
assign v1836 = ~(w3939 | w3941);
assign w4219 = v1836;
assign w4220 = (~w3950 & ~w3951) | (~w3950 & w8943) | (~w3951 & w8943);
assign w4221 = ~w4219 & w4220;
assign w4222 = w4219 & ~w4220;
assign v1837 = ~(w4221 | w4222);
assign w4223 = v1837;
assign w4224 = ~w4218 & w4223;
assign w4225 = w4218 & ~w4223;
assign v1838 = ~(w4224 | w4225);
assign w4226 = v1838;
assign w4227 = (~w3903 & ~w3905) | (~w3903 & w8739) | (~w3905 & w8739);
assign v1839 = ~(w3833 | w3836);
assign w4228 = v1839;
assign w4229 = (~w3872 & ~w3874) | (~w3872 & w9147) | (~w3874 & w9147);
assign v1840 = ~(w4228 | w4229);
assign w4230 = v1840;
assign w4231 = w4228 & w4229;
assign v1841 = ~(w4230 | w4231);
assign w4232 = v1841;
assign w4233 = ~w4232 & w4227;
assign w4234 = (w3905 & w9148) | (w3905 & w9149) | (w9148 & w9149);
assign v1842 = ~(w4233 | w4234);
assign w4235 = v1842;
assign w4236 = w4226 & w4235;
assign v1843 = ~(w4226 | w4235);
assign w4237 = v1843;
assign v1844 = ~(w4236 | w4237);
assign w4238 = v1844;
assign w4239 = w4217 & ~w4238;
assign w4240 = ~w4217 & w4238;
assign v1845 = ~(w4239 | w4240);
assign w4241 = v1845;
assign v1846 = ~(w4177 | w4241);
assign w4242 = v1846;
assign w4243 = w4177 & w4241;
assign v1847 = ~(w4242 | w4243);
assign w4244 = v1847;
assign w4245 = (~w3990 & w3987) | (~w3990 & w9150) | (w3987 & w9150);
assign w4246 = (~w3922 & w3982) | (~w3922 & w8944) | (w3982 & w8944);
assign v1848 = ~(w3917 | w3919);
assign w4247 = v1848;
assign w4248 = (~w3978 & ~w3979) | (~w3978 & w8945) | (~w3979 & w8945);
assign w4249 = w4247 & w4248;
assign v1849 = ~(w4247 | w4248);
assign w4250 = v1849;
assign v1850 = ~(w4249 | w4250);
assign w4251 = v1850;
assign w4252 = w4246 & ~w4251;
assign w4253 = ~w4246 & w4251;
assign v1851 = ~(w4252 | w4253);
assign w4254 = v1851;
assign w4255 = w4245 & ~w4254;
assign w4256 = ~w4245 & w4254;
assign v1852 = ~(w4255 | w4256);
assign w4257 = v1852;
assign w4258 = w4244 & w4257;
assign v1853 = ~(w4244 | w4257);
assign w4259 = v1853;
assign v1854 = ~(w4258 | w4259);
assign w4260 = v1854;
assign v1855 = ~(w4012 | w4260);
assign w4261 = v1855;
assign w4262 = w4012 & w4260;
assign v1856 = ~(w4261 | w4262);
assign w4263 = v1856;
assign w4264 = w4011 & ~w4263;
assign w4265 = ~w4003 & w4263;
assign w4266 = ~w4006 & w4265;
assign v1857 = ~(w4264 | w4266);
assign w4267 = v1857;
assign w4268 = pi19 & pi45;
assign w4269 = pi23 & pi41;
assign w4270 = pi24 & pi40;
assign v1858 = ~(w4042 | w4270);
assign w4271 = v1858;
assign w4272 = pi25 & pi40;
assign w4273 = w3788 & w4272;
assign v1859 = ~(w4271 | w4273);
assign w4274 = v1859;
assign w4275 = w4269 & ~w4274;
assign w4276 = ~w4269 & w4274;
assign v1860 = ~(w4275 | w4276);
assign w4277 = v1860;
assign w4278 = w4268 & ~w4277;
assign w4279 = ~w4268 & w4277;
assign v1861 = ~(w4278 | w4279);
assign w4280 = v1861;
assign w4281 = pi20 & pi44;
assign w4282 = pi21 & pi43;
assign v1862 = ~(w4054 | w4282);
assign w4283 = v1862;
assign w4284 = pi22 & pi43;
assign w4285 = w3800 & w4284;
assign v1863 = ~(w4283 | w4285);
assign w4286 = v1863;
assign w4287 = w4281 & ~w4286;
assign w4288 = ~w4281 & w4286;
assign v1864 = ~(w4287 | w4288);
assign w4289 = v1864;
assign w4290 = w4280 & ~w4289;
assign w4291 = ~w4280 & w4289;
assign v1865 = ~(w4290 | w4291);
assign w4292 = v1865;
assign w4293 = pi26 & pi38;
assign w4294 = pi30 & pi34;
assign w4295 = pi31 & pi33;
assign w4296 = ~w4294 & w4295;
assign w4297 = w4294 & ~w4295;
assign v1866 = ~(w4296 | w4297);
assign w4298 = v1866;
assign w4299 = w4293 & ~w4298;
assign w4300 = ~w4293 & w4298;
assign v1867 = ~(w4299 | w4300);
assign w4301 = v1867;
assign w4302 = pi27 & pi37;
assign w4303 = pi28 & pi36;
assign v1868 = ~(w4078 | w4303);
assign w4304 = v1868;
assign w4305 = pi29 & pi36;
assign w4306 = w3824 & w4305;
assign v1869 = ~(w4304 | w4306);
assign w4307 = v1869;
assign w4308 = w4302 & ~w4307;
assign w4309 = ~w4302 & w4307;
assign v1870 = ~(w4308 | w4309);
assign w4310 = v1870;
assign w4311 = w4301 & ~w4310;
assign w4312 = ~w4301 & w4310;
assign v1871 = ~(w4311 | w4312);
assign w4313 = v1871;
assign w4314 = w4292 & w4313;
assign v1872 = ~(w4292 | w4313);
assign w4315 = v1872;
assign v1873 = ~(w4314 | w4315);
assign w4316 = v1873;
assign w4317 = pi12 & pi52;
assign w4318 = pi16 & pi48;
assign w4319 = pi17 & pi47;
assign v1874 = ~(w4017 | w4319);
assign w4320 = v1874;
assign w4321 = pi18 & pi47;
assign w4322 = w3763 & w4321;
assign v1875 = ~(w4320 | w4322);
assign w4323 = v1875;
assign w4324 = w4318 & ~w4323;
assign w4325 = ~w4318 & w4323;
assign v1876 = ~(w4324 | w4325);
assign w4326 = v1876;
assign w4327 = w4317 & ~w4326;
assign w4328 = ~w4317 & w4326;
assign v1877 = ~(w4327 | w4328);
assign w4329 = v1877;
assign w4330 = pi13 & pi51;
assign w4331 = pi14 & pi50;
assign v1878 = ~(w4029 | w4331);
assign w4332 = v1878;
assign w4333 = pi15 & pi50;
assign w4334 = w3775 & w4333;
assign v1879 = ~(w4332 | w4334);
assign w4335 = v1879;
assign w4336 = w4330 & ~w4335;
assign w4337 = ~w4330 & w4335;
assign v1880 = ~(w4336 | w4337);
assign w4338 = v1880;
assign w4339 = w4329 & ~w4338;
assign w4340 = ~w4329 & w4338;
assign v1881 = ~(w4339 | w4340);
assign w4341 = v1881;
assign w4342 = w4316 & w4341;
assign v1882 = ~(w4316 | w4341);
assign w4343 = v1882;
assign v1883 = ~(w4342 | w4343);
assign w4344 = v1883;
assign w4345 = pi05 & pi59;
assign w4346 = pi09 & pi55;
assign w4347 = pi10 & pi54;
assign v1884 = ~(w4097 | w4347);
assign w4348 = v1884;
assign w4349 = pi11 & pi54;
assign w4350 = w3882 & w4349;
assign v1885 = ~(w4348 | w4350);
assign w4351 = v1885;
assign w4352 = w4346 & ~w4351;
assign w4353 = ~w4346 & w4351;
assign v1886 = ~(w4352 | w4353);
assign w4354 = v1886;
assign w4355 = w4345 & ~w4354;
assign w4356 = ~w4345 & w4354;
assign v1887 = ~(w4355 | w4356);
assign w4357 = v1887;
assign w4358 = pi06 & pi58;
assign w4359 = pi07 & pi57;
assign v1888 = ~(w4109 | w4359);
assign w4360 = v1888;
assign w4361 = pi08 & pi57;
assign w4362 = w3894 & w4361;
assign v1889 = ~(w4360 | w4362);
assign w4363 = v1889;
assign w4364 = w4358 & ~w4363;
assign w4365 = ~w4358 & w4363;
assign v1890 = ~(w4364 | w4365);
assign w4366 = v1890;
assign w4367 = w4357 & ~w4366;
assign w4368 = ~w4357 & w4366;
assign v1891 = ~(w4367 | w4368);
assign w4369 = v1891;
assign w4370 = (~w4103 & ~w4105) | (~w4103 & w8621) | (~w4105 & w8621);
assign w4371 = w4106 & ~w4108;
assign v1892 = ~(w4110 | w4371);
assign w4372 = v1892;
assign w4373 = w4094 & ~w4096;
assign v1893 = ~(w4098 | w4373);
assign w4374 = v1893;
assign v1894 = ~(w4372 | w4374);
assign w4375 = v1894;
assign w4376 = w4372 & w4374;
assign v1895 = ~(w4375 | w4376);
assign w4377 = v1895;
assign w4378 = ~w4370 & w4377;
assign w4379 = w4370 & ~w4377;
assign v1896 = ~(w4378 | w4379);
assign w4380 = v1896;
assign w4381 = (~w4023 & ~w4025) | (~w4023 & w8622) | (~w4025 & w8622);
assign w4382 = w4026 & ~w4028;
assign v1897 = ~(w4030 | w4382);
assign w4383 = v1897;
assign w4384 = w4014 & ~w4016;
assign v1898 = ~(w4018 | w4384);
assign w4385 = v1898;
assign v1899 = ~(w4383 | w4385);
assign w4386 = v1899;
assign w4387 = w4383 & w4385;
assign v1900 = ~(w4386 | w4387);
assign w4388 = v1900;
assign w4389 = ~w4381 & w4388;
assign w4390 = w4381 & ~w4388;
assign v1901 = ~(w4389 | w4390);
assign w4391 = v1901;
assign w4392 = w4380 & w4391;
assign v1902 = ~(w4380 | w4391);
assign w4393 = v1902;
assign v1903 = ~(w4392 | w4393);
assign w4394 = v1903;
assign v1904 = ~(w4153 | w4165);
assign w4395 = v1904;
assign w4396 = w4156 & ~w4158;
assign v1905 = ~(w4160 | w4396);
assign w4397 = v1905;
assign v1906 = ~(w4395 | w4397);
assign w4398 = v1906;
assign w4399 = w4395 & w4397;
assign v1907 = ~(w4398 | w4399);
assign w4400 = v1907;
assign w4401 = w4394 & w4400;
assign v1908 = ~(w4394 | w4400);
assign w4402 = v1908;
assign v1909 = ~(w4401 | w4402);
assign w4403 = v1909;
assign w4404 = w4369 & w4403;
assign v1910 = ~(w4369 | w4403);
assign w4405 = v1910;
assign v1911 = ~(w4404 | w4405);
assign w4406 = v1911;
assign w4407 = w4344 & w4406;
assign v1912 = ~(w4344 | w4406);
assign w4408 = v1912;
assign v1913 = ~(w4407 | w4408);
assign w4409 = v1913;
assign w4410 = pi01 & pi63;
assign w4411 = pi02 & pi62;
assign w4412 = pi03 & pi61;
assign v1914 = ~(w4159 | w4412);
assign w4413 = v1914;
assign w4414 = pi04 & pi61;
assign w4415 = w3912 & w4414;
assign v1915 = ~(w4413 | w4415);
assign w4416 = v1915;
assign w4417 = w4411 & w4416;
assign v1916 = ~(w4411 | w4416);
assign w4418 = v1916;
assign v1917 = ~(w4417 | w4418);
assign w4419 = v1917;
assign w4420 = ~w4410 & w4419;
assign w4421 = w4410 & ~w4419;
assign v1918 = ~(w4420 | w4421);
assign w4422 = v1918;
assign w4423 = (w4422 & w4224) | (w4422 & w9151) | (w4224 & w9151);
assign w4424 = ~w4224 & w9152;
assign v1919 = ~(w4423 | w4424);
assign w4425 = v1919;
assign w4426 = (~w4230 & w4227) | (~w4230 & w8946) | (w4227 & w8946);
assign w4427 = w4425 & ~w4426;
assign w4428 = ~w4425 & w4426;
assign v1920 = ~(w4427 | w4428);
assign w4429 = v1920;
assign v1921 = ~(w4409 | w4429);
assign w4430 = v1921;
assign w4431 = w4409 & w4429;
assign v1922 = ~(w4430 | w4431);
assign w4432 = v1922;
assign w4433 = (~w4072 & ~w4074) | (~w4072 & w8623) | (~w4074 & w8623);
assign w4434 = (~w4066 & ~w4068) | (~w4066 & w8947) | (~w4068 & w8947);
assign w4435 = w4075 & ~w4077;
assign v1923 = ~(w4079 | w4435);
assign w4436 = v1923;
assign v1924 = ~(w4434 | w4436);
assign w4437 = v1924;
assign w4438 = w4434 & w4436;
assign v1925 = ~(w4437 | w4438);
assign w4439 = v1925;
assign w4440 = ~w4433 & w4439;
assign w4441 = w4433 & ~w4439;
assign v1926 = ~(w4440 | w4441);
assign w4442 = v1926;
assign w4443 = (~w4134 & w4129) | (~w4134 & w9153) | (w4129 & w9153);
assign w4444 = (~w4123 & w4118) | (~w4123 & w9154) | (w4118 & w9154);
assign v1927 = ~(w4443 | w4444);
assign w4445 = v1927;
assign w4446 = w4443 & w4444;
assign v1928 = ~(w4445 | w4446);
assign w4447 = v1928;
assign w4448 = w4442 & w4447;
assign v1929 = ~(w4442 | w4447);
assign w4449 = v1929;
assign v1930 = ~(w4448 | w4449);
assign w4450 = v1930;
assign w4451 = (~w4048 & ~w4050) | (~w4048 & w8624) | (~w4050 & w8624);
assign w4452 = w4051 & ~w4053;
assign v1931 = ~(w4055 | w4452);
assign w4453 = v1931;
assign w4454 = w4039 & ~w4041;
assign v1932 = ~(w4043 | w4454);
assign w4455 = v1932;
assign v1933 = ~(w4453 | w4455);
assign w4456 = v1933;
assign w4457 = w4453 & w4455;
assign v1934 = ~(w4456 | w4457);
assign w4458 = v1934;
assign w4459 = ~w4451 & w4458;
assign w4460 = w4451 & ~w4458;
assign v1935 = ~(w4459 | w4460);
assign w4461 = v1935;
assign w4462 = (~w4201 & w4196) | (~w4201 & w9155) | (w4196 & w9155);
assign w4463 = (~w4182 & w4178) | (~w4182 & w9156) | (w4178 & w9156);
assign w4464 = w4462 & w4463;
assign v1936 = ~(w4462 | w4463);
assign w4465 = v1936;
assign v1937 = ~(w4464 | w4465);
assign w4466 = v1937;
assign w4467 = w4461 & ~w4466;
assign w4468 = ~w4461 & w4466;
assign v1938 = ~(w4467 | w4468);
assign w4469 = v1938;
assign w4470 = w4450 & w4469;
assign v1939 = ~(w4450 | w4469);
assign w4471 = v1939;
assign v1940 = ~(w4470 | w4471);
assign w4472 = v1940;
assign v1941 = ~(w4212 | w4215);
assign w4473 = v1941;
assign w4474 = (~w4190 & ~w4192) | (~w4190 & w8948) | (~w4192 & w8948);
assign v1942 = ~(w4209 | w4474);
assign w4475 = v1942;
assign w4476 = w4209 & w4474;
assign v1943 = ~(w4475 | w4476);
assign w4477 = v1943;
assign w4478 = ~w4473 & w4477;
assign w4479 = w4473 & ~w4477;
assign v1944 = ~(w4478 | w4479);
assign w4480 = v1944;
assign w4481 = (~w4146 & ~w4148) | (~w4146 & w8740) | (~w4148 & w8740);
assign w4482 = (~w4087 & ~w4089) | (~w4087 & w9157) | (~w4089 & w9157);
assign v1945 = ~(w3913 | w4140);
assign w4483 = v1945;
assign v1946 = ~(w4141 | w4483);
assign w4484 = v1946;
assign w4485 = ~w4482 & w4484;
assign w4486 = w4482 & ~w4484;
assign v1947 = ~(w4485 | w4486);
assign w4487 = v1947;
assign w4488 = (~w4148 & w8949) | (~w4148 & w8950) | (w8949 & w8950);
assign w4489 = (w4148 & w8951) | (w4148 & w8952) | (w8951 & w8952);
assign v1948 = ~(w4488 | w4489);
assign w4490 = v1948;
assign v1949 = ~(w4480 | w4490);
assign w4491 = v1949;
assign w4492 = w4480 & w4490;
assign v1950 = ~(w4491 | w4492);
assign w4493 = v1950;
assign w4494 = w4472 & ~w4493;
assign w4495 = ~w4472 & w4493;
assign v1951 = ~(w4494 | w4495);
assign w4496 = v1951;
assign w4497 = w4432 & w4496;
assign v1952 = ~(w4432 | w4496);
assign w4498 = v1952;
assign v1953 = ~(w4497 | w4498);
assign w4499 = v1953;
assign w4500 = (~w4175 & ~w4241) | (~w4175 & w8953) | (~w4241 & w8953);
assign v1954 = ~(w4168 | w4172);
assign w4501 = v1954;
assign w4502 = (~w4237 & ~w4238) | (~w4237 & w8954) | (~w4238 & w8954);
assign w4503 = ~w4501 & w4502;
assign w4504 = w4501 & ~w4502;
assign v1955 = ~(w4503 | w4504);
assign w4505 = v1955;
assign w4506 = w4500 & w4505;
assign v1956 = ~(w4500 | w4505);
assign w4507 = v1956;
assign v1957 = ~(w4506 | w4507);
assign w4508 = v1957;
assign w4509 = (~w4249 & w4246) | (~w4249 & w9158) | (w4246 & w9158);
assign w4510 = w4508 & ~w4509;
assign w4511 = ~w4508 & w4509;
assign v1958 = ~(w4510 | w4511);
assign w4512 = v1958;
assign w4513 = ~w4499 & w4512;
assign w4514 = w4499 & ~w4512;
assign v1959 = ~(w4513 | w4514);
assign w4515 = v1959;
assign w4516 = (~w4255 & ~w4257) | (~w4255 & w9159) | (~w4257 & w9159);
assign w4517 = w4515 & w4516;
assign v1960 = ~(w4515 | w4516);
assign w4518 = v1960;
assign v1961 = ~(w4517 | w4518);
assign w4519 = v1961;
assign w4520 = (w8732 & w9270) | (w8732 & w9271) | (w9270 & w9271);
assign w4521 = ~w4262 & w9298;
assign w4522 = (~w4010 & w8955) | (~w4010 & w8956) | (w8955 & w8956);
assign v1962 = ~(w4519 | w4521);
assign w4523 = v1962;
assign v1963 = ~(w4522 | w4523);
assign w4524 = v1963;
assign w4525 = (w4010 & w9040) | (w4010 & w9041) | (w9040 & w9041);
assign w4526 = (~w4510 & ~w4512) | (~w4510 & w8786) | (~w4512 & w8786);
assign w4527 = pi16 & pi49;
assign w4528 = pi17 & pi48;
assign v1964 = ~(w4527 | w4528);
assign w4529 = v1964;
assign w4530 = pi17 & pi49;
assign w4531 = w4318 & w4530;
assign v1965 = ~(w4529 | w4531);
assign w4532 = v1965;
assign w4533 = w4333 & ~w4532;
assign w4534 = ~w4333 & w4532;
assign v1966 = ~(w4533 | w4534);
assign w4535 = v1966;
assign w4536 = w4349 & ~w4535;
assign w4537 = ~w4349 & w4535;
assign v1967 = ~(w4536 | w4537);
assign w4538 = v1967;
assign w4539 = pi12 & pi53;
assign w4540 = pi13 & pi52;
assign w4541 = pi14 & pi51;
assign v1968 = ~(w4540 | w4541);
assign w4542 = v1968;
assign w4543 = pi14 & pi52;
assign w4544 = w4330 & w4543;
assign v1969 = ~(w4542 | w4544);
assign w4545 = v1969;
assign w4546 = w4539 & ~w4545;
assign w4547 = ~w4539 & w4545;
assign v1970 = ~(w4546 | w4547);
assign w4548 = v1970;
assign w4549 = w4538 & ~w4548;
assign w4550 = ~w4538 & w4548;
assign v1971 = ~(w4549 | w4550);
assign w4551 = v1971;
assign w4552 = pi23 & pi42;
assign w4553 = pi24 & pi41;
assign v1972 = ~(w4552 | w4553);
assign w4554 = v1972;
assign w4555 = pi24 & pi42;
assign w4556 = w4269 & w4555;
assign v1973 = ~(w4554 | w4556);
assign w4557 = v1973;
assign w4558 = w4284 & ~w4557;
assign w4559 = ~w4284 & w4557;
assign v1974 = ~(w4558 | w4559);
assign w4560 = v1974;
assign w4561 = w4321 & ~w4560;
assign w4562 = ~w4321 & w4560;
assign v1975 = ~(w4561 | w4562);
assign w4563 = v1975;
assign w4564 = pi19 & pi46;
assign w4565 = pi20 & pi45;
assign w4566 = pi21 & pi44;
assign v1976 = ~(w4565 | w4566);
assign w4567 = v1976;
assign w4568 = pi21 & pi45;
assign w4569 = w4281 & w4568;
assign v1977 = ~(w4567 | w4569);
assign w4570 = v1977;
assign w4571 = w4564 & ~w4570;
assign w4572 = ~w4564 & w4570;
assign v1978 = ~(w4571 | w4572);
assign w4573 = v1978;
assign w4574 = w4563 & ~w4573;
assign w4575 = ~w4563 & w4573;
assign v1979 = ~(w4574 | w4575);
assign w4576 = v1979;
assign w4577 = pi31 & pi34;
assign w4578 = pi30 & pi35;
assign w4579 = ~w4577 & w4578;
assign w4580 = w4577 & ~w4578;
assign v1980 = ~(w4579 | w4580);
assign w4581 = v1980;
assign w4582 = w4305 & w4581;
assign v1981 = ~(w4305 | w4581);
assign w4583 = v1981;
assign v1982 = ~(w4582 | w4583);
assign w4584 = v1982;
assign w4585 = w4272 & w4584;
assign v1983 = ~(w4272 | w4584);
assign w4586 = v1983;
assign v1984 = ~(w4585 | w4586);
assign w4587 = v1984;
assign w4588 = pi26 & pi39;
assign w4589 = pi27 & pi38;
assign w4590 = pi28 & pi37;
assign v1985 = ~(w4589 | w4590);
assign w4591 = v1985;
assign w4592 = pi28 & pi38;
assign w4593 = w4302 & w4592;
assign v1986 = ~(w4591 | w4593);
assign w4594 = v1986;
assign w4595 = w4588 & ~w4594;
assign w4596 = ~w4588 & w4594;
assign v1987 = ~(w4595 | w4596);
assign w4597 = v1987;
assign w4598 = w4587 & ~w4597;
assign w4599 = ~w4587 & w4597;
assign v1988 = ~(w4598 | w4599);
assign w4600 = v1988;
assign w4601 = w4576 & w4600;
assign v1989 = ~(w4576 | w4600);
assign w4602 = v1989;
assign v1990 = ~(w4601 | w4602);
assign w4603 = v1990;
assign w4604 = w4551 & w4603;
assign v1991 = ~(w4551 | w4603);
assign w4605 = v1991;
assign v1992 = ~(w4604 | w4605);
assign w4606 = v1992;
assign w4607 = pi09 & pi56;
assign w4608 = pi10 & pi55;
assign v1993 = ~(w4607 | w4608);
assign w4609 = v1993;
assign w4610 = pi10 & pi56;
assign w4611 = w4346 & w4610;
assign v1994 = ~(w4609 | w4611);
assign w4612 = v1994;
assign w4613 = w4361 & ~w4612;
assign w4614 = ~w4361 & w4612;
assign v1995 = ~(w4613 | w4614);
assign w4615 = v1995;
assign w4616 = w4414 & ~w4615;
assign w4617 = ~w4414 & w4615;
assign v1996 = ~(w4616 | w4617);
assign w4618 = v1996;
assign w4619 = pi05 & pi60;
assign w4620 = pi06 & pi59;
assign w4621 = pi07 & pi58;
assign v1997 = ~(w4620 | w4621);
assign w4622 = v1997;
assign w4623 = pi07 & pi59;
assign w4624 = w4358 & w4623;
assign v1998 = ~(w4622 | w4624);
assign w4625 = v1998;
assign w4626 = w4619 & ~w4625;
assign w4627 = ~w4619 & w4625;
assign v1999 = ~(w4626 | w4627);
assign w4628 = v1999;
assign w4629 = w4618 & ~w4628;
assign w4630 = ~w4618 & w4628;
assign v2000 = ~(w4629 | w4630);
assign w4631 = v2000;
assign w4632 = w4415 & w4420;
assign v2001 = ~(w4415 | w4420);
assign w4633 = v2001;
assign v2002 = ~(w4632 | w4633);
assign w4634 = v2002;
assign v2003 = ~(w4417 | w4634);
assign w4635 = v2003;
assign w4636 = (~w4355 & ~w4357) | (~w4355 & w8741) | (~w4357 & w8741);
assign w4637 = w4358 & ~w4360;
assign v2004 = ~(w4362 | w4637);
assign w4638 = v2004;
assign w4639 = w4346 & ~w4348;
assign v2005 = ~(w4350 | w4639);
assign w4640 = v2005;
assign v2006 = ~(w4638 | w4640);
assign w4641 = v2006;
assign w4642 = w4638 & w4640;
assign v2007 = ~(w4641 | w4642);
assign w4643 = v2007;
assign w4644 = ~w4636 & w4643;
assign w4645 = w4636 & ~w4643;
assign v2008 = ~(w4644 | w4645);
assign w4646 = v2008;
assign w4647 = (~w4327 & ~w4329) | (~w4327 & w8742) | (~w4329 & w8742);
assign w4648 = w4330 & ~w4332;
assign v2009 = ~(w4334 | w4648);
assign w4649 = v2009;
assign w4650 = w4318 & ~w4320;
assign v2010 = ~(w4322 | w4650);
assign w4651 = v2010;
assign v2011 = ~(w4649 | w4651);
assign w4652 = v2011;
assign w4653 = w4649 & w4651;
assign v2012 = ~(w4652 | w4653);
assign w4654 = v2012;
assign w4655 = ~w4647 & w4654;
assign w4656 = w4647 & ~w4654;
assign v2013 = ~(w4655 | w4656);
assign w4657 = v2013;
assign w4658 = w4646 & w4657;
assign v2014 = ~(w4646 | w4657);
assign w4659 = v2014;
assign v2015 = ~(w4658 | w4659);
assign w4660 = v2015;
assign w4661 = ~w4635 & w4660;
assign w4662 = w4635 & ~w4660;
assign v2016 = ~(w4661 | w4662);
assign w4663 = v2016;
assign v2017 = ~(w4631 | w4663);
assign w4664 = v2017;
assign w4665 = w4631 & w4663;
assign v2018 = ~(w4664 | w4665);
assign w4666 = v2018;
assign w4667 = ~w4606 & w4666;
assign w4668 = w4606 & ~w4666;
assign v2019 = ~(w4667 | w4668);
assign w4669 = v2019;
assign w4670 = pi02 & pi63;
assign w4671 = pi03 & pi62;
assign w4672 = w4670 & ~w4671;
assign w4673 = ~w4670 & w4671;
assign v2020 = ~(w4672 | w4673);
assign w4674 = v2020;
assign w4675 = (~w4674 & w8787) | (~w4674 & w4478) | (w8787 & w4478);
assign w4676 = (w8788 & w4473) | (w8788 & w8957) | (w4473 & w8957);
assign v2021 = ~(w4675 | w4676);
assign w4677 = v2021;
assign w4678 = (~w4485 & ~w4481) | (~w4485 & w8789) | (~w4481 & w8789);
assign w4679 = w4677 & ~w4678;
assign w4680 = ~w4677 & w4678;
assign v2022 = ~(w4679 | w4680);
assign w4681 = v2022;
assign w4682 = ~w4669 & w4681;
assign w4683 = w4669 & ~w4681;
assign v2023 = ~(w4682 | w4683);
assign w4684 = v2023;
assign v2024 = ~(w4299 | w4311);
assign w4685 = v2024;
assign w4686 = w4302 & ~w4304;
assign v2025 = ~(w4306 | w4686);
assign w4687 = v2025;
assign v2026 = ~(w4296 | w4687);
assign w4688 = v2026;
assign w4689 = w4296 & w4687;
assign v2027 = ~(w4688 | w4689);
assign w4690 = v2027;
assign w4691 = ~w4685 & w4690;
assign w4692 = w4685 & ~w4690;
assign v2028 = ~(w4691 | w4692);
assign w4693 = v2028;
assign w4694 = (~w4375 & w4370) | (~w4375 & w8958) | (w4370 & w8958);
assign w4695 = w4398 & ~w4694;
assign w4696 = ~w4398 & w4694;
assign v2029 = ~(w4695 | w4696);
assign w4697 = v2029;
assign w4698 = w4693 & w4697;
assign v2030 = ~(w4693 | w4697);
assign w4699 = v2030;
assign v2031 = ~(w4698 | w4699);
assign w4700 = v2031;
assign w4701 = (~w4278 & ~w4280) | (~w4278 & w8625) | (~w4280 & w8625);
assign w4702 = w4281 & ~w4283;
assign v2032 = ~(w4285 | w4702);
assign w4703 = v2032;
assign w4704 = w4269 & ~w4271;
assign v2033 = ~(w4273 | w4704);
assign w4705 = v2033;
assign v2034 = ~(w4703 | w4705);
assign w4706 = v2034;
assign w4707 = w4703 & w4705;
assign v2035 = ~(w4706 | w4707);
assign w4708 = v2035;
assign w4709 = ~w4701 & w4708;
assign w4710 = w4701 & ~w4708;
assign v2036 = ~(w4709 | w4710);
assign w4711 = v2036;
assign v2037 = ~(w4386 | w4389);
assign w4712 = v2037;
assign w4713 = (~w4437 & w4433) | (~w4437 & w8743) | (w4433 & w8743);
assign w4714 = (~w4456 & w4451) | (~w4456 & w8744) | (w4451 & w8744);
assign v2038 = ~(w4713 | w4714);
assign w4715 = v2038;
assign w4716 = w4713 & w4714;
assign v2039 = ~(w4715 | w4716);
assign w4717 = v2039;
assign w4718 = ~w4712 & w4717;
assign w4719 = w4712 & ~w4717;
assign v2040 = ~(w4718 | w4719);
assign w4720 = v2040;
assign w4721 = w4711 & w4720;
assign v2041 = ~(w4711 | w4720);
assign w4722 = v2041;
assign v2042 = ~(w4721 | w4722);
assign w4723 = v2042;
assign w4724 = w4700 & w4723;
assign v2043 = ~(w4700 | w4723);
assign w4725 = v2043;
assign v2044 = ~(w4724 | w4725);
assign w4726 = v2044;
assign v2045 = ~(w4467 | w4470);
assign w4727 = v2045;
assign w4728 = (~w4445 & ~w4447) | (~w4445 & w8790) | (~w4447 & w8790);
assign v2046 = ~(w4464 | w4728);
assign w4729 = v2046;
assign w4730 = w4464 & w4728;
assign v2047 = ~(w4729 | w4730);
assign w4731 = v2047;
assign w4732 = ~w4727 & w4731;
assign w4733 = w4727 & ~w4731;
assign v2048 = ~(w4732 | w4733);
assign w4734 = v2048;
assign w4735 = (~w4404 & ~w4406) | (~w4404 & w8745) | (~w4406 & w8745);
assign v2049 = ~(w4314 | w4342);
assign w4736 = v2049;
assign v2050 = ~(w4392 | w4401);
assign w4737 = v2050;
assign v2051 = ~(w4736 | w4737);
assign w4738 = v2051;
assign w4739 = w4736 & w4737;
assign v2052 = ~(w4738 | w4739);
assign w4740 = v2052;
assign w4741 = ~w4735 & w4740;
assign w4742 = w4735 & ~w4740;
assign v2053 = ~(w4741 | w4742);
assign w4743 = v2053;
assign w4744 = w4734 & w4743;
assign v2054 = ~(w4734 | w4743);
assign w4745 = v2054;
assign v2055 = ~(w4744 | w4745);
assign w4746 = v2055;
assign w4747 = w4726 & ~w4746;
assign w4748 = ~w4726 & w4746;
assign v2056 = ~(w4747 | w4748);
assign w4749 = v2056;
assign w4750 = w4684 & ~w4749;
assign w4751 = ~w4684 & w4749;
assign v2057 = ~(w4750 | w4751);
assign w4752 = v2057;
assign w4753 = (~w4503 & ~w4500) | (~w4503 & w9160) | (~w4500 & w9160);
assign v2058 = ~(w4430 | w4497);
assign w4754 = v2058;
assign v2059 = ~(w4423 | w4427);
assign w4755 = v2059;
assign w4756 = (~w4491 & ~w4493) | (~w4491 & w8791) | (~w4493 & w8791);
assign w4757 = ~w4755 & w4756;
assign w4758 = w4755 & ~w4756;
assign v2060 = ~(w4757 | w4758);
assign w4759 = v2060;
assign w4760 = w4754 & w4759;
assign v2061 = ~(w4754 | w4759);
assign w4761 = v2061;
assign v2062 = ~(w4760 | w4761);
assign w4762 = v2062;
assign w4763 = ~w4753 & w4762;
assign w4764 = w4753 & ~w4762;
assign v2063 = ~(w4763 | w4764);
assign w4765 = v2063;
assign w4766 = w4752 & w4765;
assign v2064 = ~(w4752 | w4765);
assign w4767 = v2064;
assign v2065 = ~(w4766 | w4767);
assign w4768 = v2065;
assign w4769 = w4526 & ~w4768;
assign w4770 = ~w4526 & w4768;
assign v2066 = ~(w4769 | w4770);
assign w4771 = v2066;
assign w4772 = w4525 & ~w4771;
assign w4773 = ~w4525 & w4771;
assign v2067 = ~(w4772 | w4773);
assign w4774 = v2067;
assign w4775 = (~w4763 & ~w4765) | (~w4763 & w8792) | (~w4765 & w8792);
assign w4776 = pi11 & pi55;
assign w4777 = pi15 & pi51;
assign w4778 = pi16 & pi50;
assign v2068 = ~(w4530 | w4778);
assign w4779 = v2068;
assign w4780 = pi17 & pi50;
assign w4781 = w4527 & w4780;
assign v2069 = ~(w4779 | w4781);
assign w4782 = v2069;
assign w4783 = w4777 & ~w4782;
assign w4784 = ~w4777 & w4782;
assign v2070 = ~(w4783 | w4784);
assign w4785 = v2070;
assign w4786 = w4776 & ~w4785;
assign w4787 = ~w4776 & w4785;
assign v2071 = ~(w4786 | w4787);
assign w4788 = v2071;
assign w4789 = pi12 & pi54;
assign w4790 = pi13 & pi53;
assign v2072 = ~(w4543 | w4790);
assign w4791 = v2072;
assign w4792 = pi14 & pi53;
assign w4793 = w4540 & w4792;
assign v2073 = ~(w4791 | w4793);
assign w4794 = v2073;
assign w4795 = w4789 & ~w4794;
assign w4796 = ~w4789 & w4794;
assign v2074 = ~(w4795 | w4796);
assign w4797 = v2074;
assign w4798 = w4788 & ~w4797;
assign w4799 = ~w4788 & w4797;
assign v2075 = ~(w4798 | w4799);
assign w4800 = v2075;
assign w4801 = pi18 & pi48;
assign w4802 = pi22 & pi44;
assign w4803 = pi23 & pi43;
assign v2076 = ~(w4555 | w4803);
assign w4804 = v2076;
assign w4805 = pi24 & pi43;
assign w4806 = w4552 & w4805;
assign v2077 = ~(w4804 | w4806);
assign w4807 = v2077;
assign w4808 = w4802 & ~w4807;
assign w4809 = ~w4802 & w4807;
assign v2078 = ~(w4808 | w4809);
assign w4810 = v2078;
assign w4811 = w4801 & ~w4810;
assign w4812 = ~w4801 & w4810;
assign v2079 = ~(w4811 | w4812);
assign w4813 = v2079;
assign w4814 = pi19 & pi47;
assign w4815 = pi20 & pi46;
assign v2080 = ~(w4568 | w4815);
assign w4816 = v2080;
assign w4817 = pi21 & pi46;
assign w4818 = w4565 & w4817;
assign v2081 = ~(w4816 | w4818);
assign w4819 = v2081;
assign w4820 = w4814 & ~w4819;
assign w4821 = ~w4814 & w4819;
assign v2082 = ~(w4820 | w4821);
assign w4822 = v2082;
assign w4823 = w4813 & ~w4822;
assign w4824 = ~w4813 & w4822;
assign v2083 = ~(w4823 | w4824);
assign w4825 = v2083;
assign w4826 = pi25 & pi41;
assign w4827 = pi29 & pi37;
assign w4828 = pi31 & pi35;
assign w4829 = pi30 & pi36;
assign w4830 = ~w4828 & w4829;
assign w4831 = w4828 & ~w4829;
assign v2084 = ~(w4830 | w4831);
assign w4832 = v2084;
assign w4833 = w4827 & w4832;
assign v2085 = ~(w4827 | w4832);
assign w4834 = v2085;
assign v2086 = ~(w4833 | w4834);
assign w4835 = v2086;
assign w4836 = w4826 & w4835;
assign v2087 = ~(w4826 | w4835);
assign w4837 = v2087;
assign v2088 = ~(w4836 | w4837);
assign w4838 = v2088;
assign w4839 = pi26 & pi40;
assign w4840 = pi27 & pi39;
assign v2089 = ~(w4592 | w4840);
assign w4841 = v2089;
assign w4842 = pi28 & pi39;
assign w4843 = w4589 & w4842;
assign v2090 = ~(w4841 | w4843);
assign w4844 = v2090;
assign w4845 = w4839 & ~w4844;
assign w4846 = ~w4839 & w4844;
assign v2091 = ~(w4845 | w4846);
assign w4847 = v2091;
assign w4848 = w4838 & ~w4847;
assign w4849 = ~w4838 & w4847;
assign v2092 = ~(w4848 | w4849);
assign w4850 = v2092;
assign w4851 = w4825 & w4850;
assign v2093 = ~(w4825 | w4850);
assign w4852 = v2093;
assign v2094 = ~(w4851 | w4852);
assign w4853 = v2094;
assign w4854 = w4800 & w4853;
assign v2095 = ~(w4800 | w4853);
assign w4855 = v2095;
assign v2096 = ~(w4854 | w4855);
assign w4856 = v2096;
assign w4857 = (~w4616 & ~w4618) | (~w4616 & w8746) | (~w4618 & w8746);
assign w4858 = w4619 & ~w4622;
assign v2097 = ~(w4624 | w4858);
assign w4859 = v2097;
assign w4860 = w4361 & ~w4609;
assign v2098 = ~(w4611 | w4860);
assign w4861 = v2098;
assign v2099 = ~(w4859 | w4861);
assign w4862 = v2099;
assign w4863 = w4859 & w4861;
assign v2100 = ~(w4862 | w4863);
assign w4864 = v2100;
assign w4865 = ~w4857 & w4864;
assign w4866 = w4857 & ~w4864;
assign v2101 = ~(w4865 | w4866);
assign w4867 = v2101;
assign w4868 = (~w4536 & ~w4538) | (~w4536 & w8626) | (~w4538 & w8626);
assign w4869 = w4539 & ~w4542;
assign v2102 = ~(w4544 | w4869);
assign w4870 = v2102;
assign w4871 = w4333 & ~w4529;
assign v2103 = ~(w4531 | w4871);
assign w4872 = v2103;
assign v2104 = ~(w4870 | w4872);
assign w4873 = v2104;
assign w4874 = w4870 & w4872;
assign v2105 = ~(w4873 | w4874);
assign w4875 = v2105;
assign w4876 = ~w4868 & w4875;
assign w4877 = w4868 & ~w4875;
assign v2106 = ~(w4876 | w4877);
assign w4878 = v2106;
assign w4879 = w4867 & w4878;
assign v2107 = ~(w4867 | w4878);
assign w4880 = v2107;
assign v2108 = ~(w4879 | w4880);
assign w4881 = v2108;
assign w4882 = ~w4672 & w4881;
assign w4883 = w4672 & ~w4881;
assign v2109 = ~(w4882 | w4883);
assign w4884 = v2109;
assign w4885 = pi04 & pi62;
assign w4886 = pi08 & pi58;
assign w4887 = pi09 & pi57;
assign v2110 = ~(w4610 | w4887);
assign w4888 = v2110;
assign w4889 = pi10 & pi57;
assign w4890 = w4607 & w4889;
assign v2111 = ~(w4888 | w4890);
assign w4891 = v2111;
assign w4892 = w4886 & ~w4891;
assign w4893 = ~w4886 & w4891;
assign v2112 = ~(w4892 | w4893);
assign w4894 = v2112;
assign w4895 = w4885 & ~w4894;
assign w4896 = ~w4885 & w4894;
assign v2113 = ~(w4895 | w4896);
assign w4897 = v2113;
assign w4898 = pi05 & pi61;
assign w4899 = pi06 & pi60;
assign v2114 = ~(w4623 | w4899);
assign w4900 = v2114;
assign w4901 = pi07 & pi60;
assign w4902 = w4620 & w4901;
assign v2115 = ~(w4900 | w4902);
assign w4903 = v2115;
assign w4904 = w4898 & ~w4903;
assign w4905 = ~w4898 & w4903;
assign v2116 = ~(w4904 | w4905);
assign w4906 = v2116;
assign w4907 = w4897 & ~w4906;
assign w4908 = ~w4897 & w4906;
assign v2117 = ~(w4907 | w4908);
assign w4909 = v2117;
assign w4910 = w4884 & w4909;
assign v2118 = ~(w4884 | w4909);
assign w4911 = v2118;
assign v2119 = ~(w4910 | w4911);
assign w4912 = v2119;
assign w4913 = w4856 & w4912;
assign v2120 = ~(w4856 | w4912);
assign w4914 = v2120;
assign v2121 = ~(w4913 | w4914);
assign w4915 = v2121;
assign w4916 = (~w4738 & w4735) | (~w4738 & w9042) | (w4735 & w9042);
assign w4917 = pi03 & pi63;
assign w4918 = (~w4729 & w4727) | (~w4729 & w8793) | (w4727 & w8793);
assign w4919 = w4917 & ~w4918;
assign w4920 = ~w4917 & w4918;
assign v2122 = ~(w4919 | w4920);
assign w4921 = v2122;
assign w4922 = ~w4916 & w4921;
assign w4923 = w4916 & ~w4921;
assign v2123 = ~(w4922 | w4923);
assign w4924 = v2123;
assign w4925 = w4915 & w4924;
assign v2124 = ~(w4915 | w4924);
assign w4926 = v2124;
assign v2125 = ~(w4925 | w4926);
assign w4927 = v2125;
assign w4928 = (~w4585 & ~w4587) | (~w4585 & w8627) | (~w4587 & w8627);
assign w4929 = (~w4579 & ~w4581) | (~w4579 & w8794) | (~w4581 & w8794);
assign w4930 = w4588 & ~w4591;
assign v2126 = ~(w4593 | w4930);
assign w4931 = v2126;
assign v2127 = ~(w4929 | w4931);
assign w4932 = v2127;
assign w4933 = w4929 & w4931;
assign v2128 = ~(w4932 | w4933);
assign w4934 = v2128;
assign w4935 = ~w4928 & w4934;
assign w4936 = w4928 & ~w4934;
assign v2129 = ~(w4935 | w4936);
assign w4937 = v2129;
assign w4938 = (~w4641 & w4636) | (~w4641 & w9043) | (w4636 & w9043);
assign w4939 = w4632 & ~w4938;
assign w4940 = ~w4632 & w4938;
assign v2130 = ~(w4939 | w4940);
assign w4941 = v2130;
assign w4942 = w4937 & w4941;
assign v2131 = ~(w4937 | w4941);
assign w4943 = v2131;
assign v2132 = ~(w4942 | w4943);
assign w4944 = v2132;
assign w4945 = (~w4561 & ~w4563) | (~w4561 & w8628) | (~w4563 & w8628);
assign w4946 = w4564 & ~w4567;
assign v2133 = ~(w4569 | w4946);
assign w4947 = v2133;
assign w4948 = w4284 & ~w4554;
assign v2134 = ~(w4556 | w4948);
assign w4949 = v2134;
assign v2135 = ~(w4947 | w4949);
assign w4950 = v2135;
assign w4951 = w4947 & w4949;
assign v2136 = ~(w4950 | w4951);
assign w4952 = v2136;
assign w4953 = ~w4945 & w4952;
assign w4954 = w4945 & ~w4952;
assign v2137 = ~(w4953 | w4954);
assign w4955 = v2137;
assign v2138 = ~(w4652 | w4655);
assign w4956 = v2138;
assign w4957 = (~w4688 & w4685) | (~w4688 & w8795) | (w4685 & w8795);
assign w4958 = (~w4706 & w4701) | (~w4706 & w8747) | (w4701 & w8747);
assign v2139 = ~(w4957 | w4958);
assign w4959 = v2139;
assign w4960 = w4957 & w4958;
assign v2140 = ~(w4959 | w4960);
assign w4961 = v2140;
assign w4962 = ~w4956 & w4961;
assign w4963 = w4956 & ~w4961;
assign v2141 = ~(w4962 | w4963);
assign w4964 = v2141;
assign w4965 = w4955 & w4964;
assign v2142 = ~(w4955 | w4964);
assign w4966 = v2142;
assign v2143 = ~(w4965 | w4966);
assign w4967 = v2143;
assign w4968 = w4944 & w4967;
assign v2144 = ~(w4944 | w4967);
assign w4969 = v2144;
assign v2145 = ~(w4968 | w4969);
assign w4970 = v2145;
assign w4971 = (~w4721 & ~w4723) | (~w4721 & w8796) | (~w4723 & w8796);
assign w4972 = (~w4695 & ~w4697) | (~w4695 & w9044) | (~w4697 & w9044);
assign w4973 = (~w4715 & ~w4717) | (~w4715 & w9045) | (~w4717 & w9045);
assign v2146 = ~(w4972 | w4973);
assign w4974 = v2146;
assign w4975 = w4972 & w4973;
assign v2147 = ~(w4974 | w4975);
assign w4976 = v2147;
assign w4977 = ~w4971 & w4976;
assign w4978 = w4971 & ~w4976;
assign v2148 = ~(w4977 | w4978);
assign w4979 = v2148;
assign w4980 = (~w4664 & ~w4666) | (~w4664 & w8797) | (~w4666 & w8797);
assign v2149 = ~(w4601 | w4604);
assign w4981 = v2149;
assign v2150 = ~(w4658 | w4661);
assign w4982 = v2150;
assign v2151 = ~(w4981 | w4982);
assign w4983 = v2151;
assign w4984 = w4981 & w4982;
assign v2152 = ~(w4983 | w4984);
assign w4985 = v2152;
assign w4986 = w4980 & w4985;
assign v2153 = ~(w4980 | w4985);
assign w4987 = v2153;
assign v2154 = ~(w4986 | w4987);
assign w4988 = v2154;
assign v2155 = ~(w4979 | w4988);
assign w4989 = v2155;
assign w4990 = w4979 & w4988;
assign v2156 = ~(w4989 | w4990);
assign w4991 = v2156;
assign w4992 = w4970 & w4991;
assign v2157 = ~(w4970 | w4991);
assign w4993 = v2157;
assign v2158 = ~(w4992 | w4993);
assign w4994 = v2158;
assign w4995 = w4927 & w4994;
assign v2159 = ~(w4927 | w4994);
assign w4996 = v2159;
assign v2160 = ~(w4995 | w4996);
assign w4997 = v2160;
assign w4998 = (~w4757 & ~w4754) | (~w4757 & w8798) | (~w4754 & w8798);
assign w4999 = (~w4682 & w4749) | (~w4682 & w8799) | (w4749 & w8799);
assign w5000 = (~w4675 & w4678) | (~w4675 & w9046) | (w4678 & w9046);
assign w5001 = ~w5000 & w9299;
assign w5002 = (w4746 & w8959) | (w4746 & w8960) | (w8959 & w8960);
assign v2161 = ~(w5001 | w5002);
assign w5003 = v2161;
assign w5004 = ~w4999 & w5003;
assign w5005 = w4999 & ~w5003;
assign v2162 = ~(w5004 | w5005);
assign w5006 = v2162;
assign w5007 = ~w4998 & w5006;
assign w5008 = w4998 & ~w5006;
assign v2163 = ~(w5007 | w5008);
assign w5009 = v2163;
assign w5010 = w4997 & w5009;
assign v2164 = ~(w4997 | w5009);
assign w5011 = v2164;
assign v2165 = ~(w5010 | w5011);
assign w5012 = v2165;
assign w5013 = ~w4775 & w5012;
assign w5014 = w4775 & ~w5012;
assign v2166 = ~(w5013 | w5014);
assign w5015 = v2166;
assign w5016 = (~w4769 & w9047) | (~w4769 & ~w4525) | (w9047 & ~w4525);
assign w5017 = (~w4010 & w9272) | (~w4010 & w9273) | (w9272 & w9273);
assign v2167 = ~(w5015 | w5016);
assign w5018 = v2167;
assign v2168 = ~(w5017 | w5018);
assign w5019 = v2168;
assign v2169 = ~(w5013 | w5017);
assign w5020 = v2169;
assign w5021 = (~w5007 & ~w5009) | (~w5007 & w8961) | (~w5009 & w8961);
assign w5022 = (~w5001 & w4999) | (~w5001 & w8962) | (w4999 & w8962);
assign v2170 = ~(w4862 | w4865);
assign w5023 = v2170;
assign w5024 = (~w4950 & w4945) | (~w4950 & w8748) | (w4945 & w8748);
assign w5025 = (~w4873 & w4868) | (~w4873 & w8749) | (w4868 & w8749);
assign v2171 = ~(w5024 | w5025);
assign w5026 = v2171;
assign w5027 = w5024 & w5025;
assign v2172 = ~(w5026 | w5027);
assign w5028 = v2172;
assign w5029 = ~w5023 & w5028;
assign w5030 = w5023 & ~w5028;
assign v2173 = ~(w5029 | w5030);
assign w5031 = v2173;
assign w5032 = (~w4836 & ~w4838) | (~w4836 & w8629) | (~w4838 & w8629);
assign v2174 = ~(w4830 | w4833);
assign w5033 = v2174;
assign w5034 = w4839 & ~w4841;
assign v2175 = ~(w4843 | w5034);
assign w5035 = v2175;
assign v2176 = ~(w5033 | w5035);
assign w5036 = v2176;
assign w5037 = w5033 & w5035;
assign v2177 = ~(w5036 | w5037);
assign w5038 = v2177;
assign w5039 = ~w5032 & w5038;
assign w5040 = w5032 & ~w5038;
assign v2178 = ~(w5039 | w5040);
assign w5041 = v2178;
assign w5042 = pi04 & pi63;
assign w5043 = (w4928 & w8801) | (w4928 & w8802) | (w8801 & w8802);
assign w5044 = ~w5042 & w9300;
assign v2179 = ~(w5043 | w5044);
assign w5045 = v2179;
assign w5046 = w5041 & ~w5045;
assign w5047 = ~w5041 & w5045;
assign v2180 = ~(w5046 | w5047);
assign w5048 = v2180;
assign w5049 = w5031 & w5048;
assign v2181 = ~(w5031 | w5048);
assign w5050 = v2181;
assign v2182 = ~(w5049 | w5050);
assign w5051 = v2182;
assign w5052 = (~w4910 & ~w4912) | (~w4910 & w8803) | (~w4912 & w8803);
assign v2183 = ~(w4851 | w4854);
assign w5053 = v2183;
assign v2184 = ~(w4879 | w4882);
assign w5054 = v2184;
assign v2185 = ~(w5053 | w5054);
assign w5055 = v2185;
assign w5056 = w5053 & w5054;
assign v2186 = ~(w5055 | w5056);
assign w5057 = v2186;
assign w5058 = ~w5052 & w5057;
assign w5059 = w5052 & ~w5057;
assign v2187 = ~(w5058 | w5059);
assign w5060 = v2187;
assign w5061 = (~w4965 & ~w4967) | (~w4965 & w8804) | (~w4967 & w8804);
assign v2188 = ~(w4939 | w4942);
assign w5062 = v2188;
assign v2189 = ~(w4959 | w4962);
assign w5063 = v2189;
assign v2190 = ~(w5062 | w5063);
assign w5064 = v2190;
assign w5065 = w5062 & w5063;
assign v2191 = ~(w5064 | w5065);
assign w5066 = v2191;
assign w5067 = ~w5061 & w5066;
assign w5068 = w5061 & ~w5066;
assign v2192 = ~(w5067 | w5068);
assign w5069 = v2192;
assign w5070 = w5060 & w5069;
assign v2193 = ~(w5060 | w5069);
assign w5071 = v2193;
assign v2194 = ~(w5070 | w5071);
assign w5072 = v2194;
assign w5073 = w5051 & w5072;
assign v2195 = ~(w5051 | w5072);
assign w5074 = v2195;
assign v2196 = ~(w5073 | w5074);
assign w5075 = v2196;
assign w5076 = pi25 & pi42;
assign w5077 = pi29 & pi38;
assign w5078 = pi31 & pi36;
assign w5079 = pi30 & pi37;
assign w5080 = ~w5078 & w5079;
assign w5081 = w5078 & ~w5079;
assign v2197 = ~(w5080 | w5081);
assign w5082 = v2197;
assign w5083 = w5077 & w5082;
assign v2198 = ~(w5077 | w5082);
assign w5084 = v2198;
assign v2199 = ~(w5083 | w5084);
assign w5085 = v2199;
assign w5086 = w5076 & w5085;
assign v2200 = ~(w5076 | w5085);
assign w5087 = v2200;
assign v2201 = ~(w5086 | w5087);
assign w5088 = v2201;
assign w5089 = pi26 & pi41;
assign w5090 = pi27 & pi40;
assign v2202 = ~(w4842 | w5090);
assign w5091 = v2202;
assign w5092 = pi28 & pi40;
assign w5093 = w4840 & w5092;
assign v2203 = ~(w5091 | w5093);
assign w5094 = v2203;
assign w5095 = w5089 & ~w5094;
assign w5096 = ~w5089 & w5094;
assign v2204 = ~(w5095 | w5096);
assign w5097 = v2204;
assign w5098 = w5088 & ~w5097;
assign w5099 = ~w5088 & w5097;
assign v2205 = ~(w5098 | w5099);
assign w5100 = v2205;
assign w5101 = ~w4917 & w5100;
assign w5102 = w4917 & ~w5100;
assign v2206 = ~(w5101 | w5102);
assign w5103 = v2206;
assign w5104 = pi18 & pi49;
assign w5105 = pi22 & pi45;
assign w5106 = pi23 & pi44;
assign v2207 = ~(w4805 | w5106);
assign w5107 = v2207;
assign w5108 = pi24 & pi44;
assign w5109 = w4803 & w5108;
assign v2208 = ~(w5107 | w5109);
assign w5110 = v2208;
assign w5111 = w5105 & ~w5110;
assign w5112 = ~w5105 & w5110;
assign v2209 = ~(w5111 | w5112);
assign w5113 = v2209;
assign w5114 = w5104 & ~w5113;
assign w5115 = ~w5104 & w5113;
assign v2210 = ~(w5114 | w5115);
assign w5116 = v2210;
assign w5117 = pi19 & pi48;
assign w5118 = pi20 & pi47;
assign v2211 = ~(w4817 | w5118);
assign w5119 = v2211;
assign w5120 = pi21 & pi47;
assign w5121 = w4815 & w5120;
assign v2212 = ~(w5119 | w5121);
assign w5122 = v2212;
assign w5123 = w5117 & ~w5122;
assign w5124 = ~w5117 & w5122;
assign v2213 = ~(w5123 | w5124);
assign w5125 = v2213;
assign w5126 = w5116 & ~w5125;
assign w5127 = ~w5116 & w5125;
assign v2214 = ~(w5126 | w5127);
assign w5128 = v2214;
assign w5129 = w5103 & w5128;
assign v2215 = ~(w5103 | w5128);
assign w5130 = v2215;
assign v2216 = ~(w5129 | w5130);
assign w5131 = v2216;
assign w5132 = pi11 & pi56;
assign w5133 = pi15 & pi52;
assign w5134 = pi16 & pi51;
assign v2217 = ~(w4780 | w5134);
assign w5135 = v2217;
assign w5136 = pi17 & pi51;
assign w5137 = w4778 & w5136;
assign v2218 = ~(w5135 | w5137);
assign w5138 = v2218;
assign w5139 = w5133 & ~w5138;
assign w5140 = ~w5133 & w5138;
assign v2219 = ~(w5139 | w5140);
assign w5141 = v2219;
assign w5142 = w5132 & ~w5141;
assign w5143 = ~w5132 & w5141;
assign v2220 = ~(w5142 | w5143);
assign w5144 = v2220;
assign w5145 = pi12 & pi55;
assign w5146 = pi13 & pi54;
assign v2221 = ~(w4792 | w5146);
assign w5147 = v2221;
assign w5148 = pi14 & pi54;
assign w5149 = w4790 & w5148;
assign v2222 = ~(w5147 | w5149);
assign w5150 = v2222;
assign w5151 = w5145 & ~w5150;
assign w5152 = ~w5145 & w5150;
assign v2223 = ~(w5151 | w5152);
assign w5153 = v2223;
assign w5154 = w5144 & ~w5153;
assign w5155 = ~w5144 & w5153;
assign v2224 = ~(w5154 | w5155);
assign w5156 = v2224;
assign v2225 = ~(w4895 | w4907);
assign w5157 = v2225;
assign w5158 = w4898 & ~w4900;
assign v2226 = ~(w4902 | w5158);
assign w5159 = v2226;
assign w5160 = w4886 & ~w4888;
assign v2227 = ~(w4890 | w5160);
assign w5161 = v2227;
assign v2228 = ~(w5159 | w5161);
assign w5162 = v2228;
assign w5163 = w5159 & w5161;
assign v2229 = ~(w5162 | w5163);
assign w5164 = v2229;
assign w5165 = ~w5157 & w5164;
assign w5166 = w5157 & ~w5164;
assign v2230 = ~(w5165 | w5166);
assign w5167 = v2230;
assign w5168 = (~w4786 & ~w4788) | (~w4786 & w8630) | (~w4788 & w8630);
assign w5169 = w4789 & ~w4791;
assign v2231 = ~(w4793 | w5169);
assign w5170 = v2231;
assign w5171 = w4777 & ~w4779;
assign v2232 = ~(w4781 | w5171);
assign w5172 = v2232;
assign v2233 = ~(w5170 | w5172);
assign w5173 = v2233;
assign w5174 = w5170 & w5172;
assign v2234 = ~(w5173 | w5174);
assign w5175 = v2234;
assign w5176 = ~w5168 & w5175;
assign w5177 = w5168 & ~w5175;
assign v2235 = ~(w5176 | w5177);
assign w5178 = v2235;
assign w5179 = (~w4811 & ~w4813) | (~w4811 & w8631) | (~w4813 & w8631);
assign w5180 = w4814 & ~w4816;
assign v2236 = ~(w4818 | w5180);
assign w5181 = v2236;
assign w5182 = w4802 & ~w4804;
assign v2237 = ~(w4806 | w5182);
assign w5183 = v2237;
assign v2238 = ~(w5181 | w5183);
assign w5184 = v2238;
assign w5185 = w5181 & w5183;
assign v2239 = ~(w5184 | w5185);
assign w5186 = v2239;
assign w5187 = ~w5179 & w5186;
assign w5188 = w5179 & ~w5186;
assign v2240 = ~(w5187 | w5188);
assign w5189 = v2240;
assign w5190 = w5178 & w5189;
assign v2241 = ~(w5178 | w5189);
assign w5191 = v2241;
assign v2242 = ~(w5190 | w5191);
assign w5192 = v2242;
assign w5193 = w5167 & w5192;
assign v2243 = ~(w5167 | w5192);
assign w5194 = v2243;
assign v2244 = ~(w5193 | w5194);
assign w5195 = v2244;
assign v2245 = ~(w5156 | w5195);
assign w5196 = v2245;
assign w5197 = w5156 & w5195;
assign v2246 = ~(w5196 | w5197);
assign w5198 = v2246;
assign w5199 = ~w5131 & w5198;
assign w5200 = w5131 & ~w5198;
assign v2247 = ~(w5199 | w5200);
assign w5201 = v2247;
assign w5202 = (~w4983 & ~w4980) | (~w4983 & w9048) | (~w4980 & w9048);
assign w5203 = pi08 & pi59;
assign w5204 = pi09 & pi58;
assign v2248 = ~(w4889 | w5204);
assign w5205 = v2248;
assign w5206 = pi10 & pi58;
assign w5207 = w4887 & w5206;
assign v2249 = ~(w5205 | w5207);
assign w5208 = v2249;
assign w5209 = w5203 & ~w5208;
assign w5210 = ~w5203 & w5208;
assign v2250 = ~(w5209 | w5210);
assign w5211 = v2250;
assign w5212 = pi05 & pi62;
assign w5213 = pi06 & pi61;
assign v2251 = ~(w4901 | w5213);
assign w5214 = v2251;
assign w5215 = pi07 & pi61;
assign w5216 = w4899 & w5215;
assign v2252 = ~(w5214 | w5216);
assign w5217 = v2252;
assign w5218 = w5212 & ~w5217;
assign w5219 = ~w5212 & w5217;
assign v2253 = ~(w5218 | w5219);
assign w5220 = v2253;
assign v2254 = ~(w5211 | w5220);
assign w5221 = v2254;
assign w5222 = w5211 & w5220;
assign v2255 = ~(w5221 | w5222);
assign w5223 = v2255;
assign w5224 = (w4971 & w9049) | (w4971 & w9050) | (w9049 & w9050);
assign w5225 = w5223 & w9301;
assign v2256 = ~(w5224 | w5225);
assign w5226 = v2256;
assign w5227 = w5202 & w5226;
assign v2257 = ~(w5202 | w5226);
assign w5228 = v2257;
assign v2258 = ~(w5227 | w5228);
assign w5229 = v2258;
assign v2259 = ~(w5201 | w5229);
assign w5230 = v2259;
assign w5231 = w5201 & w5229;
assign v2260 = ~(w5230 | w5231);
assign w5232 = v2260;
assign w5233 = w5075 & w5232;
assign v2261 = ~(w5075 | w5232);
assign w5234 = v2261;
assign v2262 = ~(w5233 | w5234);
assign w5235 = v2262;
assign w5236 = ~w5022 & w5235;
assign w5237 = w5022 & ~w5235;
assign v2263 = ~(w5236 | w5237);
assign w5238 = v2263;
assign w5239 = (~w4925 & ~w4994) | (~w4925 & w9163) | (~w4994 & w9163);
assign v2264 = ~(w4919 | w4922);
assign w5240 = v2264;
assign w5241 = (~w4990 & ~w4991) | (~w4990 & w9051) | (~w4991 & w9051);
assign v2265 = ~(w5240 | w5241);
assign w5242 = v2265;
assign w5243 = w5240 & w5241;
assign v2266 = ~(w5242 | w5243);
assign w5244 = v2266;
assign w5245 = w5239 & ~w5244;
assign w5246 = ~w5239 & w5244;
assign v2267 = ~(w5245 | w5246);
assign w5247 = v2267;
assign w5248 = w5238 & ~w5247;
assign w5249 = ~w5238 & w5247;
assign v2268 = ~(w5248 | w5249);
assign w5250 = v2268;
assign v2269 = ~(w5021 | w5250);
assign w5251 = v2269;
assign w5252 = w5021 & w5250;
assign v2270 = ~(w5251 | w5252);
assign w5253 = v2270;
assign w5254 = w5020 & ~w5253;
assign w5255 = ~w5020 & w5253;
assign v2271 = ~(w5254 | w5255);
assign w5256 = v2271;
assign w5257 = ~w5014 & w5253;
assign v2272 = ~(w4770 | w5013);
assign w5258 = v2272;
assign w5259 = w4519 & ~w4769;
assign w5260 = w5259 & w8805;
assign w5261 = w4517 & ~w4769;
assign w5262 = w5258 & ~w5261;
assign w5263 = (~w5251 & w5262) | (~w5251 & w8806) | (w5262 & w8806);
assign w5264 = (w4010 & w8964) | (w4010 & w8965) | (w8964 & w8965);
assign w5265 = pi05 & pi63;
assign w5266 = pi06 & pi62;
assign w5267 = w5265 & ~w5266;
assign w5268 = ~w5265 & w5266;
assign v2273 = ~(w5267 | w5268);
assign w5269 = v2273;
assign w5270 = (~w5269 & w5165) | (~w5269 & w8966) | (w5165 & w8966);
assign w5271 = ~w5165 & w8967;
assign v2274 = ~(w5270 | w5271);
assign w5272 = v2274;
assign v2275 = ~(w5173 | w5176);
assign w5273 = v2275;
assign w5274 = (~w5036 & w5032) | (~w5036 & w8807) | (w5032 & w8807);
assign w5275 = (~w5184 & w5179) | (~w5184 & w8808) | (w5179 & w8808);
assign v2276 = ~(w5274 | w5275);
assign w5276 = v2276;
assign w5277 = w5274 & w5275;
assign v2277 = ~(w5276 | w5277);
assign w5278 = v2277;
assign w5279 = ~w5273 & w5278;
assign w5280 = w5273 & ~w5278;
assign v2278 = ~(w5279 | w5280);
assign w5281 = v2278;
assign w5282 = w5272 & w5281;
assign v2279 = ~(w5272 | w5281);
assign w5283 = v2279;
assign v2280 = ~(w5282 | w5283);
assign w5284 = v2280;
assign w5285 = (~w5046 & ~w5031) | (~w5046 & w8809) | (~w5031 & w8809);
assign w5286 = (~w5026 & ~w5028) | (~w5026 & w8810) | (~w5028 & w8810);
assign v2281 = ~(w5043 | w5286);
assign w5287 = v2281;
assign w5288 = w5043 & w5286;
assign v2282 = ~(w5287 | w5288);
assign w5289 = v2282;
assign w5290 = ~w5285 & w5289;
assign w5291 = w5285 & ~w5289;
assign v2283 = ~(w5290 | w5291);
assign w5292 = v2283;
assign w5293 = (~w5196 & ~w5198) | (~w5196 & w8751) | (~w5198 & w8751);
assign v2284 = ~(w5101 | w5129);
assign w5294 = v2284;
assign w5295 = (~w5190 & ~w5192) | (~w5190 & w8968) | (~w5192 & w8968);
assign v2285 = ~(w5294 | w5295);
assign w5296 = v2285;
assign w5297 = w5294 & w5295;
assign v2286 = ~(w5296 | w5297);
assign w5298 = v2286;
assign w5299 = w5298 & w5293;
assign w5300 = (w5198 & w9274) | (w5198 & w9275) | (w9274 & w9275);
assign v2287 = ~(w5299 | w5300);
assign w5301 = v2287;
assign w5302 = w5292 & w5301;
assign v2288 = ~(w5292 | w5301);
assign w5303 = v2288;
assign v2289 = ~(w5302 | w5303);
assign w5304 = v2289;
assign w5305 = w5284 & w5304;
assign v2290 = ~(w5284 | w5304);
assign w5306 = v2290;
assign v2291 = ~(w5305 | w5306);
assign w5307 = v2291;
assign w5308 = pi18 & pi50;
assign w5309 = pi22 & pi46;
assign w5310 = pi23 & pi45;
assign v2292 = ~(w5108 | w5310);
assign w5311 = v2292;
assign w5312 = pi24 & pi45;
assign w5313 = w5106 & w5312;
assign v2293 = ~(w5311 | w5313);
assign w5314 = v2293;
assign w5315 = w5309 & ~w5314;
assign w5316 = ~w5309 & w5314;
assign v2294 = ~(w5315 | w5316);
assign w5317 = v2294;
assign w5318 = w5308 & ~w5317;
assign w5319 = ~w5308 & w5317;
assign v2295 = ~(w5318 | w5319);
assign w5320 = v2295;
assign w5321 = pi19 & pi49;
assign w5322 = pi20 & pi48;
assign v2296 = ~(w5120 | w5322);
assign w5323 = v2296;
assign w5324 = pi21 & pi48;
assign w5325 = w5118 & w5324;
assign v2297 = ~(w5323 | w5325);
assign w5326 = v2297;
assign w5327 = w5321 & ~w5326;
assign w5328 = ~w5321 & w5326;
assign v2298 = ~(w5327 | w5328);
assign w5329 = v2298;
assign w5330 = w5320 & ~w5329;
assign w5331 = ~w5320 & w5329;
assign v2299 = ~(w5330 | w5331);
assign w5332 = v2299;
assign w5333 = w5212 & ~w5214;
assign v2300 = ~(w5216 | w5333);
assign w5334 = v2300;
assign w5335 = w5203 & ~w5205;
assign v2301 = ~(w5207 | w5335);
assign w5336 = v2301;
assign v2302 = ~(w5334 | w5336);
assign w5337 = v2302;
assign w5338 = w5334 & w5336;
assign v2303 = ~(w5337 | w5338);
assign w5339 = v2303;
assign w5340 = w5221 & w5339;
assign v2304 = ~(w5221 | w5339);
assign w5341 = v2304;
assign v2305 = ~(w5340 | w5341);
assign w5342 = v2305;
assign w5343 = pi25 & pi43;
assign w5344 = pi29 & pi39;
assign w5345 = pi31 & pi37;
assign w5346 = pi30 & pi38;
assign w5347 = ~w5345 & w5346;
assign w5348 = w5345 & ~w5346;
assign v2306 = ~(w5347 | w5348);
assign w5349 = v2306;
assign w5350 = w5344 & w5349;
assign v2307 = ~(w5344 | w5349);
assign w5351 = v2307;
assign v2308 = ~(w5350 | w5351);
assign w5352 = v2308;
assign w5353 = w5343 & w5352;
assign v2309 = ~(w5343 | w5352);
assign w5354 = v2309;
assign v2310 = ~(w5353 | w5354);
assign w5355 = v2310;
assign w5356 = pi26 & pi42;
assign w5357 = pi27 & pi41;
assign v2311 = ~(w5092 | w5357);
assign w5358 = v2311;
assign w5359 = pi28 & pi41;
assign w5360 = w5090 & w5359;
assign v2312 = ~(w5358 | w5360);
assign w5361 = v2312;
assign w5362 = w5356 & ~w5361;
assign w5363 = ~w5356 & w5361;
assign v2313 = ~(w5362 | w5363);
assign w5364 = v2313;
assign w5365 = w5355 & ~w5364;
assign w5366 = ~w5355 & w5364;
assign v2314 = ~(w5365 | w5366);
assign w5367 = v2314;
assign w5368 = w5342 & w5367;
assign v2315 = ~(w5342 | w5367);
assign w5369 = v2315;
assign v2316 = ~(w5368 | w5369);
assign w5370 = v2316;
assign w5371 = w5332 & w5370;
assign v2317 = ~(w5332 | w5370);
assign w5372 = v2317;
assign v2318 = ~(w5371 | w5372);
assign w5373 = v2318;
assign w5374 = (~w5142 & ~w5144) | (~w5142 & w8811) | (~w5144 & w8811);
assign w5375 = w5145 & ~w5147;
assign v2319 = ~(w5149 | w5375);
assign w5376 = v2319;
assign w5377 = w5133 & ~w5135;
assign v2320 = ~(w5137 | w5377);
assign w5378 = v2320;
assign v2321 = ~(w5376 | w5378);
assign w5379 = v2321;
assign w5380 = w5376 & w5378;
assign v2322 = ~(w5379 | w5380);
assign w5381 = v2322;
assign w5382 = ~w5374 & w5381;
assign w5383 = w5374 & ~w5381;
assign v2323 = ~(w5382 | w5383);
assign w5384 = v2323;
assign w5385 = (~w5114 & ~w5116) | (~w5114 & w8632) | (~w5116 & w8632);
assign w5386 = w5117 & ~w5119;
assign v2324 = ~(w5121 | w5386);
assign w5387 = v2324;
assign w5388 = w5105 & ~w5107;
assign v2325 = ~(w5109 | w5388);
assign w5389 = v2325;
assign v2326 = ~(w5387 | w5389);
assign w5390 = v2326;
assign w5391 = w5387 & w5389;
assign v2327 = ~(w5390 | w5391);
assign w5392 = v2327;
assign w5393 = ~w5385 & w5392;
assign w5394 = w5385 & ~w5392;
assign v2328 = ~(w5393 | w5394);
assign w5395 = v2328;
assign w5396 = (~w5086 & ~w5088) | (~w5086 & w8633) | (~w5088 & w8633);
assign w5397 = (~w5080 & ~w5082) | (~w5080 & w8969) | (~w5082 & w8969);
assign w5398 = w5089 & ~w5091;
assign v2329 = ~(w5093 | w5398);
assign w5399 = v2329;
assign v2330 = ~(w5397 | w5399);
assign w5400 = v2330;
assign w5401 = w5397 & w5399;
assign v2331 = ~(w5400 | w5401);
assign w5402 = v2331;
assign w5403 = ~w5396 & w5402;
assign w5404 = w5396 & ~w5402;
assign v2332 = ~(w5403 | w5404);
assign w5405 = v2332;
assign w5406 = w5395 & w5405;
assign v2333 = ~(w5395 | w5405);
assign w5407 = v2333;
assign v2334 = ~(w5406 | w5407);
assign w5408 = v2334;
assign w5409 = w5384 & w5408;
assign v2335 = ~(w5384 | w5408);
assign w5410 = v2335;
assign v2336 = ~(w5409 | w5410);
assign w5411 = v2336;
assign w5412 = pi11 & pi57;
assign w5413 = pi15 & pi53;
assign w5414 = pi16 & pi52;
assign v2337 = ~(w5136 | w5414);
assign w5415 = v2337;
assign w5416 = pi17 & pi52;
assign w5417 = w5134 & w5416;
assign v2338 = ~(w5415 | w5417);
assign w5418 = v2338;
assign w5419 = w5413 & ~w5418;
assign w5420 = ~w5413 & w5418;
assign v2339 = ~(w5419 | w5420);
assign w5421 = v2339;
assign w5422 = w5412 & ~w5421;
assign w5423 = ~w5412 & w5421;
assign v2340 = ~(w5422 | w5423);
assign w5424 = v2340;
assign w5425 = pi12 & pi56;
assign w5426 = pi13 & pi55;
assign v2341 = ~(w5148 | w5426);
assign w5427 = v2341;
assign w5428 = pi14 & pi55;
assign w5429 = w5146 & w5428;
assign v2342 = ~(w5427 | w5429);
assign w5430 = v2342;
assign w5431 = w5425 & ~w5430;
assign w5432 = ~w5425 & w5430;
assign v2343 = ~(w5431 | w5432);
assign w5433 = v2343;
assign w5434 = w5424 & ~w5433;
assign w5435 = ~w5424 & w5433;
assign v2344 = ~(w5434 | w5435);
assign w5436 = v2344;
assign w5437 = w5411 & w5436;
assign v2345 = ~(w5411 | w5436);
assign w5438 = v2345;
assign v2346 = ~(w5437 | w5438);
assign w5439 = v2346;
assign w5440 = w5373 & w5439;
assign v2347 = ~(w5373 | w5439);
assign w5441 = v2347;
assign v2348 = ~(w5440 | w5441);
assign w5442 = v2348;
assign w5443 = (~w5055 & w5052) | (~w5055 & w9052) | (w5052 & w9052);
assign w5444 = pi08 & pi60;
assign w5445 = pi09 & pi59;
assign v2349 = ~(w5206 | w5445);
assign w5446 = v2349;
assign w5447 = pi10 & pi59;
assign w5448 = w5204 & w5447;
assign v2350 = ~(w5446 | w5448);
assign w5449 = v2350;
assign w5450 = w5444 & w5449;
assign v2351 = ~(w5444 | w5449);
assign w5451 = v2351;
assign v2352 = ~(w5450 | w5451);
assign w5452 = v2352;
assign w5453 = w5215 & w5452;
assign v2353 = ~(w5215 | w5452);
assign w5454 = v2353;
assign v2354 = ~(w5453 | w5454);
assign w5455 = v2354;
assign w5456 = (w8970 & w5061) | (w8970 & w9053) | (w5061 & w9053);
assign w5457 = (w5455 & w8971) | (w5455 & w5067) | (w8971 & w5067);
assign v2355 = ~(w5456 | w5457);
assign w5458 = v2355;
assign w5459 = w5443 & w5458;
assign v2356 = ~(w5443 | w5458);
assign w5460 = v2356;
assign v2357 = ~(w5459 | w5460);
assign w5461 = v2357;
assign w5462 = w5442 & ~w5461;
assign w5463 = ~w5442 & w5461;
assign v2358 = ~(w5462 | w5463);
assign w5464 = v2358;
assign w5465 = w5307 & w5464;
assign v2359 = ~(w5307 | w5464);
assign w5466 = v2359;
assign v2360 = ~(w5465 | w5466);
assign w5467 = v2360;
assign w5468 = (w5467 & w5246) | (w5467 & w8972) | (w5246 & w8972);
assign w5469 = ~w5246 & w8973;
assign v2361 = ~(w5468 | w5469);
assign w5470 = v2361;
assign v2362 = ~(w5230 | w5233);
assign w5471 = v2362;
assign v2363 = ~(w5224 | w5227);
assign w5472 = v2363;
assign w5473 = (~w5070 & ~w5072) | (~w5070 & w8974) | (~w5072 & w8974);
assign w5474 = w5472 & ~w5473;
assign w5475 = ~w5472 & w5473;
assign v2364 = ~(w5474 | w5475);
assign w5476 = v2364;
assign w5477 = w5471 & w5476;
assign v2365 = ~(w5471 | w5476);
assign w5478 = v2365;
assign v2366 = ~(w5477 | w5478);
assign w5479 = v2366;
assign w5480 = w5470 & w5479;
assign v2367 = ~(w5470 | w5479);
assign w5481 = v2367;
assign v2368 = ~(w5480 | w5481);
assign w5482 = v2368;
assign v2369 = ~(w5237 | w5248);
assign w5483 = v2369;
assign w5484 = ~w5482 & w5483;
assign w5485 = w5482 & ~w5483;
assign v2370 = ~(w5484 | w5485);
assign w5486 = v2370;
assign w5487 = ~w5264 & w5486;
assign w5488 = w5264 & ~w5486;
assign v2371 = ~(w5487 | w5488);
assign w5489 = v2371;
assign w5490 = (~w5484 & w5264) | (~w5484 & w9276) | (w5264 & w9276);
assign v2372 = ~(w5462 | w5465);
assign w5491 = v2372;
assign v2373 = ~(w5456 | w5459);
assign w5492 = v2373;
assign w5493 = (~w5302 & ~w5304) | (~w5302 & w8812) | (~w5304 & w8812);
assign w5494 = w5492 & ~w5493;
assign w5495 = ~w5492 & w5493;
assign v2374 = ~(w5494 | w5495);
assign w5496 = v2374;
assign w5497 = ~w5491 & w5496;
assign w5498 = w5491 & ~w5496;
assign v2375 = ~(w5497 | w5498);
assign w5499 = v2375;
assign v2376 = ~(w5230 | w5474);
assign w5500 = v2376;
assign w5501 = ~w5233 & w5500;
assign w5502 = pi18 & pi51;
assign w5503 = pi22 & pi47;
assign w5504 = pi23 & pi46;
assign v2377 = ~(w5312 | w5504);
assign w5505 = v2377;
assign w5506 = pi24 & pi46;
assign w5507 = w5310 & w5506;
assign v2378 = ~(w5505 | w5507);
assign w5508 = v2378;
assign w5509 = w5503 & ~w5508;
assign w5510 = ~w5503 & w5508;
assign v2379 = ~(w5509 | w5510);
assign w5511 = v2379;
assign w5512 = w5502 & ~w5511;
assign w5513 = ~w5502 & w5511;
assign v2380 = ~(w5512 | w5513);
assign w5514 = v2380;
assign w5515 = pi19 & pi50;
assign w5516 = pi20 & pi49;
assign v2381 = ~(w5324 | w5516);
assign w5517 = v2381;
assign w5518 = pi21 & pi49;
assign w5519 = w5322 & w5518;
assign v2382 = ~(w5517 | w5519);
assign w5520 = v2382;
assign w5521 = w5515 & ~w5520;
assign w5522 = ~w5515 & w5520;
assign v2383 = ~(w5521 | w5522);
assign w5523 = v2383;
assign w5524 = w5514 & ~w5523;
assign w5525 = ~w5514 & w5523;
assign v2384 = ~(w5524 | w5525);
assign w5526 = v2384;
assign w5527 = pi25 & pi44;
assign w5528 = pi29 & pi40;
assign w5529 = pi31 & pi38;
assign w5530 = pi30 & pi39;
assign w5531 = ~w5529 & w5530;
assign w5532 = w5529 & ~w5530;
assign v2385 = ~(w5531 | w5532);
assign w5533 = v2385;
assign w5534 = w5528 & w5533;
assign v2386 = ~(w5528 | w5533);
assign w5535 = v2386;
assign v2387 = ~(w5534 | w5535);
assign w5536 = v2387;
assign w5537 = w5527 & w5536;
assign v2388 = ~(w5527 | w5536);
assign w5538 = v2388;
assign v2389 = ~(w5537 | w5538);
assign w5539 = v2389;
assign w5540 = pi26 & pi43;
assign w5541 = pi27 & pi42;
assign v2390 = ~(w5359 | w5541);
assign w5542 = v2390;
assign w5543 = pi28 & pi42;
assign w5544 = w5357 & w5543;
assign v2391 = ~(w5542 | w5544);
assign w5545 = v2391;
assign w5546 = w5540 & ~w5545;
assign w5547 = ~w5540 & w5545;
assign v2392 = ~(w5546 | w5547);
assign w5548 = v2392;
assign w5549 = w5539 & ~w5548;
assign w5550 = ~w5539 & w5548;
assign v2393 = ~(w5549 | w5550);
assign w5551 = v2393;
assign w5552 = w5448 & w5453;
assign v2394 = ~(w5448 | w5453);
assign w5553 = v2394;
assign v2395 = ~(w5552 | w5553);
assign w5554 = v2395;
assign v2396 = ~(w5450 | w5554);
assign w5555 = v2396;
assign w5556 = w5551 & ~w5555;
assign w5557 = ~w5551 & w5555;
assign v2397 = ~(w5556 | w5557);
assign w5558 = v2397;
assign w5559 = w5526 & w5558;
assign v2398 = ~(w5526 | w5558);
assign w5560 = v2398;
assign v2399 = ~(w5559 | w5560);
assign w5561 = v2399;
assign w5562 = (~w5422 & ~w5424) | (~w5422 & w8813) | (~w5424 & w8813);
assign w5563 = w5425 & ~w5427;
assign v2400 = ~(w5429 | w5563);
assign w5564 = v2400;
assign w5565 = w5413 & ~w5415;
assign v2401 = ~(w5417 | w5565);
assign w5566 = v2401;
assign v2402 = ~(w5564 | w5566);
assign w5567 = v2402;
assign w5568 = w5564 & w5566;
assign v2403 = ~(w5567 | w5568);
assign w5569 = v2403;
assign w5570 = ~w5562 & w5569;
assign w5571 = w5562 & ~w5569;
assign v2404 = ~(w5570 | w5571);
assign w5572 = v2404;
assign w5573 = (~w5318 & ~w5320) | (~w5318 & w8634) | (~w5320 & w8634);
assign w5574 = w5321 & ~w5323;
assign v2405 = ~(w5325 | w5574);
assign w5575 = v2405;
assign w5576 = w5309 & ~w5311;
assign v2406 = ~(w5313 | w5576);
assign w5577 = v2406;
assign v2407 = ~(w5575 | w5577);
assign w5578 = v2407;
assign w5579 = w5575 & w5577;
assign v2408 = ~(w5578 | w5579);
assign w5580 = v2408;
assign w5581 = ~w5573 & w5580;
assign w5582 = w5573 & ~w5580;
assign v2409 = ~(w5581 | w5582);
assign w5583 = v2409;
assign w5584 = (~w5353 & ~w5355) | (~w5353 & w8635) | (~w5355 & w8635);
assign w5585 = (~w5347 & ~w5349) | (~w5347 & w8814) | (~w5349 & w8814);
assign w5586 = w5356 & ~w5358;
assign v2410 = ~(w5360 | w5586);
assign w5587 = v2410;
assign v2411 = ~(w5585 | w5587);
assign w5588 = v2411;
assign w5589 = w5585 & w5587;
assign v2412 = ~(w5588 | w5589);
assign w5590 = v2412;
assign w5591 = ~w5584 & w5590;
assign w5592 = w5584 & ~w5590;
assign v2413 = ~(w5591 | w5592);
assign w5593 = v2413;
assign w5594 = w5583 & w5593;
assign v2414 = ~(w5583 | w5593);
assign w5595 = v2414;
assign v2415 = ~(w5594 | w5595);
assign w5596 = v2415;
assign w5597 = w5572 & w5596;
assign v2416 = ~(w5572 | w5596);
assign w5598 = v2416;
assign v2417 = ~(w5597 | w5598);
assign w5599 = v2417;
assign w5600 = pi11 & pi58;
assign w5601 = pi15 & pi54;
assign w5602 = pi16 & pi53;
assign v2418 = ~(w5416 | w5602);
assign w5603 = v2418;
assign w5604 = pi17 & pi53;
assign w5605 = w5414 & w5604;
assign v2419 = ~(w5603 | w5605);
assign w5606 = v2419;
assign w5607 = w5601 & ~w5606;
assign w5608 = ~w5601 & w5606;
assign v2420 = ~(w5607 | w5608);
assign w5609 = v2420;
assign w5610 = w5600 & ~w5609;
assign w5611 = ~w5600 & w5609;
assign v2421 = ~(w5610 | w5611);
assign w5612 = v2421;
assign w5613 = pi12 & pi57;
assign w5614 = pi13 & pi56;
assign v2422 = ~(w5428 | w5614);
assign w5615 = v2422;
assign w5616 = pi14 & pi56;
assign w5617 = w5426 & w5616;
assign v2423 = ~(w5615 | w5617);
assign w5618 = v2423;
assign w5619 = w5613 & ~w5618;
assign w5620 = ~w5613 & w5618;
assign v2424 = ~(w5619 | w5620);
assign w5621 = v2424;
assign w5622 = w5612 & ~w5621;
assign w5623 = ~w5612 & w5621;
assign v2425 = ~(w5622 | w5623);
assign w5624 = v2425;
assign w5625 = w5599 & w5624;
assign v2426 = ~(w5599 | w5624);
assign w5626 = v2426;
assign v2427 = ~(w5625 | w5626);
assign w5627 = v2427;
assign w5628 = w5561 & w5627;
assign v2428 = ~(w5561 | w5627);
assign w5629 = v2428;
assign v2429 = ~(w5628 | w5629);
assign w5630 = v2429;
assign w5631 = (~w5296 & ~w5293) | (~w5296 & w8815) | (~w5293 & w8815);
assign w5632 = pi08 & pi61;
assign w5633 = pi09 & pi60;
assign v2430 = ~(w5447 | w5633);
assign w5634 = v2430;
assign w5635 = pi10 & pi60;
assign w5636 = w5445 & w5635;
assign v2431 = ~(w5634 | w5636);
assign w5637 = v2431;
assign w5638 = w5632 & ~w5637;
assign w5639 = ~w5632 & w5637;
assign v2432 = ~(w5638 | w5639);
assign w5640 = v2432;
assign w5641 = (~w5640 & w5290) | (~w5640 & w8975) | (w5290 & w8975);
assign w5642 = ~w5290 & w8976;
assign v2433 = ~(w5641 | w5642);
assign w5643 = v2433;
assign w5644 = ~w5631 & w5643;
assign w5645 = w5631 & ~w5643;
assign v2434 = ~(w5644 | w5645);
assign w5646 = v2434;
assign w5647 = w5630 & w5646;
assign v2435 = ~(w5630 | w5646);
assign w5648 = v2435;
assign v2436 = ~(w5647 | w5648);
assign w5649 = v2436;
assign v2437 = ~(w5337 | w5340);
assign w5650 = v2437;
assign w5651 = pi06 & pi63;
assign w5652 = pi07 & pi62;
assign w5653 = w5651 & ~w5652;
assign w5654 = ~w5651 & w5652;
assign v2438 = ~(w5653 | w5654);
assign w5655 = v2438;
assign v2439 = ~(w5650 | w5655);
assign w5656 = v2439;
assign w5657 = w5650 & w5655;
assign v2440 = ~(w5656 | w5657);
assign w5658 = v2440;
assign w5659 = (~w5379 & w5374) | (~w5379 & w8977) | (w5374 & w8977);
assign w5660 = (~w5400 & w5396) | (~w5400 & w8816) | (w5396 & w8816);
assign w5661 = (~w5390 & w5385) | (~w5390 & w8817) | (w5385 & w8817);
assign v2441 = ~(w5660 | w5661);
assign w5662 = v2441;
assign w5663 = w5660 & w5661;
assign v2442 = ~(w5662 | w5663);
assign w5664 = v2442;
assign w5665 = ~w5659 & w5664;
assign w5666 = w5659 & ~w5664;
assign v2443 = ~(w5665 | w5666);
assign w5667 = v2443;
assign w5668 = w5658 & w5667;
assign v2444 = ~(w5658 | w5667);
assign w5669 = v2444;
assign v2445 = ~(w5668 | w5669);
assign w5670 = v2445;
assign w5671 = (~w5270 & ~w5281) | (~w5270 & w8978) | (~w5281 & w8978);
assign w5672 = (~w5276 & ~w5278) | (~w5276 & w8979) | (~w5278 & w8979);
assign v2446 = ~(w5267 | w5672);
assign w5673 = v2446;
assign w5674 = w5267 & w5672;
assign v2447 = ~(w5673 | w5674);
assign w5675 = v2447;
assign w5676 = ~w5671 & w5675;
assign w5677 = w5671 & ~w5675;
assign v2448 = ~(w5676 | w5677);
assign w5678 = v2448;
assign w5679 = (~w5437 & ~w5439) | (~w5437 & w8752) | (~w5439 & w8752);
assign v2449 = ~(w5368 | w5371);
assign w5680 = v2449;
assign w5681 = (~w5406 & ~w5408) | (~w5406 & w8980) | (~w5408 & w8980);
assign v2450 = ~(w5680 | w5681);
assign w5682 = v2450;
assign w5683 = w5680 & w5681;
assign v2451 = ~(w5682 | w5683);
assign w5684 = v2451;
assign w5685 = (w5439 & w9164) | (w5439 & w9165) | (w9164 & w9165);
assign w5686 = ~w5684 & w5679;
assign v2452 = ~(w5685 | w5686);
assign w5687 = v2452;
assign w5688 = w5678 & w5687;
assign v2453 = ~(w5678 | w5687);
assign w5689 = v2453;
assign v2454 = ~(w5688 | w5689);
assign w5690 = v2454;
assign w5691 = w5670 & ~w5690;
assign w5692 = ~w5670 & w5690;
assign v2455 = ~(w5691 | w5692);
assign w5693 = v2455;
assign w5694 = w5649 & ~w5693;
assign w5695 = ~w5649 & w5693;
assign v2456 = ~(w5694 | w5695);
assign w5696 = v2456;
assign w5697 = ~w5501 & w8753;
assign w5698 = (~w5696 & w5501) | (~w5696 & w8754) | (w5501 & w8754);
assign v2457 = ~(w5697 | w5698);
assign w5699 = v2457;
assign w5700 = w5499 & ~w5699;
assign w5701 = ~w5499 & w5699;
assign v2458 = ~(w5700 | w5701);
assign w5702 = v2458;
assign w5703 = (~w5469 & ~w5470) | (~w5469 & w8755) | (~w5470 & w8755);
assign w5704 = w5702 & ~w5703;
assign w5705 = ~w5702 & w5703;
assign v2459 = ~(w5704 | w5705);
assign w5706 = v2459;
assign w5707 = w5490 & ~w5706;
assign w5708 = (w5706 & w8756) | (w5706 & w5487) | (w8756 & w5487);
assign v2460 = ~(w5707 | w5708);
assign w5709 = v2460;
assign w5710 = (~w5462 & w5493) | (~w5462 & w9054) | (w5493 & w9054);
assign w5711 = (~w5495 & w5465) | (~w5495 & w8757) | (w5465 & w8757);
assign w5712 = (~w5647 & w5693) | (~w5647 & w8818) | (w5693 & w8818);
assign v2461 = ~(w5641 | w5644);
assign w5713 = v2461;
assign w5714 = (~w5689 & ~w5690) | (~w5689 & w8758) | (~w5690 & w8758);
assign w5715 = ~w5713 & w5714;
assign w5716 = w5713 & ~w5714;
assign v2462 = ~(w5715 | w5716);
assign w5717 = v2462;
assign w5718 = ~w5712 & w5717;
assign w5719 = w5712 & ~w5717;
assign v2463 = ~(w5718 | w5719);
assign w5720 = v2463;
assign w5721 = w5720 & w9277;
assign v2464 = ~(w5567 | w5570);
assign w5722 = v2464;
assign w5723 = (~w5588 & w5584) | (~w5588 & w8759) | (w5584 & w8759);
assign w5724 = (~w5578 & w5573) | (~w5578 & w8760) | (w5573 & w8760);
assign v2465 = ~(w5723 | w5724);
assign w5725 = v2465;
assign w5726 = w5723 & w5724;
assign v2466 = ~(w5725 | w5726);
assign w5727 = v2466;
assign w5728 = ~w5722 & w5727;
assign w5729 = w5722 & ~w5727;
assign v2467 = ~(w5728 | w5729);
assign w5730 = v2467;
assign w5731 = pi07 & pi63;
assign w5732 = pi08 & pi62;
assign w5733 = w5731 & ~w5732;
assign w5734 = ~w5731 & w5732;
assign v2468 = ~(w5733 | w5734);
assign w5735 = v2468;
assign w5736 = w5552 & ~w5735;
assign w5737 = ~w5552 & w5735;
assign v2469 = ~(w5736 | w5737);
assign w5738 = v2469;
assign w5739 = w5730 & w5738;
assign v2470 = ~(w5730 | w5738);
assign w5740 = v2470;
assign v2471 = ~(w5739 | w5740);
assign w5741 = v2471;
assign w5742 = (~w5656 & ~w5667) | (~w5656 & w8761) | (~w5667 & w8761);
assign w5743 = (~w5662 & ~w5664) | (~w5662 & w8762) | (~w5664 & w8762);
assign v2472 = ~(w5653 | w5743);
assign w5744 = v2472;
assign w5745 = w5653 & w5743;
assign v2473 = ~(w5744 | w5745);
assign w5746 = v2473;
assign w5747 = ~w5742 & w5746;
assign w5748 = w5742 & ~w5746;
assign v2474 = ~(w5747 | w5748);
assign w5749 = v2474;
assign w5750 = (~w5625 & ~w5627) | (~w5625 & w8763) | (~w5627 & w8763);
assign v2475 = ~(w5556 | w5559);
assign w5751 = v2475;
assign w5752 = (~w5594 & ~w5596) | (~w5594 & w8983) | (~w5596 & w8983);
assign v2476 = ~(w5751 | w5752);
assign w5753 = v2476;
assign w5754 = w5751 & w5752;
assign v2477 = ~(w5753 | w5754);
assign w5755 = v2477;
assign w5756 = (w5627 & w9166) | (w5627 & w9167) | (w9166 & w9167);
assign w5757 = ~w5755 & w5750;
assign v2478 = ~(w5756 | w5757);
assign w5758 = v2478;
assign w5759 = w5749 & w5758;
assign v2479 = ~(w5749 | w5758);
assign w5760 = v2479;
assign v2480 = ~(w5759 | w5760);
assign w5761 = v2480;
assign w5762 = w5741 & w5761;
assign v2481 = ~(w5741 | w5761);
assign w5763 = v2481;
assign v2482 = ~(w5762 | w5763);
assign w5764 = v2482;
assign w5765 = pi25 & pi45;
assign w5766 = pi29 & pi41;
assign w5767 = pi31 & pi39;
assign w5768 = pi30 & pi40;
assign w5769 = ~w5767 & w5768;
assign w5770 = w5767 & ~w5768;
assign v2483 = ~(w5769 | w5770);
assign w5771 = v2483;
assign w5772 = w5766 & w5771;
assign v2484 = ~(w5766 | w5771);
assign w5773 = v2484;
assign v2485 = ~(w5772 | w5773);
assign w5774 = v2485;
assign w5775 = w5765 & w5774;
assign v2486 = ~(w5765 | w5774);
assign w5776 = v2486;
assign v2487 = ~(w5775 | w5776);
assign w5777 = v2487;
assign w5778 = pi26 & pi44;
assign w5779 = pi27 & pi43;
assign v2488 = ~(w5543 | w5779);
assign w5780 = v2488;
assign w5781 = pi28 & pi43;
assign w5782 = w5541 & w5781;
assign v2489 = ~(w5780 | w5782);
assign w5783 = v2489;
assign w5784 = w5778 & ~w5783;
assign w5785 = ~w5778 & w5783;
assign v2490 = ~(w5784 | w5785);
assign w5786 = v2490;
assign w5787 = w5777 & ~w5786;
assign w5788 = ~w5777 & w5786;
assign v2491 = ~(w5787 | w5788);
assign w5789 = v2491;
assign w5790 = w5632 & ~w5634;
assign v2492 = ~(w5636 | w5790);
assign w5791 = v2492;
assign w5792 = w5789 & ~w5791;
assign w5793 = ~w5789 & w5791;
assign v2493 = ~(w5792 | w5793);
assign w5794 = v2493;
assign w5795 = pi18 & pi52;
assign w5796 = pi22 & pi48;
assign w5797 = pi23 & pi47;
assign v2494 = ~(w5506 | w5797);
assign w5798 = v2494;
assign w5799 = pi24 & pi47;
assign w5800 = w5504 & w5799;
assign v2495 = ~(w5798 | w5800);
assign w5801 = v2495;
assign w5802 = w5796 & ~w5801;
assign w5803 = ~w5796 & w5801;
assign v2496 = ~(w5802 | w5803);
assign w5804 = v2496;
assign w5805 = w5795 & ~w5804;
assign w5806 = ~w5795 & w5804;
assign v2497 = ~(w5805 | w5806);
assign w5807 = v2497;
assign w5808 = pi19 & pi51;
assign w5809 = pi20 & pi50;
assign v2498 = ~(w5518 | w5809);
assign w5810 = v2498;
assign w5811 = pi21 & pi50;
assign w5812 = w5516 & w5811;
assign v2499 = ~(w5810 | w5812);
assign w5813 = v2499;
assign w5814 = w5808 & ~w5813;
assign w5815 = ~w5808 & w5813;
assign v2500 = ~(w5814 | w5815);
assign w5816 = v2500;
assign w5817 = w5807 & ~w5816;
assign w5818 = ~w5807 & w5816;
assign v2501 = ~(w5817 | w5818);
assign w5819 = v2501;
assign w5820 = w5794 & w5819;
assign v2502 = ~(w5794 | w5819);
assign w5821 = v2502;
assign v2503 = ~(w5820 | w5821);
assign w5822 = v2503;
assign w5823 = pi11 & pi59;
assign w5824 = pi15 & pi55;
assign w5825 = pi16 & pi54;
assign v2504 = ~(w5604 | w5825);
assign w5826 = v2504;
assign w5827 = pi17 & pi54;
assign w5828 = w5602 & w5827;
assign v2505 = ~(w5826 | w5828);
assign w5829 = v2505;
assign w5830 = w5824 & ~w5829;
assign w5831 = ~w5824 & w5829;
assign v2506 = ~(w5830 | w5831);
assign w5832 = v2506;
assign w5833 = w5823 & ~w5832;
assign w5834 = ~w5823 & w5832;
assign v2507 = ~(w5833 | w5834);
assign w5835 = v2507;
assign w5836 = pi12 & pi58;
assign w5837 = pi13 & pi57;
assign v2508 = ~(w5616 | w5837);
assign w5838 = v2508;
assign w5839 = pi14 & pi57;
assign w5840 = w5614 & w5839;
assign v2509 = ~(w5838 | w5840);
assign w5841 = v2509;
assign w5842 = w5836 & ~w5841;
assign w5843 = ~w5836 & w5841;
assign v2510 = ~(w5842 | w5843);
assign w5844 = v2510;
assign w5845 = w5835 & ~w5844;
assign w5846 = ~w5835 & w5844;
assign v2511 = ~(w5845 | w5846);
assign w5847 = v2511;
assign w5848 = (~w5610 & ~w5612) | (~w5610 & w8636) | (~w5612 & w8636);
assign w5849 = w5613 & ~w5615;
assign v2512 = ~(w5617 | w5849);
assign w5850 = v2512;
assign w5851 = w5601 & ~w5603;
assign v2513 = ~(w5605 | w5851);
assign w5852 = v2513;
assign v2514 = ~(w5850 | w5852);
assign w5853 = v2514;
assign w5854 = w5850 & w5852;
assign v2515 = ~(w5853 | w5854);
assign w5855 = v2515;
assign w5856 = ~w5848 & w5855;
assign w5857 = w5848 & ~w5855;
assign v2516 = ~(w5856 | w5857);
assign w5858 = v2516;
assign w5859 = (~w5512 & ~w5514) | (~w5512 & w8637) | (~w5514 & w8637);
assign w5860 = w5515 & ~w5517;
assign v2517 = ~(w5519 | w5860);
assign w5861 = v2517;
assign w5862 = w5503 & ~w5505;
assign v2518 = ~(w5507 | w5862);
assign w5863 = v2518;
assign v2519 = ~(w5861 | w5863);
assign w5864 = v2519;
assign w5865 = w5861 & w5863;
assign v2520 = ~(w5864 | w5865);
assign w5866 = v2520;
assign w5867 = ~w5859 & w5866;
assign w5868 = w5859 & ~w5866;
assign v2521 = ~(w5867 | w5868);
assign w5869 = v2521;
assign w5870 = (~w5537 & ~w5539) | (~w5537 & w8638) | (~w5539 & w8638);
assign v2522 = ~(w5531 | w5534);
assign w5871 = v2522;
assign w5872 = w5540 & ~w5542;
assign v2523 = ~(w5544 | w5872);
assign w5873 = v2523;
assign v2524 = ~(w5871 | w5873);
assign w5874 = v2524;
assign w5875 = w5871 & w5873;
assign v2525 = ~(w5874 | w5875);
assign w5876 = v2525;
assign w5877 = ~w5870 & w5876;
assign w5878 = w5870 & ~w5876;
assign v2526 = ~(w5877 | w5878);
assign w5879 = v2526;
assign w5880 = w5869 & w5879;
assign v2527 = ~(w5869 | w5879);
assign w5881 = v2527;
assign v2528 = ~(w5880 | w5881);
assign w5882 = v2528;
assign w5883 = w5858 & w5882;
assign v2529 = ~(w5858 | w5882);
assign w5884 = v2529;
assign v2530 = ~(w5883 | w5884);
assign w5885 = v2530;
assign v2531 = ~(w5847 | w5885);
assign w5886 = v2531;
assign w5887 = w5847 & w5885;
assign v2532 = ~(w5886 | w5887);
assign w5888 = v2532;
assign w5889 = ~w5822 & w5888;
assign w5890 = w5822 & ~w5888;
assign v2533 = ~(w5889 | w5890);
assign w5891 = v2533;
assign w5892 = (~w5682 & w5679) | (~w5682 & w8819) | (w5679 & w8819);
assign w5893 = pi09 & pi61;
assign v2534 = ~(w5635 | w5893);
assign w5894 = v2534;
assign w5895 = pi10 & pi61;
assign w5896 = w5633 & w5895;
assign v2535 = ~(w5894 | w5896);
assign w5897 = v2535;
assign w5898 = ~w5676 & w8764;
assign w5899 = (w5897 & w5676) | (w5897 & w8765) | (w5676 & w8765);
assign v2536 = ~(w5898 | w5899);
assign w5900 = v2536;
assign w5901 = w5892 & w5900;
assign v2537 = ~(w5892 | w5900);
assign w5902 = v2537;
assign v2538 = ~(w5901 | w5902);
assign w5903 = v2538;
assign v2539 = ~(w5891 | w5903);
assign w5904 = v2539;
assign w5905 = w5891 & w5903;
assign v2540 = ~(w5904 | w5905);
assign w5906 = v2540;
assign w5907 = w5764 & w5906;
assign v2541 = ~(w5764 | w5906);
assign w5908 = v2541;
assign v2542 = ~(w5907 | w5908);
assign w5909 = v2542;
assign w5910 = (w5909 & w5721) | (w5909 & w8766) | (w5721 & w8766);
assign w5911 = ~w5721 & w8767;
assign v2543 = ~(w5910 | w5911);
assign w5912 = v2543;
assign w5913 = (~w5698 & ~w5699) | (~w5698 & w8984) | (~w5699 & w8984);
assign w5914 = w5912 & w5913;
assign v2544 = ~(w5912 | w5913);
assign w5915 = v2544;
assign v2545 = ~(w5914 | w5915);
assign w5916 = v2545;
assign w5917 = (w5264 & w9055) | (w5264 & w9056) | (w9055 & w9056);
assign w5918 = w5916 & ~w5917;
assign w5919 = ~w5916 & w5917;
assign v2546 = ~(w5918 | w5919);
assign w5920 = v2546;
assign w5921 = (w5264 & w9278) | (w5264 & w9279) | (w9278 & w9279);
assign w5922 = w5711 & w5720;
assign v2547 = ~(w5922 | w5910);
assign w5923 = v2547;
assign w5924 = (~w5864 & w5859) | (~w5864 & w8820) | (w5859 & w8820);
assign w5925 = pi09 & pi62;
assign w5926 = pi11 & pi60;
assign v2548 = ~(w5895 | w5926);
assign w5927 = v2548;
assign w5928 = pi11 & pi61;
assign w5929 = w5635 & w5928;
assign v2549 = ~(w5927 | w5929);
assign w5930 = v2549;
assign w5931 = w5925 & ~w5930;
assign w5932 = ~w5925 & w5930;
assign v2550 = ~(w5931 | w5932);
assign w5933 = v2550;
assign v2551 = ~(w5924 | w5933);
assign w5934 = v2551;
assign w5935 = w5924 & w5933;
assign v2552 = ~(w5934 | w5935);
assign w5936 = v2552;
assign w5937 = pi08 & pi63;
assign w5938 = (~w5874 & w5870) | (~w5874 & w8821) | (w5870 & w8821);
assign w5939 = w5937 & w5938;
assign v2553 = ~(w5937 | w5938);
assign w5940 = v2553;
assign v2554 = ~(w5939 | w5940);
assign w5941 = v2554;
assign w5942 = w5936 & ~w5941;
assign w5943 = ~w5936 & w5941;
assign v2555 = ~(w5942 | w5943);
assign w5944 = v2555;
assign w5945 = (~w5736 & ~w5730) | (~w5736 & w8822) | (~w5730 & w8822);
assign w5946 = (~w5725 & ~w5727) | (~w5725 & w8823) | (~w5727 & w8823);
assign v2556 = ~(w5733 | w5946);
assign w5947 = v2556;
assign w5948 = w5733 & w5946;
assign v2557 = ~(w5947 | w5948);
assign w5949 = v2557;
assign w5950 = ~w5945 & w5949;
assign w5951 = w5945 & ~w5949;
assign v2558 = ~(w5950 | w5951);
assign w5952 = v2558;
assign w5953 = (~w5886 & ~w5888) | (~w5886 & w8768) | (~w5888 & w8768);
assign v2559 = ~(w5792 | w5820);
assign w5954 = v2559;
assign w5955 = (~w5880 & ~w5882) | (~w5880 & w8824) | (~w5882 & w8824);
assign v2560 = ~(w5954 | w5955);
assign w5956 = v2560;
assign w5957 = w5954 & w5955;
assign v2561 = ~(w5956 | w5957);
assign w5958 = v2561;
assign w5959 = w5958 & w5953;
assign w5960 = (w5888 & w9280) | (w5888 & w9281) | (w9280 & w9281);
assign v2562 = ~(w5959 | w5960);
assign w5961 = v2562;
assign w5962 = w5952 & w5961;
assign v2563 = ~(w5952 | w5961);
assign w5963 = v2563;
assign v2564 = ~(w5962 | w5963);
assign w5964 = v2564;
assign w5965 = w5944 & w5964;
assign v2565 = ~(w5944 | w5964);
assign w5966 = v2565;
assign v2566 = ~(w5965 | w5966);
assign w5967 = v2566;
assign w5968 = pi25 & pi46;
assign w5969 = pi29 & pi42;
assign w5970 = pi31 & pi40;
assign w5971 = pi30 & pi41;
assign w5972 = ~w5970 & w5971;
assign w5973 = w5970 & ~w5971;
assign v2567 = ~(w5972 | w5973);
assign w5974 = v2567;
assign w5975 = w5969 & w5974;
assign v2568 = ~(w5969 | w5974);
assign w5976 = v2568;
assign v2569 = ~(w5975 | w5976);
assign w5977 = v2569;
assign w5978 = w5968 & w5977;
assign v2570 = ~(w5968 | w5977);
assign w5979 = v2570;
assign v2571 = ~(w5978 | w5979);
assign w5980 = v2571;
assign w5981 = pi26 & pi45;
assign w5982 = pi27 & pi44;
assign v2572 = ~(w5781 | w5982);
assign w5983 = v2572;
assign w5984 = pi28 & pi44;
assign w5985 = w5779 & w5984;
assign v2573 = ~(w5983 | w5985);
assign w5986 = v2573;
assign w5987 = w5981 & ~w5986;
assign w5988 = ~w5981 & w5986;
assign v2574 = ~(w5987 | w5988);
assign w5989 = v2574;
assign w5990 = w5980 & ~w5989;
assign w5991 = ~w5980 & w5989;
assign v2575 = ~(w5990 | w5991);
assign w5992 = v2575;
assign w5993 = (~w5833 & ~w5835) | (~w5833 & w8639) | (~w5835 & w8639);
assign w5994 = w5836 & ~w5838;
assign v2576 = ~(w5840 | w5994);
assign w5995 = v2576;
assign w5996 = w5824 & ~w5826;
assign v2577 = ~(w5828 | w5996);
assign w5997 = v2577;
assign v2578 = ~(w5995 | w5997);
assign w5998 = v2578;
assign w5999 = w5995 & w5997;
assign v2579 = ~(w5998 | w5999);
assign w6000 = v2579;
assign w6001 = ~w5993 & w6000;
assign w6002 = w5993 & ~w6000;
assign v2580 = ~(w6001 | w6002);
assign w6003 = v2580;
assign w6004 = w5896 & w6003;
assign v2581 = ~(w5896 | w6003);
assign w6005 = v2581;
assign v2582 = ~(w6004 | w6005);
assign w6006 = v2582;
assign w6007 = w5992 & w6006;
assign v2583 = ~(w5992 | w6006);
assign w6008 = v2583;
assign v2584 = ~(w6007 | w6008);
assign w6009 = v2584;
assign w6010 = pi18 & pi53;
assign w6011 = pi22 & pi49;
assign w6012 = pi23 & pi48;
assign v2585 = ~(w5799 | w6012);
assign w6013 = v2585;
assign w6014 = pi24 & pi48;
assign w6015 = w5797 & w6014;
assign v2586 = ~(w6013 | w6015);
assign w6016 = v2586;
assign w6017 = w6011 & ~w6016;
assign w6018 = ~w6011 & w6016;
assign v2587 = ~(w6017 | w6018);
assign w6019 = v2587;
assign w6020 = w6010 & ~w6019;
assign w6021 = ~w6010 & w6019;
assign v2588 = ~(w6020 | w6021);
assign w6022 = v2588;
assign w6023 = pi19 & pi52;
assign w6024 = pi20 & pi51;
assign v2589 = ~(w5811 | w6024);
assign w6025 = v2589;
assign w6026 = pi21 & pi51;
assign w6027 = w5809 & w6026;
assign v2590 = ~(w6025 | w6027);
assign w6028 = v2590;
assign w6029 = w6023 & ~w6028;
assign w6030 = ~w6023 & w6028;
assign v2591 = ~(w6029 | w6030);
assign w6031 = v2591;
assign w6032 = w6022 & ~w6031;
assign w6033 = ~w6022 & w6031;
assign v2592 = ~(w6032 | w6033);
assign w6034 = v2592;
assign w6035 = (~w5805 & ~w5807) | (~w5805 & w8640) | (~w5807 & w8640);
assign w6036 = w5808 & ~w5810;
assign v2593 = ~(w5812 | w6036);
assign w6037 = v2593;
assign w6038 = w5796 & ~w5798;
assign v2594 = ~(w5800 | w6038);
assign w6039 = v2594;
assign v2595 = ~(w6037 | w6039);
assign w6040 = v2595;
assign w6041 = w6037 & w6039;
assign v2596 = ~(w6040 | w6041);
assign w6042 = v2596;
assign w6043 = ~w6035 & w6042;
assign w6044 = w6035 & ~w6042;
assign v2597 = ~(w6043 | w6044);
assign w6045 = v2597;
assign w6046 = (~w5853 & w5848) | (~w5853 & w8769) | (w5848 & w8769);
assign w6047 = (~w5775 & ~w5777) | (~w5775 & w8641) | (~w5777 & w8641);
assign v2598 = ~(w5769 | w5772);
assign w6048 = v2598;
assign w6049 = w5778 & ~w5780;
assign v2599 = ~(w5782 | w6049);
assign w6050 = v2599;
assign v2600 = ~(w6048 | w6050);
assign w6051 = v2600;
assign w6052 = w6048 & w6050;
assign v2601 = ~(w6051 | w6052);
assign w6053 = v2601;
assign w6054 = ~w6047 & w6053;
assign w6055 = w6047 & ~w6053;
assign v2602 = ~(w6054 | w6055);
assign w6056 = v2602;
assign w6057 = ~w6046 & w6056;
assign w6058 = w6046 & ~w6056;
assign v2603 = ~(w6057 | w6058);
assign w6059 = v2603;
assign w6060 = w6045 & w6059;
assign v2604 = ~(w6045 | w6059);
assign w6061 = v2604;
assign v2605 = ~(w6060 | w6061);
assign w6062 = v2605;
assign v2606 = ~(w6034 | w6062);
assign w6063 = v2606;
assign w6064 = w6034 & w6062;
assign v2607 = ~(w6063 | w6064);
assign w6065 = v2607;
assign w6066 = ~w6009 & w6065;
assign w6067 = w6009 & ~w6065;
assign v2608 = ~(w6066 | w6067);
assign w6068 = v2608;
assign w6069 = (~w5753 & w5750) | (~w5753 & w8825) | (w5750 & w8825);
assign w6070 = pi15 & pi56;
assign w6071 = pi16 & pi55;
assign v2609 = ~(w5827 | w6071);
assign w6072 = v2609;
assign w6073 = pi17 & pi55;
assign w6074 = w5825 & w6073;
assign v2610 = ~(w6072 | w6074);
assign w6075 = v2610;
assign w6076 = w6070 & ~w6075;
assign w6077 = ~w6070 & w6075;
assign v2611 = ~(w6076 | w6077);
assign w6078 = v2611;
assign w6079 = pi12 & pi59;
assign w6080 = pi13 & pi58;
assign v2612 = ~(w5839 | w6080);
assign w6081 = v2612;
assign w6082 = pi14 & pi58;
assign w6083 = w5837 & w6082;
assign v2613 = ~(w6081 | w6083);
assign w6084 = v2613;
assign w6085 = w6079 & ~w6084;
assign w6086 = ~w6079 & w6084;
assign v2614 = ~(w6085 | w6086);
assign w6087 = v2614;
assign v2615 = ~(w6078 | w6087);
assign w6088 = v2615;
assign w6089 = w6078 & w6087;
assign v2616 = ~(w6088 | w6089);
assign w6090 = v2616;
assign w6091 = ~w5747 & w8985;
assign w6092 = (w6090 & w5747) | (w6090 & w8986) | (w5747 & w8986);
assign v2617 = ~(w6091 | w6092);
assign w6093 = v2617;
assign w6094 = w6069 & w6093;
assign v2618 = ~(w6069 | w6093);
assign w6095 = v2618;
assign v2619 = ~(w6094 | w6095);
assign w6096 = v2619;
assign v2620 = ~(w6068 | w6096);
assign w6097 = v2620;
assign w6098 = w6068 & w6096;
assign v2621 = ~(w6097 | w6098);
assign w6099 = v2621;
assign w6100 = w5967 & w6099;
assign v2622 = ~(w5967 | w6099);
assign w6101 = v2622;
assign v2623 = ~(w6100 | w6101);
assign w6102 = v2623;
assign w6103 = (~w5715 & w5712) | (~w5715 & w9170) | (w5712 & w9170);
assign w6104 = (~w5904 & ~w5764) | (~w5904 & w8826) | (~w5764 & w8826);
assign v2624 = ~(w5898 | w5901);
assign w6105 = v2624;
assign w6106 = (~w5759 & ~w5761) | (~w5759 & w8827) | (~w5761 & w8827);
assign w6107 = w6105 & ~w6106;
assign w6108 = ~w6105 & w6106;
assign v2625 = ~(w6107 | w6108);
assign w6109 = v2625;
assign w6110 = ~w6104 & w6109;
assign w6111 = w6104 & ~w6109;
assign v2626 = ~(w6110 | w6111);
assign w6112 = v2626;
assign w6113 = ~w6103 & w6112;
assign w6114 = w6103 & ~w6112;
assign v2627 = ~(w6113 | w6114);
assign w6115 = v2627;
assign w6116 = w6102 & w6115;
assign v2628 = ~(w6102 | w6115);
assign w6117 = v2628;
assign v2629 = ~(w6116 | w6117);
assign w6118 = v2629;
assign w6119 = w5923 & ~w6118;
assign w6120 = ~w5923 & w6118;
assign v2630 = ~(w6119 | w6120);
assign w6121 = v2630;
assign w6122 = w5921 & ~w6121;
assign w6123 = ~w5921 & w6121;
assign v2631 = ~(w6122 | w6123);
assign w6124 = v2631;
assign v2632 = ~(w5915 | w6119);
assign w6125 = v2632;
assign w6126 = w5486 & w5706;
assign w6127 = w6125 & w6126;
assign w6128 = ~w5263 & w6127;
assign w6129 = w5484 & ~w5704;
assign v2633 = ~(w5705 | w5914);
assign w6130 = v2633;
assign w6131 = ~w6120 & w9302;
assign w6132 = ~w6128 & w6131;
assign w6133 = ~w4262 & w5916;
assign w6134 = w6121 & w6133;
assign w6135 = w6126 & w6134;
assign w6136 = w5260 & w6135;
assign w6137 = ~w4520 & w6136;
assign w6138 = w6132 & ~w6137;
assign w6139 = (~w6113 & ~w6115) | (~w6113 & w8987) | (~w6115 & w8987);
assign w6140 = pi09 & pi63;
assign w6141 = pi10 & pi62;
assign w6142 = w6140 & ~w6141;
assign w6143 = ~w6140 & w6141;
assign v2634 = ~(w6142 | w6143);
assign w6144 = v2634;
assign w6145 = (~w6051 & w6047) | (~w6051 & w8828) | (w6047 & w8828);
assign w6146 = pi13 & pi59;
assign w6147 = pi12 & pi60;
assign v2635 = ~(w6146 | w6147);
assign w6148 = v2635;
assign w6149 = pi13 & pi60;
assign w6150 = w6079 & w6149;
assign v2636 = ~(w6148 | w6150);
assign w6151 = v2636;
assign w6152 = w5928 & ~w6151;
assign w6153 = ~w5928 & w6151;
assign v2637 = ~(w6152 | w6153);
assign w6154 = v2637;
assign v2638 = ~(w6145 | w6154);
assign w6155 = v2638;
assign w6156 = w6145 & w6154;
assign v2639 = ~(w6155 | w6156);
assign w6157 = v2639;
assign w6158 = ~w6144 & w6157;
assign w6159 = w6144 & ~w6157;
assign v2640 = ~(w6158 | w6159);
assign w6160 = v2640;
assign v2641 = ~(w5934 | w5942);
assign w6161 = v2641;
assign w6162 = w5925 & ~w5927;
assign v2642 = ~(w5929 | w6162);
assign w6163 = v2642;
assign v2643 = ~(w5939 | w6163);
assign w6164 = v2643;
assign w6165 = w5939 & w6163;
assign v2644 = ~(w6164 | w6165);
assign w6166 = v2644;
assign w6167 = ~w6161 & w6166;
assign w6168 = w6161 & ~w6166;
assign v2645 = ~(w6167 | w6168);
assign w6169 = v2645;
assign w6170 = (~w6063 & ~w6065) | (~w6063 & w8771) | (~w6065 & w8771);
assign w6171 = (~w6004 & ~w6006) | (~w6004 & w8829) | (~w6006 & w8829);
assign w6172 = (~w6057 & ~w6059) | (~w6057 & w8830) | (~w6059 & w8830);
assign v2646 = ~(w6171 | w6172);
assign w6173 = v2646;
assign w6174 = w6171 & w6172;
assign v2647 = ~(w6173 | w6174);
assign w6175 = v2647;
assign w6176 = w6170 & w6175;
assign v2648 = ~(w6170 | w6175);
assign w6177 = v2648;
assign v2649 = ~(w6176 | w6177);
assign w6178 = v2649;
assign w6179 = w6169 & w6178;
assign v2650 = ~(w6169 | w6178);
assign w6180 = v2650;
assign v2651 = ~(w6179 | w6180);
assign w6181 = v2651;
assign w6182 = w6160 & w6181;
assign v2652 = ~(w6160 | w6181);
assign w6183 = v2652;
assign v2653 = ~(w6182 | w6183);
assign w6184 = v2653;
assign w6185 = pi25 & pi47;
assign w6186 = pi29 & pi43;
assign w6187 = pi31 & pi41;
assign w6188 = pi30 & pi42;
assign w6189 = ~w6187 & w6188;
assign w6190 = w6187 & ~w6188;
assign v2654 = ~(w6189 | w6190);
assign w6191 = v2654;
assign w6192 = w6186 & w6191;
assign v2655 = ~(w6186 | w6191);
assign w6193 = v2655;
assign v2656 = ~(w6192 | w6193);
assign w6194 = v2656;
assign w6195 = w6185 & w6194;
assign v2657 = ~(w6185 | w6194);
assign w6196 = v2657;
assign v2658 = ~(w6195 | w6196);
assign w6197 = v2658;
assign w6198 = pi26 & pi46;
assign w6199 = pi27 & pi45;
assign v2659 = ~(w5984 | w6199);
assign w6200 = v2659;
assign w6201 = pi28 & pi45;
assign w6202 = w5982 & w6201;
assign v2660 = ~(w6200 | w6202);
assign w6203 = v2660;
assign w6204 = w6198 & ~w6203;
assign w6205 = ~w6198 & w6203;
assign v2661 = ~(w6204 | w6205);
assign w6206 = v2661;
assign w6207 = w6197 & ~w6206;
assign w6208 = ~w6197 & w6206;
assign v2662 = ~(w6207 | w6208);
assign w6209 = v2662;
assign w6210 = w6079 & ~w6081;
assign v2663 = ~(w6083 | w6210);
assign w6211 = v2663;
assign w6212 = w6070 & ~w6072;
assign v2664 = ~(w6074 | w6212);
assign w6213 = v2664;
assign v2665 = ~(w6211 | w6213);
assign w6214 = v2665;
assign w6215 = w6211 & w6213;
assign v2666 = ~(w6214 | w6215);
assign w6216 = v2666;
assign w6217 = w6088 & w6216;
assign v2667 = ~(w6088 | w6216);
assign w6218 = v2667;
assign v2668 = ~(w6217 | w6218);
assign w6219 = v2668;
assign w6220 = (~w6020 & ~w6022) | (~w6020 & w8642) | (~w6022 & w8642);
assign w6221 = w6023 & ~w6025;
assign v2669 = ~(w6027 | w6221);
assign w6222 = v2669;
assign w6223 = w6011 & ~w6013;
assign v2670 = ~(w6015 | w6223);
assign w6224 = v2670;
assign v2671 = ~(w6222 | w6224);
assign w6225 = v2671;
assign w6226 = w6222 & w6224;
assign v2672 = ~(w6225 | w6226);
assign w6227 = v2672;
assign w6228 = ~w6220 & w6227;
assign w6229 = w6220 & ~w6227;
assign v2673 = ~(w6228 | w6229);
assign w6230 = v2673;
assign w6231 = w6219 & w6230;
assign v2674 = ~(w6219 | w6230);
assign w6232 = v2674;
assign v2675 = ~(w6231 | w6232);
assign w6233 = v2675;
assign w6234 = w6209 & w6233;
assign v2676 = ~(w6209 | w6233);
assign w6235 = v2676;
assign v2677 = ~(w6234 | w6235);
assign w6236 = v2677;
assign w6237 = pi18 & pi54;
assign w6238 = pi22 & pi50;
assign w6239 = pi23 & pi49;
assign v2678 = ~(w6014 | w6239);
assign w6240 = v2678;
assign w6241 = pi24 & pi49;
assign w6242 = w6012 & w6241;
assign v2679 = ~(w6240 | w6242);
assign w6243 = v2679;
assign w6244 = w6238 & ~w6243;
assign w6245 = ~w6238 & w6243;
assign v2680 = ~(w6244 | w6245);
assign w6246 = v2680;
assign w6247 = w6237 & ~w6246;
assign w6248 = ~w6237 & w6246;
assign v2681 = ~(w6247 | w6248);
assign w6249 = v2681;
assign w6250 = pi19 & pi53;
assign w6251 = pi20 & pi52;
assign v2682 = ~(w6026 | w6251);
assign w6252 = v2682;
assign w6253 = pi21 & pi52;
assign w6254 = w6024 & w6253;
assign v2683 = ~(w6252 | w6254);
assign w6255 = v2683;
assign w6256 = w6250 & ~w6255;
assign w6257 = ~w6250 & w6255;
assign v2684 = ~(w6256 | w6257);
assign w6258 = v2684;
assign w6259 = w6249 & ~w6258;
assign w6260 = ~w6249 & w6258;
assign v2685 = ~(w6259 | w6260);
assign w6261 = v2685;
assign w6262 = (~w5978 & ~w5980) | (~w5978 & w8772) | (~w5980 & w8772);
assign w6263 = (~w5972 & ~w5974) | (~w5972 & w8988) | (~w5974 & w8988);
assign w6264 = w5981 & ~w5983;
assign v2686 = ~(w5985 | w6264);
assign w6265 = v2686;
assign v2687 = ~(w6263 | w6265);
assign w6266 = v2687;
assign w6267 = w6263 & w6265;
assign v2688 = ~(w6266 | w6267);
assign w6268 = v2688;
assign w6269 = ~w6262 & w6268;
assign w6270 = w6262 & ~w6268;
assign v2689 = ~(w6269 | w6270);
assign w6271 = v2689;
assign w6272 = (~w6040 & w6035) | (~w6040 & w8643) | (w6035 & w8643);
assign w6273 = (~w5998 & w5993) | (~w5998 & w8644) | (w5993 & w8644);
assign v2690 = ~(w6272 | w6273);
assign w6274 = v2690;
assign w6275 = w6272 & w6273;
assign v2691 = ~(w6274 | w6275);
assign w6276 = v2691;
assign w6277 = w6271 & w6276;
assign v2692 = ~(w6271 | w6276);
assign w6278 = v2692;
assign v2693 = ~(w6277 | w6278);
assign w6279 = v2693;
assign v2694 = ~(w6261 | w6279);
assign w6280 = v2694;
assign w6281 = w6261 & w6279;
assign v2695 = ~(w6280 | w6281);
assign w6282 = v2695;
assign w6283 = ~w6236 & w6282;
assign w6284 = w6236 & ~w6282;
assign v2696 = ~(w6283 | w6284);
assign w6285 = v2696;
assign w6286 = (~w5956 & ~w5953) | (~w5956 & w8645) | (~w5953 & w8645);
assign w6287 = pi15 & pi57;
assign w6288 = pi16 & pi56;
assign v2697 = ~(w6073 | w6288);
assign w6289 = v2697;
assign w6290 = pi17 & pi56;
assign w6291 = w6071 & w6290;
assign v2698 = ~(w6289 | w6291);
assign w6292 = v2698;
assign w6293 = w6287 & w6292;
assign v2699 = ~(w6287 | w6292);
assign w6294 = v2699;
assign v2700 = ~(w6293 | w6294);
assign w6295 = v2700;
assign w6296 = w6082 & w6295;
assign v2701 = ~(w6082 | w6295);
assign w6297 = v2701;
assign v2702 = ~(w6296 | w6297);
assign w6298 = v2702;
assign w6299 = (w6298 & w5950) | (w6298 & w8646) | (w5950 & w8646);
assign w6300 = ~w5950 & w8647;
assign v2703 = ~(w6299 | w6300);
assign w6301 = v2703;
assign w6302 = ~w6286 & w6301;
assign w6303 = w6286 & ~w6301;
assign v2704 = ~(w6302 | w6303);
assign w6304 = v2704;
assign w6305 = ~w6285 & w6304;
assign w6306 = w6285 & ~w6304;
assign v2705 = ~(w6305 | w6306);
assign w6307 = v2705;
assign w6308 = w6184 & w6307;
assign v2706 = ~(w6184 | w6307);
assign w6309 = v2706;
assign v2707 = ~(w6308 | w6309);
assign w6310 = v2707;
assign w6311 = (~w6107 & w6104) | (~w6107 & w9171) | (w6104 & w9171);
assign w6312 = (~w6097 & ~w5967) | (~w6097 & w8831) | (~w5967 & w8831);
assign v2708 = ~(w6091 | w6094);
assign w6313 = v2708;
assign w6314 = (w5964 & w9172) | (w5964 & w9173) | (w9172 & w9173);
assign w6315 = ~w6313 & w9303;
assign v2709 = ~(w6314 | w6315);
assign w6316 = v2709;
assign w6317 = ~w6312 & w6316;
assign w6318 = w6312 & ~w6316;
assign v2710 = ~(w6317 | w6318);
assign w6319 = v2710;
assign w6320 = ~w6311 & w6319;
assign w6321 = w6311 & ~w6319;
assign v2711 = ~(w6320 | w6321);
assign w6322 = v2711;
assign w6323 = w6310 & w6322;
assign v2712 = ~(w6310 | w6322);
assign w6324 = v2712;
assign v2713 = ~(w6323 | w6324);
assign w6325 = v2713;
assign w6326 = ~w6139 & w6325;
assign w6327 = w6139 & ~w6325;
assign v2714 = ~(w6326 | w6327);
assign w6328 = v2714;
assign w6329 = (w6328 & w6137) | (w6328 & w8832) | (w6137 & w8832);
assign w6330 = w6138 & ~w6328;
assign v2715 = ~(w6329 | w6330);
assign w6331 = v2715;
assign w6332 = (~w6137 & w8879) | (~w6137 & w8880) | (w8879 & w8880);
assign w6333 = (~w6320 & ~w6322) | (~w6320 & w8649) | (~w6322 & w8649);
assign w6334 = pi10 & pi63;
assign w6335 = pi11 & pi62;
assign w6336 = w6334 & ~w6335;
assign w6337 = ~w6334 & w6335;
assign v2716 = ~(w6336 | w6337);
assign w6338 = v2716;
assign w6339 = pi12 & pi61;
assign w6340 = pi14 & pi59;
assign v2717 = ~(w6149 | w6340);
assign w6341 = v2717;
assign w6342 = pi14 & pi60;
assign w6343 = w6146 & w6342;
assign v2718 = ~(w6341 | w6343);
assign w6344 = v2718;
assign w6345 = w6339 & ~w6344;
assign w6346 = ~w6339 & w6344;
assign v2719 = ~(w6345 | w6346);
assign w6347 = v2719;
assign w6348 = ~w6347 & w9304;
assign w6349 = (w6262 & w8989) | (w6262 & w8990) | (w8989 & w8990);
assign v2720 = ~(w6348 | w6349);
assign w6350 = v2720;
assign w6351 = ~w6338 & w6350;
assign w6352 = w6338 & ~w6350;
assign v2721 = ~(w6351 | w6352);
assign w6353 = v2721;
assign w6354 = (~w6155 & ~w6157) | (~w6155 & w8882) | (~w6157 & w8882);
assign w6355 = w5928 & ~w6148;
assign v2722 = ~(w6150 | w6355);
assign w6356 = v2722;
assign v2723 = ~(w6142 | w6356);
assign w6357 = v2723;
assign w6358 = w6142 & w6356;
assign v2724 = ~(w6357 | w6358);
assign w6359 = v2724;
assign w6360 = ~w6354 & w6359;
assign w6361 = w6354 & ~w6359;
assign v2725 = ~(w6360 | w6361);
assign w6362 = v2725;
assign w6363 = (~w6280 & ~w6282) | (~w6280 & w8773) | (~w6282 & w8773);
assign w6364 = (~w6231 & ~w6233) | (~w6231 & w8833) | (~w6233 & w8833);
assign w6365 = (~w6274 & ~w6276) | (~w6274 & w8883) | (~w6276 & w8883);
assign v2726 = ~(w6364 | w6365);
assign w6366 = v2726;
assign w6367 = w6364 & w6365;
assign v2727 = ~(w6366 | w6367);
assign w6368 = v2727;
assign w6369 = w6363 & w6368;
assign v2728 = ~(w6363 | w6368);
assign w6370 = v2728;
assign v2729 = ~(w6369 | w6370);
assign w6371 = v2729;
assign w6372 = w6362 & w6371;
assign v2730 = ~(w6362 | w6371);
assign w6373 = v2730;
assign v2731 = ~(w6372 | w6373);
assign w6374 = v2731;
assign w6375 = w6353 & w6374;
assign v2732 = ~(w6353 | w6374);
assign w6376 = v2732;
assign v2733 = ~(w6375 | w6376);
assign w6377 = v2733;
assign w6378 = (~w6173 & ~w6170) | (~w6173 & w8650) | (~w6170 & w8650);
assign v2734 = ~(w6164 | w6167);
assign w6379 = v2734;
assign w6380 = pi15 & pi58;
assign w6381 = pi16 & pi57;
assign v2735 = ~(w6290 | w6381);
assign w6382 = v2735;
assign w6383 = pi17 & pi57;
assign w6384 = w6288 & w6383;
assign v2736 = ~(w6382 | w6384);
assign w6385 = v2736;
assign w6386 = w6380 & ~w6385;
assign w6387 = ~w6380 & w6385;
assign v2737 = ~(w6386 | w6387);
assign w6388 = v2737;
assign v2738 = ~(w6379 | w6388);
assign w6389 = v2738;
assign w6390 = w6379 & w6388;
assign v2739 = ~(w6389 | w6390);
assign w6391 = v2739;
assign w6392 = ~w6378 & w6391;
assign w6393 = w6378 & ~w6391;
assign v2740 = ~(w6392 | w6393);
assign w6394 = v2740;
assign w6395 = pi25 & pi48;
assign w6396 = pi29 & pi44;
assign w6397 = pi31 & pi42;
assign w6398 = pi30 & pi43;
assign w6399 = ~w6397 & w6398;
assign w6400 = w6397 & ~w6398;
assign v2741 = ~(w6399 | w6400);
assign w6401 = v2741;
assign w6402 = w6396 & w6401;
assign v2742 = ~(w6396 | w6401);
assign w6403 = v2742;
assign v2743 = ~(w6402 | w6403);
assign w6404 = v2743;
assign w6405 = w6395 & w6404;
assign v2744 = ~(w6395 | w6404);
assign w6406 = v2744;
assign v2745 = ~(w6405 | w6406);
assign w6407 = v2745;
assign w6408 = pi26 & pi47;
assign w6409 = pi27 & pi46;
assign v2746 = ~(w6201 | w6409);
assign w6410 = v2746;
assign w6411 = pi28 & pi46;
assign w6412 = w6199 & w6411;
assign v2747 = ~(w6410 | w6412);
assign w6413 = v2747;
assign w6414 = w6408 & ~w6413;
assign w6415 = ~w6408 & w6413;
assign v2748 = ~(w6414 | w6415);
assign w6416 = v2748;
assign w6417 = w6407 & ~w6416;
assign w6418 = ~w6407 & w6416;
assign v2749 = ~(w6417 | w6418);
assign w6419 = v2749;
assign w6420 = (~w6247 & ~w6249) | (~w6247 & w8651) | (~w6249 & w8651);
assign w6421 = w6250 & ~w6252;
assign v2750 = ~(w6254 | w6421);
assign w6422 = v2750;
assign w6423 = w6238 & ~w6240;
assign v2751 = ~(w6242 | w6423);
assign w6424 = v2751;
assign v2752 = ~(w6422 | w6424);
assign w6425 = v2752;
assign w6426 = w6422 & w6424;
assign v2753 = ~(w6425 | w6426);
assign w6427 = v2753;
assign w6428 = ~w6420 & w6427;
assign w6429 = w6420 & ~w6427;
assign v2754 = ~(w6428 | w6429);
assign w6430 = v2754;
assign v2755 = ~(w6291 | w6296);
assign w6431 = v2755;
assign w6432 = w6295 & w8884;
assign v2756 = ~(w6431 | w6432);
assign w6433 = v2756;
assign v2757 = ~(w6293 | w6433);
assign w6434 = v2757;
assign w6435 = w6430 & ~w6434;
assign w6436 = ~w6430 & w6434;
assign v2758 = ~(w6435 | w6436);
assign w6437 = v2758;
assign w6438 = w6419 & w6437;
assign v2759 = ~(w6419 | w6437);
assign w6439 = v2759;
assign v2760 = ~(w6438 | w6439);
assign w6440 = v2760;
assign w6441 = pi18 & pi55;
assign w6442 = pi22 & pi51;
assign w6443 = pi23 & pi50;
assign v2761 = ~(w6241 | w6443);
assign w6444 = v2761;
assign w6445 = pi24 & pi50;
assign w6446 = w6239 & w6445;
assign v2762 = ~(w6444 | w6446);
assign w6447 = v2762;
assign w6448 = w6442 & ~w6447;
assign w6449 = ~w6442 & w6447;
assign v2763 = ~(w6448 | w6449);
assign w6450 = v2763;
assign w6451 = w6441 & ~w6450;
assign w6452 = ~w6441 & w6450;
assign v2764 = ~(w6451 | w6452);
assign w6453 = v2764;
assign w6454 = pi19 & pi54;
assign w6455 = pi20 & pi53;
assign v2765 = ~(w6253 | w6455);
assign w6456 = v2765;
assign w6457 = pi21 & pi53;
assign w6458 = w6251 & w6457;
assign v2766 = ~(w6456 | w6458);
assign w6459 = v2766;
assign w6460 = w6454 & ~w6459;
assign w6461 = ~w6454 & w6459;
assign v2767 = ~(w6460 | w6461);
assign w6462 = v2767;
assign w6463 = w6453 & ~w6462;
assign w6464 = ~w6453 & w6462;
assign v2768 = ~(w6463 | w6464);
assign w6465 = v2768;
assign w6466 = (~w6195 & ~w6197) | (~w6195 & w8774) | (~w6197 & w8774);
assign v2769 = ~(w6189 | w6192);
assign w6467 = v2769;
assign w6468 = w6198 & ~w6200;
assign v2770 = ~(w6202 | w6468);
assign w6469 = v2770;
assign v2771 = ~(w6467 | w6469);
assign w6470 = v2771;
assign w6471 = w6467 & w6469;
assign v2772 = ~(w6470 | w6471);
assign w6472 = v2772;
assign w6473 = ~w6466 & w6472;
assign w6474 = w6466 & ~w6472;
assign v2773 = ~(w6473 | w6474);
assign w6475 = v2773;
assign w6476 = (~w6225 & w6220) | (~w6225 & w8652) | (w6220 & w8652);
assign v2774 = ~(w6214 | w6217);
assign w6477 = v2774;
assign v2775 = ~(w6476 | w6477);
assign w6478 = v2775;
assign w6479 = w6476 & w6477;
assign v2776 = ~(w6478 | w6479);
assign w6480 = v2776;
assign w6481 = w6475 & w6480;
assign v2777 = ~(w6475 | w6480);
assign w6482 = v2777;
assign v2778 = ~(w6481 | w6482);
assign w6483 = v2778;
assign v2779 = ~(w6465 | w6483);
assign w6484 = v2779;
assign w6485 = w6465 & w6483;
assign v2780 = ~(w6484 | w6485);
assign w6486 = v2780;
assign w6487 = ~w6440 & w6486;
assign w6488 = w6440 & ~w6486;
assign v2781 = ~(w6487 | w6488);
assign w6489 = v2781;
assign w6490 = w6394 & ~w6489;
assign w6491 = ~w6394 & w6489;
assign v2782 = ~(w6490 | w6491);
assign w6492 = v2782;
assign w6493 = w6377 & w6492;
assign v2783 = ~(w6377 | w6492);
assign w6494 = v2783;
assign v2784 = ~(w6493 | w6494);
assign w6495 = v2784;
assign w6496 = (~w6314 & w6312) | (~w6314 & w8653) | (w6312 & w8653);
assign w6497 = (~w6305 & ~w6184) | (~w6305 & w8654) | (~w6184 & w8654);
assign v2785 = ~(w6299 | w6302);
assign w6498 = v2785;
assign w6499 = (w6181 & w9174) | (w6181 & w9175) | (w9174 & w9175);
assign w6500 = w6498 & w9305;
assign v2786 = ~(w6499 | w6500);
assign w6501 = v2786;
assign w6502 = ~w6497 & w6501;
assign w6503 = w6497 & ~w6501;
assign v2787 = ~(w6502 | w6503);
assign w6504 = v2787;
assign w6505 = ~w6496 & w6504;
assign w6506 = w6496 & ~w6504;
assign v2788 = ~(w6505 | w6506);
assign w6507 = v2788;
assign w6508 = w6495 & w6507;
assign v2789 = ~(w6495 | w6507);
assign w6509 = v2789;
assign v2790 = ~(w6508 | w6509);
assign w6510 = v2790;
assign w6511 = w6333 & ~w6510;
assign w6512 = ~w6333 & w6510;
assign v2791 = ~(w6511 | w6512);
assign w6513 = v2791;
assign w6514 = w6332 & ~w6513;
assign w6515 = ~w6332 & w6513;
assign v2792 = ~(w6514 | w6515);
assign w6516 = v2792;
assign w6517 = (~w6505 & ~w6507) | (~w6505 & w8885) | (~w6507 & w8885);
assign w6518 = pi11 & pi63;
assign w6519 = pi12 & pi62;
assign w6520 = w6518 & ~w6519;
assign w6521 = ~w6518 & w6519;
assign v2793 = ~(w6520 | w6521);
assign w6522 = v2793;
assign w6523 = (~w6470 & w6466) | (~w6470 & w8991) | (w6466 & w8991);
assign w6524 = pi13 & pi61;
assign w6525 = pi15 & pi59;
assign v2794 = ~(w6342 | w6525);
assign w6526 = v2794;
assign w6527 = pi15 & pi60;
assign w6528 = w6340 & w6527;
assign v2795 = ~(w6526 | w6528);
assign w6529 = v2795;
assign w6530 = w6524 & ~w6529;
assign w6531 = ~w6524 & w6529;
assign v2796 = ~(w6530 | w6531);
assign w6532 = v2796;
assign v2797 = ~(w6523 | w6532);
assign w6533 = v2797;
assign w6534 = w6523 & w6532;
assign v2798 = ~(w6533 | w6534);
assign w6535 = v2798;
assign w6536 = ~w6522 & w6535;
assign w6537 = w6522 & ~w6535;
assign v2799 = ~(w6536 | w6537);
assign w6538 = v2799;
assign v2800 = ~(w6348 | w6351);
assign w6539 = v2800;
assign w6540 = w6339 & ~w6341;
assign v2801 = ~(w6343 | w6540);
assign w6541 = v2801;
assign v2802 = ~(w6336 | w6541);
assign w6542 = v2802;
assign w6543 = w6336 & w6541;
assign v2803 = ~(w6542 | w6543);
assign w6544 = v2803;
assign w6545 = ~w6539 & w6544;
assign w6546 = w6539 & ~w6544;
assign v2804 = ~(w6545 | w6546);
assign w6547 = v2804;
assign w6548 = (~w6484 & ~w6486) | (~w6484 & w8775) | (~w6486 & w8775);
assign w6549 = (~w6435 & ~w6437) | (~w6435 & w8834) | (~w6437 & w8834);
assign w6550 = (~w6478 & ~w6480) | (~w6478 & w8992) | (~w6480 & w8992);
assign v2805 = ~(w6549 | w6550);
assign w6551 = v2805;
assign w6552 = w6549 & w6550;
assign v2806 = ~(w6551 | w6552);
assign w6553 = v2806;
assign w6554 = w6548 & w6553;
assign v2807 = ~(w6548 | w6553);
assign w6555 = v2807;
assign v2808 = ~(w6554 | w6555);
assign w6556 = v2808;
assign w6557 = w6547 & w6556;
assign v2809 = ~(w6547 | w6556);
assign w6558 = v2809;
assign v2810 = ~(w6557 | w6558);
assign w6559 = v2810;
assign w6560 = w6538 & w6559;
assign v2811 = ~(w6538 | w6559);
assign w6561 = v2811;
assign v2812 = ~(w6560 | w6561);
assign w6562 = v2812;
assign w6563 = pi25 & pi49;
assign w6564 = pi29 & pi45;
assign w6565 = pi31 & pi43;
assign w6566 = pi30 & pi44;
assign w6567 = ~w6565 & w6566;
assign w6568 = w6565 & ~w6566;
assign v2813 = ~(w6567 | w6568);
assign w6569 = v2813;
assign w6570 = w6564 & w6569;
assign v2814 = ~(w6564 | w6569);
assign w6571 = v2814;
assign v2815 = ~(w6570 | w6571);
assign w6572 = v2815;
assign w6573 = w6563 & w6572;
assign v2816 = ~(w6563 | w6572);
assign w6574 = v2816;
assign v2817 = ~(w6573 | w6574);
assign w6575 = v2817;
assign w6576 = pi26 & pi48;
assign w6577 = pi27 & pi47;
assign v2818 = ~(w6411 | w6577);
assign w6578 = v2818;
assign w6579 = pi28 & pi47;
assign w6580 = w6409 & w6579;
assign v2819 = ~(w6578 | w6580);
assign w6581 = v2819;
assign w6582 = w6576 & ~w6581;
assign w6583 = ~w6576 & w6581;
assign v2820 = ~(w6582 | w6583);
assign w6584 = v2820;
assign w6585 = w6575 & ~w6584;
assign w6586 = ~w6575 & w6584;
assign v2821 = ~(w6585 | w6586);
assign w6587 = v2821;
assign w6588 = (~w6451 & ~w6453) | (~w6451 & w8835) | (~w6453 & w8835);
assign w6589 = w6454 & ~w6456;
assign v2822 = ~(w6458 | w6589);
assign w6590 = v2822;
assign w6591 = w6442 & ~w6444;
assign v2823 = ~(w6446 | w6591);
assign w6592 = v2823;
assign v2824 = ~(w6590 | w6592);
assign w6593 = v2824;
assign w6594 = w6590 & w6592;
assign v2825 = ~(w6593 | w6594);
assign w6595 = v2825;
assign w6596 = ~w6588 & w6595;
assign w6597 = w6588 & ~w6595;
assign v2826 = ~(w6596 | w6597);
assign w6598 = v2826;
assign w6599 = w6380 & ~w6382;
assign v2827 = ~(w6384 | w6599);
assign w6600 = v2827;
assign w6601 = w6598 & ~w6600;
assign w6602 = ~w6598 & w6600;
assign v2828 = ~(w6601 | w6602);
assign w6603 = v2828;
assign w6604 = w6587 & w6603;
assign v2829 = ~(w6587 | w6603);
assign w6605 = v2829;
assign v2830 = ~(w6604 | w6605);
assign w6606 = v2830;
assign w6607 = pi18 & pi56;
assign w6608 = pi22 & pi52;
assign w6609 = pi23 & pi51;
assign v2831 = ~(w6445 | w6609);
assign w6610 = v2831;
assign w6611 = pi24 & pi51;
assign w6612 = w6443 & w6611;
assign v2832 = ~(w6610 | w6612);
assign w6613 = v2832;
assign w6614 = w6608 & ~w6613;
assign w6615 = ~w6608 & w6613;
assign v2833 = ~(w6614 | w6615);
assign w6616 = v2833;
assign w6617 = w6607 & ~w6616;
assign w6618 = ~w6607 & w6616;
assign v2834 = ~(w6617 | w6618);
assign w6619 = v2834;
assign w6620 = pi19 & pi55;
assign w6621 = pi20 & pi54;
assign v2835 = ~(w6457 | w6621);
assign w6622 = v2835;
assign w6623 = pi21 & pi54;
assign w6624 = w6455 & w6623;
assign v2836 = ~(w6622 | w6624);
assign w6625 = v2836;
assign w6626 = w6620 & ~w6625;
assign w6627 = ~w6620 & w6625;
assign v2837 = ~(w6626 | w6627);
assign w6628 = v2837;
assign w6629 = w6619 & ~w6628;
assign w6630 = ~w6619 & w6628;
assign v2838 = ~(w6629 | w6630);
assign w6631 = v2838;
assign w6632 = (~w6405 & ~w6407) | (~w6405 & w8836) | (~w6407 & w8836);
assign w6633 = (~w6399 & ~w6401) | (~w6399 & w8993) | (~w6401 & w8993);
assign w6634 = w6408 & ~w6410;
assign v2839 = ~(w6412 | w6634);
assign w6635 = v2839;
assign v2840 = ~(w6633 | w6635);
assign w6636 = v2840;
assign w6637 = w6633 & w6635;
assign v2841 = ~(w6636 | w6637);
assign w6638 = v2841;
assign w6639 = ~w6632 & w6638;
assign w6640 = w6632 & ~w6638;
assign v2842 = ~(w6639 | w6640);
assign w6641 = v2842;
assign w6642 = (~w6420 & w8837) | (~w6420 & w8838) | (w8837 & w8838);
assign w6643 = (w6420 & w8839) | (w6420 & w8840) | (w8839 & w8840);
assign v2843 = ~(w6642 | w6643);
assign w6644 = v2843;
assign w6645 = w6641 & w6644;
assign v2844 = ~(w6641 | w6644);
assign w6646 = v2844;
assign v2845 = ~(w6645 | w6646);
assign w6647 = v2845;
assign w6648 = w6631 & w6647;
assign v2846 = ~(w6631 | w6647);
assign w6649 = v2846;
assign v2847 = ~(w6648 | w6649);
assign w6650 = v2847;
assign w6651 = w6606 & w6650;
assign v2848 = ~(w6606 | w6650);
assign w6652 = v2848;
assign v2849 = ~(w6651 | w6652);
assign w6653 = v2849;
assign w6654 = (~w6366 & ~w6363) | (~w6366 & w8841) | (~w6363 & w8841);
assign w6655 = pi16 & pi58;
assign v2850 = ~(w6383 | w6655);
assign w6656 = v2850;
assign w6657 = pi17 & pi58;
assign w6658 = w6381 & w6657;
assign v2851 = ~(w6656 | w6658);
assign w6659 = v2851;
assign v2852 = ~(w6357 | w6360);
assign w6660 = v2852;
assign w6661 = ~w6659 & w6660;
assign w6662 = w6659 & ~w6660;
assign v2853 = ~(w6661 | w6662);
assign w6663 = v2853;
assign w6664 = w6654 & w6663;
assign v2854 = ~(w6654 | w6663);
assign w6665 = v2854;
assign v2855 = ~(w6664 | w6665);
assign w6666 = v2855;
assign w6667 = w6653 & ~w6666;
assign w6668 = ~w6653 & w6666;
assign v2856 = ~(w6667 | w6668);
assign w6669 = v2856;
assign w6670 = w6562 & w6669;
assign v2857 = ~(w6562 | w6669);
assign w6671 = v2857;
assign v2858 = ~(w6670 | w6671);
assign w6672 = v2858;
assign w6673 = (~w6499 & w6497) | (~w6499 & w9176) | (w6497 & w9176);
assign v2859 = ~(w6490 | w6493);
assign w6674 = v2859;
assign v2860 = ~(w6389 | w6392);
assign w6675 = v2860;
assign w6676 = (~w6372 & ~w6374) | (~w6372 & w8842) | (~w6374 & w8842);
assign v2861 = ~(w6675 | w6676);
assign w6677 = v2861;
assign w6678 = w6675 & w6676;
assign v2862 = ~(w6677 | w6678);
assign w6679 = v2862;
assign w6680 = ~w6674 & w6679;
assign w6681 = w6674 & ~w6679;
assign v2863 = ~(w6680 | w6681);
assign w6682 = v2863;
assign w6683 = ~w6673 & w6682;
assign w6684 = w6673 & ~w6682;
assign v2864 = ~(w6683 | w6684);
assign w6685 = v2864;
assign w6686 = w6672 & w6685;
assign v2865 = ~(w6672 | w6685);
assign w6687 = v2865;
assign v2866 = ~(w6686 | w6687);
assign w6688 = v2866;
assign w6689 = ~w6517 & w6688;
assign w6690 = w6517 & ~w6688;
assign v2867 = ~(w6689 | w6690);
assign w6691 = v2867;
assign w6692 = (w6137 & w8994) | (w6137 & w8995) | (w8994 & w8995);
assign w6693 = w6691 & w6692;
assign v2868 = ~(w6691 | w6692);
assign w6694 = v2868;
assign v2869 = ~(w6693 | w6694);
assign w6695 = v2869;
assign w6696 = (~w6137 & w9177) | (~w6137 & w9178) | (w9177 & w9178);
assign w6697 = (~w6683 & ~w6685) | (~w6683 & w8843) | (~w6685 & w8843);
assign w6698 = pi12 & pi63;
assign w6699 = pi16 & pi59;
assign w6700 = pi18 & pi57;
assign v2870 = ~(w6657 | w6700);
assign w6701 = v2870;
assign w6702 = pi18 & pi58;
assign w6703 = w6383 & w6702;
assign v2871 = ~(w6701 | w6703);
assign w6704 = v2871;
assign w6705 = w6699 & ~w6704;
assign w6706 = ~w6699 & w6704;
assign v2872 = ~(w6705 | w6706);
assign w6707 = v2872;
assign v2873 = ~(w6698 | w6707);
assign w6708 = v2873;
assign w6709 = w6698 & w6707;
assign v2874 = ~(w6708 | w6709);
assign w6710 = v2874;
assign w6711 = pi13 & pi62;
assign w6712 = pi14 & pi61;
assign v2875 = ~(w6527 | w6712);
assign w6713 = v2875;
assign w6714 = pi15 & pi61;
assign w6715 = w6342 & w6714;
assign v2876 = ~(w6713 | w6715);
assign w6716 = v2876;
assign w6717 = w6711 & ~w6716;
assign w6718 = ~w6711 & w6716;
assign v2877 = ~(w6717 | w6718);
assign w6719 = v2877;
assign w6720 = w6710 & ~w6719;
assign w6721 = ~w6710 & w6719;
assign v2878 = ~(w6720 | w6721);
assign w6722 = v2878;
assign v2879 = ~(w6533 | w6536);
assign w6723 = v2879;
assign w6724 = w6524 & ~w6526;
assign v2880 = ~(w6528 | w6724);
assign w6725 = v2880;
assign v2881 = ~(w6520 | w6725);
assign w6726 = v2881;
assign w6727 = w6520 & w6725;
assign v2882 = ~(w6726 | w6727);
assign w6728 = v2882;
assign w6729 = ~w6723 & w6728;
assign w6730 = w6723 & ~w6728;
assign v2883 = ~(w6729 | w6730);
assign w6731 = v2883;
assign v2884 = ~(w6648 | w6651);
assign w6732 = v2884;
assign w6733 = (~w6601 & ~w6603) | (~w6601 & w8887) | (~w6603 & w8887);
assign v2885 = ~(w6642 | w6645);
assign w6734 = v2885;
assign v2886 = ~(w6733 | w6734);
assign w6735 = v2886;
assign w6736 = w6733 & w6734;
assign v2887 = ~(w6735 | w6736);
assign w6737 = v2887;
assign w6738 = ~w6732 & w6737;
assign w6739 = w6732 & ~w6737;
assign v2888 = ~(w6738 | w6739);
assign w6740 = v2888;
assign w6741 = w6731 & w6740;
assign v2889 = ~(w6731 | w6740);
assign w6742 = v2889;
assign v2890 = ~(w6741 | w6742);
assign w6743 = v2890;
assign w6744 = w6722 & w6743;
assign v2891 = ~(w6722 | w6743);
assign w6745 = v2891;
assign v2892 = ~(w6744 | w6745);
assign w6746 = v2892;
assign w6747 = pi25 & pi50;
assign w6748 = pi29 & pi46;
assign w6749 = pi31 & pi44;
assign w6750 = pi30 & pi45;
assign w6751 = ~w6749 & w6750;
assign w6752 = w6749 & ~w6750;
assign v2893 = ~(w6751 | w6752);
assign w6753 = v2893;
assign w6754 = w6748 & w6753;
assign v2894 = ~(w6748 | w6753);
assign w6755 = v2894;
assign v2895 = ~(w6754 | w6755);
assign w6756 = v2895;
assign w6757 = w6747 & w6756;
assign v2896 = ~(w6747 | w6756);
assign w6758 = v2896;
assign v2897 = ~(w6757 | w6758);
assign w6759 = v2897;
assign w6760 = pi26 & pi49;
assign w6761 = pi27 & pi48;
assign v2898 = ~(w6579 | w6761);
assign w6762 = v2898;
assign w6763 = pi28 & pi48;
assign w6764 = w6577 & w6763;
assign v2899 = ~(w6762 | w6764);
assign w6765 = v2899;
assign w6766 = w6760 & ~w6765;
assign w6767 = ~w6760 & w6765;
assign v2900 = ~(w6766 | w6767);
assign w6768 = v2900;
assign w6769 = w6759 & ~w6768;
assign w6770 = ~w6759 & w6768;
assign v2901 = ~(w6769 | w6770);
assign w6771 = v2901;
assign w6772 = (~w6593 & w6588) | (~w6593 & w8888) | (w6588 & w8888);
assign w6773 = (~w6636 & w6632) | (~w6636 & w8889) | (w6632 & w8889);
assign w6774 = w6772 & w6773;
assign v2902 = ~(w6772 | w6773);
assign w6775 = v2902;
assign v2903 = ~(w6774 | w6775);
assign w6776 = v2903;
assign w6777 = w6771 & ~w6776;
assign w6778 = ~w6771 & w6776;
assign v2904 = ~(w6777 | w6778);
assign w6779 = v2904;
assign w6780 = (~w6617 & ~w6619) | (~w6617 & w8844) | (~w6619 & w8844);
assign w6781 = w6620 & ~w6622;
assign v2905 = ~(w6624 | w6781);
assign w6782 = v2905;
assign w6783 = w6608 & ~w6610;
assign v2906 = ~(w6612 | w6783);
assign w6784 = v2906;
assign v2907 = ~(w6782 | w6784);
assign w6785 = v2907;
assign w6786 = w6782 & w6784;
assign v2908 = ~(w6785 | w6786);
assign w6787 = v2908;
assign w6788 = ~w6780 & w6787;
assign w6789 = w6780 & ~w6787;
assign v2909 = ~(w6788 | w6789);
assign w6790 = v2909;
assign w6791 = (~w6573 & ~w6575) | (~w6573 & w8845) | (~w6575 & w8845);
assign w6792 = (~w6567 & ~w6569) | (~w6567 & w8996) | (~w6569 & w8996);
assign w6793 = w6576 & ~w6578;
assign v2910 = ~(w6580 | w6793);
assign w6794 = v2910;
assign v2911 = ~(w6792 | w6794);
assign w6795 = v2911;
assign w6796 = w6792 & w6794;
assign v2912 = ~(w6795 | w6796);
assign w6797 = v2912;
assign w6798 = ~w6791 & w6797;
assign w6799 = w6791 & ~w6797;
assign v2913 = ~(w6798 | w6799);
assign w6800 = v2913;
assign w6801 = w6790 & w6800;
assign v2914 = ~(w6790 | w6800);
assign w6802 = v2914;
assign v2915 = ~(w6801 | w6802);
assign w6803 = v2915;
assign w6804 = w6658 & w6803;
assign v2916 = ~(w6658 | w6803);
assign w6805 = v2916;
assign v2917 = ~(w6804 | w6805);
assign w6806 = v2917;
assign w6807 = w6779 & w6806;
assign v2918 = ~(w6779 | w6806);
assign w6808 = v2918;
assign v2919 = ~(w6807 | w6808);
assign w6809 = v2919;
assign w6810 = (~w6551 & ~w6548) | (~w6551 & w8890) | (~w6548 & w8890);
assign v2920 = ~(w6542 | w6545);
assign w6811 = v2920;
assign w6812 = pi19 & pi56;
assign w6813 = pi20 & pi55;
assign v2921 = ~(w6623 | w6813);
assign w6814 = v2921;
assign w6815 = pi21 & pi55;
assign w6816 = w6621 & w6815;
assign v2922 = ~(w6814 | w6816);
assign w6817 = v2922;
assign w6818 = w6812 & ~w6817;
assign w6819 = ~w6812 & w6817;
assign v2923 = ~(w6818 | w6819);
assign w6820 = v2923;
assign w6821 = pi22 & pi53;
assign w6822 = pi23 & pi52;
assign v2924 = ~(w6611 | w6822);
assign w6823 = v2924;
assign w6824 = pi24 & pi52;
assign w6825 = w6609 & w6824;
assign v2925 = ~(w6823 | w6825);
assign w6826 = v2925;
assign w6827 = w6821 & ~w6826;
assign w6828 = ~w6821 & w6826;
assign v2926 = ~(w6827 | w6828);
assign w6829 = v2926;
assign v2927 = ~(w6820 | w6829);
assign w6830 = v2927;
assign w6831 = w6820 & w6829;
assign v2928 = ~(w6830 | w6831);
assign w6832 = v2928;
assign w6833 = w6811 & ~w6832;
assign w6834 = ~w6811 & w6832;
assign v2929 = ~(w6833 | w6834);
assign w6835 = v2929;
assign w6836 = w6810 & w6835;
assign v2930 = ~(w6810 | w6835);
assign w6837 = v2930;
assign v2931 = ~(w6836 | w6837);
assign w6838 = v2931;
assign w6839 = w6809 & ~w6838;
assign w6840 = ~w6809 & w6838;
assign v2932 = ~(w6839 | w6840);
assign w6841 = v2932;
assign w6842 = w6746 & w6841;
assign v2933 = ~(w6746 | w6841);
assign w6843 = v2933;
assign v2934 = ~(w6842 | w6843);
assign w6844 = v2934;
assign w6845 = (~w6677 & w6674) | (~w6677 & w8846) | (w6674 & w8846);
assign w6846 = (~w6667 & ~w6562) | (~w6667 & w8847) | (~w6562 & w8847);
assign v2935 = ~(w6661 | w6664);
assign w6847 = v2935;
assign w6848 = (w6559 & w9179) | (w6559 & w9180) | (w9179 & w9180);
assign w6849 = ~w6847 & w9306;
assign v2936 = ~(w6848 | w6849);
assign w6850 = v2936;
assign w6851 = ~w6846 & w6850;
assign w6852 = w6846 & ~w6850;
assign v2937 = ~(w6851 | w6852);
assign w6853 = v2937;
assign w6854 = ~w6845 & w6853;
assign w6855 = w6845 & ~w6853;
assign v2938 = ~(w6854 | w6855);
assign w6856 = v2938;
assign w6857 = w6844 & w6856;
assign v2939 = ~(w6844 | w6856);
assign w6858 = v2939;
assign v2940 = ~(w6857 | w6858);
assign w6859 = v2940;
assign w6860 = ~w6697 & w6859;
assign w6861 = w6697 & ~w6859;
assign v2941 = ~(w6860 | w6861);
assign w6862 = v2941;
assign w6863 = w6696 & ~w6862;
assign w6864 = ~w6696 & w6862;
assign v2942 = ~(w6863 | w6864);
assign w6865 = v2942;
assign w6866 = w6326 & ~w6511;
assign v2943 = ~(w6512 | w6689);
assign w6867 = v2943;
assign w6868 = ~w6866 & w6867;
assign w6869 = ~w6690 & w6862;
assign w6870 = (~w6860 & w6868) | (~w6860 & w8656) | (w6868 & w8656);
assign w6871 = w6328 & ~w6511;
assign w6872 = w6871 & w8891;
assign w6873 = (~w4520 & w9181) | (~w4520 & w9182) | (w9181 & w9182);
assign w6874 = (~w6854 & ~w6856) | (~w6854 & w8997) | (~w6856 & w8997);
assign w6875 = pi14 & pi62;
assign w6876 = pi20 & pi56;
assign w6877 = pi19 & pi57;
assign v2944 = ~(w6876 | w6877);
assign w6878 = v2944;
assign w6879 = pi20 & pi57;
assign w6880 = w6812 & w6879;
assign v2945 = ~(w6878 | w6880);
assign w6881 = v2945;
assign w6882 = w6702 & ~w6881;
assign w6883 = ~w6702 & w6881;
assign v2946 = ~(w6882 | w6883);
assign w6884 = v2946;
assign w6885 = w6875 & ~w6884;
assign w6886 = ~w6875 & w6884;
assign v2947 = ~(w6885 | w6886);
assign w6887 = v2947;
assign w6888 = pi17 & pi59;
assign w6889 = pi16 & pi60;
assign v2948 = ~(w6888 | w6889);
assign w6890 = v2948;
assign w6891 = pi17 & pi60;
assign w6892 = w6699 & w6891;
assign v2949 = ~(w6890 | w6892);
assign w6893 = v2949;
assign w6894 = w6714 & ~w6893;
assign w6895 = ~w6714 & w6893;
assign v2950 = ~(w6894 | w6895);
assign w6896 = v2950;
assign w6897 = w6887 & ~w6896;
assign w6898 = ~w6887 & w6896;
assign v2951 = ~(w6897 | w6898);
assign w6899 = v2951;
assign v2952 = ~(w6708 | w6720);
assign w6900 = v2952;
assign w6901 = w6711 & ~w6713;
assign v2953 = ~(w6715 | w6901);
assign w6902 = v2953;
assign w6903 = w6699 & ~w6701;
assign v2954 = ~(w6703 | w6903);
assign w6904 = v2954;
assign v2955 = ~(w6902 | w6904);
assign w6905 = v2955;
assign w6906 = w6902 & w6904;
assign v2956 = ~(w6905 | w6906);
assign w6907 = v2956;
assign w6908 = ~w6900 & w6907;
assign w6909 = w6900 & ~w6907;
assign v2957 = ~(w6908 | w6909);
assign w6910 = v2957;
assign w6911 = (~w6777 & ~w6806) | (~w6777 & w8892) | (~w6806 & w8892);
assign w6912 = (~w6801 & ~w6803) | (~w6801 & w8850) | (~w6803 & w8850);
assign v2958 = ~(w6774 | w6912);
assign w6913 = v2958;
assign w6914 = w6774 & w6912;
assign v2959 = ~(w6913 | w6914);
assign w6915 = v2959;
assign w6916 = ~w6911 & w6915;
assign w6917 = w6911 & ~w6915;
assign v2960 = ~(w6916 | w6917);
assign w6918 = v2960;
assign w6919 = w6910 & w6918;
assign v2961 = ~(w6910 | w6918);
assign w6920 = v2961;
assign v2962 = ~(w6919 | w6920);
assign w6921 = v2962;
assign w6922 = w6899 & w6921;
assign v2963 = ~(w6899 | w6921);
assign w6923 = v2963;
assign v2964 = ~(w6922 | w6923);
assign w6924 = v2964;
assign w6925 = w6812 & ~w6814;
assign v2965 = ~(w6816 | w6925);
assign w6926 = v2965;
assign w6927 = w6821 & ~w6823;
assign v2966 = ~(w6825 | w6927);
assign w6928 = v2966;
assign v2967 = ~(w6926 | w6928);
assign w6929 = v2967;
assign w6930 = w6926 & w6928;
assign v2968 = ~(w6929 | w6930);
assign w6931 = v2968;
assign w6932 = w6830 & w6931;
assign v2969 = ~(w6830 | w6931);
assign w6933 = v2969;
assign v2970 = ~(w6932 | w6933);
assign w6934 = v2970;
assign w6935 = (~w6785 & w6780) | (~w6785 & w8893) | (w6780 & w8893);
assign w6936 = (~w6757 & ~w6759) | (~w6757 & w8851) | (~w6759 & w8851);
assign w6937 = (~w6751 & ~w6753) | (~w6751 & w8998) | (~w6753 & w8998);
assign w6938 = w6760 & ~w6762;
assign v2971 = ~(w6764 | w6938);
assign w6939 = v2971;
assign v2972 = ~(w6937 | w6939);
assign w6940 = v2972;
assign w6941 = w6937 & w6939;
assign v2973 = ~(w6940 | w6941);
assign w6942 = v2973;
assign w6943 = ~w6936 & w6942;
assign w6944 = w6936 & ~w6942;
assign v2974 = ~(w6943 | w6944);
assign w6945 = v2974;
assign w6946 = ~w6935 & w6945;
assign w6947 = w6935 & ~w6945;
assign v2975 = ~(w6946 | w6947);
assign w6948 = v2975;
assign w6949 = w6934 & w6948;
assign v2976 = ~(w6934 | w6948);
assign w6950 = v2976;
assign v2977 = ~(w6949 | w6950);
assign w6951 = v2977;
assign w6952 = pi25 & pi51;
assign w6953 = pi29 & pi47;
assign w6954 = pi31 & pi45;
assign w6955 = pi30 & pi46;
assign w6956 = ~w6954 & w6955;
assign w6957 = w6954 & ~w6955;
assign v2978 = ~(w6956 | w6957);
assign w6958 = v2978;
assign w6959 = w6953 & w6958;
assign v2979 = ~(w6953 | w6958);
assign w6960 = v2979;
assign v2980 = ~(w6959 | w6960);
assign w6961 = v2980;
assign w6962 = w6952 & w6961;
assign v2981 = ~(w6952 | w6961);
assign w6963 = v2981;
assign v2982 = ~(w6962 | w6963);
assign w6964 = v2982;
assign w6965 = pi26 & pi50;
assign w6966 = pi27 & pi49;
assign v2983 = ~(w6763 | w6966);
assign w6967 = v2983;
assign w6968 = pi28 & pi49;
assign w6969 = w6761 & w6968;
assign v2984 = ~(w6967 | w6969);
assign w6970 = v2984;
assign w6971 = w6965 & ~w6970;
assign w6972 = ~w6965 & w6970;
assign v2985 = ~(w6971 | w6972);
assign w6973 = v2985;
assign w6974 = w6964 & ~w6973;
assign w6975 = ~w6964 & w6973;
assign v2986 = ~(w6974 | w6975);
assign w6976 = v2986;
assign w6977 = pi13 & pi63;
assign w6978 = (w6791 & w8999) | (w6791 & w9000) | (w8999 & w9000);
assign w6979 = ~w6977 & w9307;
assign v2987 = ~(w6978 | w6979);
assign w6980 = v2987;
assign w6981 = w6976 & ~w6980;
assign w6982 = ~w6976 & w6980;
assign v2988 = ~(w6981 | w6982);
assign w6983 = v2988;
assign w6984 = w6951 & w6983;
assign v2989 = ~(w6951 | w6983);
assign w6985 = v2989;
assign v2990 = ~(w6984 | w6985);
assign w6986 = v2990;
assign w6987 = (~w6735 & w6732) | (~w6735 & w8895) | (w6732 & w8895);
assign w6988 = (~w6726 & w6723) | (~w6726 & w8852) | (w6723 & w8852);
assign w6989 = pi22 & pi54;
assign w6990 = pi23 & pi53;
assign v2991 = ~(w6824 | w6990);
assign w6991 = v2991;
assign w6992 = pi24 & pi53;
assign w6993 = w6822 & w6992;
assign v2992 = ~(w6991 | w6993);
assign w6994 = v2992;
assign w6995 = w6989 & w6994;
assign v2993 = ~(w6989 | w6994);
assign w6996 = v2993;
assign v2994 = ~(w6995 | w6996);
assign w6997 = v2994;
assign w6998 = w6815 & w6997;
assign v2995 = ~(w6815 | w6997);
assign w6999 = v2995;
assign v2996 = ~(w6998 | w6999);
assign w7000 = v2996;
assign w7001 = ~w6988 & w7000;
assign w7002 = w6988 & ~w7000;
assign v2997 = ~(w7001 | w7002);
assign w7003 = v2997;
assign w7004 = ~w6987 & w7003;
assign w7005 = w6987 & ~w7003;
assign v2998 = ~(w7004 | w7005);
assign w7006 = v2998;
assign w7007 = w6986 & w7006;
assign v2999 = ~(w6986 | w7006);
assign w7008 = v2999;
assign v3000 = ~(w7007 | w7008);
assign w7009 = v3000;
assign w7010 = w6924 & w7009;
assign v3001 = ~(w6924 | w7009);
assign w7011 = v3001;
assign v3002 = ~(w7010 | w7011);
assign w7012 = v3002;
assign w7013 = (~w6848 & w6846) | (~w6848 & w9183) | (w6846 & w9183);
assign w7014 = (~w6839 & ~w6746) | (~w6839 & w8896) | (~w6746 & w8896);
assign v3003 = ~(w6833 | w6836);
assign w7015 = v3003;
assign w7016 = (w6743 & w9184) | (w6743 & w9185) | (w9184 & w9185);
assign w7017 = ~w7015 & w9308;
assign v3004 = ~(w7016 | w7017);
assign w7018 = v3004;
assign w7019 = ~w7014 & w7018;
assign w7020 = w7014 & ~w7018;
assign v3005 = ~(w7019 | w7020);
assign w7021 = v3005;
assign w7022 = ~w7013 & w7021;
assign w7023 = w7013 & ~w7021;
assign v3006 = ~(w7022 | w7023);
assign w7024 = v3006;
assign w7025 = w7012 & w7024;
assign v3007 = ~(w7012 | w7024);
assign w7026 = v3007;
assign v3008 = ~(w7025 | w7026);
assign w7027 = v3008;
assign w7028 = ~w6874 & w7027;
assign w7029 = w6874 & ~w7027;
assign v3009 = ~(w7028 | w7029);
assign w7030 = v3009;
assign w7031 = (w7030 & w6873) | (w7030 & w8854) | (w6873 & w8854);
assign w7032 = ~w6873 & w9282;
assign v3010 = ~(w7031 | w7032);
assign w7033 = v3010;
assign w7034 = (~w6137 & w9001) | (~w6137 & w9002) | (w9001 & w9002);
assign w7035 = (~w7022 & ~w7024) | (~w7022 & w8855) | (~w7024 & w8855);
assign w7036 = pi15 & pi62;
assign w7037 = pi19 & pi58;
assign w7038 = pi21 & pi56;
assign v3011 = ~(w6879 | w7038);
assign w7039 = v3011;
assign w7040 = pi21 & pi57;
assign w7041 = w6876 & w7040;
assign v3012 = ~(w7039 | w7041);
assign w7042 = v3012;
assign w7043 = w7037 & ~w7042;
assign w7044 = ~w7037 & w7042;
assign v3013 = ~(w7043 | w7044);
assign w7045 = v3013;
assign w7046 = w7036 & ~w7045;
assign w7047 = ~w7036 & w7045;
assign v3014 = ~(w7046 | w7047);
assign w7048 = v3014;
assign w7049 = pi16 & pi61;
assign w7050 = pi18 & pi59;
assign v3015 = ~(w6891 | w7050);
assign w7051 = v3015;
assign w7052 = pi18 & pi60;
assign w7053 = w6888 & w7052;
assign v3016 = ~(w7051 | w7053);
assign w7054 = v3016;
assign w7055 = w7049 & ~w7054;
assign w7056 = ~w7049 & w7054;
assign v3017 = ~(w7055 | w7056);
assign w7057 = v3017;
assign w7058 = w7048 & ~w7057;
assign w7059 = ~w7048 & w7057;
assign v3018 = ~(w7058 | w7059);
assign w7060 = v3018;
assign w7061 = (~w6981 & ~w6951) | (~w6981 & w8899) | (~w6951 & w8899);
assign w7062 = (~w6946 & ~w6948) | (~w6946 & w8900) | (~w6948 & w8900);
assign v3019 = ~(w6978 | w7062);
assign w7063 = v3019;
assign w7064 = w6978 & w7062;
assign v3020 = ~(w7063 | w7064);
assign w7065 = v3020;
assign w7066 = ~w7061 & w7065;
assign w7067 = w7061 & ~w7065;
assign v3021 = ~(w7066 | w7067);
assign w7068 = v3021;
assign v3022 = ~(w6885 | w6897);
assign w7069 = v3022;
assign w7070 = w6714 & ~w6890;
assign v3023 = ~(w6892 | w7070);
assign w7071 = v3023;
assign w7072 = w6702 & ~w6878;
assign v3024 = ~(w6880 | w7072);
assign w7073 = v3024;
assign v3025 = ~(w7071 | w7073);
assign w7074 = v3025;
assign w7075 = w7071 & w7073;
assign v3026 = ~(w7074 | w7075);
assign w7076 = v3026;
assign w7077 = ~w7069 & w7076;
assign w7078 = w7069 & ~w7076;
assign v3027 = ~(w7077 | w7078);
assign w7079 = v3027;
assign w7080 = w7068 & w7079;
assign v3028 = ~(w7068 | w7079);
assign w7081 = v3028;
assign v3029 = ~(w7080 | w7081);
assign w7082 = v3029;
assign w7083 = w7060 & w7082;
assign v3030 = ~(w7060 | w7082);
assign w7084 = v3030;
assign v3031 = ~(w7083 | w7084);
assign w7085 = v3031;
assign v3032 = ~(w6929 | w6932);
assign w7086 = v3032;
assign w7087 = (~w6962 & ~w6964) | (~w6962 & w8856) | (~w6964 & w8856);
assign w7088 = (~w6956 & ~w6958) | (~w6956 & w9003) | (~w6958 & w9003);
assign w7089 = w6965 & ~w6967;
assign v3033 = ~(w6969 | w7089);
assign w7090 = v3033;
assign v3034 = ~(w7088 | w7090);
assign w7091 = v3034;
assign w7092 = w7088 & w7090;
assign v3035 = ~(w7091 | w7092);
assign w7093 = v3035;
assign w7094 = ~w7087 & w7093;
assign w7095 = w7087 & ~w7093;
assign v3036 = ~(w7094 | w7095);
assign w7096 = v3036;
assign w7097 = ~w7086 & w7096;
assign w7098 = w7086 & ~w7096;
assign v3037 = ~(w7097 | w7098);
assign w7099 = v3037;
assign v3038 = ~(w6993 | w6998);
assign w7100 = v3038;
assign w7101 = w6993 & w6998;
assign v3039 = ~(w7100 | w7101);
assign w7102 = v3039;
assign v3040 = ~(w6995 | w7102);
assign w7103 = v3040;
assign w7104 = w7099 & ~w7103;
assign w7105 = ~w7099 & w7103;
assign v3041 = ~(w7104 | w7105);
assign w7106 = v3041;
assign w7107 = pi25 & pi52;
assign w7108 = pi29 & pi48;
assign w7109 = pi31 & pi46;
assign w7110 = pi30 & pi47;
assign w7111 = ~w7109 & w7110;
assign w7112 = w7109 & ~w7110;
assign v3042 = ~(w7111 | w7112);
assign w7113 = v3042;
assign w7114 = w7108 & w7113;
assign v3043 = ~(w7108 | w7113);
assign w7115 = v3043;
assign v3044 = ~(w7114 | w7115);
assign w7116 = v3044;
assign w7117 = w7107 & w7116;
assign v3045 = ~(w7107 | w7116);
assign w7118 = v3045;
assign v3046 = ~(w7117 | w7118);
assign w7119 = v3046;
assign w7120 = pi26 & pi51;
assign w7121 = pi27 & pi50;
assign v3047 = ~(w6968 | w7121);
assign w7122 = v3047;
assign w7123 = pi28 & pi50;
assign w7124 = w6966 & w7123;
assign v3048 = ~(w7122 | w7124);
assign w7125 = v3048;
assign w7126 = w7120 & ~w7125;
assign w7127 = ~w7120 & w7125;
assign v3049 = ~(w7126 | w7127);
assign w7128 = v3049;
assign w7129 = w7119 & ~w7128;
assign w7130 = ~w7119 & w7128;
assign v3050 = ~(w7129 | w7130);
assign w7131 = v3050;
assign w7132 = pi14 & pi63;
assign w7133 = (w6936 & w9004) | (w6936 & w9005) | (w9004 & w9005);
assign w7134 = ~w7132 & w9309;
assign v3051 = ~(w7133 | w7134);
assign w7135 = v3051;
assign w7136 = w7131 & ~w7135;
assign w7137 = ~w7131 & w7135;
assign v3052 = ~(w7136 | w7137);
assign w7138 = v3052;
assign w7139 = w7106 & w7138;
assign v3053 = ~(w7106 | w7138);
assign w7140 = v3053;
assign v3054 = ~(w7139 | w7140);
assign w7141 = v3054;
assign v3055 = ~(w6905 | w6908);
assign w7142 = v3055;
assign w7143 = pi22 & pi55;
assign w7144 = pi23 & pi54;
assign v3056 = ~(w6992 | w7144);
assign w7145 = v3056;
assign w7146 = pi24 & pi54;
assign w7147 = w6990 & w7146;
assign v3057 = ~(w7145 | w7147);
assign w7148 = v3057;
assign w7149 = w7143 & ~w7148;
assign w7150 = ~w7143 & w7148;
assign v3058 = ~(w7149 | w7150);
assign w7151 = v3058;
assign v3059 = ~(w7142 | w7151);
assign w7152 = v3059;
assign w7153 = w7142 & w7151;
assign v3060 = ~(w7152 | w7153);
assign w7154 = v3060;
assign w7155 = (w7154 & w6916) | (w7154 & w9006) | (w6916 & w9006);
assign w7156 = ~w6916 & w9007;
assign v3061 = ~(w7155 | w7156);
assign w7157 = v3061;
assign w7158 = w7141 & w7157;
assign v3062 = ~(w7141 | w7157);
assign w7159 = v3062;
assign v3063 = ~(w7158 | w7159);
assign w7160 = v3063;
assign w7161 = w7085 & w7160;
assign v3064 = ~(w7085 | w7160);
assign w7162 = v3064;
assign v3065 = ~(w7161 | w7162);
assign w7163 = v3065;
assign w7164 = (~w7016 & w7014) | (~w7016 & w8857) | (w7014 & w8857);
assign v3066 = ~(w7007 | w7010);
assign w7165 = v3066;
assign w7166 = (~w6919 & ~w6921) | (~w6919 & w8858) | (~w6921 & w8858);
assign v3067 = ~(w7001 | w7004);
assign w7167 = v3067;
assign v3068 = ~(w7166 | w7167);
assign w7168 = v3068;
assign w7169 = w7166 & w7167;
assign v3069 = ~(w7168 | w7169);
assign w7170 = v3069;
assign w7171 = ~w7165 & w7170;
assign w7172 = w7165 & ~w7170;
assign v3070 = ~(w7171 | w7172);
assign w7173 = v3070;
assign w7174 = ~w7164 & w7173;
assign w7175 = w7164 & ~w7173;
assign v3071 = ~(w7174 | w7175);
assign w7176 = v3071;
assign w7177 = w7163 & w7176;
assign v3072 = ~(w7163 | w7176);
assign w7178 = v3072;
assign v3073 = ~(w7177 | w7178);
assign w7179 = v3073;
assign w7180 = w7035 & ~w7179;
assign w7181 = ~w7035 & w7179;
assign v3074 = ~(w7180 | w7181);
assign w7182 = v3074;
assign w7183 = w7034 & w7182;
assign v3075 = ~(w7034 | w7182);
assign w7184 = v3075;
assign v3076 = ~(w7183 | w7184);
assign w7185 = v3076;
assign w7186 = (~w7174 & ~w7176) | (~w7174 & w9008) | (~w7176 & w9008);
assign w7187 = w7143 & ~w7145;
assign v3077 = ~(w7147 | w7187);
assign w7188 = v3077;
assign w7189 = (~w7117 & ~w7119) | (~w7117 & w8859) | (~w7119 & w8859);
assign v3078 = ~(w7111 | w7114);
assign w7190 = v3078;
assign w7191 = w7120 & ~w7122;
assign v3079 = ~(w7124 | w7191);
assign w7192 = v3079;
assign v3080 = ~(w7190 | w7192);
assign w7193 = v3080;
assign w7194 = w7190 & w7192;
assign v3081 = ~(w7193 | w7194);
assign w7195 = v3081;
assign w7196 = ~w7189 & w7195;
assign w7197 = w7189 & ~w7195;
assign v3082 = ~(w7196 | w7197);
assign w7198 = v3082;
assign w7199 = w7101 & ~w7198;
assign w7200 = ~w7101 & w7198;
assign v3083 = ~(w7199 | w7200);
assign w7201 = v3083;
assign v3084 = ~(w7188 | w7201);
assign w7202 = v3084;
assign w7203 = w7188 & w7201;
assign v3085 = ~(w7202 | w7203);
assign w7204 = v3085;
assign w7205 = pi25 & pi53;
assign w7206 = pi29 & pi49;
assign w7207 = pi31 & pi47;
assign w7208 = pi30 & pi48;
assign w7209 = ~w7207 & w7208;
assign w7210 = w7207 & ~w7208;
assign v3086 = ~(w7209 | w7210);
assign w7211 = v3086;
assign w7212 = w7206 & w7211;
assign v3087 = ~(w7206 | w7211);
assign w7213 = v3087;
assign v3088 = ~(w7212 | w7213);
assign w7214 = v3088;
assign w7215 = w7205 & w7214;
assign v3089 = ~(w7205 | w7214);
assign w7216 = v3089;
assign v3090 = ~(w7215 | w7216);
assign w7217 = v3090;
assign w7218 = pi26 & pi52;
assign w7219 = pi27 & pi51;
assign v3091 = ~(w7123 | w7219);
assign w7220 = v3091;
assign w7221 = pi28 & pi51;
assign w7222 = w7121 & w7221;
assign v3092 = ~(w7220 | w7222);
assign w7223 = v3092;
assign w7224 = w7218 & ~w7223;
assign w7225 = ~w7218 & w7223;
assign v3093 = ~(w7224 | w7225);
assign w7226 = v3093;
assign w7227 = w7217 & ~w7226;
assign w7228 = ~w7217 & w7226;
assign v3094 = ~(w7227 | w7228);
assign w7229 = v3094;
assign w7230 = pi15 & pi63;
assign w7231 = (w7087 & w9009) | (w7087 & w9010) | (w9009 & w9010);
assign w7232 = ~w7230 & w9310;
assign v3095 = ~(w7231 | w7232);
assign w7233 = v3095;
assign w7234 = w7229 & ~w7233;
assign w7235 = ~w7229 & w7233;
assign v3096 = ~(w7234 | w7235);
assign w7236 = v3096;
assign w7237 = w7204 & w7236;
assign v3097 = ~(w7204 | w7236);
assign w7238 = v3097;
assign v3098 = ~(w7237 | w7238);
assign w7239 = v3098;
assign w7240 = pi23 & pi55;
assign v3099 = ~(w7146 | w7240);
assign w7241 = v3099;
assign w7242 = pi24 & pi55;
assign w7243 = w7144 & w7242;
assign v3100 = ~(w7241 | w7243);
assign w7244 = v3100;
assign v3101 = ~(w7074 | w7077);
assign w7245 = v3101;
assign w7246 = w7244 & ~w7245;
assign w7247 = ~w7244 & w7245;
assign v3102 = ~(w7246 | w7247);
assign w7248 = v3102;
assign w7249 = (w7248 & w7066) | (w7248 & w9011) | (w7066 & w9011);
assign w7250 = ~w7066 & w9012;
assign v3103 = ~(w7249 | w7250);
assign w7251 = v3103;
assign w7252 = w7239 & w7251;
assign v3104 = ~(w7239 | w7251);
assign w7253 = v3104;
assign v3105 = ~(w7252 | w7253);
assign w7254 = v3105;
assign w7255 = pi16 & pi62;
assign w7256 = pi20 & pi58;
assign w7257 = pi22 & pi56;
assign v3106 = ~(w7040 | w7257);
assign w7258 = v3106;
assign w7259 = pi22 & pi57;
assign w7260 = w7038 & w7259;
assign v3107 = ~(w7258 | w7260);
assign w7261 = v3107;
assign w7262 = w7256 & ~w7261;
assign w7263 = ~w7256 & w7261;
assign v3108 = ~(w7262 | w7263);
assign w7264 = v3108;
assign w7265 = w7255 & ~w7264;
assign w7266 = ~w7255 & w7264;
assign v3109 = ~(w7265 | w7266);
assign w7267 = v3109;
assign w7268 = pi17 & pi61;
assign w7269 = pi19 & pi59;
assign v3110 = ~(w7052 | w7269);
assign w7270 = v3110;
assign w7271 = pi19 & pi60;
assign w7272 = w7050 & w7271;
assign v3111 = ~(w7270 | w7272);
assign w7273 = v3111;
assign w7274 = w7268 & ~w7273;
assign w7275 = ~w7268 & w7273;
assign v3112 = ~(w7274 | w7275);
assign w7276 = v3112;
assign w7277 = w7267 & ~w7276;
assign w7278 = ~w7267 & w7276;
assign v3113 = ~(w7277 | w7278);
assign w7279 = v3113;
assign w7280 = (~w7136 & ~w7106) | (~w7136 & w8903) | (~w7106 & w8903);
assign w7281 = (~w7097 & ~w7099) | (~w7097 & w8904) | (~w7099 & w8904);
assign v3114 = ~(w7133 | w7281);
assign w7282 = v3114;
assign w7283 = w7133 & w7281;
assign v3115 = ~(w7282 | w7283);
assign w7284 = v3115;
assign w7285 = ~w7280 & w7284;
assign w7286 = w7280 & ~w7284;
assign v3116 = ~(w7285 | w7286);
assign w7287 = v3116;
assign v3117 = ~(w7046 | w7058);
assign w7288 = v3117;
assign w7289 = w7049 & ~w7051;
assign v3118 = ~(w7053 | w7289);
assign w7290 = v3118;
assign w7291 = w7037 & ~w7039;
assign v3119 = ~(w7041 | w7291);
assign w7292 = v3119;
assign v3120 = ~(w7290 | w7292);
assign w7293 = v3120;
assign w7294 = w7290 & w7292;
assign v3121 = ~(w7293 | w7294);
assign w7295 = v3121;
assign w7296 = ~w7288 & w7295;
assign w7297 = w7288 & ~w7295;
assign v3122 = ~(w7296 | w7297);
assign w7298 = v3122;
assign w7299 = w7287 & w7298;
assign v3123 = ~(w7287 | w7298);
assign w7300 = v3123;
assign v3124 = ~(w7299 | w7300);
assign w7301 = v3124;
assign w7302 = w7279 & w7301;
assign v3125 = ~(w7279 | w7301);
assign w7303 = v3125;
assign v3126 = ~(w7302 | w7303);
assign w7304 = v3126;
assign w7305 = w7254 & w7304;
assign v3127 = ~(w7254 | w7304);
assign w7306 = v3127;
assign v3128 = ~(w7305 | w7306);
assign w7307 = v3128;
assign w7308 = (~w7168 & w7165) | (~w7168 & w9013) | (w7165 & w9013);
assign w7309 = (~w7158 & ~w7085) | (~w7158 & w9014) | (~w7085 & w9014);
assign v3129 = ~(w7152 | w7155);
assign w7310 = v3129;
assign w7311 = (~w7080 & ~w7082) | (~w7080 & w9015) | (~w7082 & w9015);
assign v3130 = ~(w7310 | w7311);
assign w7312 = v3130;
assign w7313 = w7310 & w7311;
assign v3131 = ~(w7312 | w7313);
assign w7314 = v3131;
assign w7315 = ~w7309 & w7314;
assign w7316 = w7309 & ~w7314;
assign v3132 = ~(w7315 | w7316);
assign w7317 = v3132;
assign w7318 = ~w7308 & w7317;
assign w7319 = w7308 & ~w7317;
assign v3133 = ~(w7318 | w7319);
assign w7320 = v3133;
assign w7321 = w7307 & w7320;
assign v3134 = ~(w7307 | w7320);
assign w7322 = v3134;
assign v3135 = ~(w7321 | w7322);
assign w7323 = v3135;
assign w7324 = ~w7186 & w7323;
assign w7325 = w7186 & ~w7323;
assign v3136 = ~(w7324 | w7325);
assign w7326 = v3136;
assign w7327 = (w6137 & w9186) | (w6137 & w9187) | (w9186 & w9187);
assign w7328 = w7326 & ~w7327;
assign w7329 = ~w7326 & w7327;
assign v3137 = ~(w7328 | w7329);
assign w7330 = v3137;
assign v3138 = ~(w7318 | w7321);
assign w7331 = v3138;
assign w7332 = pi16 & pi63;
assign w7333 = pi17 & pi62;
assign w7334 = pi18 & pi61;
assign v3139 = ~(w7333 | w7334);
assign w7335 = v3139;
assign w7336 = pi18 & pi62;
assign w7337 = w7268 & w7336;
assign v3140 = ~(w7335 | w7337);
assign w7338 = v3140;
assign w7339 = w7332 & ~w7338;
assign w7340 = ~w7332 & w7338;
assign v3141 = ~(w7339 | w7340);
assign w7341 = v3141;
assign w7342 = w7243 & w7341;
assign v3142 = ~(w7243 | w7341);
assign w7343 = v3142;
assign v3143 = ~(w7342 | w7343);
assign w7344 = v3143;
assign w7345 = (~w7193 & w7189) | (~w7193 & w9059) | (w7189 & w9059);
assign w7346 = (~w7215 & ~w7217) | (~w7215 & w9016) | (~w7217 & w9016);
assign v3144 = ~(w7209 | w7212);
assign w7347 = v3144;
assign w7348 = w7218 & ~w7220;
assign v3145 = ~(w7222 | w7348);
assign w7349 = v3145;
assign v3146 = ~(w7347 | w7349);
assign w7350 = v3146;
assign w7351 = w7347 & w7349;
assign v3147 = ~(w7350 | w7351);
assign w7352 = v3147;
assign w7353 = ~w7346 & w7352;
assign w7354 = w7346 & ~w7352;
assign v3148 = ~(w7353 | w7354);
assign w7355 = v3148;
assign w7356 = w7345 & ~w7355;
assign w7357 = ~w7345 & w7355;
assign v3149 = ~(w7356 | w7357);
assign w7358 = v3149;
assign w7359 = w7344 & ~w7358;
assign w7360 = ~w7344 & w7358;
assign v3150 = ~(w7359 | w7360);
assign w7361 = v3150;
assign v3151 = ~(w7293 | w7296);
assign w7362 = v3151;
assign w7363 = pi29 & pi50;
assign w7364 = pi31 & pi48;
assign w7365 = pi30 & pi49;
assign w7366 = ~w7364 & w7365;
assign w7367 = w7364 & ~w7365;
assign v3152 = ~(w7366 | w7367);
assign w7368 = v3152;
assign w7369 = w7363 & w7368;
assign v3153 = ~(w7363 | w7368);
assign w7370 = v3153;
assign v3154 = ~(w7369 | w7370);
assign w7371 = v3154;
assign w7372 = pi26 & pi53;
assign w7373 = pi27 & pi52;
assign v3155 = ~(w7221 | w7373);
assign w7374 = v3155;
assign w7375 = pi28 & pi52;
assign w7376 = w7219 & w7375;
assign v3156 = ~(w7374 | w7376);
assign w7377 = v3156;
assign w7378 = w7372 & ~w7377;
assign w7379 = ~w7372 & w7377;
assign v3157 = ~(w7378 | w7379);
assign w7380 = v3157;
assign w7381 = w7371 & ~w7380;
assign w7382 = ~w7371 & w7380;
assign v3158 = ~(w7381 | w7382);
assign w7383 = v3158;
assign w7384 = ~w7362 & w7383;
assign w7385 = w7362 & ~w7383;
assign v3159 = ~(w7384 | w7385);
assign w7386 = v3159;
assign w7387 = (w7386 & w7285) | (w7386 & w9017) | (w7285 & w9017);
assign w7388 = ~w7285 & w9018;
assign v3160 = ~(w7387 | w7388);
assign w7389 = v3160;
assign w7390 = w7361 & w7389;
assign v3161 = ~(w7361 | w7389);
assign w7391 = v3161;
assign v3162 = ~(w7390 | w7391);
assign w7392 = v3162;
assign w7393 = pi23 & pi56;
assign w7394 = pi25 & pi54;
assign v3163 = ~(w7242 | w7394);
assign w7395 = v3163;
assign w7396 = pi25 & pi55;
assign w7397 = w7146 & w7396;
assign v3164 = ~(w7395 | w7397);
assign w7398 = v3164;
assign w7399 = w7393 & ~w7398;
assign w7400 = ~w7393 & w7398;
assign v3165 = ~(w7399 | w7400);
assign w7401 = v3165;
assign w7402 = w7271 & ~w7401;
assign w7403 = ~w7271 & w7401;
assign v3166 = ~(w7402 | w7403);
assign w7404 = v3166;
assign w7405 = pi20 & pi59;
assign w7406 = pi21 & pi58;
assign v3167 = ~(w7259 | w7406);
assign w7407 = v3167;
assign w7408 = pi22 & pi58;
assign w7409 = w7040 & w7408;
assign v3168 = ~(w7407 | w7409);
assign w7410 = v3168;
assign w7411 = w7405 & ~w7410;
assign w7412 = ~w7405 & w7410;
assign v3169 = ~(w7411 | w7412);
assign w7413 = v3169;
assign w7414 = w7404 & ~w7413;
assign w7415 = ~w7404 & w7413;
assign v3170 = ~(w7414 | w7415);
assign w7416 = v3170;
assign v3171 = ~(w7265 | w7277);
assign w7417 = v3171;
assign w7418 = w7268 & ~w7270;
assign v3172 = ~(w7272 | w7418);
assign w7419 = v3172;
assign w7420 = w7256 & ~w7258;
assign v3173 = ~(w7260 | w7420);
assign w7421 = v3173;
assign v3174 = ~(w7419 | w7421);
assign w7422 = v3174;
assign w7423 = w7419 & w7421;
assign v3175 = ~(w7422 | w7423);
assign w7424 = v3175;
assign w7425 = ~w7417 & w7424;
assign w7426 = w7417 & ~w7424;
assign v3176 = ~(w7425 | w7426);
assign w7427 = v3176;
assign w7428 = (~w7234 & ~w7204) | (~w7234 & w8905) | (~w7204 & w8905);
assign w7429 = ~w7231 & w9311;
assign w7430 = (w7201 & w9019) | (w7201 & w9020) | (w9019 & w9020);
assign v3177 = ~(w7429 | w7430);
assign w7431 = v3177;
assign w7432 = ~w7428 & w7431;
assign w7433 = w7428 & ~w7431;
assign v3178 = ~(w7432 | w7433);
assign w7434 = v3178;
assign w7435 = w7427 & w7434;
assign v3179 = ~(w7427 | w7434);
assign w7436 = v3179;
assign v3180 = ~(w7435 | w7436);
assign w7437 = v3180;
assign w7438 = w7416 & w7437;
assign v3181 = ~(w7416 | w7437);
assign w7439 = v3181;
assign v3182 = ~(w7438 | w7439);
assign w7440 = v3182;
assign w7441 = w7392 & w7440;
assign v3183 = ~(w7392 | w7440);
assign w7442 = v3183;
assign v3184 = ~(w7441 | w7442);
assign w7443 = v3184;
assign v3185 = ~(w7312 | w7315);
assign w7444 = v3185;
assign w7445 = (~w7252 & ~w7304) | (~w7252 & w9021) | (~w7304 & w9021);
assign v3186 = ~(w7246 | w7249);
assign w7446 = v3186;
assign w7447 = (~w7299 & ~w7301) | (~w7299 & w9022) | (~w7301 & w9022);
assign v3187 = ~(w7446 | w7447);
assign w7448 = v3187;
assign w7449 = w7446 & w7447;
assign v3188 = ~(w7448 | w7449);
assign w7450 = v3188;
assign w7451 = ~w7445 & w7450;
assign w7452 = w7445 & ~w7450;
assign v3189 = ~(w7451 | w7452);
assign w7453 = v3189;
assign w7454 = ~w7444 & w7453;
assign w7455 = w7444 & ~w7453;
assign v3190 = ~(w7454 | w7455);
assign w7456 = v3190;
assign w7457 = w7443 & w7456;
assign v3191 = ~(w7443 | w7456);
assign w7458 = v3191;
assign v3192 = ~(w7457 | w7458);
assign w7459 = v3192;
assign w7460 = ~w7331 & w7459;
assign w7461 = w7331 & ~w7459;
assign v3193 = ~(w7460 | w7461);
assign w7462 = v3193;
assign w7463 = w7030 & w7182;
assign w7464 = ~w7325 & w7463;
assign w7465 = w7028 & ~w7180;
assign v3194 = ~(w7181 | w7324);
assign w7466 = v3194;
assign w7467 = ~w7465 & w7466;
assign v3195 = ~(w7325 | w7467);
assign w7468 = v3195;
assign w7469 = (~w7468 & w6870) | (~w7468 & w8907) | (w6870 & w8907);
assign w7470 = w6132 & w7469;
assign w7471 = ~w6137 & w7470;
assign w7472 = w7326 & w7463;
assign w7473 = w6872 & w7472;
assign w7474 = w7469 & ~w7473;
assign w7475 = ~w7474 & w9312;
assign w7476 = w7462 & w9313;
assign v3196 = ~(w7475 | w7476);
assign w7477 = v3196;
assign w7478 = (~w7454 & ~w7456) | (~w7454 & w9060) | (~w7456 & w9060);
assign w7479 = pi21 & pi59;
assign w7480 = pi27 & pi53;
assign w7481 = pi26 & pi54;
assign v3197 = ~(w7480 | w7481);
assign w7482 = v3197;
assign w7483 = pi27 & pi54;
assign w7484 = w7372 & w7483;
assign v3198 = ~(w7482 | w7484);
assign w7485 = v3198;
assign w7486 = w7396 & ~w7485;
assign w7487 = ~w7396 & w7485;
assign v3199 = ~(w7486 | w7487);
assign w7488 = v3199;
assign w7489 = w7479 & ~w7488;
assign w7490 = ~w7479 & w7488;
assign v3200 = ~(w7489 | w7490);
assign w7491 = v3200;
assign w7492 = pi24 & pi56;
assign w7493 = pi23 & pi57;
assign v3201 = ~(w7492 | w7493);
assign w7494 = v3201;
assign w7495 = pi24 & pi57;
assign w7496 = w7393 & w7495;
assign v3202 = ~(w7494 | w7496);
assign w7497 = v3202;
assign w7498 = w7408 & ~w7497;
assign w7499 = ~w7408 & w7497;
assign v3203 = ~(w7498 | w7499);
assign w7500 = v3203;
assign w7501 = w7491 & ~w7500;
assign w7502 = ~w7491 & w7500;
assign v3204 = ~(w7501 | w7502);
assign w7503 = v3204;
assign v3205 = ~(w7402 | w7414);
assign w7504 = v3205;
assign w7505 = w7405 & ~w7407;
assign v3206 = ~(w7409 | w7505);
assign w7506 = v3206;
assign w7507 = w7393 & ~w7395;
assign v3207 = ~(w7397 | w7507);
assign w7508 = v3207;
assign v3208 = ~(w7506 | w7508);
assign w7509 = v3208;
assign w7510 = w7506 & w7508;
assign v3209 = ~(w7509 | w7510);
assign w7511 = v3209;
assign w7512 = ~w7504 & w7511;
assign w7513 = w7504 & ~w7511;
assign v3210 = ~(w7512 | w7513);
assign w7514 = v3210;
assign w7515 = (~w7342 & w7358) | (~w7342 & w9061) | (w7358 & w9061);
assign v3211 = ~(w7337 | w7340);
assign w7516 = v3211;
assign v3212 = ~(w7356 | w7516);
assign w7517 = v3212;
assign w7518 = w7356 & w7516;
assign v3213 = ~(w7517 | w7518);
assign w7519 = v3213;
assign w7520 = ~w7515 & w7519;
assign w7521 = w7515 & ~w7519;
assign v3214 = ~(w7520 | w7521);
assign w7522 = v3214;
assign w7523 = w7514 & w7522;
assign v3215 = ~(w7514 | w7522);
assign w7524 = v3215;
assign v3216 = ~(w7523 | w7524);
assign w7525 = v3216;
assign w7526 = w7503 & w7525;
assign v3217 = ~(w7503 | w7525);
assign w7527 = v3217;
assign v3218 = ~(w7526 | w7527);
assign w7528 = v3218;
assign v3219 = ~(w7366 | w7369);
assign w7529 = v3219;
assign w7530 = w7372 & ~w7374;
assign v3220 = ~(w7376 | w7530);
assign w7531 = v3220;
assign v3221 = ~(w7529 | w7531);
assign w7532 = v3221;
assign w7533 = w7529 & w7531;
assign v3222 = ~(w7532 | w7533);
assign w7534 = v3222;
assign w7535 = w7381 & w7534;
assign v3223 = ~(w7381 | w7534);
assign w7536 = v3223;
assign v3224 = ~(w7535 | w7536);
assign w7537 = v3224;
assign w7538 = pi20 & pi60;
assign w7539 = pi19 & pi61;
assign v3225 = ~(w7538 | w7539);
assign w7540 = v3225;
assign w7541 = pi20 & pi61;
assign w7542 = w7271 & w7541;
assign v3226 = ~(w7540 | w7542);
assign w7543 = v3226;
assign w7544 = w7336 & ~w7543;
assign w7545 = ~w7336 & w7543;
assign v3227 = ~(w7544 | w7545);
assign w7546 = v3227;
assign w7547 = w7537 & ~w7546;
assign w7548 = ~w7537 & w7546;
assign v3228 = ~(w7547 | w7548);
assign w7549 = v3228;
assign w7550 = pi17 & pi63;
assign w7551 = (~w7350 & w7346) | (~w7350 & w9062) | (w7346 & w9062);
assign w7552 = w7550 & w7551;
assign v3229 = ~(w7550 | w7551);
assign w7553 = v3229;
assign v3230 = ~(w7552 | w7553);
assign w7554 = v3230;
assign w7555 = w7549 & ~w7554;
assign w7556 = ~w7549 & w7554;
assign v3231 = ~(w7555 | w7556);
assign w7557 = v3231;
assign w7558 = (~w7429 & w7428) | (~w7429 & w9023) | (w7428 & w9023);
assign v3232 = ~(w7422 | w7425);
assign w7559 = v3232;
assign w7560 = pi29 & pi51;
assign w7561 = pi31 & pi49;
assign w7562 = pi30 & pi50;
assign w7563 = ~w7561 & w7562;
assign w7564 = w7561 & ~w7562;
assign v3233 = ~(w7563 | w7564);
assign w7565 = v3233;
assign w7566 = w7560 & w7565;
assign v3234 = ~(w7560 | w7565);
assign w7567 = v3234;
assign v3235 = ~(w7566 | w7567);
assign w7568 = v3235;
assign w7569 = w7375 & w7568;
assign v3236 = ~(w7375 | w7568);
assign w7570 = v3236;
assign v3237 = ~(w7569 | w7570);
assign w7571 = v3237;
assign w7572 = ~w7559 & w7571;
assign w7573 = w7559 & ~w7571;
assign v3238 = ~(w7572 | w7573);
assign w7574 = v3238;
assign w7575 = ~w7558 & w7574;
assign w7576 = w7558 & ~w7574;
assign v3239 = ~(w7575 | w7576);
assign w7577 = v3239;
assign w7578 = w7557 & w7577;
assign v3240 = ~(w7557 | w7577);
assign w7579 = v3240;
assign v3241 = ~(w7578 | w7579);
assign w7580 = v3241;
assign w7581 = w7528 & w7580;
assign v3242 = ~(w7528 | w7580);
assign w7582 = v3242;
assign v3243 = ~(w7581 | w7582);
assign w7583 = v3243;
assign v3244 = ~(w7448 | w7451);
assign w7584 = v3244;
assign w7585 = (~w7390 & ~w7440) | (~w7390 & w9024) | (~w7440 & w9024);
assign v3245 = ~(w7384 | w7387);
assign w7586 = v3245;
assign w7587 = (~w7435 & ~w7437) | (~w7435 & w9025) | (~w7437 & w9025);
assign v3246 = ~(w7586 | w7587);
assign w7588 = v3246;
assign w7589 = w7586 & w7587;
assign v3247 = ~(w7588 | w7589);
assign w7590 = v3247;
assign w7591 = ~w7585 & w7590;
assign w7592 = w7585 & ~w7590;
assign v3248 = ~(w7591 | w7592);
assign w7593 = v3248;
assign w7594 = ~w7584 & w7593;
assign w7595 = w7584 & ~w7593;
assign v3249 = ~(w7594 | w7595);
assign w7596 = v3249;
assign w7597 = w7583 & w7596;
assign v3250 = ~(w7583 | w7596);
assign w7598 = v3250;
assign v3251 = ~(w7597 | w7598);
assign w7599 = v3251;
assign w7600 = ~w7478 & w7599;
assign w7601 = w7478 & ~w7599;
assign v3252 = ~(w7600 | w7601);
assign w7602 = v3252;
assign w7603 = (w9064 & w9284) | (w9064 & w9285) | (w9284 & w9285);
assign w7604 = ~w7461 & w7602;
assign w7605 = (w6137 & w9190) | (w6137 & w9191) | (w9190 & w9191);
assign v3253 = ~(w7603 | w7605);
assign w7606 = v3253;
assign w7607 = (~w7594 & ~w7596) | (~w7594 & w9067) | (~w7596 & w9067);
assign w7608 = pi22 & pi59;
assign w7609 = pi26 & pi55;
assign w7610 = pi28 & pi53;
assign v3254 = ~(w7483 | w7610);
assign w7611 = v3254;
assign w7612 = pi28 & pi54;
assign w7613 = w7480 & w7612;
assign v3255 = ~(w7611 | w7613);
assign w7614 = v3255;
assign w7615 = w7609 & ~w7614;
assign w7616 = ~w7609 & w7614;
assign v3256 = ~(w7615 | w7616);
assign w7617 = v3256;
assign w7618 = w7608 & ~w7617;
assign w7619 = ~w7608 & w7617;
assign v3257 = ~(w7618 | w7619);
assign w7620 = v3257;
assign w7621 = pi23 & pi58;
assign w7622 = pi25 & pi56;
assign v3258 = ~(w7495 | w7622);
assign w7623 = v3258;
assign w7624 = pi25 & pi57;
assign w7625 = w7492 & w7624;
assign v3259 = ~(w7623 | w7625);
assign w7626 = v3259;
assign w7627 = w7621 & ~w7626;
assign w7628 = ~w7621 & w7626;
assign v3260 = ~(w7627 | w7628);
assign w7629 = v3260;
assign w7630 = w7620 & ~w7629;
assign w7631 = ~w7620 & w7629;
assign v3261 = ~(w7630 | w7631);
assign w7632 = v3261;
assign v3262 = ~(w7489 | w7501);
assign w7633 = v3262;
assign w7634 = w7408 & ~w7494;
assign v3263 = ~(w7496 | w7634);
assign w7635 = v3263;
assign w7636 = w7396 & ~w7482;
assign v3264 = ~(w7484 | w7636);
assign w7637 = v3264;
assign v3265 = ~(w7635 | w7637);
assign w7638 = v3265;
assign w7639 = w7635 & w7637;
assign v3266 = ~(w7638 | w7639);
assign w7640 = v3266;
assign w7641 = ~w7633 & w7640;
assign w7642 = w7633 & ~w7640;
assign v3267 = ~(w7641 | w7642);
assign w7643 = v3267;
assign v3268 = ~(w7547 | w7555);
assign w7644 = v3268;
assign w7645 = w7336 & ~w7540;
assign v3269 = ~(w7542 | w7645);
assign w7646 = v3269;
assign v3270 = ~(w7552 | w7646);
assign w7647 = v3270;
assign w7648 = w7552 & w7646;
assign v3271 = ~(w7647 | w7648);
assign w7649 = v3271;
assign w7650 = ~w7644 & w7649;
assign w7651 = w7644 & ~w7649;
assign v3272 = ~(w7650 | w7651);
assign w7652 = v3272;
assign w7653 = w7643 & w7652;
assign v3273 = ~(w7643 | w7652);
assign w7654 = v3273;
assign v3274 = ~(w7653 | w7654);
assign w7655 = v3274;
assign w7656 = w7632 & w7655;
assign v3275 = ~(w7632 | w7655);
assign w7657 = v3275;
assign v3276 = ~(w7656 | w7657);
assign w7658 = v3276;
assign w7659 = w7563 & w7569;
assign v3277 = ~(w7563 | w7569);
assign w7660 = v3277;
assign v3278 = ~(w7659 | w7660);
assign w7661 = v3278;
assign v3279 = ~(w7566 | w7661);
assign w7662 = v3279;
assign w7663 = pi19 & pi62;
assign w7664 = pi21 & pi60;
assign v3280 = ~(w7541 | w7664);
assign w7665 = v3280;
assign w7666 = pi21 & pi61;
assign w7667 = w7538 & w7666;
assign v3281 = ~(w7665 | w7667);
assign w7668 = v3281;
assign w7669 = w7663 & ~w7668;
assign w7670 = ~w7663 & w7668;
assign v3282 = ~(w7669 | w7670);
assign w7671 = v3282;
assign v3283 = ~(w7662 | w7671);
assign w7672 = v3283;
assign w7673 = w7662 & w7671;
assign v3284 = ~(w7672 | w7673);
assign w7674 = v3284;
assign w7675 = pi18 & pi63;
assign v3285 = ~(w7532 | w7535);
assign w7676 = v3285;
assign w7677 = w7675 & w7676;
assign v3286 = ~(w7675 | w7676);
assign w7678 = v3286;
assign v3287 = ~(w7677 | w7678);
assign w7679 = v3287;
assign w7680 = w7674 & ~w7679;
assign w7681 = ~w7674 & w7679;
assign v3288 = ~(w7680 | w7681);
assign w7682 = v3288;
assign v3289 = ~(w7517 | w7520);
assign w7683 = v3289;
assign v3290 = ~(w7509 | w7512);
assign w7684 = v3290;
assign w7685 = pi29 & pi52;
assign w7686 = pi31 & pi50;
assign w7687 = pi30 & pi51;
assign w7688 = ~w7686 & w7687;
assign w7689 = w7686 & ~w7687;
assign v3291 = ~(w7688 | w7689);
assign w7690 = v3291;
assign w7691 = w7685 & w7690;
assign v3292 = ~(w7685 | w7690);
assign w7692 = v3292;
assign v3293 = ~(w7691 | w7692);
assign w7693 = v3293;
assign w7694 = ~w7684 & w7693;
assign w7695 = w7684 & ~w7693;
assign v3294 = ~(w7694 | w7695);
assign w7696 = v3294;
assign w7697 = ~w7683 & w7696;
assign w7698 = w7683 & ~w7696;
assign v3295 = ~(w7697 | w7698);
assign w7699 = v3295;
assign w7700 = w7682 & w7699;
assign v3296 = ~(w7682 | w7699);
assign w7701 = v3296;
assign v3297 = ~(w7700 | w7701);
assign w7702 = v3297;
assign w7703 = w7658 & w7702;
assign v3298 = ~(w7658 | w7702);
assign w7704 = v3298;
assign v3299 = ~(w7703 | w7704);
assign w7705 = v3299;
assign v3300 = ~(w7588 | w7591);
assign w7706 = v3300;
assign w7707 = (~w7578 & ~w7580) | (~w7578 & w9068) | (~w7580 & w9068);
assign v3301 = ~(w7523 | w7526);
assign w7708 = v3301;
assign v3302 = ~(w7572 | w7575);
assign w7709 = v3302;
assign v3303 = ~(w7708 | w7709);
assign w7710 = v3303;
assign w7711 = w7708 & w7709;
assign v3304 = ~(w7710 | w7711);
assign w7712 = v3304;
assign w7713 = ~w7707 & w7712;
assign w7714 = w7707 & ~w7712;
assign v3305 = ~(w7713 | w7714);
assign w7715 = v3305;
assign w7716 = ~w7706 & w7715;
assign w7717 = w7706 & ~w7715;
assign v3306 = ~(w7716 | w7717);
assign w7718 = v3306;
assign w7719 = w7705 & w7718;
assign v3307 = ~(w7705 | w7718);
assign w7720 = v3307;
assign v3308 = ~(w7719 | w7720);
assign w7721 = v3308;
assign w7722 = w7607 & ~w7721;
assign w7723 = ~w7607 & w7721;
assign v3309 = ~(w7722 | w7723);
assign w7724 = v3309;
assign w7725 = w8779 & ~w7605;
assign w7726 = ~w7724 & w9314;
assign v3310 = ~(w7725 | w7726);
assign w7727 = v3310;
assign w7728 = (~w7716 & ~w7718) | (~w7716 & w9069) | (~w7718 & w9069);
assign w7729 = pi23 & pi59;
assign w7730 = pi27 & pi55;
assign w7731 = pi29 & pi53;
assign v3311 = ~(w7612 | w7731);
assign w7732 = v3311;
assign w7733 = pi29 & pi54;
assign w7734 = w7610 & w7733;
assign v3312 = ~(w7732 | w7734);
assign w7735 = v3312;
assign w7736 = w7730 & ~w7735;
assign w7737 = ~w7730 & w7735;
assign v3313 = ~(w7736 | w7737);
assign w7738 = v3313;
assign w7739 = w7729 & ~w7738;
assign w7740 = ~w7729 & w7738;
assign v3314 = ~(w7739 | w7740);
assign w7741 = v3314;
assign w7742 = pi24 & pi58;
assign w7743 = pi26 & pi56;
assign v3315 = ~(w7624 | w7743);
assign w7744 = v3315;
assign w7745 = pi26 & pi57;
assign w7746 = w7622 & w7745;
assign v3316 = ~(w7744 | w7746);
assign w7747 = v3316;
assign w7748 = w7742 & ~w7747;
assign w7749 = ~w7742 & w7747;
assign v3317 = ~(w7748 | w7749);
assign w7750 = v3317;
assign w7751 = w7741 & ~w7750;
assign w7752 = ~w7741 & w7750;
assign v3318 = ~(w7751 | w7752);
assign w7753 = v3318;
assign v3319 = ~(w7618 | w7630);
assign w7754 = v3319;
assign w7755 = w7621 & ~w7623;
assign v3320 = ~(w7625 | w7755);
assign w7756 = v3320;
assign w7757 = w7609 & ~w7611;
assign v3321 = ~(w7613 | w7757);
assign w7758 = v3321;
assign v3322 = ~(w7756 | w7758);
assign w7759 = v3322;
assign w7760 = w7756 & w7758;
assign v3323 = ~(w7759 | w7760);
assign w7761 = v3323;
assign w7762 = ~w7754 & w7761;
assign w7763 = w7754 & ~w7761;
assign v3324 = ~(w7762 | w7763);
assign w7764 = v3324;
assign v3325 = ~(w7672 | w7680);
assign w7765 = v3325;
assign w7766 = w7663 & ~w7665;
assign v3326 = ~(w7667 | w7766);
assign w7767 = v3326;
assign v3327 = ~(w7677 | w7767);
assign w7768 = v3327;
assign w7769 = w7677 & w7767;
assign v3328 = ~(w7768 | w7769);
assign w7770 = v3328;
assign w7771 = ~w7765 & w7770;
assign w7772 = w7765 & ~w7770;
assign v3329 = ~(w7771 | w7772);
assign w7773 = v3329;
assign w7774 = w7764 & w7773;
assign v3330 = ~(w7764 | w7773);
assign w7775 = v3330;
assign v3331 = ~(w7774 | w7775);
assign w7776 = v3331;
assign w7777 = w7753 & w7776;
assign v3332 = ~(w7753 | w7776);
assign w7778 = v3332;
assign v3333 = ~(w7777 | w7778);
assign w7779 = v3333;
assign w7780 = pi19 & pi63;
assign w7781 = ~w7659 & w7780;
assign w7782 = w7659 & ~w7780;
assign v3334 = ~(w7781 | w7782);
assign w7783 = v3334;
assign v3335 = ~(w7688 | w7691);
assign w7784 = v3335;
assign w7785 = pi20 & pi62;
assign w7786 = pi22 & pi60;
assign v3336 = ~(w7666 | w7786);
assign w7787 = v3336;
assign w7788 = pi22 & pi61;
assign w7789 = w7664 & w7788;
assign v3337 = ~(w7787 | w7789);
assign w7790 = v3337;
assign w7791 = w7785 & ~w7790;
assign w7792 = ~w7785 & w7790;
assign v3338 = ~(w7791 | w7792);
assign w7793 = v3338;
assign v3339 = ~(w7784 | w7793);
assign w7794 = v3339;
assign w7795 = w7784 & w7793;
assign v3340 = ~(w7794 | w7795);
assign w7796 = v3340;
assign w7797 = ~w7783 & w7796;
assign w7798 = w7783 & ~w7796;
assign v3341 = ~(w7797 | w7798);
assign w7799 = v3341;
assign v3342 = ~(w7647 | w7650);
assign w7800 = v3342;
assign v3343 = ~(w7638 | w7641);
assign w7801 = v3343;
assign w7802 = pi31 & pi51;
assign w7803 = pi30 & pi52;
assign w7804 = ~w7802 & w7803;
assign w7805 = w7802 & ~w7803;
assign v3344 = ~(w7804 | w7805);
assign w7806 = v3344;
assign w7807 = ~w7801 & w7806;
assign w7808 = w7801 & ~w7806;
assign v3345 = ~(w7807 | w7808);
assign w7809 = v3345;
assign w7810 = ~w7800 & w7809;
assign w7811 = w7800 & ~w7809;
assign v3346 = ~(w7810 | w7811);
assign w7812 = v3346;
assign w7813 = w7799 & w7812;
assign v3347 = ~(w7799 | w7812);
assign w7814 = v3347;
assign v3348 = ~(w7813 | w7814);
assign w7815 = v3348;
assign w7816 = w7779 & w7815;
assign v3349 = ~(w7779 | w7815);
assign w7817 = v3349;
assign v3350 = ~(w7816 | w7817);
assign w7818 = v3350;
assign v3351 = ~(w7710 | w7713);
assign w7819 = v3351;
assign v3352 = ~(w7700 | w7703);
assign w7820 = v3352;
assign v3353 = ~(w7653 | w7656);
assign w7821 = v3353;
assign v3354 = ~(w7694 | w7697);
assign w7822 = v3354;
assign v3355 = ~(w7821 | w7822);
assign w7823 = v3355;
assign w7824 = w7821 & w7822;
assign v3356 = ~(w7823 | w7824);
assign w7825 = v3356;
assign w7826 = ~w7820 & w7825;
assign w7827 = w7820 & ~w7825;
assign v3357 = ~(w7826 | w7827);
assign w7828 = v3357;
assign w7829 = ~w7819 & w7828;
assign w7830 = w7819 & ~w7828;
assign v3358 = ~(w7829 | w7830);
assign w7831 = v3358;
assign w7832 = w7818 & w7831;
assign v3359 = ~(w7818 | w7831);
assign w7833 = v3359;
assign v3360 = ~(w7832 | w7833);
assign w7834 = v3360;
assign w7835 = ~w7728 & w7834;
assign w7836 = w7728 & ~w7834;
assign v3361 = ~(w7835 | w7836);
assign w7837 = v3361;
assign w7838 = w7837 & w9315;
assign w7839 = (w7471 & w9192) | (w7471 & w9193) | (w9192 & w9193);
assign v3362 = ~(w7838 | w7839);
assign w7840 = v3362;
assign v3363 = ~(w7829 | w7832);
assign w7841 = v3363;
assign w7842 = pi25 & pi58;
assign w7843 = pi31 & pi52;
assign w7844 = pi30 & pi53;
assign w7845 = ~w7843 & w7844;
assign w7846 = w7843 & ~w7844;
assign v3364 = ~(w7845 | w7846);
assign w7847 = v3364;
assign w7848 = w7733 & w7847;
assign v3365 = ~(w7733 | w7847);
assign w7849 = v3365;
assign v3366 = ~(w7848 | w7849);
assign w7850 = v3366;
assign w7851 = w7842 & w7850;
assign v3367 = ~(w7842 | w7850);
assign w7852 = v3367;
assign v3368 = ~(w7851 | w7852);
assign w7853 = v3368;
assign w7854 = pi27 & pi56;
assign w7855 = pi28 & pi55;
assign v3369 = ~(w7854 | w7855);
assign w7856 = v3369;
assign w7857 = pi28 & pi56;
assign w7858 = w7730 & w7857;
assign v3370 = ~(w7856 | w7858);
assign w7859 = v3370;
assign w7860 = w7745 & ~w7859;
assign w7861 = ~w7745 & w7859;
assign v3371 = ~(w7860 | w7861);
assign w7862 = v3371;
assign w7863 = w7853 & ~w7862;
assign w7864 = ~w7853 & w7862;
assign v3372 = ~(w7863 | w7864);
assign w7865 = v3372;
assign v3373 = ~(w7794 | w7797);
assign w7866 = v3373;
assign w7867 = w7785 & ~w7787;
assign v3374 = ~(w7789 | w7867);
assign w7868 = v3374;
assign v3375 = ~(w7781 | w7868);
assign w7869 = v3375;
assign w7870 = w7781 & w7868;
assign v3376 = ~(w7869 | w7870);
assign w7871 = v3376;
assign w7872 = ~w7866 & w7871;
assign w7873 = w7866 & ~w7871;
assign v3377 = ~(w7872 | w7873);
assign w7874 = v3377;
assign v3378 = ~(w7739 | w7751);
assign w7875 = v3378;
assign w7876 = w7742 & ~w7744;
assign v3379 = ~(w7746 | w7876);
assign w7877 = v3379;
assign w7878 = w7730 & ~w7732;
assign v3380 = ~(w7734 | w7878);
assign w7879 = v3380;
assign v3381 = ~(w7877 | w7879);
assign w7880 = v3381;
assign w7881 = w7877 & w7879;
assign v3382 = ~(w7880 | w7881);
assign w7882 = v3382;
assign w7883 = ~w7875 & w7882;
assign w7884 = w7875 & ~w7882;
assign v3383 = ~(w7883 | w7884);
assign w7885 = v3383;
assign w7886 = w7874 & w7885;
assign v3384 = ~(w7874 | w7885);
assign w7887 = v3384;
assign v3385 = ~(w7886 | w7887);
assign w7888 = v3385;
assign w7889 = w7865 & w7888;
assign v3386 = ~(w7865 | w7888);
assign w7890 = v3386;
assign v3387 = ~(w7889 | w7890);
assign w7891 = v3387;
assign w7892 = pi20 & pi63;
assign w7893 = pi21 & pi62;
assign w7894 = w7892 & ~w7893;
assign w7895 = ~w7892 & w7893;
assign v3388 = ~(w7894 | w7895);
assign w7896 = v3388;
assign w7897 = pi23 & pi60;
assign w7898 = pi24 & pi59;
assign v3389 = ~(w7897 | w7898);
assign w7899 = v3389;
assign w7900 = pi24 & pi60;
assign w7901 = w7729 & w7900;
assign v3390 = ~(w7899 | w7901);
assign w7902 = v3390;
assign w7903 = w7788 & ~w7902;
assign w7904 = ~w7788 & w7902;
assign v3391 = ~(w7903 | w7904);
assign w7905 = v3391;
assign v3392 = ~(w7896 | w7905);
assign w7906 = v3392;
assign w7907 = w7896 & w7905;
assign v3393 = ~(w7906 | w7907);
assign w7908 = v3393;
assign v3394 = ~(w7768 | w7771);
assign w7909 = v3394;
assign v3395 = ~(w7759 | w7762);
assign w7910 = v3395;
assign w7911 = w7804 & ~w7910;
assign w7912 = ~w7804 & w7910;
assign v3396 = ~(w7911 | w7912);
assign w7913 = v3396;
assign w7914 = ~w7909 & w7913;
assign w7915 = w7909 & ~w7913;
assign v3397 = ~(w7914 | w7915);
assign w7916 = v3397;
assign w7917 = w7908 & w7916;
assign v3398 = ~(w7908 | w7916);
assign w7918 = v3398;
assign v3399 = ~(w7917 | w7918);
assign w7919 = v3399;
assign w7920 = w7891 & w7919;
assign v3400 = ~(w7891 | w7919);
assign w7921 = v3400;
assign v3401 = ~(w7920 | w7921);
assign w7922 = v3401;
assign v3402 = ~(w7823 | w7826);
assign w7923 = v3402;
assign v3403 = ~(w7813 | w7816);
assign w7924 = v3403;
assign v3404 = ~(w7774 | w7777);
assign w7925 = v3404;
assign v3405 = ~(w7807 | w7810);
assign w7926 = v3405;
assign v3406 = ~(w7925 | w7926);
assign w7927 = v3406;
assign w7928 = w7925 & w7926;
assign v3407 = ~(w7927 | w7928);
assign w7929 = v3407;
assign w7930 = ~w7924 & w7929;
assign w7931 = w7924 & ~w7929;
assign v3408 = ~(w7930 | w7931);
assign w7932 = v3408;
assign w7933 = ~w7923 & w7932;
assign w7934 = w7923 & ~w7932;
assign v3409 = ~(w7933 | w7934);
assign w7935 = v3409;
assign w7936 = w7922 & w7935;
assign v3410 = ~(w7922 | w7935);
assign w7937 = v3410;
assign v3411 = ~(w7936 | w7937);
assign w7938 = v3411;
assign w7939 = ~w7841 & w7938;
assign w7940 = w7841 & ~w7938;
assign v3412 = ~(w7939 | w7940);
assign w7941 = v3412;
assign w7942 = (w7471 & w9194) | (w7471 & w9195) | (w9194 & w9195);
assign w7943 = (w9072 & w9073) | (w9072 & w9315) | (w9073 & w9315);
assign v3413 = ~(w7942 | w7943);
assign w7944 = v3413;
assign v3414 = ~(w7600 | w7723);
assign w7945 = v3414;
assign v3415 = ~(w7722 | w7836);
assign w7946 = v3415;
assign w7947 = ~w7945 & w7946;
assign v3416 = ~(w7835 | w7939);
assign w7948 = v3416;
assign w7949 = (~w7940 & w7947) | (~w7940 & w9074) | (w7947 & w9074);
assign w7950 = w7724 & w7837;
assign w7951 = w7941 & w7950;
assign w7952 = w7604 & w7951;
assign w7953 = (w6137 & w9196) | (w6137 & w9197) | (w9196 & w9197);
assign v3417 = ~(w7933 | w7936);
assign w7954 = v3417;
assign w7955 = pi25 & pi59;
assign w7956 = pi29 & pi55;
assign w7957 = pi31 & pi53;
assign w7958 = pi30 & pi54;
assign w7959 = ~w7957 & w7958;
assign w7960 = w7957 & ~w7958;
assign v3418 = ~(w7959 | w7960);
assign w7961 = v3418;
assign w7962 = w7956 & w7961;
assign v3419 = ~(w7956 | w7961);
assign w7963 = v3419;
assign v3420 = ~(w7962 | w7963);
assign w7964 = v3420;
assign w7965 = w7955 & w7964;
assign v3421 = ~(w7955 | w7964);
assign w7966 = v3421;
assign v3422 = ~(w7965 | w7966);
assign w7967 = v3422;
assign w7968 = pi26 & pi58;
assign w7969 = pi27 & pi57;
assign v3423 = ~(w7857 | w7969);
assign w7970 = v3423;
assign w7971 = pi28 & pi57;
assign w7972 = w7854 & w7971;
assign v3424 = ~(w7970 | w7972);
assign w7973 = v3424;
assign w7974 = w7968 & ~w7973;
assign w7975 = ~w7968 & w7973;
assign v3425 = ~(w7974 | w7975);
assign w7976 = v3425;
assign w7977 = w7967 & ~w7976;
assign w7978 = ~w7967 & w7976;
assign v3426 = ~(w7977 | w7978);
assign w7979 = v3426;
assign w7980 = w7788 & ~w7899;
assign v3427 = ~(w7901 | w7980);
assign w7981 = v3427;
assign v3428 = ~(w7894 | w7981);
assign w7982 = v3428;
assign w7983 = w7894 & w7981;
assign v3429 = ~(w7982 | w7983);
assign w7984 = v3429;
assign w7985 = w7906 & w7984;
assign v3430 = ~(w7906 | w7984);
assign w7986 = v3430;
assign v3431 = ~(w7985 | w7986);
assign w7987 = v3431;
assign v3432 = ~(w7851 | w7863);
assign w7988 = v3432;
assign v3433 = ~(w7845 | w7848);
assign w7989 = v3433;
assign w7990 = w7745 & ~w7856;
assign v3434 = ~(w7858 | w7990);
assign w7991 = v3434;
assign v3435 = ~(w7989 | w7991);
assign w7992 = v3435;
assign w7993 = w7989 & w7991;
assign v3436 = ~(w7992 | w7993);
assign w7994 = v3436;
assign w7995 = ~w7988 & w7994;
assign w7996 = w7988 & ~w7994;
assign v3437 = ~(w7995 | w7996);
assign w7997 = v3437;
assign w7998 = w7987 & w7997;
assign v3438 = ~(w7987 | w7997);
assign w7999 = v3438;
assign v3439 = ~(w7998 | w7999);
assign w8000 = v3439;
assign w8001 = w7979 & w8000;
assign v3440 = ~(w7979 | w8000);
assign w8002 = v3440;
assign v3441 = ~(w8001 | w8002);
assign w8003 = v3441;
assign w8004 = pi21 & pi63;
assign w8005 = pi22 & pi62;
assign w8006 = pi23 & pi61;
assign v3442 = ~(w7900 | w8006);
assign w8007 = v3442;
assign w8008 = pi24 & pi61;
assign w8009 = w7897 & w8008;
assign v3443 = ~(w8007 | w8009);
assign w8010 = v3443;
assign w8011 = w8005 & w8010;
assign v3444 = ~(w8005 | w8010);
assign w8012 = v3444;
assign v3445 = ~(w8011 | w8012);
assign w8013 = v3445;
assign w8014 = w8004 & ~w8013;
assign w8015 = ~w8004 & w8013;
assign v3446 = ~(w8014 | w8015);
assign w8016 = v3446;
assign v3447 = ~(w7869 | w7872);
assign w8017 = v3447;
assign v3448 = ~(w7880 | w7883);
assign w8018 = v3448;
assign w8019 = w8017 & w8018;
assign v3449 = ~(w8017 | w8018);
assign w8020 = v3449;
assign v3450 = ~(w8019 | w8020);
assign w8021 = v3450;
assign w8022 = w8016 & ~w8021;
assign w8023 = ~w8016 & w8021;
assign v3451 = ~(w8022 | w8023);
assign w8024 = v3451;
assign w8025 = w8003 & w8024;
assign v3452 = ~(w8003 | w8024);
assign w8026 = v3452;
assign v3453 = ~(w8025 | w8026);
assign w8027 = v3453;
assign v3454 = ~(w7927 | w7930);
assign w8028 = v3454;
assign v3455 = ~(w7917 | w7920);
assign w8029 = v3455;
assign v3456 = ~(w7886 | w7889);
assign w8030 = v3456;
assign v3457 = ~(w7911 | w7914);
assign w8031 = v3457;
assign v3458 = ~(w8030 | w8031);
assign w8032 = v3458;
assign w8033 = w8030 & w8031;
assign v3459 = ~(w8032 | w8033);
assign w8034 = v3459;
assign w8035 = ~w8029 & w8034;
assign w8036 = w8029 & ~w8034;
assign v3460 = ~(w8035 | w8036);
assign w8037 = v3460;
assign w8038 = ~w8028 & w8037;
assign w8039 = w8028 & ~w8037;
assign v3461 = ~(w8038 | w8039);
assign w8040 = v3461;
assign w8041 = w8027 & w8040;
assign v3462 = ~(w8027 | w8040);
assign w8042 = v3462;
assign v3463 = ~(w8041 | w8042);
assign w8043 = v3463;
assign w8044 = ~w7954 & w8043;
assign w8045 = w7954 & ~w8043;
assign v3464 = ~(w8044 | w8045);
assign w8046 = v3464;
assign w8047 = w8046 & w9316;
assign w8048 = (w7471 & w9198) | (w7471 & w9199) | (w9198 & w9199);
assign v3465 = ~(w8047 | w8048);
assign w8049 = v3465;
assign v3466 = ~(w8038 | w8041);
assign w8050 = v3466;
assign w8051 = pi22 & pi63;
assign w8052 = pi23 & pi62;
assign v3467 = ~(w8008 | w8052);
assign w8053 = v3467;
assign w8054 = pi24 & pi62;
assign w8055 = w8006 & w8054;
assign v3468 = ~(w8053 | w8055);
assign w8056 = v3468;
assign w8057 = w8051 & ~w8056;
assign w8058 = ~w8051 & w8056;
assign v3469 = ~(w8057 | w8058);
assign w8059 = v3469;
assign v3470 = ~(w7982 | w7985);
assign w8060 = v3470;
assign v3471 = ~(w7992 | w7995);
assign w8061 = v3471;
assign w8062 = w8060 & w8061;
assign v3472 = ~(w8060 | w8061);
assign w8063 = v3472;
assign v3473 = ~(w8062 | w8063);
assign w8064 = v3473;
assign w8065 = ~w8059 & w8064;
assign w8066 = w8059 & ~w8064;
assign v3474 = ~(w8065 | w8066);
assign w8067 = v3474;
assign w8068 = pi25 & pi60;
assign w8069 = pi29 & pi56;
assign w8070 = pi31 & pi54;
assign w8071 = pi30 & pi55;
assign w8072 = ~w8070 & w8071;
assign w8073 = w8070 & ~w8071;
assign v3475 = ~(w8072 | w8073);
assign w8074 = v3475;
assign w8075 = w8069 & w8074;
assign v3476 = ~(w8069 | w8074);
assign w8076 = v3476;
assign v3477 = ~(w8075 | w8076);
assign w8077 = v3477;
assign w8078 = w8068 & w8077;
assign v3478 = ~(w8068 | w8077);
assign w8079 = v3478;
assign v3479 = ~(w8078 | w8079);
assign w8080 = v3479;
assign w8081 = pi26 & pi59;
assign w8082 = pi27 & pi58;
assign v3480 = ~(w7971 | w8082);
assign w8083 = v3480;
assign w8084 = pi28 & pi58;
assign w8085 = w7969 & w8084;
assign v3481 = ~(w8083 | w8085);
assign w8086 = v3481;
assign w8087 = w8081 & ~w8086;
assign w8088 = ~w8081 & w8086;
assign v3482 = ~(w8087 | w8088);
assign w8089 = v3482;
assign w8090 = w8080 & ~w8089;
assign w8091 = ~w8080 & w8089;
assign v3483 = ~(w8090 | w8091);
assign w8092 = v3483;
assign v3484 = ~(w7965 | w7977);
assign w8093 = v3484;
assign v3485 = ~(w7959 | w7962);
assign w8094 = v3485;
assign w8095 = w7968 & ~w7970;
assign v3486 = ~(w7972 | w8095);
assign w8096 = v3486;
assign v3487 = ~(w8094 | w8096);
assign w8097 = v3487;
assign w8098 = w8094 & w8096;
assign v3488 = ~(w8097 | w8098);
assign w8099 = v3488;
assign w8100 = ~w8093 & w8099;
assign w8101 = w8093 & ~w8099;
assign v3489 = ~(w8100 | w8101);
assign w8102 = v3489;
assign w8103 = w8009 & w8015;
assign v3490 = ~(w8009 | w8015);
assign w8104 = v3490;
assign v3491 = ~(w8103 | w8104);
assign w8105 = v3491;
assign v3492 = ~(w8011 | w8105);
assign w8106 = v3492;
assign w8107 = w8102 & ~w8106;
assign w8108 = ~w8102 & w8106;
assign v3493 = ~(w8107 | w8108);
assign w8109 = v3493;
assign w8110 = w8092 & w8109;
assign v3494 = ~(w8092 | w8109);
assign w8111 = v3494;
assign v3495 = ~(w8110 | w8111);
assign w8112 = v3495;
assign w8113 = w8067 & ~w8112;
assign w8114 = ~w8067 & w8112;
assign v3496 = ~(w8113 | w8114);
assign w8115 = v3496;
assign v3497 = ~(w8032 | w8035);
assign w8116 = v3497;
assign v3498 = ~(w8022 | w8025);
assign w8117 = v3498;
assign v3499 = ~(w7998 | w8001);
assign w8118 = v3499;
assign v3500 = ~(w8019 | w8118);
assign w8119 = v3500;
assign w8120 = w8019 & w8118;
assign v3501 = ~(w8119 | w8120);
assign w8121 = v3501;
assign w8122 = ~w8117 & w8121;
assign w8123 = w8117 & ~w8121;
assign v3502 = ~(w8122 | w8123);
assign w8124 = v3502;
assign w8125 = ~w8116 & w8124;
assign w8126 = w8116 & ~w8124;
assign v3503 = ~(w8125 | w8126);
assign w8127 = v3503;
assign w8128 = ~w8115 & w8127;
assign w8129 = w8115 & ~w8127;
assign v3504 = ~(w8128 | w8129);
assign w8130 = v3504;
assign w8131 = w8050 & ~w8130;
assign w8132 = ~w8050 & w8130;
assign v3505 = ~(w8131 | w8132);
assign w8133 = v3505;
assign w8134 = (w7471 & w9200) | (w7471 & w9201) | (w9200 & w9201);
assign w8135 = (w9075 & w9076) | (w9075 & w9316) | (w9076 & w9316);
assign v3506 = ~(w8134 | w8135);
assign w8136 = v3506;
assign w8137 = w8044 & ~w8131;
assign v3507 = ~(w8132 | w8137);
assign w8138 = v3507;
assign v3508 = ~(w8045 | w8131);
assign w8139 = v3508;
assign v3509 = ~(w8132 | w8139);
assign w8140 = v3509;
assign v3510 = ~(w8125 | w8128);
assign w8141 = v3510;
assign w8142 = pi25 & pi61;
assign w8143 = pi29 & pi57;
assign w8144 = pi31 & pi55;
assign w8145 = pi30 & pi56;
assign w8146 = ~w8144 & w8145;
assign w8147 = w8144 & ~w8145;
assign v3511 = ~(w8146 | w8147);
assign w8148 = v3511;
assign w8149 = w8143 & w8148;
assign v3512 = ~(w8143 | w8148);
assign w8150 = v3512;
assign v3513 = ~(w8149 | w8150);
assign w8151 = v3513;
assign w8152 = w8142 & w8151;
assign v3514 = ~(w8142 | w8151);
assign w8153 = v3514;
assign v3515 = ~(w8152 | w8153);
assign w8154 = v3515;
assign w8155 = pi26 & pi60;
assign w8156 = pi27 & pi59;
assign v3516 = ~(w8084 | w8156);
assign w8157 = v3516;
assign w8158 = pi28 & pi59;
assign w8159 = w8082 & w8158;
assign v3517 = ~(w8157 | w8159);
assign w8160 = v3517;
assign w8161 = w8155 & ~w8160;
assign w8162 = ~w8155 & w8160;
assign v3518 = ~(w8161 | w8162);
assign w8163 = v3518;
assign w8164 = w8154 & ~w8163;
assign w8165 = ~w8154 & w8163;
assign v3519 = ~(w8164 | w8165);
assign w8166 = v3519;
assign v3520 = ~(w8078 | w8090);
assign w8167 = v3520;
assign v3521 = ~(w8072 | w8075);
assign w8168 = v3521;
assign w8169 = w8081 & ~w8083;
assign v3522 = ~(w8085 | w8169);
assign w8170 = v3522;
assign v3523 = ~(w8168 | w8170);
assign w8171 = v3523;
assign w8172 = w8168 & w8170;
assign v3524 = ~(w8171 | w8172);
assign w8173 = v3524;
assign w8174 = ~w8167 & w8173;
assign w8175 = w8167 & ~w8173;
assign v3525 = ~(w8174 | w8175);
assign w8176 = v3525;
assign v3526 = ~(w8055 | w8058);
assign w8177 = v3526;
assign w8178 = w8176 & ~w8177;
assign w8179 = ~w8176 & w8177;
assign v3527 = ~(w8178 | w8179);
assign w8180 = v3527;
assign w8181 = w8166 & w8180;
assign v3528 = ~(w8166 | w8180);
assign w8182 = v3528;
assign v3529 = ~(w8181 | w8182);
assign w8183 = v3529;
assign w8184 = pi23 & pi63;
assign w8185 = w8054 & ~w8184;
assign w8186 = ~w8054 & w8184;
assign v3530 = ~(w8185 | w8186);
assign w8187 = v3530;
assign v3531 = ~(w8097 | w8100);
assign w8188 = v3531;
assign w8189 = ~w8103 & w8188;
assign w8190 = w8103 & ~w8188;
assign v3532 = ~(w8189 | w8190);
assign w8191 = v3532;
assign w8192 = w8187 & ~w8191;
assign w8193 = ~w8187 & w8191;
assign v3533 = ~(w8192 | w8193);
assign w8194 = v3533;
assign w8195 = w8183 & w8194;
assign v3534 = ~(w8183 | w8194);
assign w8196 = v3534;
assign v3535 = ~(w8195 | w8196);
assign w8197 = v3535;
assign v3536 = ~(w8119 | w8122);
assign w8198 = v3536;
assign v3537 = ~(w8065 | w8113);
assign w8199 = v3537;
assign v3538 = ~(w8107 | w8110);
assign w8200 = v3538;
assign v3539 = ~(w8062 | w8200);
assign w8201 = v3539;
assign w8202 = w8062 & w8200;
assign v3540 = ~(w8201 | w8202);
assign w8203 = v3540;
assign w8204 = w8199 & w8203;
assign v3541 = ~(w8199 | w8203);
assign w8205 = v3541;
assign v3542 = ~(w8204 | w8205);
assign w8206 = v3542;
assign w8207 = ~w8198 & w8206;
assign w8208 = w8198 & ~w8206;
assign v3543 = ~(w8207 | w8208);
assign w8209 = v3543;
assign w8210 = w8197 & w8209;
assign v3544 = ~(w8197 | w8209);
assign w8211 = v3544;
assign v3545 = ~(w8210 | w8211);
assign w8212 = v3545;
assign w8213 = ~w8141 & w8212;
assign w8214 = w8141 & ~w8212;
assign v3546 = ~(w8213 | w8214);
assign w8215 = v3546;
assign w8216 = (w7471 & w9202) | (w7471 & w9203) | (w9202 & w9203);
assign w8217 = ~w8215 & w9317;
assign v3547 = ~(w8216 | w8217);
assign w8218 = v3547;
assign v3548 = ~(w8207 | w8210);
assign w8219 = v3548;
assign w8220 = pi29 & pi58;
assign w8221 = pi31 & pi56;
assign w8222 = pi30 & pi57;
assign w8223 = ~w8221 & w8222;
assign w8224 = w8221 & ~w8222;
assign v3549 = ~(w8223 | w8224);
assign w8225 = v3549;
assign w8226 = w8220 & w8225;
assign v3550 = ~(w8220 | w8225);
assign w8227 = v3550;
assign v3551 = ~(w8226 | w8227);
assign w8228 = v3551;
assign w8229 = pi26 & pi61;
assign w8230 = pi27 & pi60;
assign v3552 = ~(w8158 | w8230);
assign w8231 = v3552;
assign w8232 = pi28 & pi60;
assign w8233 = w8156 & w8232;
assign v3553 = ~(w8231 | w8233);
assign w8234 = v3553;
assign w8235 = w8229 & ~w8234;
assign w8236 = ~w8229 & w8234;
assign v3554 = ~(w8235 | w8236);
assign w8237 = v3554;
assign w8238 = w8228 & ~w8237;
assign w8239 = ~w8228 & w8237;
assign v3555 = ~(w8238 | w8239);
assign w8240 = v3555;
assign w8241 = pi24 & pi63;
assign w8242 = pi25 & pi62;
assign w8243 = w8241 & ~w8242;
assign w8244 = ~w8241 & w8242;
assign v3556 = ~(w8243 | w8244);
assign w8245 = v3556;
assign w8246 = w8240 & ~w8245;
assign w8247 = ~w8240 & w8245;
assign v3557 = ~(w8246 | w8247);
assign w8248 = v3557;
assign v3558 = ~(w8171 | w8174);
assign w8249 = v3558;
assign v3559 = ~(w8152 | w8164);
assign w8250 = v3559;
assign v3560 = ~(w8146 | w8149);
assign w8251 = v3560;
assign w8252 = w8155 & ~w8157;
assign v3561 = ~(w8159 | w8252);
assign w8253 = v3561;
assign v3562 = ~(w8251 | w8253);
assign w8254 = v3562;
assign w8255 = w8251 & w8253;
assign v3563 = ~(w8254 | w8255);
assign w8256 = v3563;
assign w8257 = ~w8250 & w8256;
assign w8258 = w8250 & ~w8256;
assign v3564 = ~(w8257 | w8258);
assign w8259 = v3564;
assign w8260 = ~w8249 & w8259;
assign w8261 = w8249 & ~w8259;
assign v3565 = ~(w8260 | w8261);
assign w8262 = v3565;
assign w8263 = w8185 & w8262;
assign v3566 = ~(w8185 | w8262);
assign w8264 = v3566;
assign v3567 = ~(w8263 | w8264);
assign w8265 = v3567;
assign w8266 = w8248 & w8265;
assign v3568 = ~(w8248 | w8265);
assign w8267 = v3568;
assign v3569 = ~(w8266 | w8267);
assign w8268 = v3569;
assign v3570 = ~(w8201 | w8204);
assign w8269 = v3570;
assign v3571 = ~(w8192 | w8195);
assign w8270 = v3571;
assign v3572 = ~(w8178 | w8181);
assign w8271 = v3572;
assign v3573 = ~(w8189 | w8271);
assign w8272 = v3573;
assign w8273 = w8189 & w8271;
assign v3574 = ~(w8272 | w8273);
assign w8274 = v3574;
assign w8275 = ~w8270 & w8274;
assign w8276 = w8270 & ~w8274;
assign v3575 = ~(w8275 | w8276);
assign w8277 = v3575;
assign w8278 = ~w8269 & w8277;
assign w8279 = w8269 & ~w8277;
assign v3576 = ~(w8278 | w8279);
assign w8280 = v3576;
assign w8281 = w8268 & w8280;
assign v3577 = ~(w8268 | w8280);
assign w8282 = v3577;
assign v3578 = ~(w8281 | w8282);
assign w8283 = v3578;
assign w8284 = ~w8219 & w8283;
assign w8285 = w8219 & ~w8283;
assign v3579 = ~(w8284 | w8285);
assign w8286 = v3579;
assign w8287 = (w7471 & w9204) | (w7471 & w9205) | (w9204 & w9205);
assign w8288 = ~w8214 & w8286;
assign w8289 = (w9197 & w9286) | (w9197 & w9287) | (w9286 & w9287);
assign v3580 = ~(w8287 | w8289);
assign w8290 = v3580;
assign v3581 = ~(w8278 | w8281);
assign w8291 = v3581;
assign v3582 = ~(w8272 | w8275);
assign w8292 = v3582;
assign v3583 = ~(w8246 | w8266);
assign w8293 = v3583;
assign v3584 = ~(w8260 | w8263);
assign w8294 = v3584;
assign v3585 = ~(w8243 | w8294);
assign w8295 = v3585;
assign w8296 = w8243 & w8294;
assign v3586 = ~(w8295 | w8296);
assign w8297 = v3586;
assign w8298 = ~w8293 & w8297;
assign w8299 = w8293 & ~w8297;
assign v3587 = ~(w8298 | w8299);
assign w8300 = v3587;
assign w8301 = ~w8292 & w8300;
assign w8302 = w8292 & ~w8300;
assign v3588 = ~(w8301 | w8302);
assign w8303 = v3588;
assign w8304 = pi29 & pi59;
assign w8305 = pi31 & pi57;
assign w8306 = pi30 & pi58;
assign w8307 = ~w8305 & w8306;
assign w8308 = w8305 & ~w8306;
assign v3589 = ~(w8307 | w8308);
assign w8309 = v3589;
assign w8310 = w8304 & w8309;
assign v3590 = ~(w8304 | w8309);
assign w8311 = v3590;
assign v3591 = ~(w8310 | w8311);
assign w8312 = v3591;
assign w8313 = w8232 & w8312;
assign v3592 = ~(w8232 | w8312);
assign w8314 = v3592;
assign v3593 = ~(w8313 | w8314);
assign w8315 = v3593;
assign w8316 = pi25 & pi63;
assign w8317 = pi27 & pi61;
assign w8318 = pi26 & pi62;
assign v3594 = ~(w8317 | w8318);
assign w8319 = v3594;
assign w8320 = pi27 & pi62;
assign w8321 = w8229 & w8320;
assign v3595 = ~(w8319 | w8321);
assign w8322 = v3595;
assign w8323 = w8316 & ~w8322;
assign w8324 = ~w8316 & w8322;
assign v3596 = ~(w8323 | w8324);
assign w8325 = v3596;
assign w8326 = w8315 & w8325;
assign v3597 = ~(w8315 | w8325);
assign w8327 = v3597;
assign v3598 = ~(w8326 | w8327);
assign w8328 = v3598;
assign v3599 = ~(w8254 | w8257);
assign w8329 = v3599;
assign v3600 = ~(w8223 | w8226);
assign w8330 = v3600;
assign w8331 = w8229 & ~w8231;
assign v3601 = ~(w8233 | w8331);
assign w8332 = v3601;
assign v3602 = ~(w8330 | w8332);
assign w8333 = v3602;
assign w8334 = w8330 & w8332;
assign v3603 = ~(w8333 | w8334);
assign w8335 = v3603;
assign w8336 = w8238 & w8335;
assign v3604 = ~(w8238 | w8335);
assign w8337 = v3604;
assign v3605 = ~(w8336 | w8337);
assign w8338 = v3605;
assign w8339 = w8329 & ~w8338;
assign w8340 = ~w8329 & w8338;
assign v3606 = ~(w8339 | w8340);
assign w8341 = v3606;
assign w8342 = w8328 & ~w8341;
assign w8343 = ~w8328 & w8341;
assign v3607 = ~(w8342 | w8343);
assign w8344 = v3607;
assign w8345 = w8303 & w8344;
assign v3608 = ~(w8303 | w8344);
assign w8346 = v3608;
assign v3609 = ~(w8345 | w8346);
assign w8347 = v3609;
assign w8348 = ~w8291 & w8347;
assign w8349 = w8291 & ~w8347;
assign v3610 = ~(w8348 | w8349);
assign w8350 = v3610;
assign w8351 = (w9197 & w9288) | (w9197 & w9289) | (w9288 & w9289);
assign w8352 = (w7471 & w9206) | (w7471 & w9207) | (w9206 & w9207);
assign v3611 = ~(w8351 | w8352);
assign w8353 = v3611;
assign v3612 = ~(w8301 | w8345);
assign w8354 = v3612;
assign w8355 = pi29 & pi60;
assign w8356 = pi31 & pi58;
assign w8357 = pi30 & pi59;
assign w8358 = ~w8356 & w8357;
assign w8359 = w8356 & ~w8357;
assign v3613 = ~(w8358 | w8359);
assign w8360 = v3613;
assign w8361 = w8355 & w8360;
assign v3614 = ~(w8355 | w8360);
assign w8362 = v3614;
assign v3615 = ~(w8361 | w8362);
assign w8363 = v3615;
assign w8364 = pi26 & pi63;
assign w8365 = pi28 & pi61;
assign v3616 = ~(w8320 | w8365);
assign w8366 = v3616;
assign w8367 = pi28 & pi62;
assign w8368 = w8317 & w8367;
assign v3617 = ~(w8366 | w8368);
assign w8369 = v3617;
assign w8370 = w8364 & ~w8369;
assign w8371 = ~w8364 & w8369;
assign v3618 = ~(w8370 | w8371);
assign w8372 = v3618;
assign w8373 = w8363 & w8372;
assign v3619 = ~(w8363 | w8372);
assign w8374 = v3619;
assign v3620 = ~(w8373 | w8374);
assign w8375 = v3620;
assign w8376 = w8307 & w8313;
assign v3621 = ~(w8307 | w8313);
assign w8377 = v3621;
assign v3622 = ~(w8376 | w8377);
assign w8378 = v3622;
assign v3623 = ~(w8310 | w8378);
assign w8379 = v3623;
assign v3624 = ~(w8333 | w8336);
assign w8380 = v3624;
assign w8381 = w8379 & w8380;
assign v3625 = ~(w8379 | w8380);
assign w8382 = v3625;
assign v3626 = ~(w8381 | w8382);
assign w8383 = v3626;
assign w8384 = w8375 & ~w8383;
assign w8385 = ~w8375 & w8383;
assign v3627 = ~(w8384 | w8385);
assign w8386 = v3627;
assign v3628 = ~(w8295 | w8298);
assign w8387 = v3628;
assign v3629 = ~(w8326 | w8342);
assign w8388 = v3629;
assign v3630 = ~(w8321 | w8324);
assign w8389 = v3630;
assign v3631 = ~(w8339 | w8389);
assign w8390 = v3631;
assign w8391 = w8339 & w8389;
assign v3632 = ~(w8390 | w8391);
assign w8392 = v3632;
assign w8393 = ~w8388 & w8392;
assign w8394 = w8388 & ~w8392;
assign v3633 = ~(w8393 | w8394);
assign w8395 = v3633;
assign w8396 = ~w8387 & w8395;
assign w8397 = w8387 & ~w8395;
assign v3634 = ~(w8396 | w8397);
assign w8398 = v3634;
assign w8399 = w8386 & w8398;
assign v3635 = ~(w8386 | w8398);
assign w8400 = v3635;
assign v3636 = ~(w8399 | w8400);
assign w8401 = v3636;
assign w8402 = w8354 & ~w8401;
assign w8403 = ~w8354 & w8401;
assign v3637 = ~(w8402 | w8403);
assign w8404 = v3637;
assign w8405 = (~w7953 & w9080) | (~w7953 & w9081) | (w9080 & w9081);
assign w8406 = (w7953 & w9082) | (w7953 & w9083) | (w9082 & w9083);
assign v3638 = ~(w8405 | w8406);
assign w8407 = v3638;
assign w8408 = w8350 & w8404;
assign v3639 = ~(w8348 | w8403);
assign w8409 = v3639;
assign v3640 = ~(w8402 | w8409);
assign w8410 = v3640;
assign v3641 = ~(w8408 | w8410);
assign w8411 = v3641;
assign v3642 = ~(w8284 | w8410);
assign w8412 = v3642;
assign v3643 = ~(w8396 | w8399);
assign w8413 = v3643;
assign v3644 = ~(w8358 | w8361);
assign w8414 = v3644;
assign v3645 = ~(w8376 | w8414);
assign w8415 = v3645;
assign w8416 = pi31 & pi59;
assign w8417 = pi30 & pi60;
assign w8418 = ~w8416 & w8417;
assign w8419 = w8416 & ~w8417;
assign v3646 = ~(w8418 | w8419);
assign w8420 = v3646;
assign w8421 = pi27 & pi63;
assign w8422 = pi29 & pi61;
assign v3647 = ~(w8367 | w8422);
assign w8423 = v3647;
assign w8424 = pi29 & pi62;
assign w8425 = w8365 & w8424;
assign v3648 = ~(w8423 | w8425);
assign w8426 = v3648;
assign w8427 = w8421 & ~w8426;
assign w8428 = ~w8421 & w8426;
assign v3649 = ~(w8427 | w8428);
assign w8429 = v3649;
assign w8430 = w8420 & w8429;
assign v3650 = ~(w8420 | w8429);
assign w8431 = v3650;
assign v3651 = ~(w8430 | w8431);
assign w8432 = v3651;
assign w8433 = ~w8415 & w8432;
assign w8434 = w8415 & ~w8432;
assign v3652 = ~(w8433 | w8434);
assign w8435 = v3652;
assign v3653 = ~(w8390 | w8393);
assign w8436 = v3653;
assign v3654 = ~(w8373 | w8384);
assign w8437 = v3654;
assign v3655 = ~(w8368 | w8371);
assign w8438 = v3655;
assign v3656 = ~(w8381 | w8438);
assign w8439 = v3656;
assign w8440 = w8381 & w8438;
assign v3657 = ~(w8439 | w8440);
assign w8441 = v3657;
assign w8442 = ~w8437 & w8441;
assign w8443 = w8437 & ~w8441;
assign v3658 = ~(w8442 | w8443);
assign w8444 = v3658;
assign w8445 = ~w8436 & w8444;
assign w8446 = w8436 & ~w8444;
assign v3659 = ~(w8445 | w8446);
assign w8447 = v3659;
assign w8448 = w8435 & w8447;
assign v3660 = ~(w8435 | w8447);
assign w8449 = v3660;
assign v3661 = ~(w8448 | w8449);
assign w8450 = v3661;
assign w8451 = ~w8413 & w8450;
assign w8452 = w8413 & ~w8450;
assign v3662 = ~(w8451 | w8452);
assign w8453 = v3662;
assign w8454 = (~w7471 & w9208) | (~w7471 & w9209) | (w9208 & w9209);
assign w8455 = ~w8410 & w8453;
assign w8456 = (w7471 & w9210) | (w7471 & w9211) | (w9210 & w9211);
assign v3663 = ~(w8454 | w8456);
assign w8457 = v3663;
assign v3664 = ~(w8445 | w8448);
assign w8458 = v3664;
assign w8459 = pi28 & pi63;
assign w8460 = ~w8418 & w8459;
assign w8461 = w8418 & ~w8459;
assign v3665 = ~(w8460 | w8461);
assign w8462 = v3665;
assign w8463 = pi31 & pi60;
assign w8464 = pi30 & pi61;
assign w8465 = ~w8463 & w8464;
assign w8466 = w8463 & ~w8464;
assign v3666 = ~(w8465 | w8466);
assign w8467 = v3666;
assign w8468 = w8424 & w8467;
assign v3667 = ~(w8424 | w8467);
assign w8469 = v3667;
assign v3668 = ~(w8468 | w8469);
assign w8470 = v3668;
assign w8471 = ~w8462 & w8470;
assign w8472 = w8462 & ~w8470;
assign v3669 = ~(w8471 | w8472);
assign w8473 = v3669;
assign v3670 = ~(w8439 | w8442);
assign w8474 = v3670;
assign v3671 = ~(w8430 | w8433);
assign w8475 = v3671;
assign v3672 = ~(w8425 | w8428);
assign w8476 = v3672;
assign v3673 = ~(w8414 | w8476);
assign w8477 = v3673;
assign w8478 = w8414 & w8476;
assign v3674 = ~(w8477 | w8478);
assign w8479 = v3674;
assign w8480 = ~w8475 & w8479;
assign w8481 = w8475 & ~w8479;
assign v3675 = ~(w8480 | w8481);
assign w8482 = v3675;
assign w8483 = ~w8474 & w8482;
assign w8484 = w8474 & ~w8482;
assign v3676 = ~(w8483 | w8484);
assign w8485 = v3676;
assign w8486 = w8473 & w8485;
assign v3677 = ~(w8473 | w8485);
assign w8487 = v3677;
assign v3678 = ~(w8486 | w8487);
assign w8488 = v3678;
assign w8489 = ~w8458 & w8488;
assign w8490 = w8458 & ~w8488;
assign v3679 = ~(w8489 | w8490);
assign w8491 = v3679;
assign w8492 = (w7953 & w9086) | (w7953 & w9087) | (w9086 & w9087);
assign v3680 = ~(w8451 | w8491);
assign w8493 = v3680;
assign w8494 = w8451 & w8491;
assign v3681 = ~(w8493 | w8494);
assign w8495 = v3681;
assign w8496 = (~w7953 & w9088) | (~w7953 & w9089) | (w9088 & w9089);
assign v3682 = ~(w8492 | w8496);
assign w8497 = v3682;
assign v3683 = ~(w8483 | w8486);
assign w8498 = v3683;
assign v3684 = ~(w8465 | w8468);
assign w8499 = v3684;
assign v3685 = ~(w8460 | w8499);
assign w8500 = v3685;
assign w8501 = w8460 & w8499;
assign v3686 = ~(w8500 | w8501);
assign w8502 = v3686;
assign w8503 = w8471 & w8502;
assign v3687 = ~(w8471 | w8502);
assign w8504 = v3687;
assign v3688 = ~(w8503 | w8504);
assign w8505 = v3688;
assign v3689 = ~(w8477 | w8480);
assign w8506 = v3689;
assign w8507 = w8505 & ~w8506;
assign w8508 = ~w8505 & w8506;
assign v3690 = ~(w8507 | w8508);
assign w8509 = v3690;
assign w8510 = pi29 & pi63;
assign w8511 = pi31 & pi61;
assign w8512 = pi30 & pi62;
assign w8513 = w8511 & ~w8512;
assign w8514 = ~w8511 & w8512;
assign v3691 = ~(w8513 | w8514);
assign w8515 = v3691;
assign w8516 = w8510 & ~w8515;
assign w8517 = ~w8510 & w8515;
assign v3692 = ~(w8516 | w8517);
assign w8518 = v3692;
assign w8519 = w8509 & ~w8518;
assign w8520 = ~w8509 & w8518;
assign v3693 = ~(w8519 | w8520);
assign w8521 = v3693;
assign w8522 = ~w8498 & w8521;
assign w8523 = w8498 & ~w8521;
assign v3694 = ~(w8522 | w8523);
assign w8524 = v3694;
assign v3695 = ~(w8452 | w8490);
assign w8525 = v3695;
assign w8526 = ~w8455 & w8525;
assign v3696 = ~(w8489 | w8526);
assign w8527 = v3696;
assign w8528 = ~w8284 & w8527;
assign w8529 = w8408 & w8525;
assign w8530 = w8527 & ~w8529;
assign w8531 = (w9197 & w9290) | (w9197 & w9291) | (w9290 & w9291);
assign w8532 = (w7471 & w9212) | (w7471 & w9213) | (w9212 & w9213);
assign v3697 = ~(w8531 | w8532);
assign w8533 = v3697;
assign v3698 = ~(w8507 | w8519);
assign w8534 = v3698;
assign v3699 = ~(w8500 | w8503);
assign w8535 = v3699;
assign w8536 = ~w8510 & w8514;
assign w8537 = pi31 & pi63;
assign w8538 = ~w8512 & w8537;
assign w8539 = w8422 & w8538;
assign v3700 = ~(w8536 | w8539);
assign w8540 = v3700;
assign w8541 = ~w8535 & w8540;
assign w8542 = w8535 & ~w8540;
assign v3701 = ~(w8541 | w8542);
assign w8543 = v3701;
assign w8544 = pi31 & pi62;
assign w8545 = pi30 & pi63;
assign w8546 = w8544 & ~w8545;
assign w8547 = ~w8544 & w8545;
assign v3702 = ~(w8546 | w8547);
assign w8548 = v3702;
assign w8549 = w8543 & w8548;
assign v3703 = ~(w8543 | w8548);
assign w8550 = v3703;
assign v3704 = ~(w8549 | w8550);
assign w8551 = v3704;
assign w8552 = w8534 & ~w8551;
assign w8553 = ~w8534 & w8551;
assign v3705 = ~(w8552 | w8553);
assign w8554 = v3705;
assign w8555 = w8522 & ~w8554;
assign w8556 = ~w8522 & w8554;
assign v3706 = ~(w8555 | w8556);
assign w8557 = v3706;
assign w8558 = (~w7953 & w9091) | (~w7953 & w9092) | (w9091 & w9092);
assign w8559 = w8524 & w8554;
assign w8560 = (w9197 & w9292) | (w9197 & w9293) | (w9292 & w9293);
assign v3707 = ~(w8558 | w8560);
assign w8561 = v3707;
assign v3708 = ~(w8541 | w8549);
assign w8562 = v3708;
assign v3709 = ~(w8536 | w8538);
assign w8563 = v3709;
assign w8564 = w8562 & w8563;
assign v3710 = ~(w8562 | w8563);
assign w8565 = v3710;
assign v3711 = ~(w8564 | w8565);
assign w8566 = v3711;
assign v3712 = ~(w8552 | w8556);
assign w8567 = v3712;
assign v3713 = ~(w8566 | w8567);
assign w8568 = v3713;
assign w8569 = w8566 & w8567;
assign v3714 = ~(w8568 | w8569);
assign w8570 = v3714;
assign w8571 = (~w7953 & w9093) | (~w7953 & w9094) | (w9093 & w9094);
assign w8572 = (w7953 & w9095) | (w7953 & w9096) | (w9095 & w9096);
assign v3715 = ~(w8571 | w8572);
assign w8573 = v3715;
assign v3716 = ~(w8565 | w8567);
assign w8574 = v3716;
assign w8575 = (~w7953 & w9097) | (~w7953 & w9098) | (w9097 & w9098);
assign v3717 = ~(w8564 | w8575);
assign w8576 = v3717;
assign v3718 = ~(w1 | w9);
assign w8577 = v3718;
assign w8578 = w15 & ~w29;
assign w8579 = w35 & ~w56;
assign v3719 = ~(w268 | w262);
assign w8580 = v3719;
assign v3720 = ~(w275 | w274);
assign w8581 = v3720;
assign w8582 = w310 & ~w295;
assign v3721 = ~(w349 | w382);
assign w8583 = v3721;
assign v3722 = ~(w478 | w476);
assign w8584 = v3722;
assign v3723 = ~(w448 | w446);
assign w8585 = v3723;
assign w8586 = (~w472 & ~w483) | (~w472 & w8662) | (~w483 & w8662);
assign w8587 = w440 & ~w558;
assign w8588 = w768 & ~w757;
assign v3724 = ~(w1068 | w1067);
assign w8589 = v3724;
assign v3725 = ~(w1410 | w1408);
assign w8590 = v3725;
assign w8591 = w1520 & ~w1509;
assign v3726 = ~(w1543 | w1541);
assign w8592 = v3726;
assign v3727 = ~(w1443 | w1564);
assign w8593 = v3727;
assign w8594 = w1443 & w1564;
assign w8595 = w1734 & ~w1723;
assign v3728 = ~(w1715 | w1717);
assign w8596 = v3728;
assign w8597 = (~w1889 & w1723) | (~w1889 & w8663) | (w1723 & w8663);
assign w8598 = ~w1888 & w2026;
assign v3729 = ~(w2029 | w2030);
assign w8599 = v3729;
assign w8600 = w1924 & ~w1913;
assign w8601 = w1862 & ~w1851;
assign w8602 = w2060 & ~w2049;
assign w8603 = w2087 & ~w2076;
assign w8604 = w2292 & ~w2281;
assign w8605 = w2250 & ~w2239;
assign w8606 = (~w2465 & w2281) | (~w2465 & w8664) | (w2281 & w8664);
assign v3730 = ~(w2413 | w2412);
assign w8607 = v3730;
assign w8608 = w2758 & ~w2747;
assign w8609 = w2961 & ~w2950;
assign w8610 = w2985 & ~w2974;
assign w8611 = w3093 & ~w3082;
assign w8612 = w3065 & ~w3054;
assign w8613 = w3349 & ~w3338;
assign w8614 = w3373 & ~w3362;
assign w8615 = w3723 & ~w3712;
assign w8616 = w3691 & ~w3680;
assign w8617 = w3592 & ~w3581;
assign w8618 = w3616 & ~w3605;
assign w8619 = w3899 & ~w3888;
assign w8620 = w3780 & ~w3769;
assign w8621 = w4114 & ~w4103;
assign w8622 = w4034 & ~w4023;
assign w8623 = w4083 & ~w4072;
assign w8624 = w4059 & ~w4048;
assign w8625 = w4289 & ~w4278;
assign w8626 = w4548 & ~w4536;
assign w8627 = w4597 & ~w4585;
assign w8628 = w4573 & ~w4561;
assign w8629 = w4847 & ~w4836;
assign w8630 = w4797 & ~w4786;
assign w8631 = w4822 & ~w4811;
assign w8632 = w5125 & ~w5114;
assign w8633 = w5097 & ~w5086;
assign w8634 = w5329 & ~w5318;
assign w8635 = w5364 & ~w5353;
assign w8636 = w5621 & ~w5610;
assign w8637 = w5523 & ~w5512;
assign w8638 = w5548 & ~w5537;
assign w8639 = w5844 & ~w5833;
assign w8640 = w5816 & ~w5805;
assign w8641 = w5786 & ~w5775;
assign w8642 = w6031 & ~w6020;
assign v3731 = ~(w6042 | w6040);
assign w8643 = v3731;
assign v3732 = ~(w6000 | w5998);
assign w8644 = v3732;
assign v3733 = ~(w5958 | w5956);
assign w8645 = v3733;
assign w8646 = w5947 & w6298;
assign v3734 = ~(w5947 | w6298);
assign w8647 = v3734;
assign w8648 = (~w5944 & ~w5961) | (~w5944 & w9099) | (~w5961 & w9099);
assign v3735 = ~(w6310 | w6320);
assign w8649 = v3735;
assign v3736 = ~(w6175 | w6173);
assign w8650 = v3736;
assign w8651 = w6258 & ~w6247;
assign v3737 = ~(w6227 | w6225);
assign w8652 = v3737;
assign v3738 = ~(w6316 | w6314);
assign w8653 = v3738;
assign v3739 = ~(w6307 | w6305);
assign w8654 = v3739;
assign w8655 = (~w6160 & ~w6178) | (~w6160 & w9100) | (~w6178 & w9100);
assign v3740 = ~(w6869 | w6860);
assign w8656 = v3740;
assign w8657 = w7952 & w7460;
assign w8658 = (w7952 & ~w7474) | (w7952 & w8657) | (~w7474 & w8657);
assign w8659 = (~w8140 & w7949) | (~w8140 & w9101) | (w7949 & w9101);
assign w8660 = ~w8213 & w8140;
assign v3741 = ~(w8213 | w8659);
assign w8661 = v3741;
assign v3742 = ~(w344 | w472);
assign w8662 = v3742;
assign w8663 = w1888 & ~w1889;
assign w8664 = w2464 & ~w2465;
assign w8665 = w193 & ~w162;
assign v3743 = ~(w190 | w178);
assign w8666 = v3743;
assign v3744 = ~(w158 | w156);
assign w8667 = v3744;
assign w8668 = w252 & ~w242;
assign v3745 = ~(w341 | w339);
assign w8669 = v3745;
assign v3746 = ~(w359 | w361);
assign w8670 = v3746;
assign w8671 = ~w367 & w478;
assign w8672 = w367 & ~w478;
assign w8673 = w469 & ~w458;
assign v3747 = ~(w450 | w452);
assign w8674 = v3747;
assign w8675 = w550 & w476;
assign w8676 = w550 & ~w8584;
assign v3748 = ~(w594 | w589);
assign w8677 = v3748;
assign w8678 = w525 & ~w514;
assign v3749 = ~(w506 | w508);
assign w8679 = v3749;
assign w8680 = w617 & ~w606;
assign w8681 = w722 & ~w711;
assign v3750 = ~(w932 | w927);
assign w8682 = v3750;
assign w8683 = w843 & w984;
assign w8684 = ~w845 & w986;
assign w8685 = w888 & ~w876;
assign v3751 = ~(w1038 | w1036);
assign w8686 = v3751;
assign w8687 = w969 & ~w957;
assign w8688 = w1017 & ~w1005;
assign w8689 = w1140 & ~w1129;
assign w8690 = (~w1067 & w1286) | (~w1067 & w9214) | (w1286 & w9214);
assign w8691 = ~w1287 & w8589;
assign w8692 = ~w1286 & w9215;
assign w8693 = w1287 & ~w8589;
assign v3752 = ~(w1403 | w1401);
assign w8694 = v3752;
assign w8695 = ~w1419 & w1624;
assign v3753 = ~(w1536 | w1534);
assign w8696 = v3753;
assign v3754 = ~(w1548 | w1550);
assign w8697 = v3754;
assign v3755 = ~(w1756 | w1754);
assign w8698 = v3755;
assign v3756 = ~(w1694 | w1693);
assign w8699 = v3756;
assign v3757 = ~(w1749 | w1747);
assign w8700 = v3757;
assign v3758 = ~(w1765 | w1975);
assign w8701 = v3758;
assign w8702 = w1765 & w1975;
assign v3759 = ~(w2026 | w1889);
assign w8703 = v3759;
assign w8704 = ~w2026 & w8597;
assign v3760 = ~(w1877 | w1875);
assign w8705 = v3760;
assign w8706 = (w1883 & w1893) | (w1883 & w9216) | (w1893 & w9216);
assign v3761 = ~(w2098 | w2097);
assign w8707 = v3761;
assign v3762 = ~(w2108 | w2106);
assign w8708 = v3762;
assign w8709 = w2090 & ~w2112;
assign w8710 = ~w2330 & w2429;
assign v3763 = ~(w2064 | w2328);
assign w8711 = v3763;
assign v3764 = ~(w2261 | w2259);
assign w8712 = v3764;
assign v3765 = ~(w2307 | w2305);
assign w8713 = v3765;
assign v3766 = ~(w2511 | w2509);
assign w8714 = v3766;
assign v3767 = ~(w2471 | w2465);
assign w8715 = v3767;
assign w8716 = ~w2471 & w8606;
assign w8717 = w2455 & ~w2444;
assign w8718 = w2713 & ~w2702;
assign v3768 = ~(w2739 | w2741);
assign w8719 = v3768;
assign w8720 = w2685 & ~w2674;
assign v3769 = ~(w3017 | w3030);
assign w8721 = v3769;
assign v3770 = ~(w2826 | w2824);
assign w8722 = v3770;
assign w8723 = w2926 & ~w2925;
assign v3771 = ~(w3026 | w3024);
assign w8724 = v3771;
assign w8725 = (~w3264 & w3036) | (~w3264 & w8782) | (w3036 & w8782);
assign w8726 = (~w3099 & ~w3137) | (~w3099 & w8867) | (~w3137 & w8867);
assign w8727 = (~w3386 & ~w3424) | (~w3386 & w8868) | (~w3424 & w8868);
assign v3772 = ~(w3415 | w3413);
assign w8728 = v3772;
assign v3773 = ~(w3405 | w3403);
assign w8729 = v3773;
assign v3774 = ~(w3650 | w3648);
assign w8730 = v3774;
assign w8731 = (w3631 & ~w3669) | (w3631 & w8869) | (~w3669 & w8869);
assign w8732 = ~w3753 & w4009;
assign w8733 = w3829 & ~w3818;
assign v3775 = ~(w3857 | w3855);
assign w8734 = v3775;
assign v3776 = ~(w3846 | w3844);
assign w8735 = v3776;
assign w8736 = w3805 & ~w3794;
assign v3777 = ~(w3868 | w3866);
assign w8737 = v3777;
assign v3778 = ~(w3931 | w3929);
assign w8738 = v3778;
assign w8739 = (~w3838 & ~w3877) | (~w3838 & w8870) | (~w3877 & w8870);
assign w8740 = (w4092 & ~w4145) | (w4092 & w8871) | (~w4145 & w8871);
assign w8741 = w4366 & ~w4355;
assign w8742 = w4338 & ~w4327;
assign v3779 = ~(w4439 | w4437);
assign w8743 = v3779;
assign v3780 = ~(w4458 | w4456);
assign w8744 = v3780;
assign w8745 = (~w4344 & ~w4403) | (~w4344 & w8872) | (~w4403 & w8872);
assign w8746 = w4628 & ~w4616;
assign v3781 = ~(w4708 | w4706);
assign w8747 = v3781;
assign v3782 = ~(w4952 | w4950);
assign w8748 = v3782;
assign v3783 = ~(w4875 | w4873);
assign w8749 = v3783;
assign v3784 = ~(w4934 | w4932);
assign w8750 = v3784;
assign w8751 = (w5131 & w5195) | (w5131 & w9102) | (w5195 & w9102);
assign w8752 = (~w5373 & ~w5411) | (~w5373 & w9103) | (~w5411 & w9103);
assign w8753 = ~w5475 & w5696;
assign w8754 = w5475 & ~w5696;
assign v3785 = ~(w5479 | w5469);
assign w8755 = v3785;
assign w8756 = w5484 & w5706;
assign v3786 = ~(w5710 | w5495);
assign w8757 = v3786;
assign w8758 = (w5670 & w5687) | (w5670 & w9104) | (w5687 & w9104);
assign v3787 = ~(w5590 | w5588);
assign w8759 = v3787;
assign v3788 = ~(w5580 | w5578);
assign w8760 = v3788;
assign v3789 = ~(w5658 | w5656);
assign w8761 = v3789;
assign w8762 = w5659 & ~w5662;
assign w8763 = (~w5561 & ~w5599) | (~w5561 & w9105) | (~w5599 & w9105);
assign v3790 = ~(w5673 | w5897);
assign w8764 = v3790;
assign w8765 = w5673 & w5897;
assign w8766 = ~w5720 & w9106;
assign w8767 = (~w5909 & w5720) | (~w5909 & w9107) | (w5720 & w9107);
assign w8768 = (w5822 & w5885) | (w5822 & w9217) | (w5885 & w9217);
assign v3791 = ~(w5855 | w5853);
assign w8769 = v3791;
assign w8770 = ~w6130 & w6125;
assign w8771 = w6009 & ~w6063;
assign w8772 = w5989 & ~w5978;
assign w8773 = w6236 & ~w6280;
assign w8774 = w6206 & ~w6195;
assign w8775 = w6440 & ~w6484;
assign v3792 = ~(w6427 | w6425);
assign w8776 = v3792;
assign w8777 = w7604 & w7460;
assign w8778 = (w7604 & ~w7474) | (w7604 & w8777) | (~w7474 & w8777);
assign w8779 = ~w7600 & w7724;
assign w8780 = w8288 & ~w8660;
assign w8781 = w8288 & ~w8661;
assign w8782 = w3263 & ~w3264;
assign w8783 = w4004 & ~w4261;
assign w8784 = ~w4262 & w4261;
assign v3793 = ~(w4262 | w8783);
assign w8785 = v3793;
assign w8786 = w4499 & ~w4510;
assign w8787 = w4475 & ~w4674;
assign w8788 = ~w4475 & w4674;
assign v3794 = ~(w4487 | w4485);
assign w8789 = v3794;
assign v3795 = ~(w4442 | w4445);
assign w8790 = v3795;
assign w8791 = (w4472 & w4490) | (w4472 & w8873) | (w4490 & w8873);
assign v3796 = ~(w4752 | w4763);
assign w8792 = v3796;
assign v3797 = ~(w4731 | w4729);
assign w8793 = v3797;
assign v3798 = ~(w4305 | w4579);
assign w8794 = v3798;
assign v3799 = ~(w4690 | w4688);
assign w8795 = v3799;
assign v3800 = ~(w4700 | w4721);
assign w8796 = v3800;
assign w8797 = (w4606 & w4663) | (w4606 & w9108) | (w4663 & w9108);
assign v3801 = ~(w4759 | w4757);
assign w8798 = v3801;
assign v3802 = ~(w4684 | w4682);
assign w8799 = v3802;
assign w8800 = (w4726 & w4743) | (w4726 & w8874) | (w4743 & w8874);
assign w8801 = w5042 & ~w4932;
assign w8802 = w5042 & w8750;
assign w8803 = (~w4856 & ~w4884) | (~w4856 & w9109) | (~w4884 & w9109);
assign v3803 = ~(w4944 | w4965);
assign w8804 = v3803;
assign w8805 = w5258 & w5257;
assign w8806 = (~w5251 & ~w5253) | (~w5251 & w8875) | (~w5253 & w8875);
assign v3804 = ~(w5038 | w5036);
assign w8807 = v3804;
assign v3805 = ~(w5186 | w5184);
assign w8808 = v3805;
assign v3806 = ~(w5048 | w5046);
assign w8809 = v3806;
assign w8810 = w5023 & ~w5026;
assign w8811 = w5153 & ~w5142;
assign v3807 = ~(w5284 | w5302);
assign w8812 = v3807;
assign w8813 = w5433 & ~w5422;
assign v3808 = ~(w5344 | w5347);
assign w8814 = v3808;
assign v3809 = ~(w5298 | w5296);
assign w8815 = v3809;
assign v3810 = ~(w5402 | w5400);
assign w8816 = v3810;
assign v3811 = ~(w5392 | w5390);
assign w8817 = v3811;
assign v3812 = ~(w5649 | w5647);
assign w8818 = v3812;
assign v3813 = ~(w5684 | w5682);
assign w8819 = v3813;
assign v3814 = ~(w5866 | w5864);
assign w8820 = v3814;
assign v3815 = ~(w5876 | w5874);
assign w8821 = v3815;
assign v3816 = ~(w5738 | w5736);
assign w8822 = v3816;
assign w8823 = w5722 & ~w5725;
assign v3817 = ~(w5858 | w5880);
assign w8824 = v3817;
assign v3818 = ~(w5755 | w5753);
assign w8825 = v3818;
assign v3819 = ~(w5906 | w5904);
assign w8826 = v3819;
assign w8827 = (~w5741 & ~w5758) | (~w5741 & w9110) | (~w5758 & w9110);
assign v3820 = ~(w6053 | w6051);
assign w8828 = v3820;
assign v3821 = ~(w5992 | w6004);
assign w8829 = v3821;
assign v3822 = ~(w6045 | w6057);
assign w8830 = v3822;
assign v3823 = ~(w6099 | w6097);
assign w8831 = v3823;
assign w8832 = (w6328 & w6128) | (w6328 & w8876) | (w6128 & w8876);
assign w8833 = (~w6209 & ~w6230) | (~w6209 & w9111) | (~w6230 & w9111);
assign w8834 = (~w6419 & ~w6430) | (~w6419 & w9112) | (~w6430 & w9112);
assign w8835 = w6462 & ~w6451;
assign w8836 = w6416 & ~w6405;
assign w8837 = w6432 & w6425;
assign w8838 = w6432 & ~w8776;
assign v3824 = ~(w6432 | w6425);
assign w8839 = v3824;
assign w8840 = ~w6432 & w8776;
assign v3825 = ~(w6368 | w6366);
assign w8841 = v3825;
assign w8842 = (~w6353 & ~w6371) | (~w6353 & w9113) | (~w6371 & w9113);
assign w8843 = (~w6672 & ~w6682) | (~w6672 & w9218) | (~w6682 & w9218);
assign w8844 = w6628 & ~w6617;
assign w8845 = w6584 & ~w6573;
assign v3826 = ~(w6679 | w6677);
assign w8846 = v3826;
assign v3827 = ~(w6669 | w6667);
assign w8847 = v3827;
assign w8848 = (~w6538 & ~w6556) | (~w6538 & w9114) | (~w6556 & w9114);
assign w8849 = (w6872 & w6128) | (w6872 & w9115) | (w6128 & w9115);
assign v3828 = ~(w6658 | w6801);
assign w8850 = v3828;
assign w8851 = w6768 & ~w6757;
assign v3829 = ~(w6728 | w6726);
assign w8852 = v3829;
assign w8853 = (~w6722 & ~w6740) | (~w6722 & w9116) | (~w6740 & w9116);
assign w8854 = ~w6870 & w7030;
assign v3830 = ~(w7012 | w7022);
assign w8855 = v3830;
assign w8856 = w6973 & ~w6962;
assign v3831 = ~(w7018 | w7016);
assign w8857 = v3831;
assign v3832 = ~(w6899 | w6919);
assign w8858 = v3832;
assign w8859 = w7128 & ~w7117;
assign v3833 = ~(w8779 | w7722);
assign w8860 = v3833;
assign v3834 = ~(w8284 | w8780);
assign w8861 = v3834;
assign v3835 = ~(w8284 | w8781);
assign w8862 = v3835;
assign w8863 = w8412 & ~w8780;
assign w8864 = w8412 & ~w8781;
assign w8865 = w8528 & ~w8780;
assign w8866 = w8528 & ~w8781;
assign v3836 = ~(w3162 | w3099);
assign w8867 = v3836;
assign v3837 = ~(w3449 | w3386);
assign w8868 = v3837;
assign w8869 = ~w3694 & w3631;
assign v3838 = ~(w3902 | w3838);
assign w8870 = v3838;
assign w8871 = w4117 & w4092;
assign v3839 = ~(w4369 | w4344);
assign w8872 = v3839;
assign w8873 = w4480 & w4472;
assign w8874 = w4734 & w4726;
assign w8875 = w5014 & ~w5251;
assign w8876 = ~w6131 & w6328;
assign w8877 = w5260 & w8784;
assign w8878 = w5260 & w8785;
assign v3840 = ~(w6326 | w6328);
assign w8879 = v3840;
assign v3841 = ~(w6326 | w8832);
assign w8880 = v3841;
assign v3842 = ~(w6268 | w6266);
assign w8881 = v3842;
assign w8882 = w6144 & ~w6155;
assign v3843 = ~(w6271 | w6274);
assign w8883 = v3843;
assign w8884 = w6082 & w6291;
assign v3844 = ~(w6495 | w6505);
assign w8885 = v3844;
assign w8886 = w6512 & ~w6511;
assign w8887 = (~w6587 & ~w6598) | (~w6587 & w9117) | (~w6598 & w9117);
assign v3845 = ~(w6595 | w6593);
assign w8888 = v3845;
assign v3846 = ~(w6638 | w6636);
assign w8889 = v3846;
assign v3847 = ~(w6553 | w6551);
assign w8890 = v3847;
assign w8891 = w6867 & w6869;
assign v3848 = ~(w6779 | w6777);
assign w8892 = v3848;
assign v3849 = ~(w6787 | w6785);
assign w8893 = v3849;
assign v3850 = ~(w6797 | w6795);
assign w8894 = v3850;
assign v3851 = ~(w6737 | w6735);
assign w8895 = v3851;
assign v3852 = ~(w6841 | w6839);
assign w8896 = v3852;
assign v3853 = ~(w7028 | w7030);
assign w8897 = v3853;
assign w8898 = (~w7028 & w6870) | (~w7028 & w8897) | (w6870 & w8897);
assign v3854 = ~(w6983 | w6981);
assign w8899 = v3854;
assign v3855 = ~(w6934 | w6946);
assign w8900 = v3855;
assign v3856 = ~(w6942 | w6940);
assign w8901 = v3856;
assign v3857 = ~(w7093 | w7091);
assign w8902 = v3857;
assign v3858 = ~(w7138 | w7136);
assign w8903 = v3858;
assign w8904 = w7103 & ~w7097;
assign v3859 = ~(w7236 | w7234);
assign w8905 = v3859;
assign w8906 = w7188 & ~w7101;
assign v3860 = ~(w7464 | w7468);
assign w8907 = v3860;
assign w8908 = (~w7722 & w8860) | (~w7722 & w8777) | (w8860 & w8777);
assign w8909 = (~w7722 & w8860) | (~w7722 & w8778) | (w8860 & w8778);
assign v3861 = ~(w7949 | w8657);
assign w8910 = v3861;
assign w8911 = (w7474 & w9219) | (w7474 & w8910) | (w9219 & w8910);
assign w8912 = w8350 & ~w8861;
assign w8913 = w8350 & ~w8862;
assign v3862 = ~(w8411 | w8863);
assign w8914 = v3862;
assign v3863 = ~(w8411 | w8864);
assign w8915 = v3863;
assign v3864 = ~(w8530 | w8865);
assign w8916 = v3864;
assign v3865 = ~(w8530 | w8866);
assign w8917 = v3865;
assign w8918 = w2906 & ~w2895;
assign v3866 = ~(w2966 | w2968);
assign w8919 = v3866;
assign v3867 = ~(w3216 | w2925);
assign w8920 = v3867;
assign w8921 = ~w3216 & w8723;
assign w8922 = w3293 & w3126;
assign w8923 = (w3293 & w3128) | (w3293 & w8922) | (w3128 & w8922);
assign v3868 = ~(w3293 | w3126);
assign w8924 = v3868;
assign w8925 = ~w3128 & w8924;
assign w8926 = w3159 & ~w3148;
assign v3869 = ~(w3046 | w3048);
assign w8927 = v3869;
assign w8928 = w3446 & ~w3435;
assign v3870 = ~(w3354 | w3356);
assign w8929 = v3870;
assign v3871 = ~(w3318 | w3316);
assign w8930 = v3871;
assign v3872 = ~(w3536 | w3534);
assign w8931 = v3872;
assign v3873 = ~(w3597 | w3599);
assign w8932 = v3873;
assign w8933 = w3940 & w3658;
assign w8934 = (w3940 & w3660) | (w3940 & w8933) | (w3660 & w8933);
assign v3874 = ~(w3940 | w3658);
assign w8935 = v3874;
assign w8936 = ~w3660 & w8935;
assign v3875 = ~(w3555 | w3553);
assign w8937 = v3875;
assign w8938 = w3556 & ~w3559;
assign v3876 = ~(w3735 | w3733);
assign w8939 = v3876;
assign w8940 = (~w3567 & ~w3539) | (~w3567 & w9118) | (~w3539 & w9118);
assign v3877 = ~(w3973 | w3972);
assign w8941 = v3877;
assign v3878 = ~(w3946 | w3944);
assign w8942 = v3878;
assign v3879 = ~(w3947 | w3950);
assign w8943 = v3879;
assign v3880 = ~(w3924 | w3922);
assign w8944 = v3880;
assign w8945 = (w3957 & ~w3976) | (w3957 & w9119) | (~w3976 & w9119);
assign v3881 = ~(w4232 | w4230);
assign w8946 = v3881;
assign v3882 = ~(w4064 | w4066);
assign w8947 = v3882;
assign v3883 = ~(w4187 | w4190);
assign w8948 = v3883;
assign w8949 = w4487 & w8740;
assign w8950 = w4487 & ~w4146;
assign v3884 = ~(w4487 | w8740);
assign w8951 = v3884;
assign w8952 = ~w4487 & w4146;
assign v3885 = ~(w4177 | w4175);
assign w8953 = v3885;
assign w8954 = (w4217 & w4235) | (w4217 & w9120) | (w4235 & w9120);
assign w8955 = w4519 & w8784;
assign w8956 = ~w8783 & w9121;
assign w8957 = ~w4477 & w8788;
assign v3886 = ~(w4377 | w4375);
assign w8958 = v3886;
assign w8959 = w5000 & ~w8800;
assign w8960 = w5000 & w4745;
assign w8961 = (~w4997 & ~w5006) | (~w4997 & w9122) | (~w5006 & w9122);
assign v3887 = ~(w5003 | w5001);
assign w8962 = v3887;
assign v3888 = ~(w4976 | w4974);
assign w8963 = v3888;
assign w8964 = w5263 & ~w8878;
assign w8965 = w5263 & ~w8877;
assign w8966 = w5162 & ~w5269;
assign w8967 = ~w5162 & w5269;
assign v3889 = ~(w5167 | w5190);
assign w8968 = v3889;
assign v3890 = ~(w5077 | w5080);
assign w8969 = v3890;
assign v3891 = ~(w5064 | w5455);
assign w8970 = v3891;
assign w8971 = w5064 & w5455;
assign w8972 = w5242 & w5467;
assign v3892 = ~(w5242 | w5467);
assign w8973 = v3892;
assign v3893 = ~(w5051 | w5070);
assign w8974 = v3893;
assign w8975 = w5287 & ~w5640;
assign w8976 = ~w5287 & w5640;
assign v3894 = ~(w5381 | w5379);
assign w8977 = v3894;
assign v3895 = ~(w5272 | w5270);
assign w8978 = v3895;
assign w8979 = w5273 & ~w5276;
assign v3896 = ~(w5384 | w5406);
assign w8980 = v3896;
assign w8981 = w8756 & w5706;
assign w8982 = (w5706 & w8756) | (w5706 & w5486) | (w8756 & w5486);
assign v3897 = ~(w5572 | w5594);
assign w8983 = v3897;
assign w8984 = w5499 & ~w5698;
assign v3898 = ~(w5744 | w6090);
assign w8985 = v3898;
assign w8986 = w5744 & w6090;
assign v3899 = ~(w6102 | w6113);
assign w8987 = v3899;
assign v3900 = ~(w5969 | w5972);
assign w8988 = v3900;
assign w8989 = w6347 & ~w6266;
assign w8990 = w6347 & w8881;
assign v3901 = ~(w6472 | w6470);
assign w8991 = v3901;
assign v3902 = ~(w6475 | w6478);
assign w8992 = v3902;
assign v3903 = ~(w6396 | w6399);
assign w8993 = v3903;
assign w8994 = (~w6511 & w8886) | (~w6511 & ~w8879) | (w8886 & ~w8879);
assign w8995 = (w8832 & w9123) | (w8832 & w9124) | (w9123 & w9124);
assign v3904 = ~(w6564 | w6567);
assign w8996 = v3904;
assign v3905 = ~(w6844 | w6854);
assign w8997 = v3905;
assign v3906 = ~(w6748 | w6751);
assign w8998 = v3906;
assign w8999 = w6977 & ~w6795;
assign w9000 = w6977 & w8894;
assign w9001 = (w8897 & w8898) | (w8897 & ~w6872) | (w8898 & ~w6872);
assign w9002 = (w8897 & w8898) | (w8897 & ~w8849) | (w8898 & ~w8849);
assign v3907 = ~(w6953 | w6956);
assign w9003 = v3907;
assign w9004 = w7132 & ~w6940;
assign w9005 = w7132 & w8901;
assign w9006 = w6913 & w7154;
assign v3908 = ~(w6913 | w7154);
assign w9007 = v3908;
assign v3909 = ~(w7163 | w7174);
assign w9008 = v3909;
assign w9009 = w7230 & ~w7091;
assign w9010 = w7230 & w8902;
assign w9011 = w7063 & w7248;
assign v3910 = ~(w7063 | w7248);
assign w9012 = v3910;
assign v3911 = ~(w7170 | w7168);
assign w9013 = v3911;
assign v3912 = ~(w7160 | w7158);
assign w9014 = v3912;
assign v3913 = ~(w7060 | w7080);
assign w9015 = v3913;
assign w9016 = w7226 & ~w7215;
assign w9017 = w7282 & w7386;
assign v3914 = ~(w7282 | w7386);
assign w9018 = v3914;
assign w9019 = w7231 & ~w7101;
assign w9020 = w7231 & w8906;
assign v3915 = ~(w7254 | w7252);
assign w9021 = v3915;
assign v3916 = ~(w7279 | w7299);
assign w9022 = v3916;
assign v3917 = ~(w7431 | w7429);
assign w9023 = v3917;
assign v3918 = ~(w7392 | w7390);
assign w9024 = v3918;
assign v3919 = ~(w7416 | w7435);
assign w9025 = v3919;
assign v3920 = ~(w7837 | w7835);
assign w9026 = v3920;
assign v3921 = ~(w8046 | w8044);
assign w9027 = v3921;
assign v3922 = ~(w8213 | w9077);
assign w9028 = v3922;
assign w9029 = (w7474 & w9220) | (w7474 & w9028) | (w9220 & w9028);
assign w9030 = (w8861 & w8862) | (w8861 & ~w8657) | (w8862 & ~w8657);
assign w9031 = (w7474 & w9221) | (w7474 & w9030) | (w9221 & w9030);
assign v3923 = ~(w8348 | w8912);
assign w9032 = v3923;
assign v3924 = ~(w8348 | w8913);
assign w9033 = v3924;
assign w9034 = w8453 & w8914;
assign w9035 = w8453 & w8915;
assign w9036 = w8524 & w8916;
assign w9037 = w8524 & w8917;
assign w9038 = w8559 & w8916;
assign w9039 = w8559 & w8917;
assign v3925 = ~(w4517 | w8955);
assign w9040 = v3925;
assign w9041 = (~w4517 & ~w9121) | (~w4517 & w9222) | (~w9121 & w9222);
assign v3926 = ~(w4740 | w4738);
assign w9042 = v3926;
assign v3927 = ~(w4643 | w4641);
assign w9043 = v3927;
assign v3928 = ~(w4693 | w4695);
assign w9044 = v3928;
assign w9045 = w4712 & ~w4715;
assign v3929 = ~(w4677 | w4675);
assign w9046 = v3929;
assign w9047 = w4770 & ~w4769;
assign v3930 = ~(w4985 | w4983);
assign w9048 = v3930;
assign v3931 = ~(w5223 | w4974);
assign w9049 = v3931;
assign w9050 = ~w5223 & w8963;
assign v3932 = ~(w4970 | w4990);
assign w9051 = v3932;
assign v3933 = ~(w5057 | w5055);
assign w9052 = v3933;
assign w9053 = ~w5066 & w8970;
assign v3934 = ~(w5492 | w5462);
assign w9054 = v3934;
assign v3935 = ~(w5705 | w8982);
assign w9055 = v3935;
assign v3936 = ~(w5705 | w8981);
assign w9056 = v3936;
assign v3937 = ~(w6691 | w6689);
assign w9057 = v3937;
assign w9058 = w7181 & ~w7180;
assign v3938 = ~(w7195 | w7193);
assign w9059 = v3938;
assign v3939 = ~(w7443 | w7454);
assign w9060 = v3939;
assign v3940 = ~(w7344 | w7342);
assign w9061 = v3940;
assign v3941 = ~(w7352 | w7350);
assign w9062 = v3941;
assign w9063 = w7474 & ~w7460;
assign w9064 = (~w7460 & w9063) | (~w7460 & w7470) | (w9063 & w7470);
assign v3942 = ~(w7600 | w8777);
assign w9065 = v3942;
assign w9066 = (w7474 & w9223) | (w7474 & w9065) | (w9223 & w9065);
assign v3943 = ~(w7583 | w7594);
assign w9067 = v3943;
assign v3944 = ~(w7528 | w7578);
assign w9068 = v3944;
assign v3945 = ~(w7705 | w7716);
assign w9069 = v3945;
assign v3946 = ~(w7941 | w7835);
assign w9070 = v3946;
assign w9071 = ~w7941 & w9026;
assign w9072 = w7941 & w7835;
assign w9073 = w7941 & ~w9026;
assign v3947 = ~(w7948 | w7940);
assign w9074 = v3947;
assign w9075 = w8133 & w8044;
assign w9076 = w8133 & ~w9027;
assign w9077 = (~w8140 & w8659) | (~w8140 & w8657) | (w8659 & w8657);
assign w9078 = (~w8140 & w8659) | (~w8140 & w8658) | (w8659 & w8658);
assign w9079 = w8214 & ~w8286;
assign w9080 = w8404 & w9032;
assign w9081 = w8404 & w9033;
assign v3948 = ~(w8404 | w9032);
assign w9082 = v3948;
assign v3949 = ~(w8404 | w9033);
assign w9083 = v3949;
assign w9084 = (w8914 & w8915) | (w8914 & w8657) | (w8915 & w8657);
assign w9085 = ~w8408 & w8455;
assign w9086 = ~w8491 & w9034;
assign w9087 = ~w8491 & w9035;
assign w9088 = w8495 & ~w9034;
assign w9089 = w8495 & ~w9035;
assign w9090 = (w8916 & w8917) | (w8916 & w8657) | (w8917 & w8657);
assign w9091 = w8557 & ~w9036;
assign w9092 = w8557 & ~w9037;
assign v3950 = ~(w8570 | w9038);
assign w9093 = v3950;
assign v3951 = ~(w8570 | w9039);
assign w9094 = v3951;
assign w9095 = w8566 & w9038;
assign w9096 = w8566 & w9039;
assign w9097 = w8574 & ~w9038;
assign w9098 = w8574 & ~w9039;
assign v3952 = ~(w5952 | w5944);
assign w9099 = v3952;
assign v3953 = ~(w6169 | w6160);
assign w9100 = v3953;
assign v3954 = ~(w8138 | w8140);
assign w9101 = v3954;
assign w9102 = w5156 & w5131;
assign v3955 = ~(w5436 | w5373);
assign w9103 = v3955;
assign w9104 = w5678 & w5670;
assign v3956 = ~(w5624 | w5561);
assign w9105 = v3956;
assign w9106 = w5711 & w5909;
assign v3957 = ~(w5711 | w5909);
assign w9107 = v3957;
assign w9108 = w4631 & w4606;
assign v3958 = ~(w4909 | w4856);
assign w9109 = v3958;
assign v3959 = ~(w5749 | w5741);
assign w9110 = v3959;
assign v3960 = ~(w6219 | w6209);
assign w9111 = v3960;
assign w9112 = w6434 & ~w6419;
assign v3961 = ~(w6362 | w6353);
assign w9113 = v3961;
assign v3962 = ~(w6547 | w6538);
assign w9114 = v3962;
assign w9115 = ~w6131 & w6872;
assign v3963 = ~(w6731 | w6722);
assign w9116 = v3963;
assign w9117 = w6600 & ~w6587;
assign v3964 = ~(w3530 | w3567);
assign w9118 = v3964;
assign w9119 = w3967 & w3957;
assign w9120 = w4226 & w4217;
assign w9121 = ~w4262 & w4519;
assign w9122 = w4998 & ~w4997;
assign w9123 = w8886 | ~w6511;
assign w9124 = (~w6511 & w8886) | (~w6511 & w6326) | (w8886 & w6326);
assign w9125 = w2501 & ~w2490;
assign v3965 = ~(w2996 | w2994);
assign w9126 = v3965;
assign v3966 = ~(w2917 | w2915);
assign w9127 = v3966;
assign v3967 = ~(w3107 | w3105);
assign w9128 = v3967;
assign v3968 = ~(w3118 | w3116);
assign w9129 = v3968;
assign v3969 = ~(w3214 | w3212);
assign w9130 = v3969;
assign w9131 = w3215 & ~w3217;
assign v3970 = ~(w3110 | w3132);
assign w9132 = v3970;
assign w9133 = w3318 & ~w8726;
assign w9134 = w3318 & w3163;
assign v3971 = ~(w3291 | w3289);
assign w9135 = v3971;
assign w9136 = w3292 & ~w3294;
assign v3972 = ~(w3397 | w3419);
assign w9137 = v3972;
assign w9138 = w3536 & ~w8727;
assign w9139 = w3536 & w3450;
assign v3973 = ~(w3394 | w3392);
assign w9140 = v3973;
assign v3974 = ~(w3639 | w3637);
assign w9141 = v3974;
assign v3975 = ~(w3642 | w3664);
assign w9142 = v3975;
assign v3976 = ~(w3973 | w8731);
assign w9143 = v3976;
assign w9144 = ~w3973 & w3695;
assign w9145 = w3962 & w4167;
assign v3977 = ~(w3962 | w4167);
assign w9146 = v3977;
assign v3978 = ~(w3849 | w3872);
assign w9147 = v3978;
assign w9148 = w4232 & ~w8739;
assign w9149 = w4232 & w3903;
assign v3979 = ~(w3992 | w3990);
assign w9150 = v3979;
assign w9151 = w4221 & w4422;
assign v3980 = ~(w4221 | w4422);
assign w9152 = v3980;
assign v3981 = ~(w4136 | w4134);
assign w9153 = v3981;
assign v3982 = ~(w4125 | w4123);
assign w9154 = v3982;
assign v3983 = ~(w4203 | w4201);
assign w9155 = v3983;
assign v3984 = ~(w4184 | w4182);
assign w9156 = v3984;
assign v3985 = ~(w4037 | w4087);
assign w9157 = v3985;
assign v3986 = ~(w4251 | w4249);
assign w9158 = v3986;
assign v3987 = ~(w4244 | w4255);
assign w9159 = v3987;
assign v3988 = ~(w4505 | w4503);
assign w9160 = v3988;
assign w9161 = (~w4769 & w9047) | (~w4769 & ~w9040) | (w9047 & ~w9040);
assign w9162 = (~w4769 & w9047) | (~w4769 & ~w9041) | (w9047 & ~w9041);
assign v3989 = ~(w4927 | w4925);
assign w9163 = v3989;
assign w9164 = w5684 & ~w8752;
assign w9165 = w5684 & w5437;
assign w9166 = w5755 & ~w8763;
assign w9167 = w5755 & w5625;
assign w9168 = w5916 & ~w9056;
assign w9169 = w5916 & ~w9055;
assign v3990 = ~(w5717 | w5715);
assign w9170 = v3990;
assign v3991 = ~(w6109 | w6107);
assign w9171 = v3991;
assign w9172 = w6313 & ~w8648;
assign w9173 = w6313 & w5962;
assign v3992 = ~(w6498 | w8655);
assign w9174 = v3992;
assign w9175 = ~w6498 & w6179;
assign v3993 = ~(w6501 | w6499);
assign w9176 = v3993;
assign w9177 = (~w6689 & w9057) | (~w6689 & ~w8994) | (w9057 & ~w8994);
assign w9178 = (~w8832 & w9224) | (~w8832 & w9225) | (w9224 & w9225);
assign w9179 = w6847 & ~w8848;
assign w9180 = w6847 & w6557;
assign w9181 = w8849 & w6872;
assign w9182 = (w6872 & w8849) | (w6872 & w6136) | (w8849 & w6136);
assign v3994 = ~(w6850 | w6848);
assign w9183 = v3994;
assign w9184 = w7015 & ~w8853;
assign w9185 = w7015 & w6741;
assign w9186 = (w8849 & w9226) | (w8849 & w9227) | (w9226 & w9227);
assign w9187 = (~w7180 & w9058) | (~w7180 & ~w9001) | (w9058 & ~w9001);
assign v3995 = ~(w7470 | w7474);
assign w9188 = v3995;
assign w9189 = w7461 & ~w7602;
assign w9190 = (w8777 & ~w7474) | (w8777 & w9228) | (~w7474 & w9228);
assign w9191 = (w8777 & w8778) | (w8777 & ~w7470) | (w8778 & ~w7470);
assign v3996 = ~(w7837 | w8908);
assign w9192 = v3996;
assign v3997 = ~(w7837 | w8909);
assign w9193 = v3997;
assign w9194 = ~w7941 & w9318;
assign w9195 = (w9070 & w9071) | (w9070 & ~w8909) | (w9071 & ~w8909);
assign w9196 = (w8657 & ~w7474) | (w8657 & w9229) | (~w7474 & w9229);
assign w9197 = (w8657 & w8658) | (w8657 & ~w7470) | (w8658 & ~w7470);
assign w9198 = ~w8046 & w8910;
assign w9199 = ~w8046 & w8911;
assign w9200 = ~w8133 & w9319;
assign w9201 = ~w8133 & w9320;
assign w9202 = w8215 & ~w9077;
assign w9203 = w8215 & ~w9078;
assign w9204 = (~w8286 & w9079) | (~w8286 & w9028) | (w9079 & w9028);
assign w9205 = (~w8286 & w9079) | (~w8286 & w9029) | (w9079 & w9029);
assign w9206 = ~w8350 & w9030;
assign w9207 = ~w8350 & w9031;
assign w9208 = (w8658 & w9230) | (w8658 & w9231) | (w9230 & w9231);
assign w9209 = ~w8453 & w9084;
assign w9210 = (w8455 & w9085) | (w8455 & w9030) | (w9085 & w9030);
assign w9211 = (w8455 & w9085) | (w8455 & w9031) | (w9085 & w9031);
assign w9212 = (~w8658 & w9232) | (~w8658 & w9233) | (w9232 & w9233);
assign v3998 = ~(w8524 | w9090);
assign w9213 = v3998;
assign w9214 = w1072 & ~w1067;
assign w9215 = ~w1072 & w1067;
assign w9216 = w1762 & w1883;
assign w9217 = w5847 & w5822;
assign w9218 = w6673 & ~w6672;
assign v3999 = ~(w7949 | w7952);
assign w9219 = v3999;
assign w9220 = ~w8213 & w9321;
assign w9221 = (w8861 & w8862) | (w8861 & ~w7952) | (w8862 & ~w7952);
assign w9222 = w8783 & ~w4517;
assign v4000 = ~(w7600 | w7604);
assign w9223 = v4000;
assign w9224 = (~w6689 & w9057) | (~w6689 & ~w9124) | (w9057 & ~w9124);
assign w9225 = (~w6689 & w9057) | (~w6689 & ~w9123) | (w9057 & ~w9123);
assign w9226 = (~w7180 & w9058) | (~w7180 & ~w8897) | (w9058 & ~w8897);
assign w9227 = (~w7180 & w9058) | (~w7180 & ~w8898) | (w9058 & ~w8898);
assign w9228 = w8777 | w7604;
assign w9229 = w8657 | w7952;
assign w9230 = ~w8453 & w8914;
assign w9231 = ~w8453 & w8915;
assign v4001 = ~(w8524 | w8916);
assign w9232 = v4001;
assign v4002 = ~(w8524 | w8917);
assign w9233 = v4002;
assign w9234 = w631 & ~w630;
assign v4003 = ~(w654 | w653);
assign w9235 = v4003;
assign v4004 = ~(w749 | w751);
assign w9236 = v4004;
assign v4005 = ~(w744 | w742);
assign w9237 = v4005;
assign v4006 = ~(w905 | w903);
assign w9238 = v4006;
assign v4007 = ~(w838 | w860);
assign w9239 = v4007;
assign v4008 = ~(w856 | w854);
assign w9240 = v4008;
assign v4009 = ~(w1028 | w1026);
assign w9241 = v4009;
assign w9242 = w1020 & ~w1045;
assign v4010 = ~(w1161 | w1159);
assign w9243 = v4010;
assign v4011 = ~(w1182 | w1180);
assign w9244 = v4011;
assign w9245 = w1143 & ~w1166;
assign w9246 = w1174 & ~w1186;
assign v4012 = ~(w1233 | w1231);
assign w9247 = v4012;
assign w9248 = w1223 & ~w1211;
assign v4013 = ~(w1312 | w1301);
assign w9249 = v4013;
assign v4014 = ~(w1331 | w1330);
assign w9250 = v4014;
assign w9251 = w1416 & ~w1623;
assign w9252 = w1623 & ~w1417;
assign v4015 = ~(w1501 | w1503);
assign w9253 = v4015;
assign v4016 = ~(w1871 | w1754);
assign w9254 = v4016;
assign w9255 = ~w1871 & w8698;
assign w9256 = w1781 & w1930;
assign v4017 = ~(w1781 | w1930);
assign w9257 = v4017;
assign v4018 = ~(w1825 | w1823);
assign w9258 = v4018;
assign v4019 = ~(w1990 | w2002);
assign w9259 = v4019;
assign v4020 = ~(w1936 | w1934);
assign w9260 = v4020;
assign w9261 = w1961 & ~w1983;
assign v4021 = ~(w1996 | w1994);
assign w9262 = v4021;
assign w9263 = w1976 & w2129;
assign v4022 = ~(w1976 | w2129);
assign w9264 = v4022;
assign w9265 = w2137 & ~w8706;
assign w9266 = w2137 & w1895;
assign v4023 = ~(w2008 | w1836);
assign w9267 = v4023;
assign w9268 = ~w2202 & w2403;
assign w9269 = w3752 & w2405;
assign w9270 = w8783 & ~w4261;
assign w9271 = (~w4261 & w8783) | (~w4261 & ~w3754) | (w8783 & ~w3754);
assign w9272 = w5015 & w9162;
assign w9273 = w5015 & w9161;
assign v4024 = ~(w5298 | w8751);
assign w9274 = v4024;
assign w9275 = ~w5298 & w5196;
assign v4025 = ~(w5486 | w5484);
assign w9276 = v4025;
assign v4026 = ~(w5494 | w5497);
assign w9277 = v4026;
assign v4027 = ~(w5914 | w9169);
assign w9278 = v4027;
assign v4028 = ~(w5914 | w9168);
assign w9279 = v4028;
assign v4029 = ~(w5958 | w8768);
assign w9280 = v4029;
assign w9281 = ~w5958 & w5886;
assign w9282 = w6870 & ~w7030;
assign w9283 = ~w7462 & w6137;
assign w9284 = (~w7602 & w9189) | (~w7602 & ~w6137) | (w9189 & ~w6137);
assign w9285 = (~w7602 & w9189) | (~w7602 & w9063) | (w9189 & w9063);
assign w9286 = w8288 & w9322;
assign w9287 = w8288 & w9323;
assign w9288 = w8350 & w9324;
assign w9289 = w8350 & w9325;
assign w9290 = (w9036 & w9037) | (w9036 & w6137) | (w9037 & w6137);
assign w9291 = (w9036 & w9037) | (w9036 & w9196) | (w9037 & w9196);
assign w9292 = (w9038 & w9039) | (w9038 & w6137) | (w9039 & w6137);
assign w9293 = (w9038 & w9039) | (w9038 & w9196) | (w9039 & w9196);
assign w9294 = (~w476 & w8584) | (~w476 & ~w480) | (w8584 & ~w480);
assign w9295 = (w1754 & ~w8698) | (w1754 & ~w1750) | (~w8698 & ~w1750);
assign w9296 = (w8706 & ~w1895) | (w8706 & ~w1896) | (~w1895 & ~w1896);
assign w9297 = (w2925 & ~w8723) | (w2925 & ~w2921) | (~w8723 & ~w2921);
assign w9298 = (w4261 & ~w8783) | (w4261 & ~w4010) | (~w8783 & ~w4010);
assign w9299 = (w8800 & ~w4745) | (w8800 & ~w4746) | (~w4745 & ~w4746);
assign w9300 = (w4932 & ~w8750) | (w4932 & ~w4928) | (~w8750 & ~w4928);
assign w9301 = (w4974 & ~w8963) | (w4974 & ~w4971) | (~w8963 & ~w4971);
assign w9302 = (~w6125 & ~w6129) | (~w6125 & ~w8770) | (~w6129 & ~w8770);
assign w9303 = (w8648 & ~w5962) | (w8648 & ~w5964) | (~w5962 & ~w5964);
assign w9304 = (w6266 & ~w8881) | (w6266 & ~w6262) | (~w8881 & ~w6262);
assign w9305 = (w8655 & ~w6179) | (w8655 & ~w6181) | (~w6179 & ~w6181);
assign w9306 = (w8848 & ~w6557) | (w8848 & ~w6559) | (~w6557 & ~w6559);
assign w9307 = (w6795 & ~w8894) | (w6795 & ~w6791) | (~w8894 & ~w6791);
assign w9308 = (w8853 & ~w6741) | (w8853 & ~w6743) | (~w6741 & ~w6743);
assign w9309 = (w6940 & ~w8901) | (w6940 & ~w6936) | (~w8901 & ~w6936);
assign w9310 = (w7091 & ~w8902) | (w7091 & ~w7087) | (~w8902 & ~w7087);
assign w9311 = (w7101 & ~w8906) | (w7101 & ~w7201) | (~w8906 & ~w7201);
assign w9312 = (~w7470 & ~w7462) | (~w7470 & w9283) | (~w7462 & w9283);
assign w9313 = (w7474 & ~w6137) | (w7474 & ~w9188) | (~w6137 & ~w9188);
assign w9314 = (~w9065 & ~w9066) | (~w9065 & ~w7471) | (~w9066 & ~w7471);
assign w9315 = (w8908 & w8909) | (w8908 & ~w7471) | (w8909 & ~w7471);
assign w9316 = (~w8910 & ~w8911) | (~w8910 & ~w7471) | (~w8911 & ~w7471);
assign w9317 = (w9077 & w9078) | (w9077 & ~w7471) | (w9078 & ~w7471);
assign w9318 = (~w7835 & w9026) | (~w7835 & ~w8908) | (w9026 & ~w8908);
assign w9319 = (~w8044 & w9027) | (~w8044 & w8910) | (w9027 & w8910);
assign w9320 = (~w8044 & w9027) | (~w8044 & w8911) | (w9027 & w8911);
assign w9321 = (w8140 & ~w8659) | (w8140 & ~w7952) | (~w8659 & ~w7952);
assign w9322 = (~w8660 & ~w8661) | (~w8660 & w6137) | (~w8661 & w6137);
assign w9323 = (~w8660 & ~w8661) | (~w8660 & w9196) | (~w8661 & w9196);
assign w9324 = (~w8861 & ~w8862) | (~w8861 & w6137) | (~w8862 & w6137);
assign w9325 = (~w8861 & ~w8862) | (~w8861 & w9196) | (~w8862 & w9196);
assign one = 1;
assign po00 = w3;// level 3
assign po01 = w14;// level 7
assign po02 = w34;// level 9
assign po03 = w61;// level 11
assign po04 = w97;// level 13
assign po05 = ~w150;// level 16
assign po06 = ~w205;// level 17
assign po07 = w267;// level 19
assign po08 = w337;// level 19
assign po09 = ~w412;// level 21
assign po10 = w501;// level 22
assign po11 = ~w593;// level 24
assign po12 = ~w698;// level 25
assign po13 = w812;// level 27
assign po14 = w931;// level 28
assign po15 = ~w1061;// level 28
assign po16 = w1200;// level 30
assign po17 = ~w1344;// level 32
assign po18 = w1498;// level 34
assign po19 = w1661;// level 36
assign po20 = w1840;// level 31
assign po21 = ~w2014;// level 33
assign po22 = w2206;// level 35
assign po23 = ~w2402;// level 34
assign po24 = w2608;// level 34
assign po25 = w2819;// level 36
assign po26 = w3042;// level 38
assign po27 = ~w3268;// level 40
assign po28 = w3509;// level 37
assign po29 = w3751;// level 39
assign po30 = w4008;// level 38
assign po31 = ~w4267;// level 39
assign po32 = w4524;// level 40
assign po33 = w4774;// level 39
assign po34 = w5019;// level 40
assign po35 = w5256;// level 41
assign po36 = w5489;// level 40
assign po37 = w5709;// level 41
assign po38 = w5920;// level 41
assign po39 = w6124;// level 41
assign po40 = w6331;// level 40
assign po41 = w6516;// level 41
assign po42 = w6695;// level 41
assign po43 = w6865;// level 41
assign po44 = w7033;// level 41
assign po45 = ~w7185;// level 41
assign po46 = ~w7330;// level 41
assign po47 = ~w7477;// level 41
assign po48 = w7606;// level 40
assign po49 = ~w7727;// level 41
assign po50 = w7840;// level 41
assign po51 = w7944;// level 41
assign po52 = w8049;// level 41
assign po53 = w8136;// level 41
assign po54 = ~w8218;// level 41
assign po55 = w8290;// level 41
assign po56 = w8353;// level 41
assign po57 = ~w8407;// level 41
assign po58 = ~w8457;// level 41
assign po59 = ~w8497;// level 41
assign po60 = w8533;// level 41
assign po61 = w8561;// level 41
assign po62 = w8573;// level 41
assign po63 = ~w8576;// level 41
assign po64 = ~w8576;// level 41
endmodule
