//Written by the Majority Logic Package Thu Apr 30 23:48:42 2015
module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, v802, v803, v804, v805, v806, v807, v808, v809, v810, v811, v812, v813, v814, v815, v816, v817, v818, v819, v820, v821, v822, v823, v824, v825, v826, v827, v828, v829, v830, v831, v832, v833, v834, v835, v836, v837, v838, v839, v840, v841, v842, v843, v844, v845, v846, v847, v848, v849, v850, v851, v852, v853, v854, v855, v856, v857, v858, v859, v860, v861, v862, v863, v864, v865, v866, v867, v868, v869, v870, v871, v872, v873, v874, v875, v876, v877, v878, v879, v880, v881, v882, v883, v884, v885, v886, v887, v888, v889, v890, v891, v892, v893, v894, v895, v896, v897, v898, v899, v900, v901, v902, v903, v904, v905, v906, v907, v908, v909, v910, v911, v912, v913, v914, v915, v916, v917, v918, v919, v920, v921, v922, v923, v924, v925, v926, v927, v928, v929, v930, v931, v932, v933, v934, v935, v936, v937, v938, v939, v940, v941, v942, v943, v944, v945, v946, v947, v948, v949, v950, v951, v952, v953, v954, v955, v956, v957, v958, v959, v960, v961, v962, v963, v964, v965, v966, v967, v968, v969, v970, v971, v972, v973, v974, v975, v976, v977, v978, v979, v980, v981, v982, v983, v984, v985, v986, v987, v988, v989, v990, v991, v992, v993, v994, v995, v996, v997, v998, v999, v1000, v1001, v1002, v1003, v1004, v1005, v1006, v1007, v1008, v1009, v1010, v1011, v1012, v1013, v1014, v1015, v1016, v1017, v1018, v1019, v1020, v1021, v1022, v1023, v1024, v1025, v1026, v1027, v1028, v1029, v1030, v1031, v1032, v1033, v1034, v1035, v1036, v1037, v1038, v1039, v1040, v1041, v1042, v1043, v1044, v1045, v1046, v1047, v1048, v1049, v1050, v1051, v1052, v1053, v1054, v1055, v1056, v1057, v1058, v1059, v1060, v1061, v1062, v1063, v1064, v1065, v1066, v1067, v1068, v1069, v1070, v1071, v1072, v1073, v1074, v1075, v1076, v1077, v1078, v1079, v1080, v1081, v1082, v1083, v1084, v1085, v1086, v1087, v1088, v1089, v1090, v1091, v1092, v1093, v1094, v1095, v1096, v1097, v1098, v1099, v1100, v1101, v1102, v1103, v1104, v1105, v1106, v1107, v1108, v1109, v1110, v1111, v1112, v1113, v1114, v1115, v1116, v1117, v1118, v1119, v1120, v1121, v1122, v1123, v1124, v1125, v1126, v1127, v1128, v1129, v1130, v1131, v1132, v1133, v1134, v1135, v1136, v1137, v1138, v1139, v1140, v1141, v1142, v1143, v1144, v1145, v1146, v1147, v1148, v1149, v1150, v1151, v1152, v1153, v1154, v1155, v1156, v1157, v1158, v1159, v1160, v1161, v1162, v1163, v1164, v1165, v1166, v1167, v1168, v1169, v1170, v1171, v1172, v1173, v1174, v1175, v1176, v1177, v1178, v1179, v1180, v1181, v1182, v1183, v1184, v1185, v1186, v1187, v1188, v1189, v1190, v1191, v1192, v1193, v1194, v1195, v1196, v1197, v1198, v1199, v1200, v1201, v1202, v1203, v1204, v1205, v1206, v1207, v1208, v1209, v1210, v1211, v1212, v1213, v1214, v1215, v1216, v1217, v1218, v1219, v1220, v1221, v1222, v1223, v1224, v1225, v1226, v1227, v1228, v1229, v1230, v1231, v1232, v1233, v1234, v1235, v1236, v1237, v1238, v1239, v1240, v1241, v1242, v1243, v1244, v1245, v1246, v1247, v1248, v1249, v1250, v1251, v1252, v1253, v1254, v1255, v1256, v1257, v1258, v1259, v1260, v1261, v1262, v1263, v1264, v1265, v1266, v1267, v1268, v1269, v1270, v1271, v1272, v1273, v1274, v1275, v1276, v1277, v1278, v1279, v1280, v1281, v1282, v1283, v1284, v1285, v1286, v1287, v1288, v1289, v1290, v1291, v1292, v1293, v1294, v1295, v1296, v1297, v1298, v1299, v1300, v1301, v1302, v1303, v1304, v1305, v1306, v1307, v1308, v1309, v1310, v1311, v1312, v1313, v1314, v1315, v1316, v1317, v1318, v1319, v1320, v1321, v1322, v1323, v1324, v1325, v1326, v1327, v1328, v1329, v1330, v1331, v1332, v1333, v1334, v1335, v1336, v1337, v1338, v1339, v1340, v1341, v1342, v1343, v1344, v1345, v1346, v1347, v1348, v1349, v1350, v1351, v1352, v1353, v1354, v1355, v1356, v1357, v1358, v1359, v1360, v1361, v1362, v1363, v1364, v1365, v1366, v1367, v1368, v1369, v1370, v1371, v1372, v1373, v1374, v1375, v1376, v1377, v1378, v1379, v1380, v1381, v1382, v1383, v1384, v1385, v1386, v1387, v1388, v1389, v1390, v1391, v1392, v1393, v1394, v1395, v1396, v1397, v1398, v1399, v1400, v1401, v1402, v1403, v1404, v1405, v1406, v1407, v1408, v1409, v1410, v1411, v1412, v1413, v1414, v1415, v1416, v1417, v1418, v1419, v1420, v1421, v1422, v1423, v1424, v1425, v1426, v1427, v1428, v1429, v1430, v1431, v1432, v1433, v1434, v1435, v1436, v1437, v1438, v1439, v1440, v1441, v1442, v1443, v1444, v1445, v1446, v1447, v1448, v1449, v1450, v1451, v1452, v1453, v1454, v1455, v1456, v1457, v1458, v1459, v1460, v1461, v1462, v1463, v1464, v1465, v1466, v1467, v1468, v1469, v1470, v1471, v1472, v1473, v1474, v1475, v1476, v1477, v1478, v1479, v1480, v1481, v1482, v1483, v1484, v1485, v1486, v1487, v1488, v1489, v1490, v1491, v1492, v1493, v1494, v1495, v1496, v1497, v1498, v1499, v1500, v1501, v1502, v1503, v1504, v1505, v1506, v1507, v1508, v1509, v1510, v1511, v1512, v1513, v1514, v1515, v1516, v1517, v1518, v1519, v1520, v1521, v1522, v1523, v1524, v1525, v1526, v1527, v1528, v1529, v1530, v1531, v1532, v1533, v1534, v1535, v1536, v1537, v1538, v1539, v1540, v1541, v1542, v1543, v1544, v1545, v1546, v1547, v1548, v1549, v1550, v1551, v1552, v1553, v1554, v1555, v1556, v1557, v1558, v1559, v1560, v1561, v1562, v1563, v1564, v1565, v1566, v1567, v1568, v1569, v1570, v1571, v1572, v1573, v1574, v1575, v1576, v1577, v1578, v1579, v1580, v1581, v1582, v1583, v1584, v1585, v1586, v1587, v1588, v1589, v1590, v1591, v1592, v1593, v1594, v1595, v1596, v1597, v1598, v1599, v1600, v1601, v1602, v1603, v1604, v1605, v1606, v1607, v1608, v1609, v1610, v1611, v1612, v1613, v1614, v1615, v1616, v1617, v1618, v1619, v1620, v1621, v1622, v1623, v1624, v1625, v1626, v1627, v1628, v1629, v1630, v1631, v1632, v1633, v1634, v1635, v1636, v1637, v1638, v1639, v1640, v1641, v1642, v1643, v1644, v1645, v1646, v1647, v1648, v1649, v1650, v1651, v1652, v1653, v1654, v1655, v1656, v1657, v1658, v1659, v1660, v1661, v1662, v1663, v1664, v1665, v1666, v1667, v1668, v1669, v1670, v1671, v1672, v1673, v1674, v1675, v1676, v1677, v1678, v1679, v1680, v1681, v1682, v1683, v1684, v1685, v1686, v1687, v1688, v1689, v1690, v1691, v1692, v1693, v1694, v1695, v1696, v1697, v1698, v1699, v1700, v1701, v1702, v1703, v1704, v1705, v1706, v1707, v1708, v1709, v1710, v1711, v1712, v1713, v1714, v1715, v1716, v1717, v1718, v1719, v1720, v1721, v1722, v1723, v1724, v1725, v1726, v1727, v1728, v1729, v1730, v1731, v1732, v1733, v1734, v1735, v1736, v1737, v1738, v1739, v1740, v1741, v1742, v1743, v1744, v1745, v1746, v1747, v1748, v1749, v1750, v1751, v1752, v1753, v1754, v1755, v1756, v1757, v1758, v1759, v1760, v1761, v1762, v1763, v1764, v1765, v1766, v1767, v1768, v1769, v1770, v1771, v1772, v1773, v1774, v1775, v1776, v1777, v1778, v1779, v1780, v1781, v1782, v1783, v1784, v1785, v1786, v1787, v1788, v1789, v1790, v1791, v1792, v1793, v1794, v1795, v1796, v1797, v1798, v1799, v1800, v1801, v1802, v1803, v1804, v1805, v1806, v1807, v1808, v1809, v1810, v1811, v1812, v1813, v1814, v1815, v1816, v1817, v1818, v1819, v1820, v1821, v1822, v1823, v1824, v1825, v1826, v1827, v1828, v1829, v1830, v1831, v1832, v1833, v1834, v1835, v1836, v1837, v1838, v1839, v1840, v1841, v1842, v1843, v1844, v1845, v1846, v1847, v1848, v1849, v1850, v1851, v1852, v1853, v1854, v1855, v1856, v1857, v1858, v1859, v1860, v1861, v1862, v1863, v1864, v1865, v1866, v1867, v1868, v1869, v1870, v1871, v1872, v1873, v1874, v1875, v1876, v1877, v1878, v1879, v1880, v1881, v1882, v1883, v1884, v1885, v1886, v1887, v1888, v1889, v1890, v1891, v1892, v1893, v1894, v1895, v1896, v1897, v1898, v1899, v1900, v1901, v1902, v1903, v1904, v1905, v1906, v1907, v1908, v1909, v1910, v1911, v1912, v1913, v1914, v1915, v1916, v1917, v1918, v1919, v1920, v1921, v1922, v1923, v1924, v1925, v1926, v1927, v1928, v1929, v1930, v1931, v1932, v1933, v1934, v1935, v1936, v1937, v1938, v1939, v1940, v1941, v1942, v1943, v1944, v1945, v1946, v1947, v1948, v1949, v1950, v1951, v1952, v1953, v1954, v1955, v1956, v1957, v1958, v1959, v1960, v1961, v1962, v1963, v1964, v1965, v1966, v1967, v1968, v1969, v1970, v1971, v1972, v1973, v1974, v1975, v1976, v1977, v1978, v1979, v1980, v1981, v1982, v1983, v1984, v1985, v1986, v1987, v1988, v1989, v1990, v1991, v1992, v1993, v1994, v1995, v1996, v1997, v1998, v1999, v2000, v2001, v2002, v2003, v2004, v2005, v2006, v2007, v2008, v2009, v2010, v2011, v2012, v2013, v2014, v2015, v2016, v2017, v2018, v2019, v2020, v2021, v2022, v2023, v2024, v2025, v2026, v2027, v2028, v2029, v2030, v2031, v2032, v2033, v2034, v2035, v2036, v2037, v2038, v2039, v2040, v2041, v2042, v2043, v2044, v2045, v2046, v2047, v2048, v2049, v2050, v2051, v2052, v2053, v2054, v2055, v2056, v2057, v2058, v2059, v2060, v2061, v2062, v2063, v2064, v2065, v2066, v2067, v2068, v2069, v2070, v2071, v2072, v2073, v2074, v2075, v2076, v2077, v2078, v2079, v2080, v2081, v2082, v2083, v2084, v2085, v2086, v2087, v2088, v2089, v2090, v2091, v2092, v2093, v2094, v2095, v2096, v2097, v2098, v2099, v2100, v2101, v2102, v2103, v2104, v2105, v2106, v2107, v2108, v2109, v2110, v2111, v2112, v2113, v2114, v2115, v2116, v2117, v2118, v2119, v2120, v2121, v2122, v2123, v2124, v2125, v2126, v2127, v2128, v2129, v2130, v2131, v2132, v2133, v2134, v2135, v2136, v2137, v2138, v2139, v2140, v2141, v2142, v2143, v2144, v2145, v2146, v2147, v2148, v2149, v2150, v2151, v2152, v2153, v2154, v2155, v2156, v2157, v2158, v2159, v2160, v2161, v2162, v2163, v2164, v2165, v2166, v2167, v2168, v2169, v2170, v2171, v2172, v2173, v2174, v2175, v2176, v2177, v2178, v2179, v2180, v2181, v2182, v2183, v2184, v2185, v2186, v2187, v2188, v2189, v2190, v2191, v2192, v2193, v2194, v2195, v2196, v2197, v2198, v2199, v2200, v2201, v2202, v2203, v2204, v2205, v2206, v2207, v2208, v2209, v2210, v2211, v2212, v2213, v2214, v2215, v2216, v2217, v2218, v2219, v2220, v2221, v2222, v2223, v2224, v2225, v2226, v2227, v2228, v2229, v2230, v2231, v2232, v2233, v2234, v2235, v2236, v2237, v2238, v2239, v2240, v2241, v2242, v2243, v2244, v2245, v2246, v2247, v2248, v2249, v2250, v2251, v2252, v2253, v2254, v2255, v2256, v2257, v2258, v2259, v2260, v2261, v2262, v2263, v2264, v2265, v2266, v2267, v2268, v2269, v2270, v2271, v2272, v2273, v2274, v2275, v2276, v2277, v2278, v2279, v2280, v2281, v2282, v2283, v2284, v2285, v2286, v2287, v2288, v2289, v2290, v2291, v2292, v2293, v2294, v2295, v2296, v2297, v2298, v2299, v2300, v2301, v2302, v2303, v2304, v2305, v2306, v2307, v2308, v2309, v2310, v2311, v2312, v2313, v2314, v2315, v2316, v2317, v2318, v2319, v2320, v2321, v2322, v2323, v2324, v2325, v2326, v2327, v2328, v2329, v2330, v2331, v2332, v2333, v2334, v2335, v2336, v2337, v2338, v2339, v2340, v2341, v2342, v2343, v2344, v2345, v2346, v2347, v2348, v2349, v2350, v2351, v2352, v2353, v2354, v2355, v2356, v2357, v2358, v2359, v2360, v2361, v2362, v2363, v2364, v2365, v2366, v2367, v2368, v2369, v2370, v2371, v2372, v2373, v2374, v2375, v2376, v2377, v2378, v2379, v2380, v2381, v2382, v2383, v2384, v2385, v2386, v2387, v2388, v2389, v2390, v2391, v2392, v2393, v2394, v2395, v2396, v2397, v2398, v2399, v2400, v2401, v2402, v2403, v2404, v2405, v2406, v2407, v2408, v2409, v2410, v2411, v2412, v2413, v2414, v2415, v2416, v2417, v2418, v2419, v2420, v2421, v2422, v2423, v2424, v2425, v2426, v2427, v2428, v2429, v2430, v2431, v2432, v2433, v2434, v2435, v2436, v2437, v2438, v2439, v2440, v2441, v2442, v2443, v2444, v2445, v2446, v2447, v2448, v2449, v2450, v2451, v2452, v2453, v2454, v2455, v2456, v2457, v2458, v2459, v2460, v2461, v2462, v2463, v2464, v2465, v2466, v2467, v2468, v2469, v2470, v2471, v2472, v2473, v2474, v2475, v2476, v2477, v2478, v2479, v2480, v2481, v2482, v2483, v2484, v2485, v2486, v2487, v2488, v2489, v2490, v2491, v2492, v2493, v2494, v2495, v2496, v2497, v2498, v2499, v2500, v2501, v2502, v2503, v2504, v2505, v2506, v2507, v2508, v2509, v2510, v2511, v2512, v2513, v2514, v2515, v2516, v2517, v2518, v2519, v2520, v2521, v2522, v2523, v2524, v2525, v2526, v2527, v2528, v2529, v2530, v2531, v2532, v2533, v2534, v2535, v2536, v2537, v2538, v2539, v2540, v2541, v2542, v2543, v2544, v2545, v2546, v2547, v2548, v2549, v2550, v2551, v2552, v2553, v2554, v2555, v2556, v2557, v2558, v2559, v2560, v2561, v2562, v2563, v2564, v2565, v2566, v2567, v2568, v2569, v2570, v2571, v2572, v2573, v2574, v2575, v2576, v2577, v2578, v2579, v2580, v2581, v2582, v2583, v2584, v2585, v2586, v2587, v2588, v2589, v2590, v2591, v2592, v2593, v2594, v2595, v2596, v2597, v2598, v2599, v2600, v2601, v2602, v2603, v2604, v2605, v2606, v2607, v2608, v2609, v2610, v2611, v2612, v2613, v2614, v2615, v2616, v2617, v2618, v2619, v2620, v2621, v2622, v2623, v2624, v2625, v2626, v2627, v2628, v2629, v2630, v2631, v2632, v2633, v2634, v2635, v2636, v2637, v2638, v2639, v2640, v2641, v2642, v2643, v2644, v2645, v2646, v2647, v2648, v2649, v2650, v2651, v2652, v2653, v2654, v2655, v2656, v2657, v2658, v2659, v2660, v2661, v2662, v2663, v2664, v2665, v2666, v2667, v2668, v2669, v2670, v2671, v2672, v2673, v2674, v2675, v2676, v2677, v2678, v2679, v2680, v2681, v2682, v2683, v2684, v2685, v2686, v2687, v2688, v2689, v2690, v2691, v2692, v2693, v2694, v2695, v2696, v2697, v2698, v2699, v2700, v2701, v2702, v2703, v2704, v2705, v2706, v2707, v2708, v2709, v2710, v2711, v2712, v2713, v2714, v2715, v2716, v2717, v2718, v2719, v2720, v2721, v2722, v2723, v2724, v2725, v2726, v2727, v2728, v2729, v2730, v2731, v2732, v2733, v2734, v2735, v2736, v2737, v2738, v2739, v2740, v2741, v2742, v2743, v2744, v2745, v2746, v2747, v2748, v2749, v2750, v2751, v2752, v2753, v2754, v2755, v2756, v2757, v2758, v2759, v2760, v2761, v2762, v2763, v2764, v2765, v2766, v2767, v2768, v2769, v2770, v2771, v2772, v2773, v2774, v2775, v2776, v2777, v2778, v2779, v2780, v2781, v2782, v2783, v2784, v2785, v2786, v2787, v2788, v2789, v2790, v2791, v2792, v2793, v2794, v2795, v2796, v2797, v2798, v2799, v2800, v2801, v2802, v2803, v2804, v2805, v2806, v2807, v2808, v2809, v2810, v2811, v2812, v2813, v2814, v2815, v2816, v2817, v2818, v2819, v2820, v2821, v2822, v2823, v2824, v2825, v2826, v2827, v2828, v2829, v2830, v2831, v2832, v2833, v2834, v2835, v2836, v2837, v2838, v2839, v2840, v2841, v2842, v2843, v2844, v2845, v2846, v2847, v2848, v2849, v2850, v2851, v2852, v2853, v2854, v2855, v2856, v2857, v2858, v2859, v2860, v2861, v2862, v2863, v2864, v2865, v2866, v2867, v2868, v2869, v2870, v2871, v2872, v2873, v2874, v2875, v2876, v2877, v2878, v2879, v2880, v2881, v2882, v2883, v2884, v2885, v2886, v2887, v2888, v2889, v2890, v2891, v2892, v2893, v2894, v2895, v2896, v2897, v2898, v2899, v2900, v2901, v2902, v2903, v2904, v2905, v2906, v2907, v2908, v2909, v2910, v2911, v2912, v2913, v2914, v2915, v2916, v2917, v2918, v2919, v2920, v2921, v2922, v2923, v2924, v2925, v2926, v2927, v2928, v2929, v2930, v2931, v2932, v2933, v2934, v2935, v2936, v2937, v2938, v2939, v2940, v2941, v2942, v2943, v2944, v2945, v2946, v2947, v2948, v2949, v2950, v2951, v2952, v2953, v2954, v2955, v2956, v2957, v2958, v2959, v2960, v2961, v2962, v2963, v2964, v2965, v2966, v2967, v2968, v2969, v2970, v2971, v2972, v2973, v2974, v2975, v2976, v2977, v2978, v2979, v2980, v2981, v2982, v2983, v2984, v2985, v2986, v2987, v2988, v2989, v2990, v2991, v2992, v2993, v2994, v2995, v2996, v2997, v2998, v2999, v3000, v3001, v3002, v3003, v3004, v3005, v3006, v3007, v3008, v3009, v3010, v3011, v3012, v3013, v3014, v3015, v3016, v3017, v3018, v3019, v3020, v3021, v3022, v3023, v3024, v3025, v3026, v3027, v3028, v3029, v3030, v3031, v3032, v3033, v3034, v3035, v3036, v3037, v3038, v3039, v3040, v3041, v3042, v3043, v3044, v3045, v3046, v3047, v3048, v3049, v3050, v3051, v3052, v3053, v3054, v3055, v3056, v3057, v3058, v3059, v3060, v3061, v3062, v3063, v3064, v3065, v3066, v3067, v3068, v3069, v3070, v3071, v3072, v3073, v3074, v3075, v3076, v3077, v3078, v3079, v3080, v3081, v3082, v3083, v3084, v3085, v3086, v3087, v3088, v3089, v3090, v3091, v3092, v3093, v3094, v3095, v3096, v3097, v3098, v3099, v3100, v3101, v3102, v3103, v3104, v3105, v3106, v3107, v3108, v3109, v3110, v3111, v3112, v3113, v3114, v3115, v3116, v3117, v3118, v3119, v3120, v3121, v3122, v3123, v3124, v3125, v3126, v3127, v3128, v3129, v3130, v3131, v3132, v3133, v3134, v3135, v3136, v3137, v3138, v3139, v3140, v3141, v3142, v3143, v3144, v3145, v3146, v3147, v3148, v3149, v3150, v3151, v3152, v3153, v3154, v3155, v3156, v3157, v3158, v3159, v3160, v3161, v3162, v3163, v3164, v3165, v3166, v3167, v3168, v3169, v3170, v3171, v3172, v3173, v3174, v3175, v3176, v3177, v3178, v3179, v3180, v3181, v3182, v3183, v3184, v3185, v3186, v3187, v3188, v3189, v3190, v3191, v3192, v3193, v3194, v3195, v3196, v3197, v3198, v3199, v3200, v3201, v3202, v3203, v3204, v3205, v3206, v3207, v3208, v3209, v3210, v3211, v3212, v3213, v3214, v3215, v3216, v3217, v3218, v3219, v3220, v3221, v3222, v3223, v3224, v3225, v3226, v3227, v3228, v3229, v3230, v3231, v3232, v3233, v3234, v3235, v3236, v3237, v3238, v3239, v3240, v3241, v3242, v3243, v3244, v3245, v3246, v3247, v3248, v3249, v3250, v3251, v3252, v3253, v3254, v3255, v3256, v3257, v3258, v3259, v3260, v3261, v3262, v3263, v3264, v3265, v3266, v3267, v3268, v3269, v3270, v3271, v3272, v3273, v3274, v3275, v3276, v3277, v3278, v3279, v3280, v3281, v3282, v3283, v3284, v3285, v3286, v3287, v3288, v3289, v3290, v3291, v3292, v3293, v3294, v3295, v3296, v3297, v3298, v3299, v3300, v3301, v3302, v3303, v3304, v3305, v3306, v3307, v3308, v3309, v3310, v3311, v3312, v3313, v3314, v3315, v3316, v3317, v3318, v3319, v3320, v3321, v3322, v3323, v3324, v3325, v3326, v3327, v3328, v3329, v3330, v3331, v3332, v3333, v3334, v3335, v3336, v3337, v3338, v3339, v3340, v3341, v3342, v3343, v3344, v3345, v3346, v3347, v3348, v3349, v3350, v3351, v3352, v3353, v3354, v3355, v3356, v3357, v3358, v3359, v3360, v3361, v3362, v3363, v3364, v3365, v3366, v3367, v3368, v3369, v3370, v3371, v3372, v3373, v3374, v3375, v3376, v3377, v3378, v3379, v3380, v3381, v3382, v3383, v3384, v3385, v3386, v3387, v3388, v3389, v3390, v3391, v3392, v3393, v3394, v3395, v3396, v3397, v3398, v3399, v3400, v3401, v3402, v3403, v3404, v3405, v3406, v3407, v3408, v3409, v3410, v3411, v3412, v3413, v3414, v3415, v3416, v3417, v3418, v3419, v3420, v3421, v3422, v3423, v3424, v3425, v3426, v3427, v3428, v3429, v3430, v3431, v3432, v3433, v3434, v3435, v3436, v3437, v3438, v3439, v3440, v3441, v3442, v3443, v3444, v3445, v3446, v3447, v3448, v3449, v3450, v3451, v3452, v3453, v3454, v3455, v3456, v3457, v3458, v3459, v3460, v3461, v3462, v3463, v3464, v3465, v3466, v3467, v3468, v3469, v3470, v3471, v3472, v3473, v3474, v3475, v3476, v3477, v3478, v3479, v3480, v3481, v3482, v3483, v3484, v3485, v3486, v3487, v3488, v3489, v3490, v3491, v3492, v3493, v3494, v3495, v3496, v3497, v3498, v3499, v3500, v3501, v3502, v3503, v3504, v3505, v3506, v3507, v3508, v3509, v3510, v3511, v3512, v3513, v3514, v3515, v3516, v3517, v3518, v3519, v3520, v3521, v3522, v3523, v3524, v3525, v3526, v3527, v3528, v3529, v3530, v3531, v3532, v3533, v3534, v3535, v3536, v3537, v3538, v3539, v3540, v3541, v3542, v3543, v3544, v3545, v3546, v3547, v3548, v3549, v3550, v3551, v3552, v3553, v3554, v3555, v3556, v3557, v3558, v3559, v3560, v3561, v3562, v3563, v3564, v3565, v3566, v3567, v3568, v3569, v3570, v3571, v3572, v3573, v3574, v3575, v3576, v3577, v3578, v3579, v3580, v3581, v3582, v3583, v3584, v3585, v3586, v3587, v3588, v3589, v3590, v3591, v3592, v3593, v3594, v3595, v3596, v3597, v3598, v3599, v3600, v3601, v3602, v3603, v3604, v3605, v3606, v3607, v3608, v3609, v3610, v3611, v3612, v3613, v3614, v3615, v3616, v3617, v3618, v3619, v3620, v3621, v3622, v3623, v3624, v3625, v3626, v3627, v3628, v3629, v3630, v3631, v3632, v3633, v3634, v3635, v3636, v3637, v3638, v3639, v3640, v3641, v3642, v3643, v3644, v3645, v3646, v3647, v3648, v3649, v3650, v3651, v3652, v3653, v3654, v3655, v3656, v3657, v3658, v3659, v3660, v3661, v3662, v3663, v3664, v3665, v3666, v3667, v3668, v3669, v3670, v3671, v3672, v3673, v3674, v3675, v3676, v3677, v3678, v3679, v3680, v3681, v3682, v3683, v3684, v3685, v3686, v3687, v3688, v3689, v3690, v3691, v3692, v3693, v3694, v3695, v3696, v3697, v3698, v3699, v3700, v3701, v3702, v3703, v3704, v3705, v3706, v3707, v3708, v3709, v3710, v3711, v3712, v3713, v3714, v3715, v3716, v3717, v3718, v3719, v3720, v3721, v3722, v3723, v3724, v3725, v3726, v3727, v3728, v3729, v3730, v3731, v3732, v3733, v3734, v3735, v3736, v3737, v3738, v3739, v3740, v3741, v3742, v3743, v3744, v3745, v3746, v3747, v3748, v3749, v3750, v3751, v3752, v3753, v3754, v3755, v3756, v3757, v3758, v3759, v3760, v3761, v3762, v3763, v3764, v3765, v3766, v3767, v3768, v3769, v3770, v3771, v3772, v3773, v3774, v3775, v3776, v3777, v3778, v3779, v3780, v3781, v3782, v3783, v3784, v3785, v3786, v3787, v3788, v3789, v3790, v3791, v3792, v3793, v3794, v3795, v3796, v3797, v3798, v3799, v3800, v3801, v3802, v3803, v3804, v3805, v3806, v3807, v3808, v3809, v3810, v3811, v3812, v3813, v3814, v3815, v3816, v3817, v3818, v3819, v3820, v3821, v3822, v3823, v3824, v3825, v3826, v3827, v3828, v3829, v3830, v3831, v3832, v3833, v3834, v3835, v3836, v3837, v3838, v3839, v3840, v3841, v3842, v3843, v3844, v3845, v3846, v3847, v3848, v3849, v3850, v3851, v3852, v3853, v3854, v3855, v3856, v3857, v3858, v3859, v3860, v3861, v3862, v3863, v3864, v3865, v3866, v3867, v3868, v3869, v3870, v3871, v3872, v3873, v3874, v3875, v3876, v3877, v3878, v3879, v3880, v3881, v3882, v3883, v3884, v3885, v3886, v3887, v3888, v3889, v3890, v3891, v3892, v3893, v3894, v3895, v3896, v3897, v3898, v3899, v3900, v3901, v3902, v3903, v3904, v3905, v3906, v3907, v3908, v3909, v3910, v3911, v3912, v3913, v3914, v3915, v3916, v3917, v3918, v3919, v3920, v3921, v3922, v3923, v3924, v3925, v3926, v3927, v3928, v3929, v3930, v3931, v3932, v3933, v3934, v3935, v3936, v3937, v3938, v3939, v3940, v3941, v3942, v3943, v3944, v3945, v3946, v3947, v3948, v3949, v3950, v3951, v3952, v3953, v3954, v3955, v3956, v3957, v3958, v3959, v3960, v3961, v3962, v3963, v3964, v3965, v3966, v3967, v3968, v3969, v3970, v3971, v3972, v3973, v3974, v3975, v3976, v3977, v3978, v3979, v3980, v3981, v3982, v3983, v3984, v3985, v3986, v3987, v3988, v3989, v3990, v3991, v3992, v3993, v3994, v3995, v3996, v3997, v3998, v3999, v4000, v4001, v4002, v4003, v4004, v4005, v4006, v4007, v4008, v4009, v4010, v4011, v4012, v4013, v4014, v4015, v4016, v4017, v4018, v4019, v4020, v4021, v4022, v4023, v4024, v4025, v4026, v4027, v4028, v4029, v4030, v4031, v4032, v4033, v4034, v4035, v4036, v4037, v4038, v4039, v4040, v4041, v4042, v4043, v4044, v4045, v4046, v4047, v4048, v4049, v4050, v4051, v4052, v4053, v4054, v4055, v4056, v4057, v4058, v4059, v4060, v4061, v4062, v4063, v4064, v4065, v4066, v4067, v4068, v4069, v4070, v4071, v4072, v4073, v4074, v4075, v4076, v4077, v4078, v4079, v4080, v4081, v4082, v4083, v4084, v4085, v4086, v4087, v4088, v4089, v4090, v4091, v4092, v4093, v4094, v4095, v4096, v4097, v4098, v4099, v4100, v4101, v4102, v4103, v4104, v4105, v4106, v4107, v4108, v4109, v4110, v4111, v4112, v4113, v4114, v4115, v4116, v4117, v4118, v4119, v4120, v4121, v4122, v4123, v4124, v4125, v4126, v4127, v4128, v4129, v4130, v4131, v4132, v4133, v4134, v4135, v4136, v4137, v4138, v4139, v4140, v4141, v4142, v4143, v4144, v4145, v4146, v4147, v4148, v4149, v4150, v4151, v4152, v4153, v4154, v4155, v4156, v4157, v4158, v4159, v4160, v4161, v4162, v4163, v4164, v4165, v4166, v4167, v4168, v4169, v4170, v4171, v4172, v4173, v4174, v4175, v4176, v4177, v4178, v4179, v4180, v4181, v4182, v4183, v4184, v4185, v4186, v4187, v4188, v4189, v4190, v4191, v4192, v4193, v4194, v4195, v4196, v4197, v4198, v4199, v4200, v4201, v4202, v4203, v4204, v4205, v4206, v4207, v4208, v4209, v4210, v4211, v4212, v4213, v4214, v4215, v4216, v4217, v4218, v4219, v4220, v4221, v4222, v4223, v4224, v4225, v4226, v4227, v4228, v4229, v4230, v4231, v4232, v4233, v4234, v4235, v4236, v4237, v4238, v4239, v4240, v4241, v4242, v4243, v4244, v4245, v4246, v4247, v4248, v4249, v4250, v4251, v4252, v4253, v4254, v4255, v4256, v4257, v4258, v4259, v4260, v4261, v4262, v4263, v4264, v4265, v4266, v4267, v4268, v4269, v4270, v4271, v4272, v4273, v4274, v4275, v4276, v4277, v4278, v4279, v4280, v4281, v4282, v4283, v4284, v4285, v4286, v4287, v4288, v4289, v4290, v4291, v4292, v4293, v4294, v4295, v4296, v4297, v4298, v4299, v4300, v4301, v4302, v4303, v4304, v4305, v4306, v4307, v4308, v4309, v4310, v4311, v4312, v4313, v4314, v4315, v4316, v4317, v4318, v4319, v4320, v4321, v4322, v4323, v4324, v4325, v4326, v4327, v4328, v4329, v4330, v4331, v4332, v4333, v4334, v4335, v4336, v4337, v4338, v4339, v4340, v4341, v4342, v4343, v4344, v4345, v4346, v4347, v4348, v4349, v4350, v4351, v4352, v4353, v4354, v4355, v4356, v4357, v4358, v4359, v4360, v4361, v4362, v4363, v4364, v4365, v4366, v4367, v4368, v4369, v4370, v4371, v4372, v4373, v4374, v4375, v4376, v4377, v4378, v4379, v4380, v4381, v4382, v4383, v4384, v4385, v4386, v4387, v4388, v4389, v4390, v4391, v4392, v4393, v4394, v4395, v4396, v4397, v4398, v4399, v4400, v4401, v4402, v4403, v4404, v4405, v4406, v4407, v4408, v4409, v4410, v4411, v4412, v4413, v4414, v4415, v4416, v4417, v4418, v4419, v4420, v4421, v4422, v4423, v4424, v4425, v4426, v4427, v4428, v4429, v4430, v4431, v4432, v4433, v4434, v4435, v4436, v4437, v4438, v4439, v4440, v4441, v4442, v4443, v4444, v4445, v4446, v4447, v4448, v4449, v4450, v4451, v4452, v4453, v4454, v4455, v4456, v4457, v4458, v4459, v4460, v4461, v4462, v4463, v4464, v4465, v4466, v4467, v4468, v4469, v4470, v4471, v4472, v4473, v4474, v4475, v4476, v4477, v4478, v4479, v4480, v4481, v4482, v4483, v4484, v4485, v4486, v4487, v4488, v4489, v4490, v4491, v4492, v4493, v4494, v4495, v4496, v4497, v4498, v4499, v4500, v4501, v4502, v4503, v4504, v4505, v4506, v4507, v4508, v4509, v4510, v4511, v4512, v4513, v4514, v4515, v4516, v4517, v4518, v4519, v4520, v4521, v4522, v4523, v4524, v4525, v4526, v4527, v4528, v4529, v4530, v4531, v4532, v4533, v4534, v4535, v4536, v4537, v4538, v4539, v4540, v4541, v4542, v4543, v4544, v4545, v4546, v4547, v4548, v4549, v4550, v4551, v4552, v4553, v4554, v4555, v4556, v4557, v4558, v4559, v4560, v4561, v4562, v4563, v4564, v4565, v4566, v4567, v4568, v4569, v4570, v4571, v4572, v4573, v4574, v4575, v4576, v4577, v4578, v4579, v4580, v4581, v4582, v4583, v4584, v4585, v4586, v4587, v4588, v4589, v4590, v4591, v4592, v4593, v4594, v4595, v4596, v4597, v4598, v4599, v4600, v4601, v4602, v4603, v4604, v4605, v4606, v4607, v4608, v4609, v4610, v4611, v4612, v4613, v4614, v4615, v4616, v4617, v4618, v4619, v4620, v4621, v4622, v4623, v4624, v4625, v4626, v4627, v4628, v4629, v4630, v4631, v4632, v4633, v4634, v4635, v4636, v4637, v4638, v4639, v4640, v4641, v4642, v4643, v4644, v4645, v4646, v4647, v4648, v4649, v4650, v4651, v4652, v4653, v4654, v4655, v4656, v4657, v4658, v4659, v4660, v4661, v4662, v4663, v4664, v4665, v4666, v4667, v4668, v4669, v4670, v4671, v4672, v4673, v4674, v4675, v4676, v4677, v4678, v4679, v4680, v4681, v4682, v4683, v4684, v4685, v4686, v4687, v4688, v4689, v4690, v4691, v4692, v4693, v4694, v4695, v4696, v4697, v4698, v4699, v4700, v4701, v4702, v4703, v4704, v4705, v4706, v4707, v4708, v4709, v4710, v4711, v4712, v4713, v4714, v4715, v4716, v4717, v4718, v4719, v4720, v4721, v4722, v4723, v4724, v4725, v4726, v4727, v4728, v4729, v4730, v4731, v4732, v4733, v4734, v4735, v4736, v4737, v4738, v4739, v4740, v4741, v4742, v4743, v4744, v4745, v4746, v4747, v4748, v4749, v4750, v4751, v4752, v4753, v4754, v4755, v4756, v4757, v4758, v4759, v4760, v4761, v4762, v4763, v4764, v4765, v4766, v4767, v4768, v4769, v4770, v4771, v4772, v4773, v4774, v4775, v4776, v4777, v4778, v4779, v4780, v4781, v4782, v4783, v4784, v4785, v4786, v4787, v4788, v4789, v4790, v4791, v4792, v4793, v4794, v4795, v4796, v4797, v4798, v4799, v4800, v4801, v4802, v4803, v4804, v4805, v4806, v4807, v4808, v4809, v4810, v4811, v4812, v4813, v4814, v4815, v4816, v4817, v4818, v4819, v4820, v4821, v4822, v4823, v4824, v4825, v4826, v4827, v4828, v4829, v4830, v4831, v4832, v4833, v4834, v4835, v4836, v4837, v4838, v4839, v4840, v4841, v4842, v4843, v4844, v4845, v4846, v4847, v4848, v4849, v4850, v4851, v4852, v4853, v4854, v4855, v4856, v4857, v4858, v4859, v4860, v4861, v4862, v4863, v4864, v4865, v4866, v4867, v4868, v4869, v4870, v4871, v4872, v4873, v4874, v4875, v4876, v4877, v4878, v4879, v4880, v4881, v4882, v4883, v4884, v4885, v4886, v4887, v4888, v4889, v4890, v4891, v4892, v4893, v4894, v4895, v4896, v4897, v4898, v4899, v4900, v4901, v4902, v4903, v4904, v4905, v4906, v4907, v4908, v4909, v4910, v4911, v4912, v4913, v4914, v4915, v4916, v4917, v4918, v4919, v4920, v4921, v4922, v4923, v4924, v4925, v4926, v4927, v4928, v4929, v4930, v4931, v4932, v4933, v4934, v4935, v4936, v4937, v4938, v4939, v4940, v4941, v4942, v4943, v4944, v4945, v4946, v4947, v4948, v4949, v4950, v4951, v4952, v4953, v4954, v4955, v4956, v4957, v4958, v4959, v4960, v4961, v4962, v4963, v4964, v4965, v4966, v4967, v4968, v4969, v4970, v4971, v4972, v4973, v4974, v4975, v4976, v4977, v4978, v4979, v4980, v4981, v4982, v4983, v4984, v4985, v4986, v4987, v4988, v4989, v4990, v4991, v4992, v4993, v4994, v4995, v4996, v4997, v4998, v4999, v5000, v5001, v5002, v5003, v5004, v5005, v5006, v5007, v5008, v5009, v5010, v5011, v5012, v5013, v5014, v5015, v5016, v5017, v5018, v5019, v5020, v5021, v5022, v5023, v5024, v5025, v5026, v5027, v5028, v5029, v5030, v5031, v5032, v5033, v5034, v5035, v5036, v5037, v5038, v5039, v5040, v5041, v5042, v5043, v5044, v5045, v5046, v5047, v5048, v5049, v5050, v5051, v5052, v5053, v5054, v5055, v5056, v5057, v5058, v5059, v5060, v5061, v5062, v5063, v5064, v5065, v5066, v5067, v5068, v5069, v5070, v5071, v5072, v5073, v5074, v5075, v5076, v5077, v5078, v5079, v5080, v5081, v5082, v5083, v5084, v5085, v5086, v5087, v5088, v5089, v5090, v5091, v5092, v5093, v5094, v5095, v5096, v5097, v5098, v5099, v5100, v5101, v5102, v5103, v5104, v5105, v5106, v5107, v5108, v5109, v5110, v5111, v5112, v5113, v5114, v5115, v5116, v5117, v5118, v5119, v5120, v5121, v5122, v5123, v5124, v5125, v5126, v5127, v5128, v5129, v5130, v5131, v5132, v5133, v5134, v5135, v5136, v5137, v5138, v5139, v5140, v5141, v5142, v5143, v5144, v5145, v5146, v5147, v5148, v5149, v5150, v5151, v5152, v5153, v5154, v5155, v5156, v5157, v5158, v5159, v5160, v5161, v5162, v5163, v5164, v5165, v5166, v5167, v5168, v5169, v5170, v5171, v5172, v5173, v5174, v5175, v5176, v5177, v5178, v5179, v5180, v5181, v5182, v5183, v5184, v5185, v5186, v5187, v5188, v5189, v5190, v5191, v5192, v5193, v5194, v5195, v5196, v5197, v5198, v5199, v5200, v5201, v5202, v5203, v5204, v5205, v5206, v5207, v5208, v5209, v5210, v5211, v5212, v5213, v5214, v5215, v5216, v5217, v5218, v5219, v5220, v5221, v5222, v5223, v5224, v5225, v5226, v5227, v5228, v5229, v5230, v5231, v5232, v5233, v5234, v5235, v5236, v5237, v5238, v5239, v5240, v5241, v5242, v5243, v5244, v5245, v5246, v5247, v5248, v5249, v5250, v5251, v5252, v5253, v5254, v5255, v5256, v5257, v5258, v5259, v5260, v5261, v5262, v5263, v5264, v5265, v5266, v5267, v5268, v5269, v5270, v5271, v5272, v5273, v5274, v5275, v5276, v5277, v5278, v5279, v5280, v5281, v5282, v5283, v5284, v5285, v5286, v5287, v5288, v5289, v5290, v5291, v5292, v5293, v5294, v5295, v5296, v5297, v5298, v5299, v5300, v5301, v5302, v5303, v5304, v5305, v5306, v5307, v5308, v5309, v5310, v5311, v5312, v5313, v5314, v5315, v5316, v5317, v5318, v5319, v5320, v5321, v5322, v5323, v5324, v5325, v5326, v5327, v5328, v5329, v5330, v5331, v5332, v5333, v5334, v5335, v5336, v5337, v5338, v5339, v5340, v5341, v5342, v5343, v5344, v5345, v5346, v5347, v5348, v5349, v5350, v5351, v5352, v5353, v5354, v5355, v5356, v5357, v5358, v5359, v5360, v5361, v5362, v5363, v5364, v5365, v5366, v5367, v5368, v5369, v5370, v5371, v5372, v5373, v5374, v5375, v5376, v5377, v5378, v5379, v5380, v5381, v5382, v5383, v5384, v5385, v5386, v5387, v5388, v5389, v5390, v5391, v5392, v5393, v5394, v5395, v5396, v5397, v5398, v5399, v5400, v5401, v5402, v5403, v5404, v5405, v5406, v5407, v5408, v5409, v5410, v5411, v5412, v5413, v5414, v5415, v5416, v5417, v5418, v5419, v5420, v5421, v5422, v5423, v5424, v5425, v5426, v5427, v5428, v5429, v5430, v5431, v5432, v5433, v5434, v5435, v5436, v5437, v5438, v5439, v5440, v5441, v5442, v5443, v5444, v5445, v5446, v5447, v5448, v5449, v5450, v5451, v5452, v5453, v5454, v5455, v5456, v5457, v5458, v5459, v5460, v5461, v5462, v5463, v5464, v5465, v5466, v5467, v5468, v5469, v5470, v5471, v5472, v5473, v5474, v5475, v5476, v5477, v5478, v5479, v5480, v5481, v5482, v5483, v5484, v5485, v5486, v5487, v5488, v5489, v5490, v5491, v5492, v5493, v5494, v5495, v5496, v5497, v5498, v5499, v5500, v5501, v5502, v5503, v5504, v5505, v5506, v5507, v5508, v5509, v5510, v5511, v5512, v5513, v5514, v5515, v5516, v5517, v5518, v5519, v5520, v5521, v5522, v5523, v5524, v5525, v5526, v5527, v5528, v5529, v5530, v5531, v5532, v5533, v5534, v5535, v5536, v5537, v5538, v5539, v5540, v5541, v5542, v5543, v5544, v5545, v5546, v5547, v5548, v5549, v5550, v5551, v5552, v5553, v5554, v5555, v5556, v5557, v5558, v5559, v5560, v5561, v5562, v5563, v5564, v5565, v5566, v5567, v5568, v5569, v5570, v5571, v5572, v5573, v5574, v5575, v5576, v5577, v5578, v5579, v5580, v5581, v5582, v5583, v5584, v5585, v5586, v5587, v5588, v5589, v5590, v5591, v5592, v5593, v5594, v5595, v5596, v5597, v5598, v5599, v5600, v5601, v5602, v5603, v5604, v5605, v5606, v5607, v5608, v5609, v5610, v5611, v5612, v5613, v5614, v5615, v5616, v5617, v5618, v5619, v5620, v5621, v5622, v5623, v5624, v5625, v5626, v5627, v5628, v5629, v5630, v5631, v5632, v5633, v5634, v5635, v5636, v5637, v5638, v5639, v5640, v5641, v5642, v5643, v5644, v5645, v5646, v5647, v5648, v5649, v5650, v5651, v5652, v5653, v5654, v5655, v5656, v5657, v5658, v5659, v5660, v5661, v5662, v5663, v5664, v5665, v5666, v5667, v5668, v5669, v5670, v5671, v5672, v5673, v5674, v5675, v5676, v5677, v5678, v5679, v5680, v5681, v5682, v5683, v5684, v5685, v5686, v5687, v5688, v5689, v5690, v5691, v5692, v5693, v5694, v5695, v5696, v5697, v5698, v5699, v5700, v5701, v5702, v5703, v5704, v5705, v5706, v5707, v5708, v5709, v5710, v5711, v5712, v5713, v5714, v5715, v5716, v5717, v5718, v5719, v5720, v5721, v5722, v5723, v5724, v5725, v5726, v5727, v5728, v5729, v5730, v5731, v5732, v5733, v5734, v5735, v5736, v5737, v5738, v5739, v5740, v5741, v5742, v5743, v5744, v5745, v5746, v5747, v5748, v5749, v5750, v5751, v5752, v5753, v5754, v5755, v5756, v5757, v5758, v5759, v5760, v5761, v5762, v5763, v5764, v5765, v5766, v5767, v5768, v5769, v5770, v5771, v5772, v5773, v5774, v5775, v5776, v5777, v5778, v5779, v5780, v5781, v5782, v5783, v5784, v5785, v5786, v5787, v5788, v5789, v5790, v5791, v5792, v5793, v5794, v5795, v5796, v5797, v5798, v5799, v5800, v5801, v5802, v5803, v5804, v5805, v5806, v5807, v5808, v5809, v5810, v5811, v5812, v5813, v5814, v5815, v5816, v5817, v5818, v5819, v5820, v5821, v5822, v5823, v5824, v5825, v5826, v5827, v5828, v5829, v5830, v5831, v5832, v5833, v5834, v5835, v5836, v5837, v5838, v5839, v5840, v5841, v5842, v5843, v5844, v5845, v5846, v5847, v5848, v5849, v5850, v5851, v5852, v5853, v5854, v5855, v5856, v5857, v5858, v5859, v5860, v5861, v5862, v5863, v5864, v5865, v5866, v5867, v5868, v5869, v5870, v5871, v5872, v5873, v5874, v5875, v5876, v5877, v5878, v5879, v5880, v5881, v5882, v5883, v5884, v5885, v5886, v5887, v5888, v5889, v5890, v5891, v5892, v5893, v5894, v5895, v5896, v5897, v5898, v5899, v5900, v5901, v5902, v5903, v5904, v5905, v5906, v5907, v5908, v5909, v5910, v5911, v5912, v5913, v5914, v5915, v5916, v5917, v5918, v5919, v5920, v5921, v5922, v5923, v5924, v5925, v5926, v5927, v5928, v5929, v5930, v5931, v5932, v5933, v5934, v5935, v5936, v5937, v5938, v5939, v5940, v5941, v5942, v5943, v5944, v5945, v5946, v5947, v5948, v5949, v5950, v5951, v5952, v5953, v5954, v5955, v5956, v5957, v5958, v5959, v5960, v5961, v5962, v5963, v5964, v5965, v5966, v5967, v5968, v5969, v5970, v5971, v5972, v5973, v5974, v5975, v5976, v5977, v5978, v5979, v5980, v5981, v5982, v5983, v5984, v5985, v5986, v5987, v5988, v5989, v5990, v5991, v5992, v5993, v5994, v5995, v5996, v5997, v5998, v5999, v6000, v6001, v6002, v6003, v6004, v6005, v6006, v6007, v6008, v6009, v6010, v6011, v6012, v6013, v6014, v6015, v6016, v6017, v6018, v6019, v6020, v6021, v6022, v6023, v6024, v6025, v6026, v6027, v6028, v6029, v6030, v6031, v6032, v6033, v6034, v6035, v6036, v6037, v6038, v6039, v6040, v6041, v6042, v6043, v6044, v6045, v6046, v6047, v6048, v6049, v6050, v6051, v6052, v6053, v6054, v6055, v6056, v6057, v6058, v6059, v6060, v6061, v6062, v6063, v6064, v6065, v6066, v6067, v6068, v6069, v6070, v6071, v6072, v6073, v6074, v6075, v6076, v6077, v6078, v6079, v6080, v6081, v6082, v6083, v6084, v6085, v6086, v6087, v6088, v6089, v6090, v6091, v6092, v6093, v6094, v6095, v6096, v6097, v6098, v6099, v6100, v6101, v6102, v6103, v6104, v6105, v6106, v6107, v6108, v6109, v6110, v6111, v6112, v6113, v6114, v6115, v6116, v6117, v6118, v6119, v6120, v6121, v6122, v6123, v6124, v6125, v6126, v6127, v6128, v6129, v6130, v6131, v6132, v6133, v6134, v6135, v6136, v6137, v6138, v6139, v6140, v6141, v6142, v6143, v6144, v6145, v6146, v6147, v6148, v6149, v6150, v6151, v6152, v6153, v6154, v6155, v6156, v6157, v6158, v6159, v6160, v6161, v6162, v6163, v6164, v6165, v6166, v6167, v6168, v6169, v6170, v6171, v6172, v6173, v6174, v6175, v6176, v6177, v6178, v6179, v6180, v6181, v6182, v6183, v6184, v6185, v6186, v6187, v6188, v6189, v6190, v6191, v6192, v6193, v6194, v6195, v6196, v6197, v6198, v6199, v6200, v6201, v6202, v6203, v6204, v6205, v6206, v6207, v6208, v6209, v6210, v6211, v6212, v6213, v6214, v6215, v6216, v6217, v6218, v6219, v6220, v6221, v6222, v6223, v6224, v6225, v6226, v6227, v6228, v6229, v6230, v6231, v6232, v6233, v6234, v6235, v6236, v6237, v6238, v6239, v6240, v6241, v6242, v6243, v6244, v6245, v6246, v6247, v6248, v6249, v6250, v6251, v6252, v6253, v6254, v6255, v6256, v6257, v6258, v6259, v6260, v6261, v6262, v6263, v6264, v6265, v6266, v6267, v6268, v6269, v6270, v6271, v6272, v6273, v6274, v6275, v6276, v6277, v6278, v6279, v6280, v6281, v6282, v6283, v6284, v6285, v6286, v6287, v6288, v6289, v6290, v6291, v6292, v6293, v6294, v6295, v6296, v6297, v6298, v6299, v6300, v6301, v6302, v6303, v6304, v6305, v6306, v6307, v6308, v6309, v6310, v6311, v6312, v6313, v6314, v6315, v6316, v6317, v6318, v6319, v6320, v6321, v6322, v6323, v6324, v6325, v6326, v6327, v6328, v6329, v6330, v6331, v6332, v6333, v6334, v6335, v6336, v6337, v6338, v6339, v6340, v6341, v6342, v6343, v6344, v6345, v6346, v6347, v6348, v6349, v6350, v6351, v6352, v6353, v6354, v6355, v6356, v6357, v6358, v6359, v6360, v6361, v6362, v6363, v6364, v6365, v6366, v6367, v6368, v6369, v6370, v6371, v6372, v6373, v6374, v6375, v6376, v6377, v6378, v6379, v6380, v6381, v6382, v6383, v6384, v6385, v6386, v6387, v6388, v6389, v6390, v6391, v6392, v6393, v6394, v6395, v6396, v6397, v6398, v6399, v6400, v6401, v6402, v6403, v6404, v6405, v6406, v6407, v6408, v6409, v6410, v6411, v6412, v6413, v6414, v6415, v6416, v6417, v6418, v6419, v6420, v6421, v6422, v6423, v6424, v6425, v6426, v6427, v6428, v6429, v6430, v6431, v6432, v6433, v6434, v6435, v6436, v6437, v6438, v6439, v6440, v6441, v6442, v6443, v6444, v6445, v6446, v6447, v6448, v6449, v6450, v6451, v6452, v6453, v6454, v6455, v6456, v6457, v6458, v6459, v6460, v6461, v6462, v6463, v6464, v6465, v6466, v6467, v6468, v6469, v6470, v6471, v6472, v6473, v6474, v6475, v6476, v6477, v6478, v6479, v6480, v6481, v6482, v6483, v6484, v6485, v6486, v6487, v6488, v6489, v6490, v6491, v6492, v6493, v6494, v6495, v6496, v6497, v6498, v6499, v6500, v6501, v6502, v6503, v6504, v6505, v6506, v6507, v6508, v6509, v6510, v6511, v6512, v6513, v6514, v6515, v6516, v6517, v6518, v6519, v6520, v6521, v6522, v6523, v6524, v6525, v6526, v6527, v6528, v6529, v6530, v6531, v6532, v6533, v6534, v6535, v6536, v6537, v6538, v6539, v6540, v6541, v6542, v6543, v6544, v6545, v6546, v6547, v6548, v6549, v6550, v6551, v6552, v6553, v6554, v6555, v6556, v6557, v6558, v6559, v6560, v6561, v6562, v6563, v6564, v6565, v6566, v6567, v6568, v6569, v6570, v6571, v6572, v6573, v6574, v6575, v6576, v6577, v6578, v6579, v6580, v6581, v6582, v6583, v6584, v6585, v6586, v6587, v6588, v6589, v6590, v6591, v6592, v6593, v6594, v6595, v6596, v6597, v6598, v6599, v6600, v6601, v6602, v6603, v6604, v6605, v6606, v6607, v6608, v6609, v6610, v6611, v6612, v6613, v6614, v6615, v6616, v6617, v6618, v6619, v6620, v6621, v6622, v6623, v6624, v6625, v6626, v6627, v6628, v6629, v6630, v6631, v6632, v6633, v6634, v6635, v6636, v6637, v6638, v6639, v6640, v6641, v6642, v6643, v6644, v6645, v6646, v6647, v6648, v6649, v6650, v6651, v6652, v6653, v6654, v6655, v6656, v6657, v6658, v6659, v6660, v6661, v6662, v6663, v6664, v6665, v6666, v6667, v6668, v6669, v6670, v6671, v6672, v6673, v6674, v6675, v6676, v6677, v6678, v6679, v6680, v6681, v6682, v6683, v6684, v6685, v6686, v6687, v6688, v6689, v6690, v6691, v6692, v6693, v6694, v6695, v6696, v6697, v6698, v6699, v6700, v6701, v6702, v6703, v6704, v6705, v6706, v6707, v6708, v6709, v6710, v6711, v6712, v6713, v6714, v6715, v6716, v6717, v6718, v6719, v6720, v6721, v6722, v6723, v6724, v6725, v6726, v6727, v6728, v6729, v6730, v6731, v6732, v6733, v6734, v6735, v6736, v6737, v6738, v6739, v6740, v6741, v6742, v6743, v6744, v6745, v6746, v6747, v6748, v6749, v6750, v6751, v6752, v6753, v6754, v6755, v6756, v6757, v6758, v6759, v6760, v6761, v6762, v6763, v6764, v6765, v6766, v6767, v6768, v6769, v6770, v6771, v6772, v6773, v6774, v6775, v6776, v6777, v6778, v6779, v6780, v6781, v6782, v6783, v6784, v6785, v6786, v6787, v6788, v6789, v6790, v6791, v6792, v6793, v6794, v6795, v6796, v6797, v6798, v6799, v6800, v6801, v6802, v6803, v6804, v6805, v6806, v6807, v6808, v6809, v6810, v6811, v6812, v6813, v6814, v6815, v6816, v6817, v6818, v6819, v6820, v6821, v6822, v6823, v6824, v6825, v6826, v6827, v6828, v6829, v6830, v6831, v6832, v6833, v6834, v6835, v6836, v6837, v6838, v6839, v6840, v6841, v6842, v6843, v6844, v6845, v6846, v6847, v6848, v6849, v6850, v6851, v6852, v6853, v6854, v6855, v6856, v6857, v6858, v6859, v6860, v6861, v6862, v6863, v6864, v6865, v6866, v6867, v6868, v6869, v6870, v6871, v6872, v6873, v6874, v6875, v6876, v6877, v6878, v6879, v6880, v6881, v6882, v6883, v6884, v6885, v6886, v6887, v6888, v6889, v6890, v6891, v6892, v6893, v6894, v6895, v6896, v6897, v6898, v6899, v6900, v6901, v6902, v6903, v6904, v6905, v6906, v6907, v6908, v6909, v6910, v6911, v6912, v6913, v6914, v6915, v6916, v6917, v6918, v6919, v6920, v6921, v6922, v6923, v6924, v6925, v6926, v6927, v6928, v6929, v6930, v6931, v6932, v6933, v6934, v6935, v6936, v6937, v6938, v6939, v6940, v6941, v6942, v6943, v6944, v6945, v6946, v6947, v6948, v6949, v6950, v6951, v6952, v6953, v6954, v6955, v6956, v6957, v6958, v6959, v6960, v6961, v6962, v6963, v6964, v6965, v6966, v6967, v6968, v6969, v6970, v6971, v6972, v6973, v6974, v6975, v6976, v6977, v6978, v6979, v6980, v6981, v6982, v6983, v6984, v6985, v6986, v6987, v6988, v6989, v6990, v6991, v6992, v6993, v6994, v6995, v6996, v6997, v6998, v6999, v7000, v7001, v7002, v7003, v7004, v7005, v7006, v7007, v7008, v7009, v7010, v7011, v7012, v7013, v7014, v7015, v7016, v7017, v7018, v7019, v7020, v7021, v7022, v7023, v7024, v7025, v7026, v7027, v7028, v7029, v7030, v7031, v7032, v7033, v7034, v7035, v7036, v7037, v7038, v7039, v7040, v7041, v7042, v7043, v7044, v7045, v7046, v7047, v7048, v7049, v7050, v7051, v7052, v7053, v7054, v7055, v7056, v7057, v7058, v7059, v7060, v7061, v7062, v7063, v7064, v7065, v7066, v7067, v7068, v7069, v7070, v7071, v7072, v7073, v7074, v7075, v7076, v7077, v7078, v7079, v7080, v7081, v7082, v7083, v7084, v7085, v7086, v7087, v7088, v7089, v7090, v7091, v7092, v7093, v7094, v7095, v7096, v7097, v7098, v7099, v7100, v7101, v7102, v7103, v7104, v7105, v7106, v7107, v7108, v7109, v7110, v7111, v7112, v7113, v7114, v7115, v7116, v7117, v7118, v7119, v7120, v7121, v7122, v7123, v7124, v7125, v7126, v7127, v7128, v7129, v7130, v7131, v7132, v7133, v7134, v7135, v7136, v7137, v7138, v7139, v7140, v7141, v7142, v7143, v7144, v7145, v7146, v7147, v7148, v7149, v7150, v7151, v7152, v7153, v7154, v7155, v7156, v7157, v7158, v7159, v7160, v7161, v7162, v7163, v7164, v7165, v7166, v7167, v7168, v7169, v7170, v7171, v7172, v7173, v7174, v7175, v7176, v7177, v7178, v7179, v7180, v7181, v7182, v7183, v7184, v7185, v7186, v7187, v7188, v7189, v7190, v7191, v7192, v7193, v7194, v7195, v7196, v7197, v7198, v7199, v7200, v7201, v7202, v7203, v7204, v7205, v7206, v7207, v7208, v7209, v7210, v7211, v7212, v7213, v7214, v7215, v7216, v7217, v7218, v7219, v7220, v7221, v7222, v7223, v7224, v7225, v7226, v7227, v7228, v7229, v7230, v7231, v7232, v7233, v7234, v7235, v7236, v7237, v7238, v7239, v7240, v7241, v7242, v7243, v7244, v7245, v7246, v7247, v7248, v7249, v7250, v7251, v7252, v7253, v7254, v7255, v7256, v7257, v7258, v7259, v7260, v7261, v7262, v7263, v7264, v7265, v7266, v7267, v7268, v7269, v7270, v7271, v7272, v7273, v7274, v7275, v7276, v7277, v7278, v7279, v7280, v7281, v7282, v7283, v7284, v7285, v7286, v7287, v7288, v7289, v7290, v7291, v7292, v7293, v7294, v7295, v7296, v7297, v7298, v7299, v7300, v7301, v7302, v7303, v7304, v7305, v7306, v7307, v7308, v7309, v7310, v7311, v7312, v7313, v7314, v7315, v7316, v7317, v7318, v7319, v7320, v7321, v7322, v7323, v7324, v7325, v7326, v7327, v7328, v7329, v7330, v7331, v7332, v7333, v7334, v7335, v7336, v7337, v7338, v7339, v7340, v7341, v7342, v7343, v7344, v7345, v7346, v7347, v7348, v7349, v7350, v7351, v7352, v7353, v7354, v7355, v7356, v7357, v7358, v7359, v7360, v7361, v7362, v7363, v7364, v7365, v7366, v7367, v7368, v7369, v7370, v7371, v7372, v7373, v7374, v7375, v7376, v7377, v7378, v7379, v7380, v7381, v7382, v7383, v7384, v7385, v7386, v7387, v7388, v7389, v7390, v7391, v7392, v7393, v7394, v7395, v7396, v7397, v7398, v7399, v7400, v7401, v7402, v7403, v7404, v7405, v7406, v7407, v7408, v7409, v7410, v7411, v7412, v7413, v7414, v7415, v7416, v7417, v7418, v7419, v7420, v7421, v7422, v7423, v7424, v7425, v7426, v7427, v7428, v7429, v7430, v7431, v7432, v7433, v7434, v7435, v7436, v7437, v7438, v7439, v7440, v7441, v7442, v7443, v7444, v7445, v7446, v7447, v7448, v7449, v7450, v7451, v7452, v7453, v7454, v7455, v7456, v7457, v7458, v7459, v7460, v7461, v7462, v7463, v7464, v7465, v7466, v7467, v7468, v7469, v7470, v7471, v7472, v7473, v7474, v7475, v7476, v7477, v7478, v7479, v7480, v7481, v7482, v7483, v7484, v7485, v7486, v7487, v7488, v7489, v7490, v7491, v7492, v7493, v7494, v7495, v7496, v7497, v7498, v7499, v7500, v7501, v7502, v7503, v7504, v7505, v7506, v7507, v7508, v7509, v7510, v7511, v7512, v7513, v7514, v7515, v7516, v7517, v7518, v7519, v7520, v7521, v7522, v7523, v7524, v7525, v7526, v7527, v7528, v7529, v7530, v7531, v7532, v7533, v7534, v7535, v7536, v7537, v7538, v7539, v7540, v7541, v7542, v7543, v7544, v7545, v7546, v7547, v7548, v7549, v7550, v7551, v7552, v7553, v7554, v7555, v7556, v7557, v7558, v7559, v7560, v7561, v7562, v7563, v7564, v7565, v7566, v7567, v7568, v7569, v7570, v7571, v7572, v7573, v7574, v7575, v7576, v7577, v7578, v7579, v7580, v7581, v7582, v7583, v7584, v7585, v7586, v7587, v7588, v7589, v7590, v7591, v7592, v7593, v7594, v7595, v7596, v7597, v7598, v7599, v7600, v7601, v7602, v7603, v7604, v7605, v7606, v7607, v7608, v7609, v7610, v7611, v7612, v7613, v7614, v7615, v7616, v7617, v7618, v7619, v7620, v7621, v7622, v7623, v7624, v7625, v7626, v7627, v7628, v7629, v7630, v7631, v7632, v7633, v7634, v7635, v7636, v7637, v7638, v7639, v7640, v7641, v7642, v7643, v7644, v7645, v7646, v7647, v7648, v7649, v7650, v7651, v7652, v7653, v7654, v7655, v7656, v7657, v7658, v7659, v7660, v7661, v7662, v7663, v7664, v7665, v7666, v7667, v7668, v7669, v7670, v7671, v7672, v7673, v7674, v7675, v7676, v7677, v7678, v7679, v7680, v7681, v7682, v7683, v7684, v7685, v7686, v7687, v7688, v7689, v7690, v7691, v7692, v7693, v7694, v7695, v7696, v7697, v7698, v7699, v7700, v7701, v7702, v7703, v7704, v7705, v7706, v7707, v7708, v7709, v7710, v7711, v7712, v7713, v7714, v7715, v7716, v7717, v7718, v7719, v7720, v7721, v7722, v7723, v7724, v7725, v7726, v7727, v7728, v7729, v7730, v7731, v7732, v7733, v7734, v7735, v7736, v7737, v7738, v7739, v7740, v7741, v7742, v7743, v7744, v7745, v7746, v7747, v7748, v7749, v7750, v7751, v7752, v7753, v7754, v7755, v7756, v7757, v7758, v7759, v7760, v7761, v7762, v7763, v7764, v7765, v7766, v7767, v7768, v7769, v7770, v7771, v7772, v7773, v7774, v7775, v7776, v7777, v7778, v7779, v7780, v7781, v7782, v7783, v7784, v7785, v7786, v7787, v7788, v7789, v7790, v7791, v7792, v7793, v7794, v7795, v7796, v7797, v7798, v7799, v7800, v7801, v7802, v7803, v7804, v7805, v7806, v7807, v7808, v7809, v7810, v7811, v7812, v7813, v7814, v7815, v7816, v7817, v7818, v7819, v7820, v7821, v7822, v7823, v7824, v7825, v7826, v7827, v7828, v7829, v7830, v7831, v7832, v7833, v7834, v7835, v7836, v7837, v7838, v7839, v7840, v7841, v7842, v7843, v7844, v7845, v7846, v7847, v7848, v7849, v7850, v7851, v7852, v7853, v7854, v7855, v7856, v7857, v7858, v7859, v7860, v7861, v7862, v7863, v7864, v7865, v7866, v7867, v7868, v7869, v7870, v7871, v7872, v7873, v7874, v7875, v7876, v7877, v7878, v7879, v7880, v7881, v7882, v7883, v7884, v7885, v7886, v7887, v7888, v7889, v7890, v7891, v7892, v7893, v7894, v7895, v7896, v7897, v7898, v7899, v7900, v7901, v7902, v7903, v7904, v7905, v7906, v7907, v7908, v7909, v7910, v7911, v7912, v7913, v7914, v7915, v7916, v7917, v7918, v7919, v7920, v7921, v7922, v7923, v7924, v7925, v7926, v7927, v7928, v7929, v7930, v7931, v7932, v7933, v7934, v7935, v7936, v7937, v7938, v7939, v7940, v7941, v7942, v7943, v7944, v7945, v7946, v7947, v7948, v7949, v7950, v7951, v7952, v7953, v7954, v7955, v7956, v7957, v7958, v7959, v7960, v7961, v7962, v7963, v7964, v7965, v7966, v7967, v7968, v7969, v7970, v7971, v7972, v7973, v7974, v7975, v7976, v7977, v7978, v7979, v7980, v7981, v7982, v7983, v7984, v7985, v7986, v7987, v7988, v7989, v7990, v7991, v7992, v7993, v7994, v7995, v7996, v7997, v7998, v7999, v8000, v8001, v8002, v8003, v8004, v8005, v8006, v8007, v8008, v8009, v8010, v8011, v8012, v8013, v8014, v8015, v8016, v8017, v8018, v8019, v8020, v8021, v8022, v8023, v8024, v8025, v8026, v8027, v8028, v8029, v8030, v8031, v8032, v8033, v8034, v8035, v8036, v8037, v8038, v8039, v8040, v8041, v8042, v8043, v8044, v8045, v8046, v8047, v8048, v8049, v8050, v8051, v8052, v8053, v8054, v8055, v8056, v8057, v8058, v8059, v8060, v8061, v8062, v8063, v8064, v8065, v8066, v8067, v8068, v8069, v8070, v8071, v8072, v8073, v8074, v8075, v8076, v8077, v8078, v8079, v8080, v8081, v8082, v8083, v8084, v8085, v8086, v8087, v8088, v8089, v8090, v8091, v8092, v8093, v8094, v8095, v8096, v8097, v8098, v8099, v8100, v8101, v8102, v8103, v8104, v8105, v8106, v8107, v8108, v8109, v8110, v8111, v8112, v8113, v8114, v8115, v8116, v8117, v8118, v8119, v8120, v8121, v8122, v8123, v8124, v8125, v8126, v8127, v8128, v8129, v8130, v8131, v8132, v8133, v8134, v8135, v8136, v8137, v8138, v8139, v8140, v8141, v8142, v8143, v8144, v8145, v8146, v8147, v8148, v8149, v8150, v8151, v8152, v8153, v8154, v8155, v8156, v8157, v8158, v8159, v8160, v8161, v8162, v8163, v8164, v8165, v8166, v8167, v8168, v8169, v8170, v8171, v8172, v8173, v8174, v8175, v8176, v8177, v8178, v8179, v8180, v8181, v8182, v8183, v8184, v8185, v8186, v8187, v8188, v8189, v8190, v8191, v8192, v8193, v8194, v8195, v8196, v8197, v8198, v8199, v8200, v8201, v8202, v8203, v8204, v8205, v8206, v8207, v8208, v8209, v8210, v8211, v8212, v8213, v8214, v8215, v8216, v8217, v8218, v8219, v8220, v8221, v8222, v8223, v8224, v8225, v8226, v8227, v8228, v8229, v8230, v8231, v8232, v8233, v8234, v8235, v8236, v8237, v8238, v8239, v8240, v8241, v8242, v8243, v8244, v8245, v8246, v8247, v8248, v8249, v8250, v8251, v8252, v8253, v8254, v8255, v8256, v8257, v8258, v8259, v8260, v8261, v8262, v8263, v8264, v8265, v8266, v8267, v8268, v8269, v8270, v8271, v8272, v8273, v8274, v8275, v8276, v8277, v8278, v8279, v8280, v8281, v8282, v8283, v8284, v8285, v8286, v8287, v8288, v8289, v8290, v8291, v8292, v8293, v8294, v8295, v8296, v8297, v8298, v8299, v8300, v8301, v8302, v8303, v8304, v8305, v8306, v8307, v8308, v8309, v8310, v8311, v8312, v8313, v8314, v8315, v8316, v8317, v8318, v8319, v8320, v8321, v8322, v8323, v8324, v8325, v8326, v8327, v8328, v8329, v8330, v8331, v8332, v8333, v8334, v8335, v8336, v8337, v8338, v8339, v8340, v8341, v8342, v8343, v8344, v8345, v8346, v8347, v8348, v8349, v8350, v8351, v8352, v8353, v8354, v8355, v8356, v8357, v8358, v8359, v8360, v8361, v8362, v8363, v8364, v8365, v8366, v8367, v8368, v8369, v8370, v8371, v8372, v8373, v8374, v8375, v8376, v8377, v8378, v8379, v8380, v8381, v8382, v8383, v8384, v8385, v8386, v8387, v8388, v8389, v8390, v8391, v8392, v8393, v8394, v8395, v8396, v8397, v8398, v8399, v8400, v8401, v8402, v8403, v8404, v8405, v8406, v8407, v8408, v8409, v8410, v8411, v8412, v8413, v8414, v8415, v8416, v8417, v8418, v8419, v8420, v8421, v8422, v8423, v8424, v8425, v8426, v8427, v8428, v8429, v8430, v8431, v8432, v8433, v8434, v8435, v8436, v8437, v8438, v8439, v8440, v8441, v8442, v8443, v8444, v8445, v8446, v8447, v8448, v8449, v8450, v8451, v8452, v8453, v8454, v8455, v8456, v8457, v8458, v8459, v8460, v8461, v8462, v8463, v8464, v8465, v8466, v8467, v8468, v8469, v8470, v8471, v8472, v8473, v8474, v8475, v8476, v8477, v8478, v8479, v8480, v8481, v8482, v8483, v8484, v8485, v8486, v8487, v8488, v8489, v8490, v8491, v8492, v8493, v8494, v8495, v8496, v8497, v8498, v8499, v8500, v8501, v8502, v8503, v8504, v8505, v8506, v8507, v8508, v8509, v8510, v8511, v8512, v8513, v8514, v8515, v8516, v8517, v8518, v8519, v8520, v8521, v8522, v8523, v8524, v8525, v8526, v8527, v8528, v8529, v8530, v8531, v8532, v8533, v8534, v8535, v8536, v8537, v8538, v8539, v8540, v8541, v8542, v8543, v8544, v8545, v8546, v8547, v8548, v8549, v8550, v8551, v8552, v8553, v8554, v8555, v8556, v8557, v8558, v8559, v8560, v8561, v8562, v8563, v8564, v8565, v8566, v8567, v8568, v8569, v8570, v8571, v8572, v8573, v8574, v8575, v8576, v8577, v8578, v8579, v8580, v8581, v8582, v8583, v8584, v8585, v8586, v8587, v8588, v8589, v8590, v8591, v8592, v8593, v8594, v8595, v8596, v8597, v8598, v8599, v8600, v8601, v8602, v8603, v8604, v8605, v8606, v8607, v8608, v8609, v8610, v8611, v8612, v8613, v8614, v8615, v8616, v8617, v8618, v8619, v8620, v8621, v8622, v8623, v8624, v8625, v8626, v8627, v8628, v8629, v8630, v8631, v8632, v8633, v8634, v8635, v8636, v8637, v8638, v8639, v8640, v8641, v8642, v8643, v8644, v8645, v8646, v8647, v8648, v8649, v8650, v8651, v8652, v8653, v8654, v8655, v8656, v8657, v8658, v8659, v8660, v8661, v8662, v8663, v8664, v8665, v8666, v8667, v8668, v8669, v8670, v8671, v8672, v8673, v8674, v8675, v8676, v8677, v8678, v8679, v8680, v8681, v8682, v8683, v8684, v8685, v8686, v8687, v8688, v8689, v8690, v8691, v8692, v8693, v8694, v8695, v8696, v8697, v8698, v8699, v8700, v8701, v8702, v8703, v8704, v8705, v8706, v8707, v8708, v8709, v8710, v8711, v8712, v8713, v8714, v8715, v8716, v8717, v8718, v8719, v8720, v8721, v8722, v8723, v8724, v8725, v8726, v8727, v8728, v8729, v8730, v8731, v8732, v8733, v8734, v8735, v8736, v8737, v8738, v8739, v8740, v8741, v8742, v8743, v8744, v8745, v8746, v8747, v8748, v8749, v8750, v8751, v8752, v8753, v8754, v8755, v8756, v8757, v8758, v8759, v8760, v8761, v8762, v8763, v8764, v8765, v8766, v8767, v8768, v8769, v8770, v8771, v8772, v8773, v8774, v8775, v8776, v8777, v8778, v8779, v8780, v8781, v8782, v8783, v8784, v8785, v8786, v8787, v8788, v8789, v8790, v8791, v8792, v8793, v8794, v8795, v8796, v8797, v8798, v8799, v8800, v8801, v8802, v8803, v8804, v8805, v8806, v8807, v8808, v8809, v8810, v8811, v8812, v8813, v8814, v8815, v8816, v8817, v8818, v8819, v8820, v8821, v8822, v8823, v8824, v8825, v8826, v8827, v8828, v8829, v8830, v8831, v8832, v8833, v8834, v8835, v8836, v8837, v8838, v8839, v8840, v8841, v8842, v8843, v8844, v8845, v8846, v8847, v8848, v8849, v8850, v8851, v8852, v8853, v8854, v8855, v8856, v8857, v8858, v8859, v8860, v8861, v8862, v8863, v8864, v8865, v8866, v8867, v8868, v8869, v8870, v8871, v8872, v8873, v8874, v8875, v8876, v8877, v8878, v8879, v8880, v8881, v8882, v8883, v8884, v8885, v8886, v8887, v8888, v8889, v8890, v8891, v8892, v8893, v8894, v8895, v8896, v8897, v8898, v8899, v8900, v8901, v8902, v8903, v8904, v8905, v8906, v8907, v8908, v8909, v8910, v8911, v8912, v8913, v8914, v8915, v8916, v8917, v8918, v8919, v8920, v8921, v8922, v8923, v8924, v8925, v8926, v8927, v8928, v8929, v8930, v8931, v8932, v8933, v8934, v8935, v8936, v8937, v8938, v8939, v8940, v8941, v8942, v8943, v8944, v8945, v8946, v8947, v8948, v8949, v8950, v8951, v8952, v8953, v8954, v8955, v8956, v8957, v8958, v8959, v8960, v8961, v8962, v8963, v8964, v8965, v8966, v8967, v8968, v8969, v8970, v8971, v8972, v8973, v8974, v8975, v8976, v8977, v8978, v8979, v8980, v8981, v8982, v8983, v8984, v8985, v8986, v8987, v8988, v8989, v8990, v8991, v8992, v8993, v8994, v8995, v8996, v8997, v8998, v8999, v9000, v9001, v9002, v9003, v9004, v9005, v9006, v9007, v9008, v9009, v9010, v9011, v9012, v9013, v9014, v9015, v9016, v9017, v9018, v9019, v9020, v9021, v9022, v9023, v9024, v9025, v9026, v9027, v9028, v9029, v9030, v9031, v9032, v9033, v9034, v9035, v9036, v9037, v9038, v9039, v9040, v9041, v9042, v9043, v9044, v9045, v9046, v9047, v9048, v9049, v9050, v9051, v9052, v9053, v9054, v9055, v9056, v9057, v9058, v9059, v9060, v9061, v9062, v9063, v9064, v9065, v9066, v9067, v9068, v9069, v9070, v9071, v9072, v9073, v9074, v9075, v9076, v9077, v9078, v9079, v9080, v9081, v9082, v9083, v9084, v9085, v9086, v9087, v9088, v9089, v9090, v9091, v9092, v9093, v9094, v9095, v9096, v9097, v9098, v9099, v9100, v9101, v9102, v9103, v9104, v9105, v9106, v9107, v9108, v9109, v9110, v9111, v9112, v9113, v9114, v9115, v9116, v9117, v9118, v9119, v9120, v9121, v9122, v9123, v9124, v9125, v9126, v9127, v9128, v9129, v9130, v9131, v9132, v9133, v9134, v9135, v9136, v9137, v9138, v9139, v9140, v9141, v9142, v9143, v9144, v9145, v9146, v9147, v9148, v9149, v9150, v9151, v9152, v9153, v9154, v9155, v9156, v9157, v9158, v9159, v9160, v9161, v9162, v9163, v9164, v9165, v9166, v9167, v9168, v9169, v9170, v9171, v9172, v9173, v9174, v9175, v9176, v9177, v9178, v9179, v9180, v9181, v9182, v9183, v9184, v9185, v9186, v9187, v9188, v9189, v9190, v9191, v9192, v9193, v9194, v9195, v9196, v9197, v9198, v9199, v9200, v9201, v9202, v9203, v9204, v9205, v9206, v9207, v9208, v9209, v9210, v9211, v9212, v9213, v9214, v9215, v9216, v9217, v9218, v9219, v9220, v9221, v9222, v9223, v9224, v9225, v9226, v9227, v9228, v9229, v9230, v9231, v9232, v9233, v9234, v9235, v9236, v9237, v9238, v9239, v9240, v9241, v9242, v9243, v9244, v9245, v9246, v9247, v9248, v9249, v9250, v9251, v9252, v9253, v9254, v9255, v9256, v9257, v9258, v9259, v9260, v9261, v9262, v9263, v9264, v9265, v9266, v9267, v9268, v9269, v9270, v9271, v9272, v9273, v9274, v9275, v9276, v9277, v9278, v9279, v9280, v9281, v9282, v9283, v9284, v9285, v9286, v9287, v9288, v9289, v9290, v9291, v9292, v9293, v9294, v9295, v9296, v9297, v9298, v9299, v9300, v9301, v9302, v9303, v9304, v9305, v9306, v9307, v9308, v9309, v9310, v9311, v9312, v9313, v9314, v9315, v9316, v9317, v9318, v9319, v9320, v9321, v9322, v9323, v9324, v9325, v9326, v9327, v9328, v9329, v9330, v9331, v9332, v9333, v9334, v9335, v9336, v9337, v9338, v9339, v9340, v9341, v9342, v9343, v9344, v9345, v9346, v9347, v9348, v9349, v9350, v9351, v9352, v9353, v9354, v9355, v9356, v9357, v9358, v9359, v9360, v9361, v9362, v9363, v9364, v9365, v9366, v9367, v9368, v9369, v9370, v9371, v9372, v9373, v9374, v9375, v9376, v9377, v9378, v9379, v9380, v9381, v9382, v9383, v9384, v9385, v9386, v9387, v9388, v9389, v9390, v9391, v9392, v9393, v9394, v9395, v9396, v9397, v9398, v9399, v9400, v9401, v9402, v9403, v9404, v9405, v9406, v9407, v9408, v9409, v9410, v9411, v9412, v9413, v9414, v9415, v9416, v9417, v9418, v9419, v9420, v9421, v9422, v9423, v9424, v9425, v9426, v9427, v9428, v9429, v9430, v9431, v9432, v9433, v9434, v9435, v9436, v9437, v9438, v9439, v9440, v9441, v9442, v9443, v9444, v9445, v9446, v9447, v9448, v9449, v9450, v9451, v9452, v9453, v9454, v9455, v9456, v9457, v9458, v9459, v9460, v9461, v9462, v9463, v9464, v9465, v9466, v9467, v9468, v9469, v9470, v9471, v9472, v9473, v9474, v9475, v9476, v9477, v9478, v9479, v9480, v9481, v9482, v9483, v9484, v9485, v9486, v9487, v9488, v9489, v9490, v9491, v9492, v9493, v9494, v9495, v9496, v9497, v9498, v9499, v9500, v9501, v9502, v9503, v9504, v9505, v9506, v9507, v9508, v9509, v9510, v9511, v9512, v9513, v9514, v9515, v9516, v9517, v9518, v9519, v9520, v9521, v9522, v9523, v9524, v9525, v9526, v9527, v9528, v9529, v9530, v9531, v9532, v9533, v9534, v9535, v9536, v9537, v9538, v9539, v9540, v9541, v9542, v9543, v9544, v9545, v9546, v9547, v9548, v9549, v9550, v9551, v9552, v9553, v9554, v9555, v9556, v9557, v9558, v9559, v9560, v9561, v9562, v9563, v9564, v9565, v9566, v9567, v9568, v9569, v9570, v9571, v9572, v9573, v9574, v9575, v9576, v9577, v9578, v9579, v9580, v9581, v9582, v9583, v9584, v9585, v9586, v9587, v9588, v9589, v9590, v9591, v9592, v9593, v9594, v9595, v9596, v9597, v9598, v9599, v9600, v9601, v9602, v9603, v9604, v9605, v9606, v9607, v9608, v9609, v9610, v9611, v9612, v9613, v9614, v9615, v9616, v9617, v9618, v9619, v9620, v9621, v9622, v9623, v9624, v9625, v9626, v9627, v9628, v9629, v9630, v9631, v9632, v9633, v9634, v9635, v9636, v9637, v9638, v9639, v9640, v9641, v9642, v9643, v9644, v9645, v9646, v9647, v9648, v9649, v9650, v9651, v9652, v9653, v9654, v9655, v9656, v9657, v9658, v9659, v9660, v9661, v9662, v9663, v9664, v9665, v9666, v9667, v9668, v9669, v9670, v9671, v9672, v9673, v9674, v9675, v9676, v9677, v9678, v9679, v9680, v9681, v9682, v9683, v9684, v9685, v9686, v9687, v9688, v9689, v9690, v9691, v9692, v9693, v9694, v9695, v9696, v9697, v9698, v9699, v9700, v9701, v9702, v9703, v9704, v9705, v9706, v9707, v9708, v9709, v9710, v9711, v9712, v9713, v9714, v9715, v9716, v9717, v9718, v9719, v9720, v9721, v9722, v9723, v9724, v9725, v9726, v9727, v9728, v9729, v9730, v9731, v9732, v9733, v9734, v9735, v9736, v9737, v9738, v9739, v9740, v9741, v9742, v9743, v9744, v9745, v9746, v9747, v9748, v9749, v9750, v9751, v9752, v9753, v9754, v9755, v9756, v9757, v9758, v9759, v9760, v9761, v9762, v9763, v9764, v9765, v9766, v9767, v9768, v9769, v9770, v9771, v9772, v9773, v9774, v9775, v9776, v9777, v9778, v9779, v9780, v9781, v9782, v9783, v9784, v9785, v9786, v9787, v9788, v9789, v9790, v9791, v9792, v9793, v9794, v9795, v9796, v9797, v9798, v9799, v9800, v9801, v9802, v9803, v9804, v9805, v9806, v9807, v9808, v9809, v9810, v9811, v9812, v9813, v9814, v9815, v9816, v9817, v9818, v9819, v9820, v9821, v9822, v9823, v9824, v9825, v9826, v9827, v9828, v9829, v9830, v9831, v9832, v9833, v9834, v9835, v9836, v9837, v9838, v9839, v9840, v9841, v9842, v9843, v9844, v9845, v9846, v9847, v9848, v9849, v9850, v9851, v9852, v9853, v9854, v9855, v9856, v9857, v9858, v9859, v9860, v9861, v9862, v9863, v9864, v9865, v9866, v9867, v9868, v9869, v9870, v9871, v9872, v9873,
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325;
assign w0 = ~pi01 & pi02;
assign w1 = pi00 & w0;
assign w2 = pi01 & ~pi02;
assign w3 = pi00 & w2;
assign v0 = ~(w1 | w3);
assign w4 = v0;
assign v1 = ~(pi21 | pi22);
assign w5 = v1;
assign w6 = pi21 & pi22;
assign v2 = ~(w5 | w6);
assign w7 = v2;
assign v3 = ~(pi20 | pi21);
assign w8 = v3;
assign w9 = pi20 & pi21;
assign v4 = ~(w8 | w9);
assign w10 = v4;
assign v5 = ~(w7 | w10);
assign w11 = v5;
assign w12 = pi23 & ~w11;
assign w13 = ~pi22 & w8;
assign v6 = ~(w12 | w13);
assign w14 = v6;
assign v7 = ~(pi23 | pi26);
assign w15 = v7;
assign w16 = ~pi24 & pi25;
assign w17 = w15 & w16;
assign w18 = pi29 & pi30;
assign w19 = pi27 & pi28;
assign w20 = w18 & w19;
assign w21 = w17 & w20;
assign w22 = pi23 & pi26;
assign w23 = pi24 & ~pi25;
assign w24 = w22 & w23;
assign w25 = pi27 & ~pi28;
assign w26 = w18 & w25;
assign w27 = w24 & w26;
assign w28 = w15 & w23;
assign w29 = pi29 & ~pi30;
assign w30 = w25 & w29;
assign w31 = w28 & w30;
assign v8 = ~(pi29 | pi30);
assign w32 = v8;
assign w33 = ~pi27 & pi28;
assign w34 = w32 & w33;
assign w35 = pi23 & ~pi26;
assign w36 = w23 & w35;
assign w37 = w34 & w36;
assign v9 = ~(pi24 | pi25);
assign w38 = v9;
assign w39 = w35 & w38;
assign v10 = ~(pi27 | pi28);
assign w40 = v10;
assign w41 = w18 & w40;
assign w42 = w39 & w41;
assign v11 = ~(w37 | w42);
assign w43 = v11;
assign w44 = ~w31 & w43;
assign w45 = ~pi29 & pi30;
assign w46 = w40 & w45;
assign w47 = pi24 & pi25;
assign w48 = w22 & w47;
assign w49 = w46 & w48;
assign w50 = w19 & w32;
assign w51 = w17 & w50;
assign v12 = ~(w49 | w51);
assign w52 = v12;
assign w53 = w30 & w48;
assign w54 = w15 & w38;
assign w55 = w18 & w33;
assign w56 = w54 & w55;
assign v13 = ~(w53 | w56);
assign w57 = v13;
assign w58 = w52 & w57;
assign w59 = w44 & w58;
assign w60 = ~w27 & w59;
assign w61 = ~pi23 & pi26;
assign w62 = w47 & w61;
assign w63 = w46 & w62;
assign w64 = w22 & w38;
assign w65 = w26 & w64;
assign v14 = ~(w63 | w65);
assign w66 = v14;
assign w67 = w25 & w45;
assign w68 = w36 & w67;
assign w69 = w16 & w35;
assign w70 = w20 & w69;
assign w71 = w19 & w29;
assign w72 = pi25 & w61;
assign w73 = w71 & w72;
assign w74 = pi24 & w73;
assign v15 = ~(w70 | w74);
assign w75 = v15;
assign w76 = ~w68 & w75;
assign w77 = w69 & w71;
assign w78 = w34 & w54;
assign v16 = ~(w77 | w78);
assign w79 = v16;
assign w80 = w16 & w22;
assign w81 = w33 & w45;
assign w82 = w80 & w81;
assign w83 = w79 & ~w82;
assign w84 = w76 & w83;
assign w85 = w66 & w84;
assign w86 = w60 & w85;
assign w87 = w38 & w61;
assign w88 = w67 & w87;
assign w89 = w32 & w40;
assign w90 = w24 & w89;
assign v17 = ~(w88 | w90);
assign w91 = v17;
assign w92 = w16 & w61;
assign w93 = w34 & w92;
assign w94 = w23 & w61;
assign w95 = w71 & w94;
assign v18 = ~(w93 | w95);
assign w96 = v18;
assign w97 = w91 & w96;
assign w98 = w28 & w71;
assign w99 = w69 & w89;
assign w100 = w34 & w80;
assign v19 = ~(w99 | w100);
assign w101 = v19;
assign w102 = w29 & w40;
assign w103 = w69 & w102;
assign w104 = w101 & ~w103;
assign w105 = ~w98 & w104;
assign w106 = w35 & w47;
assign w107 = w46 & w106;
assign w108 = w17 & w67;
assign v20 = ~(w107 | w108);
assign w109 = v20;
assign w110 = w28 & w46;
assign w111 = w24 & w46;
assign w112 = w71 & w80;
assign v21 = ~(w111 | w112);
assign w113 = v21;
assign w114 = ~w110 & w113;
assign w115 = w109 & w114;
assign w116 = w105 & w115;
assign w117 = w97 & w116;
assign w118 = w19 & w45;
assign w119 = w28 & w118;
assign w120 = w50 & w94;
assign v22 = ~(w119 | w120);
assign w121 = v22;
assign w122 = w25 & w32;
assign w123 = w94 & w122;
assign w124 = w15 & w47;
assign w125 = w71 & w124;
assign v23 = ~(w123 | w125);
assign w126 = v23;
assign w127 = w39 & w71;
assign w128 = w26 & w48;
assign v24 = ~(w127 | w128);
assign w129 = v24;
assign w130 = w126 & w129;
assign w131 = w67 & w92;
assign w132 = w41 & w92;
assign v25 = ~(w131 | w132);
assign w133 = v25;
assign w134 = w92 & w118;
assign w135 = w17 & w26;
assign v26 = ~(w134 | w135);
assign w136 = v26;
assign w137 = w133 & w136;
assign w138 = w130 & w137;
assign w139 = w121 & w138;
assign w140 = w39 & w81;
assign w141 = w87 & w102;
assign v27 = ~(w140 | w141);
assign w142 = v27;
assign w143 = w26 & w94;
assign w144 = w41 & w106;
assign w145 = w34 & w94;
assign v28 = ~(w144 | w145);
assign w146 = v28;
assign w147 = ~w143 & w146;
assign w148 = w142 & w147;
assign w149 = w29 & w33;
assign w150 = w62 & w149;
assign w151 = w30 & w124;
assign v29 = ~(w150 | w151);
assign w152 = v29;
assign w153 = w148 & w152;
assign w154 = w139 & w153;
assign w155 = w117 & w154;
assign w156 = w86 & w155;
assign w157 = ~w21 & w156;
assign w158 = w36 & w89;
assign w159 = w54 & w118;
assign w160 = w55 & w80;
assign v30 = ~(w159 | w160);
assign w161 = v30;
assign w162 = w39 & w122;
assign w163 = w161 & ~w162;
assign w164 = ~w158 & w163;
assign w165 = w62 & w122;
assign w166 = w164 & ~w165;
assign w167 = w54 & w149;
assign w168 = w64 & w67;
assign w169 = w34 & w87;
assign v31 = ~(w168 | w169);
assign w170 = v31;
assign w171 = ~w167 & w170;
assign w172 = w54 & w67;
assign w173 = w28 & w102;
assign v32 = ~(w172 | w173);
assign w174 = v32;
assign w175 = w171 & w174;
assign w176 = w39 & w89;
assign w177 = w54 & w102;
assign v33 = ~(w176 | w177);
assign w178 = v33;
assign w179 = w92 & w102;
assign w180 = w39 & w55;
assign v34 = ~(w179 | w180);
assign w181 = v34;
assign w182 = w178 & w181;
assign w183 = w55 & w87;
assign w184 = w41 & w80;
assign v35 = ~(w183 | w184);
assign w185 = v35;
assign w186 = w124 & w149;
assign w187 = w34 & w106;
assign v36 = ~(w186 | w187);
assign w188 = v36;
assign w189 = w185 & w188;
assign w190 = w182 & w189;
assign w191 = w39 & w118;
assign w192 = w55 & w92;
assign v37 = ~(w191 | w192);
assign w193 = v37;
assign w194 = w30 & w69;
assign w195 = w46 & w94;
assign v38 = ~(w194 | w195);
assign w196 = v38;
assign w197 = w193 & w196;
assign w198 = ~pi26 & w47;
assign w199 = w50 & w198;
assign w200 = pi23 & w199;
assign w201 = w28 & w50;
assign w202 = w48 & w89;
assign v39 = ~(w201 | w202);
assign w203 = v39;
assign w204 = ~w200 & w203;
assign w205 = w197 & w204;
assign w206 = w190 & w205;
assign w207 = w175 & w206;
assign w208 = w24 & w102;
assign w209 = w106 & w149;
assign v40 = ~(w208 | w209);
assign w210 = v40;
assign w211 = w94 & w149;
assign w212 = w36 & w149;
assign v41 = ~(w211 | w212);
assign w213 = v41;
assign w214 = w69 & w122;
assign w215 = w20 & w80;
assign w216 = w36 & w81;
assign v42 = ~(w215 | w216);
assign w217 = v42;
assign w218 = ~w214 & w217;
assign w219 = w213 & w218;
assign w220 = w26 & w69;
assign w221 = w24 & w149;
assign v43 = ~(w220 | w221);
assign w222 = v43;
assign w223 = w64 & w122;
assign w224 = w102 & w124;
assign v44 = ~(w223 | w224);
assign w225 = v44;
assign w226 = w222 & w225;
assign w227 = w219 & w226;
assign w228 = w210 & w227;
assign w229 = w207 & w228;
assign w230 = w166 & w229;
assign w231 = w67 & w80;
assign w232 = w30 & w92;
assign v45 = ~(w231 | w232);
assign w233 = v45;
assign w234 = w62 & w67;
assign w235 = w20 & w92;
assign v46 = ~(w234 | w235);
assign w236 = v46;
assign w237 = w233 & w236;
assign w238 = w28 & w81;
assign w239 = w106 & w118;
assign v47 = ~(w238 | w239);
assign w240 = v47;
assign w241 = w81 & w106;
assign w242 = w240 & ~w241;
assign w243 = w237 & w242;
assign w244 = w34 & w69;
assign w245 = w64 & w71;
assign v48 = ~(w244 | w245);
assign w246 = v48;
assign w247 = w41 & w87;
assign w248 = w118 & w124;
assign v49 = ~(w247 | w248);
assign w249 = v49;
assign w250 = w246 & w249;
assign w251 = w48 & w55;
assign w252 = w62 & w102;
assign w253 = w20 & w36;
assign v50 = ~(w252 | w253);
assign w254 = v50;
assign w255 = ~w251 & w254;
assign w256 = w250 & w255;
assign w257 = w243 & w256;
assign w258 = w20 & w124;
assign w259 = w92 & w122;
assign w260 = w55 & w106;
assign v51 = ~(w259 | w260);
assign w261 = v51;
assign w262 = ~w258 & w261;
assign w263 = w41 & w62;
assign w264 = w48 & w102;
assign v52 = ~(w263 | w264);
assign w265 = v52;
assign w266 = w64 & w89;
assign w267 = w50 & w80;
assign v53 = ~(w266 | w267);
assign w268 = v53;
assign w269 = w265 & w268;
assign w270 = w262 & w269;
assign w271 = w64 & w102;
assign w272 = w36 & w102;
assign v54 = ~(w271 | w272);
assign w273 = v54;
assign w274 = w24 & w81;
assign w275 = w273 & ~w274;
assign w276 = w270 & w275;
assign w277 = w89 & w106;
assign w278 = w30 & w64;
assign v55 = ~(w277 | w278);
assign w279 = v55;
assign w280 = w39 & w46;
assign w281 = w81 & w92;
assign w282 = w46 & w124;
assign v56 = ~(w281 | w282);
assign w283 = v56;
assign w284 = ~w280 & w283;
assign w285 = w279 & w284;
assign w286 = w80 & w89;
assign w287 = w30 & w87;
assign w288 = w81 & w124;
assign v57 = ~(w287 | w288);
assign w289 = v57;
assign w290 = ~w286 & w289;
assign w291 = w20 & w24;
assign w292 = w106 & w122;
assign v58 = ~(w291 | w292);
assign w293 = v58;
assign w294 = w290 & w293;
assign w295 = w285 & w294;
assign w296 = w276 & w295;
assign w297 = w257 & w296;
assign w298 = w81 & w87;
assign w299 = w28 & w41;
assign w300 = w24 & w118;
assign v59 = ~(w299 | w300);
assign w301 = v59;
assign w302 = w48 & w50;
assign w303 = w80 & w118;
assign v60 = ~(w302 | w303);
assign w304 = v60;
assign w305 = w301 & w304;
assign w306 = ~w298 & w305;
assign w307 = w26 & w36;
assign w308 = w50 & w69;
assign w309 = w55 & w62;
assign v61 = ~(w308 | w309);
assign w310 = v61;
assign w311 = w36 & w41;
assign w312 = w55 & w124;
assign v62 = ~(w311 | w312);
assign w313 = v62;
assign w314 = w310 & w313;
assign w315 = ~w307 & w314;
assign w316 = w34 & w48;
assign w317 = w36 & w122;
assign v63 = ~(w316 | w317);
assign w318 = v63;
assign w319 = w315 & w318;
assign w320 = w306 & w319;
assign w321 = w297 & w320;
assign w322 = w230 & w321;
assign w323 = w157 & w322;
assign w324 = w89 & w94;
assign v64 = ~(w214 | w324);
assign w325 = v64;
assign w326 = w122 & w124;
assign v65 = ~(w169 | w326);
assign w327 = v65;
assign w328 = w325 & w327;
assign w329 = w36 & w71;
assign v66 = ~(w127 | w329);
assign w330 = v66;
assign w331 = w24 & w71;
assign v67 = ~(w99 | w331);
assign w332 = v67;
assign w333 = w330 & w332;
assign w334 = w328 & w333;
assign v68 = ~(w56 | w95);
assign w335 = v68;
assign v69 = ~(w241 | w264);
assign w336 = v69;
assign w337 = w20 & w39;
assign w338 = w69 & w118;
assign v70 = ~(w337 | w338);
assign w339 = v70;
assign w340 = w336 & w339;
assign w341 = w335 & w340;
assign w342 = w334 & w341;
assign w343 = w50 & w87;
assign v71 = ~(w251 | w343);
assign w344 = v71;
assign v72 = ~(w110 | w131);
assign w345 = v72;
assign w346 = ~w187 & w345;
assign w347 = w344 & w346;
assign v73 = ~(w200 | w234);
assign w348 = v73;
assign w349 = ~w123 & w348;
assign w350 = w347 & w349;
assign w351 = w342 & w350;
assign w352 = pi25 & w35;
assign w353 = w30 & w352;
assign v74 = ~(w307 | w353);
assign w354 = v74;
assign v75 = ~(w220 | w271);
assign w355 = v75;
assign w356 = w354 & w355;
assign w357 = w351 & w356;
assign v76 = ~(w141 | w221);
assign w358 = v76;
assign w359 = w26 & w124;
assign v77 = ~(w195 | w359);
assign w360 = v77;
assign w361 = w358 & w360;
assign v78 = ~(w235 | w288);
assign w362 = v78;
assign w363 = ~w245 & w362;
assign w364 = w361 & w363;
assign w365 = w357 & w364;
assign v79 = ~(w144 | w303);
assign w366 = v79;
assign w367 = ~w291 & w366;
assign w368 = ~w232 & w367;
assign w369 = w50 & w64;
assign w370 = w17 & w149;
assign v80 = ~(w369 | w370);
assign w371 = v80;
assign w372 = w67 & w198;
assign w373 = ~pi23 & w372;
assign w374 = w67 & w69;
assign v81 = ~(w373 | w374);
assign w375 = v81;
assign w376 = w371 & w375;
assign w377 = w368 & w376;
assign w378 = w30 & w62;
assign w379 = w17 & w55;
assign v82 = ~(w378 | w379);
assign w380 = v82;
assign w381 = w17 & w71;
assign v83 = ~(w212 | w381);
assign w382 = v83;
assign w383 = w380 & w382;
assign w384 = w30 & w80;
assign w385 = w17 & w118;
assign v84 = ~(w384 | w385);
assign w386 = v84;
assign w387 = w36 & w55;
assign w388 = w48 & w122;
assign v85 = ~(w387 | w388);
assign w389 = v85;
assign w390 = w36 & w50;
assign v86 = ~(w180 | w390);
assign w391 = v86;
assign w392 = w389 & w391;
assign w393 = w386 & w392;
assign w394 = w383 & w393;
assign w395 = w377 & w394;
assign v87 = ~(w68 | w108);
assign w396 = v87;
assign w397 = ~w231 & w396;
assign w398 = w62 & w118;
assign v88 = ~(w266 | w398);
assign w399 = v88;
assign w400 = w41 & w94;
assign v89 = ~(w215 | w400);
assign w401 = v89;
assign w402 = w399 & w401;
assign w403 = w397 & w402;
assign w404 = w71 & w92;
assign w405 = w55 & w69;
assign v90 = ~(w404 | w405);
assign w406 = v90;
assign w407 = w403 & w406;
assign w408 = w395 & w407;
assign w409 = w26 & w106;
assign w410 = w24 & w122;
assign v91 = ~(w409 | w410);
assign w411 = v91;
assign v92 = ~(w100 | w191);
assign w412 = v92;
assign w413 = w411 & w412;
assign w414 = w46 & w80;
assign v93 = ~(w165 | w252);
assign w415 = v93;
assign w416 = ~w414 & w415;
assign w417 = w413 & w416;
assign w418 = w28 & w122;
assign v94 = ~(w173 | w418);
assign w419 = v94;
assign w420 = w36 & w118;
assign w421 = w419 & ~w420;
assign w422 = w34 & w62;
assign w423 = w421 & ~w422;
assign w424 = w417 & w423;
assign w425 = w20 & w28;
assign v95 = ~(w160 | w425);
assign w426 = v95;
assign w427 = w28 & w89;
assign w428 = w54 & w81;
assign v96 = ~(w151 | w428);
assign w429 = v96;
assign w430 = w50 & w62;
assign w431 = w80 & w149;
assign v97 = ~(w430 | w431);
assign w432 = v97;
assign w433 = w429 & w432;
assign w434 = ~w427 & w433;
assign w435 = w426 & w434;
assign w436 = w424 & w435;
assign w437 = w34 & w64;
assign w438 = w94 & w102;
assign v98 = ~(w437 | w438);
assign w439 = v98;
assign v99 = ~(w135 | w159);
assign w440 = v99;
assign w441 = w81 & w94;
assign v100 = ~(w98 | w441);
assign w442 = v100;
assign w443 = w440 & w442;
assign w444 = w439 & w443;
assign w445 = w436 & w444;
assign w446 = w408 & w445;
assign w447 = w69 & w149;
assign w448 = w46 & w92;
assign v101 = ~(w447 | w448);
assign w449 = v101;
assign v102 = ~(w286 | w300);
assign w450 = v102;
assign w451 = w20 & w62;
assign v103 = ~(w192 | w451);
assign w452 = v103;
assign w453 = w450 & w452;
assign w454 = w92 & w149;
assign v104 = ~(w247 | w454);
assign w455 = v104;
assign w456 = w89 & w124;
assign w457 = w20 & w48;
assign v105 = ~(w456 | w457);
assign w458 = v105;
assign w459 = w455 & w458;
assign w460 = w453 & w459;
assign w461 = w449 & w460;
assign w462 = w41 & w54;
assign w463 = w26 & w87;
assign v106 = ~(w462 | w463);
assign w464 = v106;
assign w465 = w36 & w46;
assign w466 = w62 & w89;
assign v107 = ~(w176 | w466);
assign w467 = v107;
assign w468 = ~w465 & w467;
assign w469 = w24 & w41;
assign v108 = ~(w223 | w469);
assign w470 = v108;
assign w471 = w468 & w470;
assign w472 = w464 & w471;
assign w473 = w461 & w472;
assign w474 = w17 & w102;
assign w475 = pi23 & w372;
assign v109 = ~(w474 | w475);
assign w476 = v109;
assign w477 = ~w128 & w476;
assign v110 = ~(w37 | w201);
assign w478 = v110;
assign w479 = w41 & w64;
assign w480 = w478 & ~w479;
assign w481 = w48 & w118;
assign w482 = w20 & w54;
assign v111 = ~(w481 | w482);
assign w483 = v111;
assign w484 = w30 & w39;
assign w485 = w483 & ~w484;
assign w486 = w480 & w485;
assign w487 = w477 & w486;
assign w488 = w30 & w54;
assign v112 = ~(w267 | w488);
assign w489 = v112;
assign v113 = ~(w272 | w309);
assign w490 = v113;
assign w491 = ~w111 & w490;
assign w492 = w489 & w491;
assign w493 = w17 & w34;
assign w494 = w28 & w55;
assign v114 = ~(w493 | w494);
assign w495 = v114;
assign w496 = ~w93 & w495;
assign w497 = w17 & w46;
assign v115 = ~(w119 | w497);
assign w498 = v115;
assign w499 = w46 & w69;
assign v116 = ~(w280 | w499);
assign w500 = v116;
assign w501 = w498 & w500;
assign w502 = w496 & w501;
assign w503 = w64 & w81;
assign v117 = ~(w211 | w503);
assign w504 = v117;
assign w505 = w48 & w67;
assign v118 = ~(w298 | w505);
assign w506 = v118;
assign v119 = ~(w134 | w162);
assign w507 = v119;
assign w508 = w506 & w507;
assign w509 = w504 & w508;
assign w510 = w502 & w509;
assign w511 = w492 & w510;
assign w512 = w487 & w511;
assign w513 = w473 & w512;
assign w514 = w446 & w513;
assign w515 = w365 & w514;
assign v120 = ~(w323 | w515);
assign w516 = v120;
assign w517 = w323 & w515;
assign v121 = ~(w516 | w517);
assign w518 = v121;
assign w519 = ~w14 & w518;
assign w520 = w14 & ~w518;
assign v122 = ~(w519 | w520);
assign w521 = v122;
assign w522 = w87 & w118;
assign v123 = ~(w370 | w522);
assign w523 = v123;
assign v124 = ~(w214 | w448);
assign w524 = v124;
assign w525 = w46 & w87;
assign v125 = ~(w187 | w525);
assign w526 = v125;
assign w527 = w524 & w526;
assign w528 = w523 & w527;
assign w529 = w196 & w528;
assign w530 = w34 & w39;
assign w531 = w39 & w149;
assign v126 = ~(w530 | w531);
assign w532 = v126;
assign w533 = w39 & w102;
assign v127 = ~(w384 | w533);
assign w534 = v127;
assign w535 = ~w93 & w534;
assign w536 = w532 & w535;
assign v128 = ~(w337 | w438);
assign w537 = v128;
assign w538 = w536 & w537;
assign w539 = w529 & w538;
assign v129 = ~(w208 | w454);
assign w540 = v129;
assign w541 = w26 & w80;
assign v130 = ~(w145 | w541);
assign w542 = v130;
assign w543 = w540 & w542;
assign v131 = ~(w184 | w388);
assign w544 = v131;
assign v132 = ~(w420 | w479);
assign w545 = v132;
assign w546 = w544 & w545;
assign w547 = w543 & w546;
assign w548 = w30 & w36;
assign v133 = ~(w223 | w548);
assign w549 = v133;
assign w550 = w50 & w54;
assign v134 = ~(w505 | w550);
assign w551 = v134;
assign w552 = w549 & w551;
assign v135 = ~(w173 | w312);
assign w553 = v135;
assign v136 = ~(w132 | w387);
assign w554 = v136;
assign w555 = w553 & w554;
assign w556 = w552 & w555;
assign w557 = w547 & w556;
assign w558 = w20 & w106;
assign w559 = w20 & w87;
assign v137 = ~(w253 | w559);
assign w560 = v137;
assign w561 = ~w558 & w560;
assign w562 = w246 & w561;
assign w563 = w87 & w122;
assign w564 = w17 & w81;
assign v138 = ~(w563 | w564);
assign w565 = v138;
assign w566 = w26 & w92;
assign v139 = ~(w134 | w566);
assign w567 = v139;
assign w568 = w565 & w567;
assign w569 = w562 & w568;
assign w570 = w330 & w569;
assign w571 = w557 & w570;
assign w572 = w539 & w571;
assign v140 = ~(w465 | w497);
assign w573 = v140;
assign v141 = ~(w53 | w252);
assign w574 = v141;
assign w575 = w573 & w574;
assign v142 = ~(w128 | w430);
assign w576 = v142;
assign v143 = ~(w211 | w374);
assign w577 = v143;
assign w578 = w576 & w577;
assign w579 = w575 & w578;
assign v144 = ~(w51 | w331);
assign w580 = v144;
assign w581 = w26 & w54;
assign v145 = ~(w300 | w581);
assign w582 = v145;
assign w583 = w580 & w582;
assign w584 = w48 & w149;
assign v146 = ~(w160 | w584);
assign w585 = v146;
assign w586 = w583 & w585;
assign w587 = ~w131 & w293;
assign w588 = w39 & w67;
assign v147 = ~(w503 | w588);
assign w589 = v147;
assign w590 = ~w280 & w589;
assign w591 = w587 & w590;
assign w592 = w586 & w591;
assign w593 = w17 & w41;
assign v148 = ~(w56 | w593);
assign w594 = v148;
assign w595 = w41 & w48;
assign v149 = ~(w400 | w595);
assign w596 = v149;
assign v150 = ~(w88 | w326);
assign w597 = v150;
assign w598 = w596 & w597;
assign w599 = w594 & w598;
assign v151 = ~(w21 | w248);
assign w600 = v151;
assign w601 = w193 & w600;
assign w602 = w599 & w601;
assign w603 = w592 & w602;
assign w604 = w579 & w603;
assign w605 = w24 & w50;
assign w606 = w66 & ~w605;
assign v152 = ~(w78 | w488);
assign w607 = v152;
assign w608 = ~w140 & w607;
assign w609 = w71 & w352;
assign v153 = ~(w359 | w609);
assign w610 = v153;
assign w611 = w608 & w610;
assign w612 = w606 & w611;
assign w613 = w24 & w34;
assign v154 = ~(w287 | w613);
assign w614 = v154;
assign v155 = ~(w141 | w474);
assign w615 = v155;
assign w616 = ~w112 & w615;
assign w617 = w614 & w616;
assign w618 = w612 & w617;
assign w619 = w604 & w618;
assign w620 = w572 & w619;
assign v156 = ~(w49 | w302);
assign w621 = v156;
assign v157 = ~(w68 | w186);
assign w622 = v157;
assign w623 = w621 & w622;
assign w624 = w64 & w118;
assign v158 = ~(w316 | w624);
assign w625 = v158;
assign v159 = ~(w200 | w451);
assign w626 = v159;
assign w627 = w625 & w626;
assign w628 = w623 & w627;
assign w629 = w48 & w71;
assign w630 = w87 & w149;
assign v160 = ~(w165 | w630);
assign w631 = v160;
assign w632 = ~w629 & w631;
assign w633 = w67 & w94;
assign v161 = ~(w307 | w633);
assign w634 = v161;
assign w635 = w102 & w352;
assign v162 = ~(w343 | w635);
assign w636 = v162;
assign w637 = w634 & w636;
assign w638 = w632 & w637;
assign w639 = w62 & w81;
assign w640 = w30 & w94;
assign v163 = ~(w639 | w640);
assign w641 = v163;
assign w642 = w80 & w102;
assign w643 = w55 & w64;
assign v164 = ~(w642 | w643);
assign w644 = v164;
assign w645 = ~w398 & w644;
assign w646 = w641 & w645;
assign w647 = w638 & w646;
assign w648 = w628 & w647;
assign v165 = ~(w42 | w274);
assign w649 = v165;
assign v166 = ~(w282 | w457);
assign w650 = v166;
assign w651 = ~w159 & w650;
assign w652 = w34 & w124;
assign v167 = ~(w144 | w652);
assign w653 = v167;
assign w654 = ~w390 & w653;
assign w655 = w651 & w654;
assign w656 = w55 & w94;
assign v168 = ~(w494 | w656);
assign w657 = v168;
assign v169 = ~(w288 | w482);
assign w658 = v169;
assign w659 = w657 & w658;
assign w660 = w655 & w659;
assign w661 = w649 & w660;
assign w662 = w648 & w661;
assign w663 = w620 & w662;
assign w664 = ~w323 & w663;
assign w665 = w380 & ~w558;
assign w666 = w30 & w106;
assign v170 = ~(w390 | w666);
assign w667 = v170;
assign w668 = ~w482 & w667;
assign w669 = w665 & w668;
assign v171 = ~(w373 | w463);
assign w670 = v171;
assign w671 = ~w338 & w670;
assign w672 = w669 & w671;
assign w673 = w26 & w39;
assign w674 = w69 & w81;
assign v172 = ~(w125 | w674);
assign w675 = v172;
assign v173 = ~(w359 | w639);
assign w676 = v173;
assign w677 = w594 & w676;
assign w678 = w675 & w677;
assign w679 = ~w673 & w678;
assign w680 = w17 & w122;
assign v174 = ~(w533 | w680);
assign w681 = v174;
assign v175 = ~(w324 | w656);
assign w682 = v175;
assign w683 = ~w140 & w682;
assign v176 = ~(w481 | w530);
assign w684 = v176;
assign w685 = w17 & w89;
assign v177 = ~(w119 | w685);
assign w686 = v177;
assign w687 = w684 & w686;
assign w688 = w683 & w687;
assign w689 = w681 & w688;
assign w690 = w679 & w689;
assign w691 = w672 & w690;
assign w692 = w28 & w34;
assign v178 = ~(w120 | w692);
assign w693 = v178;
assign v179 = ~(w93 | w488);
assign w694 = v179;
assign w695 = w693 & w694;
assign w696 = ~w187 & w695;
assign w697 = w87 & w89;
assign v180 = ~(w462 | w697);
assign w698 = v180;
assign w699 = w71 & w87;
assign v181 = ~(w211 | w699);
assign w700 = v181;
assign w701 = w698 & w700;
assign v182 = ~(w479 | w624);
assign w702 = v182;
assign v183 = ~(w68 | w643);
assign w703 = v183;
assign w704 = w702 & w703;
assign w705 = w701 & w704;
assign w706 = w696 & w705;
assign v184 = ~(w110 | w201);
assign w707 = v184;
assign v185 = ~(w465 | w548);
assign w708 = v185;
assign w709 = w707 & w708;
assign w710 = ~w103 & w709;
assign w711 = w89 & w92;
assign v186 = ~(w95 | w711);
assign w712 = v186;
assign w713 = w709 & w28468;
assign w714 = w706 & w713;
assign w715 = w26 & w62;
assign v187 = ~(w302 | w715);
assign w716 = v187;
assign w717 = ~w369 & w716;
assign w718 = w706 & w28469;
assign w719 = w91 & w161;
assign w720 = ~w212 & w719;
assign v188 = ~(w221 | w595);
assign w721 = v188;
assign w722 = w412 & ~w418;
assign w723 = w721 & w722;
assign w724 = w720 & w723;
assign v189 = ~(w308 | w469);
assign w725 = v189;
assign v190 = ~(w143 | w566);
assign w726 = v190;
assign w727 = w48 & w81;
assign v191 = ~(w51 | w727);
assign w728 = v191;
assign w729 = w726 & w728;
assign w730 = w725 & w729;
assign w731 = w54 & w122;
assign v192 = ~(w192 | w374);
assign w732 = v192;
assign w733 = ~w731 & w732;
assign w734 = w732 & w28470;
assign w735 = w730 & w734;
assign w736 = w724 & w735;
assign v193 = ~(w398 | w584);
assign w737 = v193;
assign w738 = ~w427 & w737;
assign w739 = w24 & w67;
assign v194 = ~(w53 | w385);
assign w740 = v194;
assign w741 = ~w739 & w740;
assign w742 = w41 & w69;
assign v195 = ~(w494 | w742);
assign w743 = v195;
assign w744 = w449 & w743;
assign w745 = w741 & w744;
assign w746 = w738 & w745;
assign w747 = w736 & w746;
assign w748 = w718 & w747;
assign w749 = w46 & w64;
assign v196 = ~(w420 | w749);
assign w750 = v196;
assign w751 = ~w588 & w750;
assign v197 = ~(w63 | w82);
assign w752 = v197;
assign w753 = w54 & w89;
assign v198 = ~(w150 | w753);
assign w754 = v198;
assign w755 = ~w630 & w754;
assign w756 = w752 & w755;
assign w757 = w751 & w756;
assign w758 = w39 & w50;
assign v199 = ~(w633 | w758);
assign w759 = v199;
assign w760 = ~w331 & w759;
assign v200 = ~(w141 | w381);
assign w761 = v200;
assign v201 = ~(w31 | w135);
assign w762 = v201;
assign w763 = w761 & w762;
assign w764 = ~w404 & w763;
assign v202 = ~(w326 | w531);
assign w765 = v202;
assign w766 = ~w132 & w765;
assign v203 = ~(w425 | w522);
assign w767 = v203;
assign v204 = ~(w437 | w484);
assign w768 = v204;
assign w769 = w767 & w768;
assign w770 = w766 & w769;
assign w771 = w764 & w770;
assign w772 = w760 & w771;
assign w773 = w757 & w772;
assign w774 = w297 & w773;
assign w775 = w748 & w774;
assign w776 = w691 & w775;
assign v205 = ~(w108 | w481);
assign w777 = v205;
assign w778 = w710 & w777;
assign v206 = ~(w264 | w673);
assign w779 = v206;
assign v207 = ~(w195 | w629);
assign w780 = v207;
assign w781 = w779 & w780;
assign w782 = w778 & w781;
assign v208 = ~(w245 | w378);
assign w783 = v208;
assign w784 = w495 & w783;
assign w785 = ~w427 & w784;
assign v209 = ~(w312 | w374);
assign w786 = v209;
assign v210 = ~(w111 | w563);
assign w787 = v210;
assign w788 = w786 & w787;
assign v211 = ~(w93 | w180);
assign w789 = v211;
assign v212 = ~(w287 | w522);
assign w790 = v212;
assign w791 = w789 & w790;
assign w792 = w788 & w791;
assign w793 = w785 & w792;
assign v213 = ~(w131 | w299);
assign w794 = v213;
assign w795 = ~w65 & w794;
assign w796 = ~w558 & w795;
assign v214 = ~(w51 | w135);
assign w797 = v214;
assign w798 = ~w209 & w797;
assign w799 = ~w73 & w798;
assign w800 = w796 & w799;
assign v215 = ~(w120 | w263);
assign w801 = v215;
assign v216 = ~(w150 | w302);
assign w802 = v216;
assign w803 = w801 & w802;
assign w804 = w800 & w803;
assign w805 = w793 & w804;
assign w806 = w782 & w805;
assign v217 = ~(w176 | w418);
assign w807 = v217;
assign w808 = ~w441 & w807;
assign v218 = ~(w125 | w652);
assign w809 = v218;
assign w810 = ~w252 & w809;
assign w811 = w808 & w810;
assign w812 = w17 & w30;
assign v219 = ~(w159 | w595);
assign w813 = v219;
assign w814 = ~w428 & w813;
assign w815 = w813 & w31148;
assign w816 = w811 & w815;
assign v220 = ~(w187 | w223);
assign w817 = v220;
assign v221 = ~(w78 | w241);
assign w818 = v221;
assign v222 = ~(w112 | w317);
assign w819 = v222;
assign w820 = w818 & w819;
assign w821 = w817 & w820;
assign w822 = w94 & w118;
assign v223 = ~(w482 | w822);
assign w823 = v223;
assign w824 = ~w186 & w823;
assign w825 = w821 & w824;
assign w826 = w816 & w825;
assign w827 = ~w479 & w726;
assign v224 = ~(w31 | w331);
assign w828 = v224;
assign w829 = ~w605 & w828;
assign w830 = w827 & w829;
assign v225 = ~(w409 | w727);
assign w831 = v225;
assign w832 = ~w469 & w831;
assign w833 = w362 & w832;
assign w834 = w830 & w833;
assign v226 = ~(w128 | w370);
assign w835 = v226;
assign w836 = w649 & w835;
assign v227 = ~(w70 | w739);
assign w837 = v227;
assign v228 = ~(w381 | w451);
assign w838 = v228;
assign w839 = ~w753 & w838;
assign w840 = w837 & w839;
assign w841 = w836 & w840;
assign w842 = w834 & w841;
assign w843 = w826 & w842;
assign v229 = ~(w132 | w158);
assign w844 = v229;
assign w845 = ~w77 & w844;
assign v230 = ~(w127 | w530);
assign w846 = v230;
assign w847 = w845 & w846;
assign v231 = ~(w231 | w267);
assign w848 = v231;
assign v232 = ~(w398 | w422);
assign w849 = v232;
assign w850 = ~w253 & w849;
assign w851 = w848 & w850;
assign v233 = ~(w95 | w239);
assign w852 = v233;
assign w853 = ~w212 & w852;
assign w854 = w851 & w853;
assign w855 = w847 & w854;
assign w856 = w843 & w855;
assign v234 = ~(w300 | w613);
assign w857 = v234;
assign w858 = ~w281 & w857;
assign v235 = ~(w179 | w208);
assign w859 = v235;
assign w860 = ~w238 & w859;
assign v236 = ~(w247 | w584);
assign w861 = v236;
assign w862 = ~w385 & w861;
assign w863 = w860 & w862;
assign v237 = ~(w140 | w232);
assign w864 = v237;
assign v238 = ~(w37 | w329);
assign w865 = v238;
assign w866 = w864 & w865;
assign w867 = w449 & w866;
assign w868 = w863 & w867;
assign w869 = w858 & w868;
assign w870 = w24 & w55;
assign v239 = ~(w162 | w870);
assign w871 = v239;
assign w872 = ~w666 & w871;
assign w873 = ~w742 & w872;
assign w874 = w20 & w64;
assign v240 = ~(w379 | w874);
assign w875 = v240;
assign w876 = ~w680 & w875;
assign w877 = w80 & w122;
assign v241 = ~(w437 | w550);
assign w878 = v241;
assign w879 = ~w877 & w878;
assign w880 = w876 & w879;
assign w881 = w873 & w880;
assign w882 = ~w384 & w881;
assign v242 = ~(w98 | w177);
assign w883 = v242;
assign v243 = ~(w280 | w414);
assign w884 = v243;
assign w885 = w883 & w884;
assign w886 = w54 & w71;
assign v244 = ~(w192 | w886);
assign w887 = v244;
assign w888 = w46 & w54;
assign v245 = ~(w173 | w888);
assign w889 = v245;
assign w890 = w887 & w889;
assign w891 = w885 & w890;
assign w892 = w50 & w124;
assign v246 = ~(w63 | w892);
assign w893 = v246;
assign v247 = ~(w260 | w699);
assign w894 = v247;
assign w895 = ~w420 & w894;
assign w896 = w893 & w895;
assign w897 = w891 & w896;
assign v248 = ~(w343 | w373);
assign w898 = v248;
assign w899 = w71 & w106;
assign v249 = ~(w309 | w643);
assign w900 = v249;
assign w901 = ~w141 & w900;
assign w902 = ~w899 & w901;
assign w903 = w898 & w902;
assign w904 = w897 & w903;
assign w905 = w882 & w904;
assign w906 = w869 & w905;
assign w907 = w856 & w906;
assign w908 = w806 & w907;
assign v250 = ~(w776 | w908);
assign w909 = v250;
assign v251 = ~(pi17 | pi18);
assign w910 = v251;
assign w911 = pi17 & pi18;
assign v252 = ~(w910 | w911);
assign w912 = v252;
assign v253 = ~(pi18 | pi19);
assign w913 = v253;
assign w914 = pi18 & pi19;
assign v254 = ~(w913 | w914);
assign w915 = v254;
assign v255 = ~(w912 | w915);
assign w916 = v255;
assign w917 = pi20 & ~w916;
assign w918 = ~pi17 & w913;
assign v256 = ~(w917 | w918);
assign w919 = v256;
assign w920 = w776 & w908;
assign v257 = ~(w909 | w920);
assign w921 = v257;
assign w922 = ~w919 & w921;
assign v258 = ~(w909 | w922);
assign w923 = v258;
assign w924 = w663 & ~w923;
assign w925 = ~w663 & w923;
assign v259 = ~(w924 | w925);
assign w926 = v259;
assign w927 = pi31 & ~w32;
assign w928 = ~w18 & w927;
assign v260 = ~(w151 | w447);
assign w929 = v260;
assign v261 = ~(w88 | w593);
assign w930 = v261;
assign w931 = ~w134 & w930;
assign w932 = w929 & w931;
assign v262 = ~(w140 | w215);
assign w933 = v262;
assign v263 = ~(w82 | w531);
assign w934 = v263;
assign w935 = w933 & w934;
assign w936 = w932 & w935;
assign v264 = ~(w180 | w499);
assign w937 = v264;
assign v265 = ~(w150 | w282);
assign w938 = v265;
assign w939 = w937 & w938;
assign w940 = w936 & w939;
assign v266 = ~(w374 | w886);
assign w941 = v266;
assign w942 = ~w248 & w941;
assign v267 = ~(w253 | w715);
assign w943 = v267;
assign w944 = w942 & w943;
assign w945 = w41 & w124;
assign v268 = ~(w160 | w945);
assign w946 = v268;
assign w947 = ~w550 & w946;
assign v269 = ~(w343 | w387);
assign w948 = v269;
assign w949 = ~w172 & w948;
assign w950 = w947 & w949;
assign w951 = w944 & w950;
assign v270 = ~(w231 | w414);
assign w952 = v270;
assign v271 = ~(w187 | w216);
assign w953 = v271;
assign w954 = ~w331 & w953;
assign v272 = ~(w37 | w533);
assign w955 = v272;
assign w956 = w954 & w955;
assign w957 = w952 & w956;
assign w958 = w951 & w957;
assign v273 = ~(w441 | w753);
assign w959 = v273;
assign v274 = ~(w234 | w870);
assign w960 = v274;
assign w961 = w959 & w960;
assign w962 = w958 & w961;
assign w963 = w940 & w962;
assign v275 = ~(w131 | w409);
assign w964 = v275;
assign v276 = ~(w454 | w630);
assign w965 = v276;
assign w966 = ~w159 & w965;
assign v277 = ~(w27 | w359);
assign w967 = v277;
assign w968 = w966 & w967;
assign w969 = w964 & w968;
assign v278 = ~(w77 | w428);
assign w970 = v278;
assign w971 = ~w70 & w970;
assign v279 = ~(w31 | w493);
assign w972 = v279;
assign w973 = ~w522 & w972;
assign w974 = w971 & w973;
assign w975 = ~w308 & w974;
assign w976 = w969 & w975;
assign v280 = ~(w143 | w505);
assign w977 = v280;
assign w978 = w20 & w94;
assign v281 = ~(w451 | w978);
assign w979 = v281;
assign w980 = w857 & w979;
assign v282 = ~(w280 | w431);
assign w981 = v282;
assign w982 = ~w398 & w981;
assign v283 = ~(w326 | w643);
assign w983 = v283;
assign w984 = ~w584 & w983;
assign w985 = w982 & w984;
assign w986 = w980 & w985;
assign w987 = w977 & w986;
assign w988 = w976 & w987;
assign w989 = w102 & w106;
assign v284 = ~(w264 | w989);
assign w990 = v284;
assign w991 = ~w317 & w990;
assign w992 = w675 & w991;
assign v285 = ~(w307 | w892);
assign w993 = v285;
assign v286 = ~(w194 | w425);
assign w994 = v286;
assign w995 = ~w427 & w994;
assign w996 = w993 & w995;
assign w997 = w64 & w149;
assign v287 = ~(w111 | w997);
assign w998 = v287;
assign w999 = w28 & w67;
assign v288 = ~(w260 | w999);
assign w1000 = v288;
assign w1001 = ~w888 & w1000;
assign w1002 = ~w564 & w1001;
assign w1003 = w998 & w1002;
assign w1004 = w996 & w1003;
assign w1005 = w992 & w1004;
assign w1006 = w988 & w1005;
assign v289 = ~(w463 | w497);
assign w1007 = v289;
assign v290 = ~(w93 | w503);
assign w1008 = v290;
assign w1009 = w1007 & w1008;
assign w1010 = ~w742 & w1009;
assign v291 = ~(w53 | w711);
assign w1011 = v291;
assign v292 = ~(w311 | w874);
assign w1012 = v292;
assign w1013 = w1011 & w1012;
assign v293 = ~(w673 | w758);
assign w1014 = v293;
assign w1015 = ~w224 & w1014;
assign w1016 = w1013 & w1015;
assign w1017 = w1010 & w1016;
assign v294 = ~(w110 | w581);
assign w1018 = v294;
assign w1019 = ~w202 & w1018;
assign v295 = ~(w378 | w481);
assign w1020 = v295;
assign w1021 = w1019 & w1020;
assign v296 = ~(w221 | w474);
assign w1022 = v296;
assign w1023 = w406 & w1022;
assign w1024 = w1021 & w1023;
assign w1025 = w1017 & w1024;
assign v297 = ~(w258 | w329);
assign w1026 = v297;
assign w1027 = w213 & w1026;
assign v298 = ~(w162 | w685);
assign w1028 = v298;
assign v299 = ~(w245 | w385);
assign w1029 = v299;
assign w1030 = ~w195 & w1029;
assign v300 = ~(w165 | w176);
assign w1031 = v300;
assign w1032 = w26 & w28;
assign v301 = ~(w119 | w1032);
assign w1033 = v301;
assign w1034 = w1031 & w1033;
assign w1035 = w1030 & w1034;
assign w1036 = w1028 & w1035;
assign w1037 = w1027 & w1036;
assign w1038 = w1025 & w1037;
assign w1039 = ~w56 & w419;
assign w1040 = ~w266 & w1039;
assign v302 = ~(w168 | w457);
assign w1041 = v302;
assign v303 = ~(w238 | w422);
assign w1042 = v303;
assign w1043 = ~w629 & w1042;
assign v304 = ~(w465 | w624);
assign w1044 = v304;
assign w1045 = w1043 & w1044;
assign w1046 = w1041 & w1045;
assign w1047 = w1040 & w1046;
assign v305 = ~(w292 | w482);
assign w1048 = v305;
assign v306 = ~(w259 | w652);
assign w1049 = v306;
assign w1050 = w1048 & w1049;
assign w1051 = ~w120 & w1050;
assign w1052 = w1047 & w1051;
assign w1053 = w1038 & w1052;
assign w1054 = w1006 & w1053;
assign w1055 = w963 & w1054;
assign v307 = ~(w381 | w699);
assign w1056 = v307;
assign w1057 = ~w739 & w1056;
assign w1058 = ~w248 & w1026;
assign w1059 = w1057 & w1058;
assign w1060 = ~w42 & w929;
assign w1061 = w57 & w1060;
assign w1062 = w1059 & w1061;
assign v308 = ~(w167 | w302);
assign w1063 = v308;
assign v309 = ~(w120 | w749);
assign w1064 = v309;
assign w1065 = w1063 & w1064;
assign v310 = ~(w165 | w369);
assign w1066 = v310;
assign w1067 = ~w160 & w1066;
assign w1068 = ~w311 & w1067;
assign w1069 = w1065 & w1068;
assign w1070 = w1062 & w1069;
assign v311 = ~(w107 | w110);
assign w1071 = v311;
assign w1072 = ~w822 & w1071;
assign v312 = ~(w140 | w244);
assign w1073 = v312;
assign v313 = ~(w550 | w692);
assign w1074 = v313;
assign w1075 = w1073 & w1074;
assign w1076 = w1072 & w1075;
assign v314 = ~(w202 | w494);
assign w1077 = v314;
assign v315 = ~(w208 | w488);
assign w1078 = v315;
assign w1079 = w1077 & w1078;
assign v316 = ~(w51 | w475);
assign w1080 = v316;
assign v317 = ~(w267 | w656);
assign w1081 = v317;
assign w1082 = w1080 & w1081;
assign w1083 = w1079 & w1082;
assign w1084 = w1076 & w1083;
assign w1085 = w1070 & w1084;
assign v318 = ~(w128 | w168);
assign w1086 = v318;
assign v319 = ~(w378 | w441);
assign w1087 = v319;
assign w1088 = w1086 & w1087;
assign w1089 = w539 & w1088;
assign w1090 = w1085 & w1089;
assign v320 = ~(w286 | w870);
assign w1091 = v320;
assign w1092 = ~w211 & w1091;
assign v321 = ~(w251 | w999);
assign w1093 = v321;
assign w1094 = w1044 & w1093;
assign w1095 = w1092 & w1094;
assign v322 = ~(w247 | w359);
assign w1096 = v322;
assign v323 = ~(w90 | w271);
assign w1097 = v323;
assign w1098 = w1096 & w1097;
assign v324 = ~(w99 | w409);
assign w1099 = v324;
assign w1100 = ~w172 & w1099;
assign w1101 = w1098 & w1100;
assign w1102 = w1095 & w1101;
assign v325 = ~(w70 | w989);
assign w1103 = v325;
assign w1104 = ~w742 & w1103;
assign w1105 = w1102 & w1104;
assign v326 = ~(w674 | w758);
assign w1106 = v326;
assign w1107 = ~w277 & w937;
assign w1108 = w50 & w92;
assign v327 = ~(w466 | w1108);
assign w1109 = v327;
assign v328 = ~(w191 | w287);
assign w1110 = v328;
assign w1111 = w1109 & w1110;
assign w1112 = w1107 & w1111;
assign w1113 = w1106 & w1112;
assign v329 = ~(w274 | w945);
assign w1114 = v329;
assign w1115 = w615 & w1114;
assign w1116 = w1113 & w1115;
assign w1117 = w1105 & w1116;
assign v330 = ~(w324 | w584);
assign w1118 = v330;
assign w1119 = w931 & w1118;
assign v331 = ~(w309 | w563);
assign w1120 = v331;
assign v332 = ~(w145 | w292);
assign w1121 = v332;
assign w1122 = ~w425 & w1121;
assign w1123 = w1120 & w1122;
assign w1124 = w1119 & w1123;
assign w1125 = w626 & w1124;
assign w1126 = w1117 & w1125;
assign v333 = ~(w150 | w731);
assign w1127 = v333;
assign v334 = ~(w212 | w379);
assign w1128 = v334;
assign w1129 = w1127 & w1128;
assign w1130 = ~w159 & w589;
assign v335 = ~(w410 | w613);
assign w1131 = v335;
assign v336 = ~(w135 | w263);
assign w1132 = v336;
assign w1133 = ~w997 & w1132;
assign w1134 = w24 & w30;
assign v337 = ~(w201 | w1134);
assign w1135 = v337;
assign w1136 = ~w317 & w1135;
assign w1137 = w1133 & w1136;
assign w1138 = w1131 & w1137;
assign w1139 = w1130 & w1138;
assign w1140 = w1129 & w1139;
assign v338 = ~(w143 | w326);
assign w1141 = v338;
assign v339 = ~(w119 | w390);
assign w1142 = v339;
assign w1143 = w970 & w1142;
assign w1144 = w236 & w752;
assign w1145 = ~w715 & w1144;
assign w1146 = w1143 & w1145;
assign v340 = ~(w177 | w298);
assign w1147 = v340;
assign w1148 = ~w316 & w1147;
assign w1149 = w1146 & w1148;
assign w1150 = w1141 & w1149;
assign w1151 = w1140 & w1150;
assign w1152 = w1126 & w1151;
assign w1153 = w1090 & w1152;
assign v341 = ~(w223 | w739);
assign w1154 = v341;
assign w1155 = ~w74 & w1154;
assign w1156 = ~w370 & w1155;
assign v342 = ~(w559 | w945);
assign w1157 = v342;
assign v343 = ~(w176 | w414);
assign w1158 = v343;
assign w1159 = w1157 & w1158;
assign w1160 = w1156 & w1159;
assign v344 = ~(w235 | w978);
assign w1161 = v344;
assign v345 = ~(w287 | w531);
assign w1162 = v345;
assign w1163 = w1161 & w1162;
assign v346 = ~(w187 | w624);
assign w1164 = v346;
assign v347 = ~(w308 | w673);
assign w1165 = v347;
assign w1166 = w1041 & w1165;
assign w1167 = w1164 & w1166;
assign v348 = ~(w288 | w566);
assign w1168 = v348;
assign w1169 = ~w359 & w1168;
assign v349 = ~(w216 | w272);
assign w1170 = v349;
assign v350 = ~(w135 | w456);
assign w1171 = v350;
assign w1172 = w1170 & w1171;
assign w1173 = w1169 & w1172;
assign w1174 = w1167 & w1173;
assign w1175 = w1163 & w1174;
assign w1176 = w476 & w1128;
assign v351 = ~(w123 | w387);
assign w1177 = v351;
assign v352 = ~(w266 | w274);
assign w1178 = v352;
assign v353 = ~(w299 | w405);
assign w1179 = v353;
assign w1180 = w1178 & w1179;
assign w1181 = w1177 & w1180;
assign w1182 = w1176 & w1181;
assign w1183 = w1042 & w1182;
assign w1184 = w1175 & w1183;
assign w1185 = w1160 & w1184;
assign v354 = ~(w134 | w656);
assign w1186 = v354;
assign w1187 = ~w128 & w1186;
assign v355 = ~(w63 | w525);
assign w1188 = v355;
assign v356 = ~(w286 | w503);
assign w1189 = v356;
assign w1190 = w1188 & w1189;
assign w1191 = ~w639 & w1190;
assign w1192 = w1187 & w1191;
assign w1193 = w30 & w72;
assign v357 = ~(w258 | w1193);
assign w1194 = v357;
assign v358 = ~(w259 | w303);
assign w1195 = v358;
assign v359 = ~(w21 | w404);
assign w1196 = v359;
assign w1197 = w1195 & w1196;
assign w1198 = w1194 & w1197;
assign w1199 = w1192 & w1198;
assign v360 = ~(w192 | w280);
assign w1200 = v360;
assign v361 = ~(w195 | w211);
assign w1201 = v361;
assign v362 = ~(w642 | w742);
assign w1202 = v362;
assign w1203 = ~w253 & w1202;
assign w1204 = w1201 & w1203;
assign v363 = ~(w267 | w381);
assign w1205 = v363;
assign w1206 = ~w481 & w1205;
assign w1207 = w28 & w149;
assign v364 = ~(w271 | w1207);
assign w1208 = v364;
assign w1209 = w1206 & w1208;
assign w1210 = w1204 & w1209;
assign w1211 = w1200 & w1210;
assign w1212 = w1199 & w1211;
assign w1213 = w1185 & w1212;
assign v365 = ~(w343 | w430);
assign w1214 = v365;
assign v366 = ~(w56 | w643);
assign w1215 = v366;
assign w1216 = w1214 & w1215;
assign w1217 = ~w90 & w1216;
assign v367 = ~(w277 | w338);
assign w1218 = v367;
assign w1219 = w802 & w977;
assign v368 = ~(w140 | w497);
assign w1220 = v368;
assign w1221 = w1219 & w1220;
assign w1222 = w1218 & w1221;
assign w1223 = w895 & w1222;
assign w1224 = w1217 & w1223;
assign v369 = ~(w454 | w613);
assign w1225 = v369;
assign v370 = ~(w374 | w581);
assign w1226 = v370;
assign w1227 = w1225 & w1226;
assign v371 = ~(w202 | w680);
assign w1228 = v371;
assign w1229 = w1029 & w1228;
assign w1230 = ~w316 & w1229;
assign w1231 = w1227 & w1230;
assign v372 = ~(w640 | w870);
assign w1232 = v372;
assign v373 = ~(w241 | w488);
assign w1233 = v373;
assign w1234 = ~w158 & w1233;
assign w1235 = ~w465 & w1234;
assign w1236 = w1232 & w1235;
assign w1237 = w1231 & w1236;
assign v374 = ~(w251 | w482);
assign w1238 = v374;
assign v375 = ~(w151 | w1134);
assign w1239 = v375;
assign v376 = ~(w209 | w877);
assign w1240 = v376;
assign w1241 = ~w685 & w1240;
assign v377 = ~(w428 | w758);
assign w1242 = v377;
assign w1243 = w109 & w1242;
assign w1244 = w1241 & w1243;
assign w1245 = w1239 & w1244;
assign w1246 = w1238 & w1245;
assign w1247 = w1237 & w1246;
assign w1248 = w1224 & w1247;
assign v378 = ~(w264 | w635);
assign w1249 = v378;
assign w1250 = ~w37 & w1249;
assign w1251 = ~w221 & w1250;
assign v379 = ~(w369 | w431);
assign w1252 = v379;
assign v380 = ~(w95 | w100);
assign w1253 = v380;
assign w1254 = w1252 & w1253;
assign w1255 = w1251 & w1254;
assign v381 = ~(w183 | w438);
assign w1256 = v381;
assign w1257 = w1255 & w1256;
assign v382 = ~(w110 | w127);
assign w1258 = v382;
assign v383 = ~(w812 | w822);
assign w1259 = v383;
assign w1260 = ~w312 & w1259;
assign w1261 = w859 & w1260;
assign v384 = ~(w200 | w292);
assign w1262 = v384;
assign v385 = ~(w65 | w278);
assign w1263 = v385;
assign v386 = ~(w77 | w533);
assign w1264 = v386;
assign w1265 = w1263 & w1264;
assign w1266 = w1262 & w1265;
assign w1267 = w1261 & w1266;
assign w1268 = w1258 & w1267;
assign w1269 = w1257 & w1268;
assign w1270 = w1248 & w1269;
assign w1271 = w1213 & w1270;
assign w1272 = w1153 & w1271;
assign v387 = ~(w1153 | w1271);
assign w1273 = v387;
assign v388 = ~(w1272 | w1273);
assign w1274 = v388;
assign w1275 = pi20 & w1274;
assign v389 = ~(w1272 | w1275);
assign w1276 = v389;
assign w1277 = w1055 & w1276;
assign v390 = ~(w1055 | w1276);
assign w1278 = v390;
assign v391 = ~(w1277 | w1278);
assign w1279 = v391;
assign v392 = ~(w216 | w258);
assign w1280 = v392;
assign w1281 = ~w192 & w1280;
assign w1282 = ~w605 & w1281;
assign v393 = ~(w374 | w465);
assign w1283 = v393;
assign v394 = ~(w200 | w652);
assign w1284 = v394;
assign w1285 = w1283 & w1284;
assign w1286 = w1282 & w1285;
assign v395 = ~(w291 | w548);
assign w1287 = v395;
assign v396 = ~(w337 | w541);
assign w1288 = v396;
assign w1289 = w1287 & w1288;
assign w1290 = ~w288 & w1289;
assign w1291 = w1286 & w1290;
assign v397 = ~(w37 | w666);
assign w1292 = v397;
assign v398 = ~(w277 | w400);
assign w1293 = v398;
assign w1294 = ~w418 & w1293;
assign w1295 = w1292 & w1294;
assign v399 = ~(w209 | w474);
assign w1296 = v399;
assign w1297 = w1064 & w1296;
assign v400 = ~(w140 | w758);
assign w1298 = v400;
assign w1299 = w1297 & w1298;
assign w1300 = w1295 & w1299;
assign v401 = ~(w329 | w978);
assign w1301 = v401;
assign w1302 = ~w251 & w1301;
assign v402 = ~(w593 | w886);
assign w1303 = v402;
assign w1304 = w91 & w1303;
assign w1305 = w1302 & w1304;
assign v403 = ~(w633 | w888);
assign w1306 = v403;
assign w1307 = ~w100 & w1306;
assign v404 = ~(w431 | w437);
assign w1308 = v404;
assign w1309 = ~w381 & w1308;
assign w1310 = w1307 & w1309;
assign w1311 = ~w281 & w1310;
assign w1312 = w1305 & w1311;
assign w1313 = w1300 & w1312;
assign w1314 = w1291 & w1313;
assign w1315 = w366 & ~w378;
assign v405 = ~(w73 | w274);
assign w1316 = v405;
assign w1317 = ~w692 & w1316;
assign w1318 = w1315 & w1317;
assign v406 = ~(w613 | w673);
assign w1319 = v406;
assign v407 = ~(w125 | w141);
assign w1320 = v407;
assign w1321 = w1319 & w1320;
assign v408 = ~(w21 | w388);
assign w1322 = v408;
assign v409 = ~(w531 | w588);
assign w1323 = v409;
assign w1324 = w1322 & w1323;
assign v410 = ~(w65 | w1207);
assign w1325 = v410;
assign v411 = ~(w176 | w753);
assign w1326 = v411;
assign w1327 = w1325 & w1326;
assign w1328 = w1324 & w1327;
assign w1329 = w1321 & w1328;
assign v412 = ~(w715 | w870);
assign w1330 = v412;
assign w1331 = ~w260 & w1330;
assign w1332 = ~w494 & w1331;
assign w1333 = w1329 & w1332;
assign w1334 = w1318 & w1333;
assign w1335 = w1314 & w1334;
assign v413 = ~(w499 | w812);
assign w1336 = v413;
assign v414 = ~(w131 | w384);
assign w1337 = v414;
assign w1338 = w1336 & w1337;
assign w1339 = w580 & w1338;
assign v415 = ~(w466 | w685);
assign w1340 = v415;
assign w1341 = ~w165 & w1340;
assign v416 = ~(w31 | w103);
assign w1342 = v416;
assign w1343 = w313 & w1342;
assign w1344 = w1341 & w1343;
assign v417 = ~(w220 | w385);
assign w1345 = v417;
assign w1346 = w152 & w1345;
assign w1347 = w1344 & w1346;
assign w1348 = w1339 & w1347;
assign v418 = ~(w49 | w111);
assign w1349 = v418;
assign w1350 = w1071 & w1349;
assign v419 = ~(w245 | w302);
assign w1351 = v419;
assign w1352 = ~w239 & w1351;
assign w1353 = w1350 & w1352;
assign w1354 = w977 & ~w989;
assign v420 = ~(w127 | w224);
assign w1355 = v420;
assign w1356 = w1354 & w1355;
assign w1357 = w1353 & w1356;
assign v421 = ~(w70 | w162);
assign w1358 = v421;
assign v422 = ~(w414 | w503);
assign w1359 = v422;
assign w1360 = w1358 & w1359;
assign w1361 = w676 & w1360;
assign w1362 = w1357 & w1361;
assign v423 = ~(w232 | w469);
assign w1363 = v423;
assign v424 = ~(w263 | w1032);
assign w1364 = v424;
assign w1365 = w318 & w1364;
assign v425 = ~(w430 | w482);
assign w1366 = v425;
assign w1367 = ~w194 & w1366;
assign w1368 = w1365 & w1367;
assign w1369 = w1363 & w1368;
assign v426 = ~(w822 | w877);
assign w1370 = v426;
assign v427 = ~(w186 | w266);
assign w1371 = v427;
assign v428 = ~(w387 | w564);
assign w1372 = v428;
assign w1373 = w1371 & w1372;
assign w1374 = w1370 & w1373;
assign w1375 = w213 & w1374;
assign w1376 = w1369 & w1375;
assign w1377 = w1362 & w1376;
assign v429 = ~(w462 | w945);
assign w1378 = v429;
assign w1379 = ~w68 & w1378;
assign w1380 = ~w191 & w1379;
assign v430 = ~(w248 | w892);
assign w1381 = v430;
assign w1382 = w1380 & w1381;
assign v431 = ~(w457 | w874);
assign w1383 = v431;
assign w1384 = w1382 & w1383;
assign w1385 = w1377 & w1384;
assign w1386 = w1348 & w1385;
assign w1387 = w1335 & w1386;
assign w1388 = w113 & ~w183;
assign w1389 = w801 & w1388;
assign v432 = ~(w373 | w414);
assign w1390 = v432;
assign w1391 = w534 & w1381;
assign w1392 = w1390 & w1391;
assign v433 = ~(w63 | w74);
assign w1393 = v433;
assign w1394 = w129 & w1393;
assign w1395 = w1392 & w1394;
assign v434 = ~(w220 | w488);
assign w1396 = v434;
assign w1397 = w641 & w1396;
assign v435 = ~(w410 | w711);
assign w1398 = v435;
assign w1399 = ~w595 & w1398;
assign w1400 = w767 & w1399;
assign w1401 = w1397 & w1400;
assign w1402 = w1395 & w1401;
assign w1403 = w1389 & w1402;
assign v436 = ~(w307 | w666);
assign w1404 = v436;
assign w1405 = ~w158 & w1404;
assign v437 = ~(w77 | w727);
assign w1406 = v437;
assign w1407 = w754 & w1406;
assign w1408 = w1405 & w1407;
assign v438 = ~(w68 | w241);
assign w1409 = v438;
assign w1410 = ~w541 & w1202;
assign w1411 = w1409 & w1410;
assign w1412 = w1408 & w1411;
assign v439 = ~(w271 | w874);
assign w1413 = v439;
assign v440 = ~(w448 | w749);
assign w1414 = v440;
assign v441 = ~(w282 | w494);
assign w1415 = v441;
assign w1416 = w1414 & w1415;
assign w1417 = w1413 & w1416;
assign v442 = ~(w169 | w558);
assign w1418 = v442;
assign w1419 = ~w252 & w1418;
assign w1420 = ~w21 & w1419;
assign w1421 = w1417 & w1420;
assign w1422 = w1412 & w1421;
assign v443 = ~(w103 | w277);
assign w1423 = v443;
assign v444 = ~(w37 | w530);
assign w1424 = v444;
assign v445 = ~(w274 | w465);
assign w1425 = v445;
assign w1426 = w1424 & w1425;
assign w1427 = w860 & w1426;
assign w1428 = ~w462 & w1427;
assign w1429 = w1423 & w1428;
assign w1430 = w1422 & w1429;
assign w1431 = w1403 & w1430;
assign v446 = ~(w259 | w1108);
assign w1432 = v446;
assign w1433 = ~w430 & w1432;
assign w1434 = w947 & w1433;
assign v447 = ~(w398 | w447);
assign w1435 = v447;
assign v448 = ~(w145 | w739);
assign w1436 = v448;
assign v449 = ~(w316 | w588);
assign w1437 = v449;
assign w1438 = w1436 & w1437;
assign w1439 = w1435 & w1438;
assign w1440 = w1434 & w1439;
assign w1441 = ~w131 & w1440;
assign v450 = ~(w132 | w300);
assign w1442 = v450;
assign w1443 = ~w343 & w1442;
assign v451 = ~(w27 | w247);
assign w1444 = v451;
assign w1445 = ~w201 & w1444;
assign w1446 = w1444 & w30772;
assign v452 = ~(w244 | w438);
assign w1447 = v452;
assign v453 = ~(w308 | w978);
assign w1448 = v453;
assign w1449 = w1447 & w1448;
assign w1450 = ~w497 & w1449;
assign w1451 = w1450 & w30773;
assign w1452 = ~w404 & w1228;
assign v454 = ~(w216 | w231);
assign w1453 = v454;
assign w1454 = ~w119 & w1453;
assign w1455 = w1452 & w1454;
assign w1456 = ~w999 & w1455;
assign w1457 = ~w870 & w1239;
assign w1458 = ~w400 & w1457;
assign w1459 = w1456 & w1458;
assign w1460 = w1451 & w1459;
assign w1461 = w1441 & w1460;
assign v455 = ~(w409 | w499);
assign w1462 = v455;
assign v456 = ~(w167 | w437);
assign w1463 = v456;
assign w1464 = w1462 & w1463;
assign v457 = ~(w49 | w209);
assign w1465 = v457;
assign v458 = ~(w311 | w484);
assign w1466 = v458;
assign w1467 = w1465 & w1466;
assign w1468 = w1464 & w1467;
assign w1469 = w109 & ~w264;
assign v459 = ~(w214 | w454);
assign w1470 = v459;
assign v460 = ~(w65 | w177);
assign w1471 = v460;
assign w1472 = w1470 & w1471;
assign w1473 = w1469 & w1472;
assign w1474 = w1468 & w1473;
assign v461 = ~(w42 | w456);
assign w1475 = v461;
assign v462 = ~(w176 | w195);
assign w1476 = v462;
assign w1477 = w1475 & w1476;
assign w1478 = w363 & w1477;
assign w1479 = w1298 & w1319;
assign w1480 = w1358 & w1479;
assign w1481 = w1478 & w1480;
assign w1482 = w1474 & w1481;
assign v463 = ~(w482 | w699);
assign w1483 = v463;
assign v464 = ~(w338 | w474);
assign w1484 = v464;
assign v465 = ~(w172 | w525);
assign w1485 = v465;
assign w1486 = w1484 & w1485;
assign w1487 = w383 & w1486;
assign v466 = ~(w251 | w457);
assign w1488 = v466;
assign w1489 = w786 & w1488;
assign v467 = ~(w388 | w997);
assign w1490 = v467;
assign w1491 = w1489 & w1490;
assign w1492 = w1487 & w1491;
assign w1493 = w1483 & w1492;
assign w1494 = w1482 & w1493;
assign w1495 = w1461 & w1494;
assign w1496 = w1431 & w1495;
assign v468 = ~(w1387 | w1496);
assign w1497 = v468;
assign w1498 = w1387 & w1496;
assign v469 = ~(w1497 | w1498);
assign w1499 = v469;
assign v470 = ~(w82 | w253);
assign w1500 = v470;
assign w1501 = ~w463 & w1500;
assign v471 = ~(w143 | w169);
assign w1502 = v471;
assign v472 = ~(w191 | w251);
assign w1503 = v472;
assign w1504 = w1502 & w1503;
assign w1505 = w1501 & w1504;
assign v473 = ~(w474 | w945);
assign w1506 = v473;
assign w1507 = w1226 & w1506;
assign v474 = ~(w42 | w135);
assign w1508 = v474;
assign w1509 = w336 & w1508;
assign w1510 = w1507 & w1509;
assign w1511 = w1505 & w1510;
assign v475 = ~(w428 | w888);
assign w1512 = v475;
assign w1513 = ~w209 & w1512;
assign w1514 = ~w220 & w1513;
assign w1515 = ~w215 & w1228;
assign w1516 = w1514 & w1515;
assign w1517 = w1511 & w1516;
assign w1518 = w632 & w1517;
assign w1519 = ~w248 & w1049;
assign v476 = ~(w112 | w231);
assign w1520 = v476;
assign v477 = ~(w326 | w409);
assign w1521 = v477;
assign w1522 = w1520 & w1521;
assign w1523 = w1120 & w1522;
assign w1524 = w1519 & w1523;
assign w1525 = ~w711 & w1524;
assign w1526 = ~w93 & w1040;
assign w1527 = w1355 & w1526;
assign w1528 = w1525 & w1527;
assign v478 = ~(w422 | w892);
assign w1529 = v478;
assign v479 = ~(w235 | w497);
assign w1530 = v479;
assign w1531 = w1529 & w1530;
assign w1532 = w1528 & w1531;
assign w1533 = w1518 & w1532;
assign v480 = ~(w566 | w643);
assign w1534 = v480;
assign v481 = ~(w239 | w1207);
assign w1535 = v481;
assign v482 = ~(w437 | w874);
assign w1536 = v482;
assign w1537 = ~w447 & w1536;
assign w1538 = ~w997 & w1537;
assign w1539 = w1535 & w1538;
assign w1540 = w1534 & w1539;
assign v483 = ~(w484 | w584);
assign w1541 = v483;
assign v484 = ~(w385 | w465);
assign w1542 = v484;
assign w1543 = w1541 & w1542;
assign w1544 = w313 & w894;
assign w1545 = w1543 & w1544;
assign v485 = ~(w21 | w541);
assign w1546 = v485;
assign v486 = ~(w208 | w595);
assign w1547 = v486;
assign w1548 = w1546 & w1547;
assign w1549 = w1545 & w1548;
assign v487 = ~(w65 | w1032);
assign w1550 = v487;
assign w1551 = ~w68 & w1550;
assign v488 = ~(w247 | w398);
assign w1552 = v488;
assign w1553 = w1551 & w1552;
assign w1554 = ~w292 & w1553;
assign w1555 = w1549 & w1554;
assign w1556 = w1540 & w1555;
assign v489 = ~(w378 | w812);
assign w1557 = v489;
assign w1558 = w213 & w1557;
assign v490 = ~(w158 | w427);
assign w1559 = v490;
assign w1560 = ~w697 & w1559;
assign w1561 = ~w456 & w1560;
assign w1562 = ~w271 & w1561;
assign v491 = ~(w39 | w48);
assign w1563 = v491;
assign w1564 = w50 & ~w1563;
assign w1565 = w1086 & ~w1564;
assign w1566 = w1562 & w1565;
assign w1567 = w1558 & w1566;
assign w1568 = w1556 & w1567;
assign w1569 = w126 & w1135;
assign w1570 = ~w95 & w1569;
assign v492 = ~(w51 | w216);
assign w1571 = v492;
assign w1572 = w1570 & w1571;
assign w1573 = ~w223 & w634;
assign v493 = ~(w186 | w479);
assign w1574 = v493;
assign v494 = ~(w108 | w441);
assign w1575 = v494;
assign w1576 = w1574 & w1575;
assign w1577 = w1573 & w1576;
assign w1578 = w1127 & w1577;
assign w1579 = w1572 & w1578;
assign w1580 = ~w499 & w1340;
assign v495 = ~(w162 | w673);
assign w1581 = v495;
assign v496 = ~(w278 | w488);
assign w1582 = v496;
assign w1583 = w1581 & w1582;
assign w1584 = w1580 & w1583;
assign w1585 = ~w373 & w1584;
assign v497 = ~(w98 | w381);
assign w1586 = v497;
assign v498 = ~(w183 | w200);
assign w1587 = v498;
assign v499 = ~(w177 | w559);
assign w1588 = v499;
assign w1589 = w366 & w1588;
assign w1590 = w1587 & w1589;
assign w1591 = w1586 & w1590;
assign w1592 = w1585 & w1591;
assign w1593 = ~w404 & w1447;
assign v500 = ~(w359 | w715);
assign w1594 = v500;
assign v501 = ~(w176 | w822);
assign w1595 = v501;
assign w1596 = w1594 & w1595;
assign v502 = ~(w100 | w353);
assign w1597 = v502;
assign w1598 = w1596 & w1597;
assign w1599 = w1593 & w1598;
assign v503 = ~(w299 | w727);
assign w1600 = v503;
assign w1601 = ~w674 & w1600;
assign w1602 = ~w370 & w1601;
assign v504 = ~(w27 | w324);
assign w1603 = v504;
assign w1604 = w1602 & w1603;
assign w1605 = w1599 & w1604;
assign w1606 = w1592 & w1605;
assign w1607 = w1579 & w1606;
assign w1608 = w1568 & w1607;
assign w1609 = w1533 & w1608;
assign v505 = ~(w1496 | w1609);
assign w1610 = v505;
assign w1611 = w1496 & w1609;
assign w1612 = ~w73 & w1093;
assign v506 = ~(w493 | w652);
assign w1613 = v506;
assign w1614 = w1529 & w1613;
assign v507 = ~(w267 | w505);
assign w1615 = v507;
assign w1616 = ~w271 & w1615;
assign w1617 = w1614 & w1616;
assign v508 = ~(w212 | w484);
assign w1618 = v508;
assign v509 = ~(w42 | w874);
assign w1619 = v509;
assign v510 = ~(w194 | w541);
assign w1620 = v510;
assign w1621 = w1619 & w1620;
assign w1622 = w1618 & w1621;
assign w1623 = w1617 & w1622;
assign w1624 = ~w522 & w1418;
assign v511 = ~(w100 | w303);
assign w1625 = v511;
assign w1626 = ~w697 & w1625;
assign w1627 = w1624 & w1626;
assign w1628 = w898 & w1627;
assign w1629 = w1623 & w1628;
assign w1630 = w1612 & w1629;
assign w1631 = ~w93 & w725;
assign v512 = ~(w232 | w425);
assign w1632 = v512;
assign w1633 = ~w642 & w1632;
assign w1634 = w1631 & w1633;
assign w1635 = w1114 & w1634;
assign v513 = ~(w215 | w643);
assign w1636 = v513;
assign w1637 = ~w151 & w1636;
assign w1638 = w953 & w1637;
assign w1639 = w1490 & w1638;
assign w1640 = w1635 & w1639;
assign v514 = ~(w379 | w525);
assign w1641 = v514;
assign v515 = ~(w457 | w1134);
assign w1642 = v515;
assign w1643 = w1641 & w1642;
assign w1644 = w1142 & w1643;
assign w1645 = w1640 & w1644;
assign w1646 = w1630 & w1645;
assign v516 = ~(w176 | w266);
assign w1647 = v516;
assign w1648 = w883 & w1252;
assign w1649 = w1647 & w1648;
assign v517 = ~(w629 | w715);
assign w1650 = v517;
assign w1651 = ~w338 & w1650;
assign w1652 = w1649 & w1651;
assign v518 = ~(w633 | w673);
assign w1653 = v518;
assign v519 = ~(w466 | w548);
assign w1654 = v519;
assign w1655 = ~w282 & w1654;
assign w1656 = w1653 & w1655;
assign v520 = ~(w329 | w441);
assign w1657 = v520;
assign w1658 = ~w405 & w1657;
assign w1659 = w1656 & w1658;
assign v521 = ~(w123 | w1207);
assign w1660 = v521;
assign v522 = ~(w481 | w989);
assign w1661 = v522;
assign w1662 = ~w107 & w1661;
assign w1663 = w1660 & w1662;
assign v523 = ~(w324 | w1032);
assign w1664 = v523;
assign w1665 = w146 & w1664;
assign v524 = ~(w179 | w238);
assign w1666 = v524;
assign v525 = ~(w201 | w418);
assign w1667 = v525;
assign w1668 = w1666 & w1667;
assign w1669 = w1665 & w1668;
assign w1670 = w1663 & w1669;
assign w1671 = w1659 & w1670;
assign w1672 = w1652 & w1671;
assign w1673 = w604 & w1672;
assign w1674 = w1646 & w1673;
assign v526 = ~(w1609 | w1674);
assign w1675 = v526;
assign w1676 = w1609 & w1674;
assign v527 = ~(w629 | w666);
assign w1677 = v527;
assign w1678 = w982 & w1677;
assign v528 = ~(w88 | w989);
assign w1679 = v528;
assign w1680 = ~w53 & w1679;
assign v529 = ~(w299 | w400);
assign w1681 = v529;
assign v530 = ~(w131 | w195);
assign w1682 = v530;
assign w1683 = w1681 & w1682;
assign v531 = ~(w425 | w892);
assign w1684 = v531;
assign w1685 = w1177 & w1684;
assign w1686 = w1683 & w1685;
assign w1687 = w1680 & w1686;
assign w1688 = w1678 & w1687;
assign v532 = ~(w303 | w410);
assign w1689 = v532;
assign v533 = ~(w258 | w462);
assign w1690 = v533;
assign w1691 = w1689 & w1690;
assign w1692 = w965 & w1691;
assign v534 = ~(w183 | w211);
assign w1693 = v534;
assign w1694 = w1041 & w1693;
assign w1695 = w1692 & w1694;
assign w1696 = w328 & ~w385;
assign w1697 = w1695 & w1696;
assign w1698 = w1688 & w1697;
assign v535 = ~(w108 | w372);
assign w1699 = v535;
assign w1700 = w900 & w1699;
assign w1701 = w1352 & w1700;
assign w1702 = ~w200 & w1701;
assign w1703 = ~w888 & w1702;
assign w1704 = w1698 & w1703;
assign w1705 = ~w287 & w1704;
assign v536 = ~(w132 | w674);
assign w1706 = v536;
assign w1707 = ~w558 & w1706;
assign v537 = ~(w162 | w422);
assign w1708 = v537;
assign w1709 = w967 & w1708;
assign v538 = ~(w266 | w378);
assign w1710 = v538;
assign v539 = ~(w247 | w749);
assign w1711 = v539;
assign w1712 = w1710 & w1711;
assign w1713 = w1709 & w1712;
assign w1714 = w1707 & w1713;
assign w1715 = w335 & ~w343;
assign v540 = ~(w134 | w300);
assign w1716 = v540;
assign w1717 = ~w165 & w1716;
assign v541 = ~(w605 | w1108);
assign w1718 = v541;
assign w1719 = w1717 & w1718;
assign w1720 = w1715 & w1719;
assign w1721 = w1714 & w1720;
assign v542 = ~(w430 | w533);
assign w1722 = v542;
assign w1723 = ~w870 & w1722;
assign w1724 = ~w337 & w1396;
assign w1725 = w1723 & w1724;
assign v543 = ~(w307 | w317);
assign w1726 = v543;
assign w1727 = w1425 & w1726;
assign w1728 = ~w822 & w1727;
assign v544 = ~(w223 | w277);
assign w1729 = v544;
assign v545 = ~(w232 | w564);
assign w1730 = v545;
assign w1731 = w1161 & w1730;
assign w1732 = w1729 & w1731;
assign w1733 = w1728 & w1732;
assign w1734 = w1725 & w1733;
assign w1735 = w1721 & w1734;
assign v546 = ~(w77 | w248);
assign w1736 = v546;
assign w1737 = ~w103 & w1325;
assign v547 = ~(w405 | w697);
assign w1738 = v547;
assign w1739 = w835 & w1738;
assign w1740 = w1737 & w1739;
assign v548 = ~(w93 | w685);
assign w1741 = v548;
assign w1742 = ~w150 & w1741;
assign v549 = ~(w438 | w550);
assign w1743 = v549;
assign w1744 = ~w499 & w1743;
assign w1745 = w1742 & w1744;
assign w1746 = w1740 & w1745;
assign w1747 = w1736 & w1746;
assign w1748 = w1228 & w29637;
assign w1749 = ~w640 & w1748;
assign w1750 = w1747 & w1749;
assign w1751 = w1735 & w1750;
assign w1752 = ~w503 & w814;
assign w1753 = ~w282 & w1752;
assign v550 = ~(w42 | w291);
assign w1754 = v550;
assign w1755 = ~w110 & w1754;
assign w1756 = w1753 & w1755;
assign w1757 = w1751 & w1756;
assign w1758 = w1705 & w1757;
assign v551 = ~(w563 | w999);
assign w1759 = v551;
assign w1760 = ~w90 & w1759;
assign v552 = ~(w278 | w886);
assign w1761 = v552;
assign w1762 = w1760 & w1761;
assign w1763 = ~w404 & w1762;
assign v553 = ~(w100 | w224);
assign w1764 = v553;
assign v554 = ~(w177 | w874);
assign w1765 = v554;
assign w1766 = w839 & w1765;
assign v555 = ~(w135 | w271);
assign w1767 = v555;
assign v556 = ~(w409 | w559);
assign w1768 = v556;
assign w1769 = w1767 & w1768;
assign w1770 = w1766 & w1769;
assign v557 = ~(w441 | w727);
assign w1771 = v557;
assign v558 = ~(w49 | w172);
assign w1772 = v558;
assign w1773 = w121 & w1772;
assign w1774 = w1771 & w1773;
assign w1775 = w1770 & w1774;
assign w1776 = ~w231 & w1202;
assign w1777 = w1666 & w1776;
assign w1778 = w1775 & w1777;
assign w1779 = w1764 & w1778;
assign v559 = ~(w194 | w481);
assign w1780 = v559;
assign v560 = ~(w447 | w711);
assign w1781 = v560;
assign w1782 = ~w652 & w1781;
assign w1783 = w726 & ~w945;
assign w1784 = w1782 & w1783;
assign w1785 = w1780 & w1784;
assign v561 = ~(w286 | w739);
assign w1786 = v561;
assign w1787 = ~w252 & w1786;
assign v562 = ~(w98 | w463);
assign w1788 = v562;
assign w1789 = ~w209 & w585;
assign w1790 = w1788 & w1789;
assign w1791 = w1787 & w1790;
assign w1792 = w1785 & w1791;
assign w1793 = w1779 & w1792;
assign w1794 = w1763 & w1793;
assign w1795 = w1758 & w1794;
assign v563 = ~(w1674 | w1795);
assign w1796 = v563;
assign w1797 = w1674 & w1795;
assign v564 = ~(w1796 | w1797);
assign w1798 = v564;
assign v565 = ~(w78 | w186);
assign w1799 = v565;
assign w1800 = w1340 & w1388;
assign w1801 = w1799 & w1800;
assign v566 = ~(w438 | w749);
assign w1802 = v566;
assign w1803 = ~w564 & w1802;
assign w1804 = w1445 & w1803;
assign v567 = ~(w90 | w324);
assign w1805 = v567;
assign w1806 = ~w326 & w1805;
assign v568 = ~(w454 | w558);
assign w1807 = v568;
assign w1808 = w1806 & w1807;
assign w1809 = w1804 & w1808;
assign w1810 = w1801 & w1809;
assign v569 = ~(w373 | w451);
assign w1811 = v569;
assign w1812 = ~w132 & w1811;
assign w1813 = ~w167 & w1812;
assign v570 = ~(w484 | w639);
assign w1814 = v570;
assign w1815 = w1018 & w1814;
assign v571 = ~(w370 | w404);
assign w1816 = v571;
assign w1817 = w1815 & w1816;
assign w1818 = w893 & w1817;
assign w1819 = w1813 & w1818;
assign w1820 = w1810 & w1819;
assign v572 = ~(w422 | w448);
assign w1821 = v572;
assign w1822 = w1727 & w28151;
assign v573 = ~(w251 | w258);
assign w1823 = v573;
assign w1824 = w1560 & w1823;
assign w1825 = w1822 & w1824;
assign v574 = ~(w457 | w563);
assign w1826 = v574;
assign w1827 = ~w593 & w1826;
assign v575 = ~(w95 | w299);
assign w1828 = v575;
assign w1829 = ~w469 & w1828;
assign w1830 = w1827 & w1829;
assign v576 = ~(w629 | w633);
assign w1831 = v576;
assign v577 = ~(w144 | w272);
assign w1832 = v577;
assign w1833 = w1831 & w1832;
assign w1834 = w1830 & w1833;
assign w1835 = w1753 & w1834;
assign w1836 = w1825 & w1835;
assign w1837 = w544 & w1087;
assign w1838 = w193 & ~w522;
assign w1839 = w1837 & w1838;
assign v578 = ~(w214 | w252);
assign w1840 = v578;
assign w1841 = w225 & w1840;
assign w1842 = w859 & w894;
assign w1843 = w1039 & w1842;
assign w1844 = w1841 & w1843;
assign w1845 = w1320 & w1844;
assign w1846 = w1839 & w1845;
assign w1847 = w1836 & w1846;
assign v579 = ~(w337 | w505);
assign w1848 = v579;
assign w1849 = w1168 & w1848;
assign v580 = ~(w308 | w899);
assign w1850 = v580;
assign w1851 = w1484 & w1850;
assign w1852 = w1849 & w1851;
assign v581 = ~(w642 | w731);
assign w1853 = v581;
assign v582 = ~(w53 | w494);
assign w1854 = v582;
assign w1855 = w1853 & w1854;
assign w1856 = ~w107 & w1855;
assign w1857 = w1852 & w1856;
assign w1858 = w958 & w1857;
assign w1859 = w1847 & w1858;
assign w1860 = w1820 & w1859;
assign v583 = ~(w1795 | w1860);
assign w1861 = v583;
assign w1862 = w1795 & w1860;
assign v584 = ~(w1861 | w1862);
assign w1863 = v584;
assign v585 = ~(w291 | w457);
assign w1864 = v585;
assign w1865 = w1284 & w1864;
assign w1866 = w779 & w1865;
assign w1867 = w881 & w1866;
assign v586 = ~(w187 | w258);
assign w1868 = v586;
assign v587 = ~(w186 | w564);
assign w1869 = v587;
assign v588 = ~(w378 | w390);
assign w1870 = v588;
assign w1871 = w1869 & w1870;
assign w1872 = w1542 & w1871;
assign w1873 = w1868 & w1872;
assign w1874 = w1867 & w1873;
assign v589 = ~(w179 | w945);
assign w1875 = v589;
assign w1876 = ~w430 & w1875;
assign v590 = ~(w400 | w503);
assign w1877 = v590;
assign v591 = ~(w280 | w282);
assign w1878 = v591;
assign w1879 = w1877 & w1878;
assign w1880 = w1876 & w1879;
assign w1881 = w1397 & w1880;
assign w1882 = w1600 & w1881;
assign w1883 = w1874 & w1882;
assign w1884 = w109 & ~w274;
assign w1885 = w1841 & w1884;
assign v592 = ~(w260 | w505);
assign w1886 = v592;
assign w1887 = ~w497 & w1886;
assign v593 = ~(w259 | w410);
assign w1888 = v593;
assign w1889 = ~w316 & w1888;
assign w1890 = w1887 & w1889;
assign w1891 = w1885 & w1890;
assign v594 = ~(w184 | w241);
assign w1892 = v594;
assign v595 = ~(w82 | w99);
assign w1893 = v595;
assign w1894 = ~w21 & w1893;
assign w1895 = w1892 & w1894;
assign v596 = ~(w373 | w494);
assign w1896 = v596;
assign w1897 = ~w120 & w1896;
assign w1898 = w1895 & w1897;
assign w1899 = w585 & w1898;
assign w1900 = w1891 & w1899;
assign w1901 = w1883 & w1900;
assign v597 = ~(w37 | w531);
assign w1902 = v597;
assign v598 = ~(w53 | w630);
assign w1903 = v598;
assign w1904 = w1902 & w1903;
assign v599 = ~(w431 | w581);
assign w1905 = v599;
assign v600 = ~(w78 | w441);
assign w1906 = v600;
assign w1907 = w545 & w1906;
assign w1908 = w1905 & w1907;
assign w1909 = w1904 & w1908;
assign w1910 = w1908 & w30774;
assign v601 = ~(w131 | w633);
assign w1911 = v601;
assign v602 = ~(w183 | w215);
assign w1912 = v602;
assign v603 = ~(w63 | w119);
assign w1913 = v603;
assign w1914 = ~w127 & w1913;
assign w1915 = w1912 & w1914;
assign v604 = ~(w135 | w559);
assign w1916 = v604;
assign w1917 = w1914 & w30775;
assign w1918 = w1911 & w1917;
assign w1919 = w1910 & w1918;
assign v605 = ~(w123 | w475);
assign w1920 = v605;
assign w1921 = ~w201 & w1920;
assign w1922 = w1502 & w1805;
assign w1923 = w1161 & w1922;
assign w1924 = ~w238 & w857;
assign w1925 = w1923 & w1924;
assign w1926 = w1921 & w1925;
assign w1927 = w1919 & w1926;
assign v606 = ~(w42 | w1108);
assign w1928 = v606;
assign w1929 = w142 & w1928;
assign v607 = ~(w286 | w812);
assign w1930 = v607;
assign w1931 = ~w566 & w1930;
assign w1932 = w1056 & w1931;
assign w1933 = w1929 & w1932;
assign v608 = ~(w167 | w888);
assign w1934 = v608;
assign v609 = ~(w159 | w588);
assign w1935 = v609;
assign w1936 = w419 & w1935;
assign w1937 = w1934 & w1936;
assign w1938 = w96 & w1937;
assign w1939 = ~w244 & w1938;
assign w1940 = w1933 & w1939;
assign w1941 = w1927 & w1940;
assign w1942 = w1901 & w1941;
assign v610 = ~(w1860 | w1942);
assign w1943 = v610;
assign w1944 = w1860 & w1942;
assign v611 = ~(w167 | w531);
assign w1945 = v611;
assign w1946 = w1853 & w1945;
assign v612 = ~(w329 | w530);
assign w1947 = v612;
assign w1948 = w1878 & w1947;
assign w1949 = w1946 & w1948;
assign w1950 = w1138 & w1949;
assign v613 = ~(w886 | w1207);
assign w1951 = v613;
assign w1952 = w972 & w1951;
assign v614 = ~(w274 | w479);
assign w1953 = v614;
assign w1954 = w1952 & w1953;
assign v615 = ~(w134 | w588);
assign w1955 = v615;
assign w1956 = ~w287 & w1955;
assign w1957 = ~w822 & w1956;
assign w1958 = w1954 & w1957;
assign w1959 = ~w656 & w1500;
assign v616 = ~(w159 | w208);
assign w1960 = v616;
assign w1961 = w1959 & w1960;
assign w1962 = w348 & w1961;
assign w1963 = w1958 & w1962;
assign w1964 = w1950 & w1963;
assign v617 = ~(w42 | w369);
assign w1965 = v617;
assign v618 = ~(w93 | w633);
assign w1966 = v618;
assign w1967 = w1965 & w1966;
assign w1968 = ~w316 & w783;
assign w1969 = ~w311 & w1968;
assign w1970 = w1967 & w1969;
assign v619 = ~(w307 | w593);
assign w1971 = v619;
assign w1972 = w675 & w1971;
assign w1973 = w1666 & w1972;
assign v620 = ~(w462 | w989);
assign w1974 = v620;
assign w1975 = w933 & w1974;
assign w1976 = ~w90 & w358;
assign w1977 = w1975 & w1976;
assign w1978 = w1973 & w1977;
assign w1979 = w1080 & w1978;
assign v621 = ~(w308 | w630);
assign w1980 = v621;
assign w1981 = ~w673 & w1980;
assign w1982 = w1001 & w1981;
assign w1983 = w1801 & w1982;
assign w1984 = w1979 & w1983;
assign w1985 = w1970 & w1984;
assign v622 = ~(w231 | w278);
assign w1986 = v622;
assign w1987 = w325 & w1986;
assign w1988 = ~w427 & w1987;
assign v623 = ~(w758 | w812);
assign w1989 = v623;
assign w1990 = ~w666 & w1989;
assign v624 = ~(w180 | w456);
assign w1991 = v624;
assign w1992 = w1588 & w1991;
assign w1993 = w1990 & w1992;
assign w1994 = w1988 & w1993;
assign v625 = ~(w187 | w373);
assign w1995 = v625;
assign v626 = ~(w68 | w212);
assign w1996 = v626;
assign w1997 = ~w150 & w1996;
assign w1998 = w1995 & w1997;
assign w1999 = w419 & w1447;
assign w2000 = ~w414 & w1999;
assign w2001 = w1998 & w2000;
assign w2002 = w1994 & w2001;
assign v627 = ~(w281 | w384);
assign w2003 = v627;
assign v628 = ~(w88 | w400);
assign w2004 = v628;
assign w2005 = w2003 & w2004;
assign v629 = ~(w288 | w550);
assign w2006 = v629;
assign w2007 = ~w132 & w2006;
assign w2008 = w2005 & w2007;
assign v630 = ~(w385 | w541);
assign w2009 = v630;
assign v631 = ~(w640 | w1108);
assign w2010 = v631;
assign w2011 = w2009 & w2010;
assign w2012 = w2008 & w2011;
assign v632 = ~(w144 | w381);
assign w2013 = v632;
assign w2014 = ~w420 & w2013;
assign v633 = ~(w581 | w899);
assign w2015 = v633;
assign v634 = ~(w191 | w259);
assign w2016 = v634;
assign w2017 = w2015 & w2016;
assign w2018 = w2014 & w2017;
assign w2019 = ~w945 & w2018;
assign w2020 = w2012 & w2019;
assign w2021 = w2002 & w2020;
assign v635 = ~(w176 | w629);
assign w2022 = v635;
assign w2023 = ~w309 & w2022;
assign v636 = ~(w100 | w202);
assign w2024 = v636;
assign w2025 = ~w605 & w2024;
assign w2026 = ~w107 & w2025;
assign v637 = ~(w264 | w266);
assign w2027 = v637;
assign v638 = ~(w65 | w277);
assign w2028 = v638;
assign w2029 = w225 & w2028;
assign w2030 = w2027 & w2029;
assign w2031 = w2026 & w2030;
assign w2032 = w2023 & w2031;
assign v639 = ~(w359 | w503);
assign w2033 = v639;
assign w2034 = w1773 & w2033;
assign w2035 = w2032 & w2034;
assign w2036 = w2021 & w2035;
assign w2037 = w1985 & w2036;
assign w2038 = w1964 & w2037;
assign v640 = ~(w1942 | w2038);
assign w2039 = v640;
assign w2040 = w1942 & w2038;
assign v641 = ~(w2039 | w2040);
assign w2041 = v641;
assign w2042 = ~w267 & w872;
assign v642 = ~(w292 | w497);
assign w2043 = v642;
assign w2044 = w72 & w122;
assign v643 = ~(w437 | w2044);
assign w2045 = v643;
assign w2046 = ~w533 & w2045;
assign w2047 = w2043 & w2046;
assign w2048 = w2042 & w2047;
assign v644 = ~(w251 | w692);
assign w2049 = v644;
assign v645 = ~(w212 | w1032);
assign w2050 = v645;
assign w2051 = ~w899 & w2050;
assign v646 = ~(w173 | w877);
assign w2052 = v646;
assign v647 = ~(w425 | w474);
assign w2053 = v647;
assign w2054 = w2052 & w2053;
assign w2055 = w2051 & w2054;
assign w2056 = w2049 & w2055;
assign w2057 = w708 & w2056;
assign w2058 = w2048 & w2057;
assign w2059 = w1807 & w2058;
assign v648 = ~(w324 | w405);
assign w2060 = v648;
assign w2061 = ~w74 & w2060;
assign w2062 = w1322 & w1995;
assign w2063 = w582 & w2062;
assign w2064 = ~w239 & w2063;
assign w2065 = w2061 & w2064;
assign w2066 = ~w151 & w1792;
assign w2067 = w2065 & w2066;
assign w2068 = w2059 & w2067;
assign v649 = ~(w274 | w288);
assign w2069 = v649;
assign w2070 = w1731 & w27992;
assign w2071 = ~w216 & w1853;
assign w2072 = w641 & w2071;
assign w2073 = w1667 & w1892;
assign w2074 = w2072 & w2073;
assign w2075 = w2070 & w2074;
assign v650 = ~(w144 | w479);
assign w2076 = v650;
assign w2077 = ~w63 & w2076;
assign v651 = ~(w525 | w699);
assign w2078 = v651;
assign v652 = ~(w329 | w493);
assign w2079 = v652;
assign w2080 = w2078 & w2079;
assign w2081 = w2077 & w2080;
assign v653 = ~(w550 | w697);
assign w2082 = v653;
assign v654 = ~(w430 | w448);
assign w2083 = v654;
assign w2084 = w2082 & w2083;
assign w2085 = w2081 & w27993;
assign w2086 = w2075 & w2085;
assign w2087 = w1775 & w2086;
assign w2088 = w1985 & w2087;
assign w2089 = w2068 & w2088;
assign w2090 = w2038 & w2089;
assign v655 = ~(w2038 | w2089);
assign w2091 = v655;
assign v656 = ~(w119 | w271);
assign w2092 = v656;
assign w2093 = w1738 & w2092;
assign v657 = ~(w169 | w291);
assign w2094 = v657;
assign v658 = ~(w186 | w202);
assign w2095 = v658;
assign w2096 = w2094 & w2095;
assign w2097 = ~w715 & w2096;
assign w2098 = w2093 & w2097;
assign v659 = ~(w331 | w874);
assign w2099 = v659;
assign v660 = ~(w385 | w699);
assign w2100 = v660;
assign v661 = ~(w179 | w613);
assign w2101 = v661;
assign w2102 = w2100 & w2101;
assign w2103 = ~w267 & w2102;
assign w2104 = w2099 & w2103;
assign w2105 = w2098 & w2104;
assign w2106 = w752 & w2105;
assign v662 = ~(w428 | w475);
assign w2107 = v662;
assign v663 = ~(w160 | w324);
assign w2108 = v663;
assign v664 = ~(w563 | w581);
assign w2109 = v664;
assign w2110 = w2108 & w2109;
assign w2111 = w2107 & w2110;
assign w2112 = w1692 & w2111;
assign w2113 = w2071 & w2112;
assign w2114 = w2106 & w2113;
assign w2115 = w362 & ~w369;
assign w2116 = w681 & w2115;
assign v665 = ~(w300 | w643);
assign w2117 = v665;
assign w2118 = w657 & w759;
assign v666 = ~(w78 | w624);
assign w2119 = v666;
assign w2120 = ~w674 & w2119;
assign w2121 = w2118 & w2120;
assign w2122 = w2117 & w2121;
assign w2123 = w2116 & w2122;
assign v667 = ~(w184 | w525);
assign w2124 = v667;
assign w2125 = w442 & w2124;
assign w2126 = ~w176 & w2125;
assign v668 = ~(w191 | w503);
assign w2127 = v668;
assign w2128 = w213 & w2127;
assign w2129 = w1388 & w2128;
assign w2130 = w2126 & w2129;
assign v669 = ~(w70 | w173);
assign w2131 = v669;
assign w2132 = w2130 & w2131;
assign w2133 = w2123 & w2132;
assign v670 = ~(w158 | w886);
assign w2134 = v670;
assign w2135 = w802 & w2134;
assign w2136 = ~w1207 & w1680;
assign w2137 = w2135 & w2136;
assign v671 = ~(w414 | w629);
assign w2138 = v671;
assign v672 = ~(w99 | w266);
assign w2139 = v672;
assign w2140 = w2138 & w2139;
assign v673 = ~(w214 | w309);
assign w2141 = v673;
assign v674 = ~(w127 | w277);
assign w2142 = v674;
assign w2143 = w2141 & w2142;
assign w2144 = w2140 & w2143;
assign w2145 = w1743 & w2144;
assign w2146 = w2137 & w2145;
assign v675 = ~(w145 | w427);
assign w2147 = v675;
assign v676 = ~(w252 | w877);
assign w2148 = v676;
assign w2149 = w2147 & w2148;
assign w2150 = w1381 & w2149;
assign w2151 = w348 & w360;
assign w2152 = w2150 & w2151;
assign w2153 = w2146 & w2152;
assign w2154 = w2133 & w2153;
assign w2155 = ~w231 & w2154;
assign v677 = ~(w159 | w272);
assign w2156 = v677;
assign w2157 = ~w640 & w2156;
assign v678 = ~(w93 | w278);
assign w2158 = v678;
assign w2159 = ~w463 & w2158;
assign v679 = ~(w167 | w605);
assign w2160 = v679;
assign w2161 = w1165 & w2160;
assign w2162 = w2159 & w2161;
assign v680 = ~(w379 | w381);
assign w2163 = v680;
assign v681 = ~(w326 | w338);
assign w2164 = v681;
assign w2165 = w2163 & w2164;
assign w2166 = ~w27 & w2165;
assign w2167 = w2162 & w2166;
assign w2168 = w2157 & w2167;
assign v682 = ~(w68 | w374);
assign w2169 = v682;
assign w2170 = w1060 & w2169;
assign w2171 = ~w107 & w2170;
assign w2172 = w2168 & w2171;
assign v683 = ~(w253 | w685);
assign w2173 = v683;
assign w2174 = ~w390 & w2173;
assign w2175 = ~w245 & w2174;
assign v684 = ~(w192 | w298);
assign w2176 = v684;
assign v685 = ~(w388 | w409);
assign w2177 = v685;
assign w2178 = w2176 & w2177;
assign w2179 = w2175 & w2178;
assign v686 = ~(w125 | w548);
assign w2180 = v686;
assign v687 = ~(w194 | w244);
assign w2181 = v687;
assign v688 = ~(w239 | w418);
assign w2182 = v688;
assign w2183 = w2181 & w2182;
assign w2184 = w2180 & w2183;
assign v689 = ~(w400 | w505);
assign w2185 = v689;
assign v690 = ~(w263 | w564);
assign w2186 = v690;
assign w2187 = ~w220 & w2186;
assign v691 = ~(w56 | w343);
assign w2188 = v691;
assign w2189 = w2187 & w30776;
assign w2190 = w2184 & w2189;
assign w2191 = w2179 & w2190;
assign w2192 = w2172 & w2191;
assign v692 = ~(w448 | w742);
assign w2193 = v692;
assign w2194 = ~w100 & w2193;
assign w2195 = w1971 & w2194;
assign v693 = ~(w172 | w812);
assign w2196 = v693;
assign w2197 = w800 & w2196;
assign w2198 = ~w666 & w2197;
assign w2199 = w2195 & w2198;
assign w2200 = w2192 & w2199;
assign w2201 = w2155 & w2200;
assign w2202 = w2114 & w2201;
assign v694 = ~(w2089 | w2202);
assign w2203 = v694;
assign w2204 = ~w95 & w864;
assign w2205 = ~w390 & w2204;
assign w2206 = ~w112 & w887;
assign v695 = ~(w309 | w1108);
assign w2207 = v695;
assign w2208 = w1157 & w2207;
assign w2209 = w2206 & w2208;
assign v696 = ~(w21 | w1032);
assign w2210 = v696;
assign w2211 = w2046 & w2210;
assign w2212 = w2209 & w2211;
assign w2213 = w2205 & w2212;
assign v697 = ~(w88 | w103);
assign w2214 = v697;
assign w2215 = w2014 & w2214;
assign w2216 = w225 & w551;
assign w2217 = ~w425 & w752;
assign w2218 = w2216 & w2217;
assign w2219 = w1165 & w1613;
assign w2220 = w794 & w937;
assign w2221 = w2219 & w2220;
assign v698 = ~(w56 | w253);
assign w2222 = v698;
assign w2223 = ~w258 & w2222;
assign w2224 = w966 & w2223;
assign w2225 = w2221 & w2224;
assign w2226 = w2225 & w29239;
assign w2227 = w2213 & w2226;
assign w2228 = w2227 & w29638;
assign v699 = ~(w53 | w595);
assign w2229 = v699;
assign w2230 = ~w1207 & w2229;
assign w2231 = w1777 & w2230;
assign w2232 = w528 & w2231;
assign v700 = ~(w111 | w298);
assign w2233 = v700;
assign w2234 = w442 & w2233;
assign v701 = ~(w169 | w311);
assign w2235 = v701;
assign w2236 = w1259 & w2235;
assign w2237 = w2234 & w2236;
assign w2238 = w2232 & w2237;
assign v702 = ~(w78 | w388);
assign w2239 = v702;
assign w2240 = w358 & w708;
assign v703 = ~(w338 | w753);
assign w2241 = v703;
assign w2242 = ~w286 & w2241;
assign w2243 = ~w475 & w2242;
assign v704 = ~(w143 | w234);
assign w2244 = v704;
assign w2245 = ~w151 & w2244;
assign w2246 = ~w280 & w1330;
assign w2247 = w2245 & w2246;
assign w2248 = w2243 & w2247;
assign w2249 = w2240 & w2248;
assign w2250 = w2239 & w2249;
assign w2251 = w2238 & w2250;
assign v705 = ~(w266 | w497);
assign w2252 = v705;
assign w2253 = ~w447 & w2252;
assign w2254 = ~w135 & w489;
assign w2255 = w2253 & w2254;
assign v706 = ~(w400 | w428);
assign w2256 = v706;
assign w2257 = w1366 & w2256;
assign w2258 = w2255 & w2257;
assign w2259 = ~w451 & w2258;
assign w2260 = w2251 & w2259;
assign v707 = ~(w369 | w563);
assign w2261 = v707;
assign v708 = ~(w252 | w307);
assign w2262 = v708;
assign w2263 = w2261 & w2262;
assign v709 = ~(w385 | w530);
assign w2264 = v709;
assign w2265 = w2263 & w2264;
assign v710 = ~(w194 | w457);
assign w2266 = v710;
assign w2267 = w1288 & w2266;
assign v711 = ~(w134 | w481);
assign w2268 = v711;
assign w2269 = w332 & w2268;
assign w2270 = w2267 & w2269;
assign v712 = ~(w49 | w343);
assign w2271 = v712;
assign v713 = ~(w215 | w431);
assign w2272 = v713;
assign v714 = ~(w177 | w277);
assign w2273 = v714;
assign w2274 = w2272 & w2273;
assign w2275 = w2271 & w2274;
assign w2276 = w2270 & w2275;
assign v715 = ~(w287 | w410);
assign w2277 = v715;
assign w2278 = ~w65 & w2277;
assign w2279 = ~w260 & w2278;
assign w2280 = ~w484 & w1077;
assign w2281 = w1892 & w2280;
assign v716 = ~(w145 | w613);
assign w2282 = v716;
assign w2283 = ~w247 & w2282;
assign w2284 = ~w235 & w2283;
assign w2285 = w2281 & w2284;
assign w2286 = w2279 & w2285;
assign w2287 = w2276 & w2286;
assign w2288 = w2265 & w2287;
assign w2289 = w2260 & w2288;
assign w2290 = w2228 & w2289;
assign v717 = ~(w2202 | w2290);
assign w2291 = v717;
assign v718 = ~(w177 | w822);
assign w2292 = v718;
assign w2293 = ~w95 & w1358;
assign w2294 = w2292 & w2293;
assign w2295 = w808 & w2294;
assign v719 = ~(w241 | w373);
assign w2296 = v719;
assign w2297 = w1245 & w2296;
assign w2298 = w2295 & w2297;
assign v720 = ~(w298 | w812);
assign w2299 = v720;
assign w2300 = w579 & w2299;
assign v721 = ~(w308 | w427);
assign w2301 = v721;
assign w2302 = w1466 & w2301;
assign v722 = ~(w238 | w945);
assign w2303 = v722;
assign w2304 = ~w886 & w2303;
assign w2305 = w2302 & w2304;
assign v723 = ~(w120 | w447);
assign w2306 = v723;
assign w2307 = w345 & w1292;
assign w2308 = w728 & w2307;
assign w2309 = w2306 & w2308;
assign w2310 = w2305 & w2309;
assign w2311 = w998 & w1823;
assign w2312 = w2310 & w2311;
assign w2313 = w2300 & w2312;
assign w2314 = w2298 & w2313;
assign v724 = ~(w259 | w493);
assign w2315 = v724;
assign v725 = ~(w27 | w309);
assign w2316 = v725;
assign w2317 = w2315 & w2316;
assign w2318 = ~w224 & w2317;
assign v726 = ~(w400 | w456);
assign w2319 = v726;
assign w2320 = w2318 & w2319;
assign w2321 = w992 & w1096;
assign w2322 = w2320 & w2321;
assign w2323 = w2105 & w2322;
assign w2324 = ~w73 & w864;
assign v727 = ~(w595 | w629);
assign w2325 = v727;
assign w2326 = w1127 & w2325;
assign w2327 = w2324 & w2326;
assign w2328 = ~w379 & w1463;
assign w2329 = w2157 & w2328;
assign w2330 = w650 & w1788;
assign v728 = ~(w292 | w584);
assign w2331 = v728;
assign w2332 = w2330 & w2331;
assign w2333 = w2329 & w2332;
assign v729 = ~(w31 | w1207);
assign w2334 = v729;
assign w2335 = w2333 & w2334;
assign w2336 = w2327 & w2335;
assign w2337 = w2323 & w2336;
assign w2338 = w572 & w2337;
assign w2339 = w2314 & w2338;
assign v730 = ~(w2290 | w2339);
assign w2340 = v730;
assign w2341 = ~w595 & w2138;
assign w2342 = ~w388 & w2341;
assign v731 = ~(w533 | w558);
assign w2343 = v731;
assign w2344 = w52 & w2343;
assign w2345 = w2176 & w2344;
assign w2346 = w2342 & w2345;
assign v732 = ~(w177 | w266);
assign w2347 = v732;
assign v733 = ~(w425 | w451);
assign w2348 = v733;
assign v734 = ~(w639 | w945);
assign w2349 = v734;
assign v735 = ~(w31 | w656);
assign w2350 = v735;
assign w2351 = w2349 & w2350;
assign w2352 = w2348 & w2351;
assign w2353 = w2347 & w2352;
assign w2354 = w2346 & w2353;
assign v736 = ~(w457 | w999);
assign w2355 = v736;
assign w2356 = w1201 & w2355;
assign w2357 = w1413 & w2356;
assign w2358 = w1603 & w2357;
assign w2359 = w2354 & w2358;
assign w2360 = ~w379 & w614;
assign w2361 = ~w441 & w2360;
assign w2362 = ~w162 & w2361;
assign v737 = ~(w145 | w172);
assign w2363 = v737;
assign w2364 = w2362 & w2363;
assign w2365 = w1747 & w2364;
assign v738 = ~(w418 | w494);
assign w2366 = v738;
assign w2367 = w2365 & w2366;
assign w2368 = w2359 & w2367;
assign w2369 = ~w466 & w1761;
assign v739 = ~(w201 | w503);
assign w2370 = v739;
assign v740 = ~(w183 | w252);
assign w2371 = v740;
assign w2372 = w2370 & w2371;
assign w2373 = w114 & w2372;
assign v741 = ~(w311 | w692);
assign w2374 = v741;
assign w2375 = w2043 & w2374;
assign w2376 = ~w484 & w2375;
assign w2377 = w2373 & w2376;
assign w2378 = w2369 & w2377;
assign w2379 = w2377 & w30777;
assign v742 = ~(w1134 | w1564);
assign w2380 = v742;
assign v743 = ~(w90 | w605);
assign w2381 = v743;
assign w2382 = ~w56 & w2381;
assign w2383 = w2380 & w2382;
assign v744 = ~(w88 | w588);
assign w2384 = v744;
assign w2385 = ~w70 & w2384;
assign w2386 = w1443 & w2385;
assign w2387 = w2383 & w2386;
assign w2388 = w330 & w1202;
assign w2389 = ~w373 & w2388;
assign w2390 = w2205 & w2389;
assign w2391 = w2387 & w2390;
assign w2392 = w2379 & w2391;
assign v745 = ~(w251 | w731);
assign w2393 = v745;
assign v746 = ~(w593 | w624);
assign w2394 = v746;
assign w2395 = w765 & w2394;
assign w2396 = w2393 & w2395;
assign v747 = ~(w108 | w119);
assign w2397 = v747;
assign v748 = ~(w21 | w264);
assign w2398 = v748;
assign v749 = ~(w410 | w673);
assign w2399 = v749;
assign w2400 = w2398 & w2399;
assign v750 = ~(w420 | w493);
assign w2401 = v750;
assign w2402 = w2109 & w2401;
assign w2403 = w2400 & w2402;
assign w2404 = w2397 & w2403;
assign v751 = ~(w288 | w715);
assign w2405 = v751;
assign w2406 = w1764 & w2405;
assign w2407 = ~w482 & w2406;
assign w2408 = ~w53 & w449;
assign w2409 = w2407 & w2408;
assign w2410 = w2404 & w2409;
assign v752 = ~(w158 | w559);
assign w2411 = v752;
assign v753 = ~(w241 | w267);
assign w2412 = v753;
assign w2413 = ~w431 & w2412;
assign w2414 = ~w209 & w2413;
assign w2415 = w2411 & w2414;
assign v754 = ~(w280 | w525);
assign w2416 = v754;
assign w2417 = w1586 & w2416;
assign w2418 = ~w877 & w2417;
assign w2419 = ~w428 & w2418;
assign w2420 = w2415 & w2419;
assign w2421 = w2410 & w2420;
assign w2422 = w2396 & w2421;
assign w2423 = w2392 & w2422;
assign w2424 = w2368 & w2423;
assign v755 = ~(w2339 | w2424);
assign w2425 = v755;
assign v756 = ~(w123 | w224);
assign w2426 = v756;
assign v757 = ~(w216 | w758);
assign w2427 = v757;
assign w2428 = ~w635 & w2427;
assign w2429 = w2426 & w2428;
assign w2430 = ~w215 & w2397;
assign w2431 = ~w533 & w2430;
assign w2432 = w2429 & w2431;
assign w2433 = ~w656 & w1396;
assign w2434 = ~w266 & w2433;
assign v758 = ~(w141 | w541);
assign w2435 = v758;
assign w2436 = w946 & w2435;
assign w2437 = w2434 & w2436;
assign w2438 = w2432 & w2437;
assign w2439 = ~w633 & w2438;
assign v759 = ~(w82 | w316);
assign w2440 = v759;
assign w2441 = ~w98 & w283;
assign w2442 = w2440 & w2441;
assign v760 = ~(w309 | w642);
assign w2443 = v760;
assign v761 = ~(w593 | w892);
assign w2444 = v761;
assign w2445 = w2443 & w2444;
assign w2446 = w2442 & w2445;
assign v762 = ~(w425 | w588);
assign w2447 = v762;
assign w2448 = ~w338 & w2447;
assign w2449 = w2279 & w2448;
assign w2450 = w2446 & w2449;
assign w2451 = w2439 & w2450;
assign v763 = ~(w200 | w697);
assign w2452 = v763;
assign v764 = ~(w27 | w711);
assign w2453 = v764;
assign w2454 = w2452 & w2453;
assign w2455 = ~w497 & w2024;
assign w2456 = w537 & w2455;
assign w2457 = w2454 & w2456;
assign w2458 = ~w978 & w2185;
assign w2459 = ~w499 & w2458;
assign w2460 = w2457 & w2459;
assign w2461 = w843 & w31149;
assign v765 = ~(w165 | w581);
assign w2462 = v765;
assign w2463 = ~w73 & w1767;
assign w2464 = w2462 & w2463;
assign v766 = ~(w51 | w390);
assign w2465 = v766;
assign w2466 = ~w63 & w2465;
assign w2467 = ~w674 & w2466;
assign w2468 = w2078 & w2467;
assign w2469 = w621 & w2468;
assign w2470 = w2464 & w2469;
assign v767 = ~(w134 | w183);
assign w2471 = v767;
assign w2472 = ~w286 & w2471;
assign v768 = ~(w329 | w431);
assign w2473 = v768;
assign w2474 = ~w201 & w2473;
assign w2475 = w2472 & w2474;
assign v769 = ~(w430 | w474);
assign w2476 = v769;
assign w2477 = w2475 & w2476;
assign v770 = ~(w465 | w899);
assign w2478 = v770;
assign w2479 = ~w111 & w898;
assign w2480 = w2478 & w2479;
assign w2481 = w2477 & w2480;
assign v771 = ~(w151 | w1207);
assign w2482 = v771;
assign w2483 = ~w466 & w2482;
assign w2484 = w2094 & w2483;
assign v772 = ~(w238 | w613);
assign w2485 = v772;
assign w2486 = ~w624 & w2485;
assign w2487 = ~w749 & w2486;
assign w2488 = w2484 & w2487;
assign w2489 = w2481 & w2488;
assign w2490 = w2470 & w2489;
assign w2491 = w2461 & w2490;
assign w2492 = w2451 & w2491;
assign v773 = ~(w2424 | w2492);
assign w2493 = v773;
assign v774 = ~(w159 | w326);
assign w2494 = v774;
assign v775 = ~(w150 | w409);
assign w2495 = v775;
assign v776 = ~(w292 | w656);
assign w2496 = v776;
assign w2497 = w2495 & w2496;
assign v777 = ~(w180 | w220);
assign w2498 = v777;
assign w2499 = w2497 & w2498;
assign w2500 = w626 & w2499;
assign w2501 = w217 & ~w381;
assign v778 = ~(w173 | w812);
assign w2502 = v778;
assign w2503 = w2501 & w31150;
assign w2504 = w2500 & w2503;
assign v779 = ~(w475 | w525);
assign w2505 = v779;
assign w2506 = w2382 & w2505;
assign v780 = ~(w112 | w302);
assign w2507 = v780;
assign v781 = ~(w151 | w309);
assign w2508 = v781;
assign w2509 = w2507 & w2508;
assign w2510 = w977 & w2509;
assign w2511 = w2506 & w2510;
assign v782 = ~(w131 | w749);
assign w2512 = v782;
assign v783 = ~(w144 | w493);
assign w2513 = v783;
assign w2514 = w2512 & w2513;
assign w2515 = w698 & w1893;
assign w2516 = w2514 & w2515;
assign v784 = ~(w179 | w438);
assign w2517 = v784;
assign w2518 = w1689 & w2517;
assign w2519 = w2516 & w30778;
assign w2520 = w2511 & w2519;
assign w2521 = w2504 & w2520;
assign w2522 = w2521 & w31151;
assign v785 = ~(w494 | w595);
assign w2523 = v785;
assign w2524 = ~w77 & w2523;
assign w2525 = w1534 & w2524;
assign v786 = ~(w272 | w404);
assign w2526 = v786;
assign v787 = ~(w274 | w758);
assign w2527 = v787;
assign w2528 = w2526 & w2527;
assign w2529 = w1536 & w2528;
assign w2530 = w2525 & w2529;
assign w2531 = w1909 & w2530;
assign w2532 = ~w588 & w1288;
assign v788 = ~(w299 | w680);
assign w2533 = v788;
assign w2534 = w1049 & w2533;
assign v789 = ~(w202 | w214);
assign w2535 = v789;
assign w2536 = w2534 & w2535;
assign w2537 = w2532 & w2536;
assign w2538 = w733 & w2537;
assign w2539 = w2531 & w2538;
assign v790 = ~(w316 | w692);
assign w2540 = v790;
assign v791 = ~(w260 | w1032);
assign w2541 = v791;
assign w2542 = w2471 & w2541;
assign w2543 = w233 & ~w390;
assign w2544 = w2542 & w2543;
assign v792 = ~(w42 | w300);
assign w2545 = v792;
assign w2546 = ~w234 & w2545;
assign v793 = ~(w359 | w388);
assign w2547 = v793;
assign w2548 = w225 & w2547;
assign w2549 = w2546 & w2548;
assign w2550 = w2544 & w2549;
assign w2551 = w2540 & w2550;
assign w2552 = w2550 & w30779;
assign w2553 = w1934 & w30780;
assign w2554 = w1027 & w2553;
assign w2555 = w2554 & w31152;
assign w2556 = w2552 & w2555;
assign w2557 = ~w88 & w1471;
assign v794 = ~(w674 | w870);
assign w2558 = v794;
assign w2559 = ~w899 & w2558;
assign w2560 = w2557 & w2559;
assign w2561 = ~w307 & w523;
assign w2562 = w1503 & w2561;
assign w2563 = ~w497 & w1772;
assign w2564 = w2562 & w2563;
assign w2565 = w2564 & w31153;
assign w2566 = w2556 & w2565;
assign w2567 = w2539 & w2566;
assign w2568 = w2522 & w2567;
assign v795 = ~(w2492 | w2568);
assign w2569 = v795;
assign w2570 = ~w247 & w589;
assign w2571 = w777 & w2570;
assign w2572 = w1113 & w2571;
assign v796 = ~(w184 | w387);
assign w2573 = v796;
assign v797 = ~(w49 | w711);
assign w2574 = v797;
assign w2575 = w2573 & w2574;
assign v798 = ~(w176 | w208);
assign w2576 = v798;
assign w2577 = ~w451 & w2576;
assign w2578 = w2575 & w2577;
assign w2579 = w845 & w2578;
assign w2580 = w2056 & w2579;
assign w2581 = w2572 & w2580;
assign w2582 = w998 & w2349;
assign w2583 = w1363 & w2582;
assign w2584 = w2581 & w2583;
assign w2585 = w1927 & w2584;
assign v799 = ~(w264 | w438);
assign w2586 = v799;
assign w2587 = ~w168 & w2586;
assign v800 = ~(w234 | w337);
assign w2588 = v800;
assign w2589 = w2587 & w2588;
assign v801 = ~(w274 | w1134);
assign w2590 = v801;
assign w2591 = ~w70 & w2590;
assign w2592 = ~w456 & w2591;
assign w2593 = w2589 & w2592;
assign w2594 = ~w144 & w2593;
assign w2595 = w2172 & w30781;
assign w2596 = w2585 & w2595;
assign v802 = ~(w2568 | w2596);
assign w2597 = v802;
assign v803 = ~(w462 | w652);
assign w2598 = v803;
assign w2599 = w1460 & w30782;
assign v804 = ~(w633 | w715);
assign w2600 = v804;
assign w2601 = w1381 & w2600;
assign w2602 = ~w753 & w2601;
assign w2603 = ~w88 & w1296;
assign w2604 = w864 & w1814;
assign w2605 = w2603 & w2604;
assign v805 = ~(w379 | w643);
assign w2606 = v805;
assign w2607 = ~w613 & w2606;
assign w2608 = w2292 & w2607;
assign w2609 = w2605 & w2608;
assign w2610 = w2602 & w2609;
assign w2611 = w2609 & w30783;
assign w2612 = ~w95 & w1559;
assign w2613 = w44 & w2612;
assign v806 = ~(w184 | w288);
assign w2614 = v806;
assign w2615 = ~w558 & w2614;
assign v807 = ~(w699 | w742);
assign w2616 = v807;
assign v808 = ~(w176 | w531);
assign w2617 = v808;
assign w2618 = w2616 & w2617;
assign w2619 = w2615 & w2618;
assign w2620 = w2613 & w2619;
assign v809 = ~(w93 | w286);
assign w2621 = v809;
assign w2622 = w693 & w2621;
assign w2623 = w188 & w2622;
assign v810 = ~(w111 | w369);
assign w2624 = v810;
assign w2625 = ~w234 & w2624;
assign w2626 = ~w134 & w2625;
assign w2627 = w2623 & w2626;
assign w2628 = w2620 & w2627;
assign w2629 = w2611 & w2628;
assign v811 = ~(w291 | w674);
assign w2630 = v811;
assign v812 = ~(w253 | w503);
assign w2631 = v812;
assign w2632 = w225 & w2631;
assign w2633 = w2630 & w2632;
assign v813 = ~(w307 | w584);
assign w2634 = v813;
assign w2635 = w1086 & w2076;
assign v814 = ~(w271 | w642);
assign w2636 = v814;
assign w2637 = w1761 & w2636;
assign w2638 = w2635 & w2637;
assign w2639 = w2634 & w2638;
assign w2640 = w2633 & w2639;
assign w2641 = ~w103 & w1600;
assign w2642 = w657 & w2641;
assign w2643 = ~w53 & w1201;
assign v815 = ~(w108 | w559);
assign w2644 = v815;
assign v816 = ~(w51 | w428);
assign w2645 = v816;
assign w2646 = w2644 & w2645;
assign w2647 = w2643 & w2646;
assign w2648 = w2642 & w2647;
assign w2649 = w1654 & w2648;
assign v817 = ~(w167 | w317);
assign w2650 = v817;
assign v818 = ~(w235 | w530);
assign w2651 = v818;
assign w2652 = w2650 & w2651;
assign v819 = ~(w110 | w387);
assign w2653 = v819;
assign w2654 = w2003 & w2653;
assign w2655 = ~w525 & w2654;
assign w2656 = w2652 & w2655;
assign w2657 = w265 & ~w1032;
assign w2658 = w265 & w30472;
assign w2659 = ~w245 & w339;
assign w2660 = w122 & w352;
assign v820 = ~(w63 | w812);
assign w2661 = v820;
assign w2662 = ~w2660 & w2661;
assign w2663 = w2659 & w2662;
assign w2664 = w2658 & w2663;
assign w2665 = w2656 & w2664;
assign w2666 = w2649 & w2665;
assign w2667 = w2666 & w30473;
assign w2668 = w2629 & w2667;
assign w2669 = w2599 & w2668;
assign v821 = ~(w2596 | w2669);
assign w2670 = v821;
assign v822 = ~(w74 | w731);
assign w2671 = v822;
assign v823 = ~(w324 | w727);
assign w2672 = v823;
assign w2673 = ~w666 & w2672;
assign w2674 = w2458 & w2673;
assign w2675 = w2671 & w2674;
assign w2676 = w851 & w2675;
assign v824 = ~(w100 | w173);
assign w2677 = v824;
assign w2678 = w2156 & w2677;
assign w2679 = ~w192 & w318;
assign w2680 = w2678 & w2679;
assign v825 = ~(w103 | w564);
assign w2681 = v825;
assign w2682 = w824 & w2681;
assign w2683 = w2680 & w2682;
assign w2684 = w1550 & w28471;
assign w2685 = w1337 & w2684;
assign w2686 = w2683 & w2685;
assign w2687 = w2676 & w2686;
assign w2688 = w2392 & w2687;
assign v826 = ~(w202 | w224);
assign w2689 = v826;
assign w2690 = w1850 & w2689;
assign w2691 = w1781 & w2690;
assign v827 = ~(w82 | w739);
assign w2692 = v827;
assign w2693 = ~w187 & w2692;
assign w2694 = ~w221 & w2693;
assign w2695 = w2691 & w2694;
assign w2696 = w236 & w1470;
assign w2697 = ~w656 & w2696;
assign w2698 = w2587 & w2697;
assign w2699 = w2695 & w2698;
assign w2700 = w1723 & w2495;
assign v828 = ~(w194 | w643);
assign w2701 = v828;
assign w2702 = ~w21 & w2701;
assign w2703 = w2700 & w2702;
assign v829 = ~(w326 | w427);
assign w2704 = v829;
assign v830 = ~(w37 | w481);
assign w2705 = v830;
assign w2706 = ~w359 & w2705;
assign w2707 = w2704 & w2706;
assign v831 = ~(w120 | w1108);
assign w2708 = v831;
assign v832 = ~(w212 | w420);
assign w2709 = v832;
assign w2710 = w2708 & w2709;
assign w2711 = ~w685 & w2334;
assign w2712 = w2710 & w2711;
assign w2713 = w2707 & w2712;
assign w2714 = w2076 & w2645;
assign w2715 = w2713 & w2714;
assign w2716 = w2703 & w2715;
assign w2717 = w786 & w1878;
assign w2718 = ~w753 & w2717;
assign v833 = ~(w385 | w494);
assign w2719 = v833;
assign w2720 = w1711 & w2719;
assign w2721 = w2718 & w2720;
assign w2722 = w780 & w2721;
assign w2723 = w2716 & w30784;
assign w2724 = w2688 & w2723;
assign v834 = ~(w2669 | w2724);
assign w2725 = v834;
assign w2726 = w2669 & w2724;
assign v835 = ~(w2725 | w2726);
assign w2727 = v835;
assign v836 = ~(w563 | w697);
assign w2728 = v836;
assign v837 = ~(w111 | w331);
assign w2729 = v837;
assign w2730 = w2728 & w2729;
assign w2731 = w2501 & w2730;
assign v838 = ~(w201 | w456);
assign w2732 = v838;
assign v839 = ~(w387 | w405);
assign w2733 = v839;
assign w2734 = w498 & w2733;
assign w2735 = w2732 & w2734;
assign w2736 = w2731 & w2735;
assign w2737 = w2546 & w2736;
assign w2738 = ~w475 & w942;
assign w2739 = w942 & w29993;
assign v840 = ~(w51 | w267);
assign w2740 = v840;
assign w2741 = w1681 & w1989;
assign w2742 = w2740 & w2741;
assign w2743 = ~w224 & w802;
assign v841 = ~(w414 | w499);
assign w2744 = v841;
assign w2745 = w657 & w2744;
assign w2746 = w2743 & w2745;
assign w2747 = w2742 & w2746;
assign w2748 = w2739 & w2747;
assign v842 = ~(w398 | w593);
assign w2749 = v842;
assign w2750 = w2749 & w29994;
assign w2751 = ~w888 & w2750;
assign w2752 = ~w463 & w1536;
assign w2753 = ~w144 & w2752;
assign w2754 = w2751 & w2753;
assign w2755 = w2748 & w2754;
assign w2756 = w2737 & w2755;
assign v843 = ~(w479 | w715);
assign w2757 = v843;
assign v844 = ~(w173 | w642);
assign w2758 = v844;
assign w2759 = w2757 & w2758;
assign w2760 = ~w239 & w2709;
assign w2761 = w865 & w2760;
assign w2762 = w2116 & w2761;
assign w2763 = w2759 & w2762;
assign v845 = ~(w82 | w1032);
assign w2764 = v845;
assign w2765 = w1710 & w2764;
assign w2766 = w1011 & w2765;
assign w2767 = ~w742 & w1816;
assign v846 = ~(w180 | w566);
assign w2768 = v846;
assign w2769 = w2355 & w2768;
assign w2770 = w2767 & w2769;
assign w2771 = w844 & w2770;
assign w2772 = w2766 & w2771;
assign w2773 = w2763 & w2772;
assign w2774 = w2756 & w2773;
assign v847 = ~(w145 | w522);
assign w2775 = v847;
assign v848 = ~(w481 | w505);
assign w2776 = v848;
assign w2777 = w2775 & w2776;
assign v849 = ~(w312 | w633);
assign w2778 = v849;
assign v850 = ~(w68 | w410);
assign w2779 = v850;
assign w2780 = w2778 & w2779;
assign w2781 = w2777 & w2780;
assign w2782 = w1109 & w1905;
assign w2783 = w2781 & w2782;
assign w2784 = w1157 & w1546;
assign w2785 = w318 & w2784;
assign w2786 = w2783 & w2785;
assign w2787 = ~w870 & w1345;
assign v851 = ~(w110 | w643);
assign w2788 = v851;
assign w2789 = ~w469 & w2788;
assign w2790 = w2787 & w2789;
assign w2791 = w2361 & w2790;
assign w2792 = ~w27 & w358;
assign w2793 = ~w281 & w2792;
assign w2794 = ~w70 & w2793;
assign w2795 = w2791 & w2794;
assign w2796 = w2786 & w2795;
assign w2797 = w675 & ~w727;
assign w2798 = w91 & ~w422;
assign w2799 = w2797 & w2798;
assign w2800 = w970 & w2124;
assign w2801 = w2799 & w2800;
assign v852 = ~(w131 | w430);
assign w2802 = v852;
assign v853 = ~(w584 | w753);
assign w2803 = v853;
assign w2804 = w261 & w2803;
assign v854 = ~(w277 | w595);
assign w2805 = v854;
assign w2806 = w2804 & w2805;
assign w2807 = w2802 & w2806;
assign w2808 = w2801 & w2807;
assign w2809 = w1414 & w2808;
assign w2810 = w2796 & w2809;
assign w2811 = w2774 & w2810;
assign w2812 = w2724 & w2811;
assign v855 = ~(w2724 | w2811);
assign w2813 = v855;
assign v856 = ~(w2812 | w2813);
assign w2814 = v856;
assign w2815 = w1442 & w2592;
assign w2816 = ~w160 & w2815;
assign v857 = ~(w110 | w482);
assign w2817 = v857;
assign w2818 = w313 & w984;
assign w2819 = w2817 & w2818;
assign w2820 = ~w892 & w1603;
assign w2821 = w1106 & w2820;
assign w2822 = w2819 & w2821;
assign w2823 = w2816 & w2822;
assign v858 = ~(w281 | w742);
assign w2824 = v858;
assign w2825 = w2749 & w2824;
assign w2826 = w2299 & w2825;
assign w2827 = w2184 & w2826;
assign w2828 = w702 & w1128;
assign w2829 = w1976 & w2828;
assign v859 = ~(w216 | w475);
assign w2830 = v859;
assign w2831 = w1765 & w2830;
assign w2832 = w2829 & w2831;
assign w2833 = w2578 & w2832;
assign w2834 = w2827 & w2833;
assign v860 = ~(w422 | w877);
assign w2835 = v860;
assign w2836 = w1414 & w2835;
assign w2837 = ~w359 & w2836;
assign w2838 = w783 & w1161;
assign w2839 = w121 & w2838;
assign w2840 = w2838 & w29639;
assign w2841 = w2837 & w2840;
assign w2842 = w1663 & w1749;
assign w2843 = w2841 & w2842;
assign w2844 = w2834 & w2843;
assign w2845 = w2823 & w2844;
assign w2846 = w2228 & w2845;
assign w2847 = w2811 & w2846;
assign v861 = ~(w2811 | w2846);
assign w2848 = v861;
assign v862 = ~(w267 | w563);
assign w2849 = v862;
assign w2850 = w725 & w2453;
assign w2851 = ~w613 & w2850;
assign v863 = ~(w307 | w448);
assign w2852 = v863;
assign w2853 = ~w475 & w2852;
assign v864 = ~(w162 | w260);
assign w2854 = v864;
assign w2855 = w2805 & w2854;
assign w2856 = w2853 & w2855;
assign w2857 = w2018 & w2856;
assign w2858 = w2851 & w2857;
assign w2859 = w236 & w29640;
assign w2860 = w2857 & w29240;
assign w2861 = w676 & w1741;
assign w2862 = w2615 & w2861;
assign v865 = ~(w231 | w299);
assign w2863 = v865;
assign w2864 = w1424 & w2863;
assign w2865 = ~w134 & w2864;
assign w2866 = w2862 & w2865;
assign w2867 = w1178 & w1409;
assign v866 = ~(w303 | w316);
assign w2868 = v866;
assign v867 = ~(w292 | w494);
assign w2869 = v867;
assign w2870 = w2868 & w2869;
assign w2871 = w2867 & w2870;
assign w2872 = w2866 & w2871;
assign v868 = ~(w87 | w106);
assign w2873 = v868;
assign w2874 = w1563 & w2873;
assign w2875 = w26 & ~w2874;
assign w2876 = w328 & ~w2875;
assign v869 = ~(w165 | w541);
assign w2877 = v869;
assign w2878 = w1330 & w2877;
assign w2879 = w1281 & w2878;
assign w2880 = w2876 & w2879;
assign w2881 = w2467 & w2880;
assign w2882 = w2872 & w2881;
assign w2883 = w2860 & w2882;
assign w2884 = w2882 & w29241;
assign v870 = ~(w150 | w370);
assign w2885 = v870;
assign w2886 = w1541 & w2885;
assign w2887 = ~w640 & w2886;
assign w2888 = w2886 & w29242;
assign v871 = ~(w431 | w447);
assign w2889 = v871;
assign w2890 = w1239 & w2889;
assign v872 = ~(w53 | w287);
assign w2891 = v872;
assign w2892 = ~w186 & w2891;
assign w2893 = w2890 & w2892;
assign w2894 = w1558 & w2893;
assign w2895 = w2888 & w2894;
assign w2896 = w2894 & w29243;
assign w2897 = ~w438 & w2896;
assign w2898 = w2896 & w29641;
assign w2899 = w2884 & w2898;
assign w2900 = w1073 & w1242;
assign v873 = ~(w201 | w656);
assign w2901 = v873;
assign w2902 = w551 & w2901;
assign w2903 = w2900 & w2902;
assign v874 = ~(w119 | w462);
assign w2904 = v874;
assign v875 = ~(w49 | w143);
assign w2905 = v875;
assign w2906 = w2904 & w2905;
assign w2907 = ~w311 & w2906;
assign w2908 = w2903 & w2907;
assign w2909 = w2825 & w2908;
assign w2910 = w1372 & w2150;
assign w2911 = w2909 & w2910;
assign v876 = ~(w497 | w749);
assign w2912 = v876;
assign w2913 = w1406 & w2912;
assign w2914 = w1413 & w2913;
assign w2915 = ~w272 & w1722;
assign v877 = ~(w177 | w302);
assign w2916 = v877;
assign w2917 = w1249 & w2916;
assign w2918 = w2915 & w2917;
assign w2919 = ~w200 & w29244;
assign v878 = ~(w95 | w263);
assign w2920 = v878;
assign w2921 = w589 & w2920;
assign w2922 = w2919 & w2921;
assign w2923 = w2918 & w2922;
assign v879 = ~(w317 | w629);
assign w2924 = v879;
assign w2925 = w1306 & w2924;
assign w2926 = ~w56 & w2925;
assign v880 = ~(w99 | w605);
assign w2927 = v880;
assign w2928 = ~w425 & w2927;
assign v881 = ~(w247 | w680);
assign w2929 = v881;
assign w2930 = ~w107 & w2929;
assign w2931 = w2928 & w2930;
assign w2932 = w2926 & w2931;
assign w2933 = w2923 & w2932;
assign w2934 = w2914 & w2933;
assign w2935 = w2911 & w2934;
assign w2936 = w1542 & w2935;
assign w2937 = w2899 & w2936;
assign v882 = ~(w2846 | w2937);
assign w2938 = v882;
assign w2939 = w2846 & w2937;
assign v883 = ~(w2938 | w2939);
assign w2940 = v883;
assign w2941 = ~w298 & w2435;
assign w2942 = ~w51 & w2941;
assign w2943 = ~w370 & w2049;
assign w2944 = w2942 & w2943;
assign w2945 = ~w469 & w1067;
assign v884 = ~(w123 | w234);
assign w2946 = v884;
assign w2947 = w101 & w2946;
assign w2948 = w1164 & w2947;
assign w2949 = w2945 & w2948;
assign w2950 = w2944 & w2949;
assign v885 = ~(w90 | w482);
assign w2951 = v885;
assign v886 = ~(w239 | w271);
assign w2952 = v886;
assign w2953 = ~w247 & w2952;
assign w2954 = w2951 & w2953;
assign v887 = ~(w211 | w235);
assign w2955 = v887;
assign v888 = ~(w107 | w652);
assign w2956 = v888;
assign w2957 = ~w899 & w2956;
assign w2958 = w2955 & w2957;
assign w2959 = w2954 & w2958;
assign v889 = ~(w65 | w244);
assign w2960 = v889;
assign w2961 = w1914 & w2960;
assign w2962 = w1781 & w2961;
assign w2963 = w2959 & w2962;
assign w2964 = w2950 & w2963;
assign v890 = ~(w266 | w311);
assign w2965 = v890;
assign w2966 = ~w588 & w2965;
assign v891 = ~(w673 | w680);
assign w2967 = v891;
assign w2968 = w2966 & w2967;
assign w2969 = w2083 & w2644;
assign w2970 = w2968 & w2969;
assign w2971 = w875 & w1574;
assign v892 = ~(w404 | w548);
assign w2972 = v892;
assign w2973 = ~w288 & w2972;
assign w2974 = w2971 & w2973;
assign w2975 = w641 & w2974;
assign w2976 = w2970 & w2975;
assign w2977 = ~w388 & w1831;
assign w2978 = w1206 & w2977;
assign v893 = ~(w132 | w282);
assign w2979 = v893;
assign w2980 = w225 & w2979;
assign w2981 = w2978 & w2980;
assign v894 = ~(w221 | w384);
assign w2982 = v894;
assign w2983 = w1195 & w2982;
assign w2984 = w600 & w2983;
assign w2985 = w2981 & w2984;
assign w2986 = w2976 & w2985;
assign w2987 = w1463 & w1853;
assign v895 = ~(w530 | w822);
assign w2988 = v895;
assign w2989 = ~w474 & w2988;
assign w2990 = w2987 & w2989;
assign v896 = ~(w112 | w337);
assign w2991 = v896;
assign w2992 = w174 & w2991;
assign w2993 = w803 & w2992;
assign w2994 = w2990 & w2993;
assign v897 = ~(w272 | w286);
assign w2995 = v897;
assign w2996 = w698 & w2995;
assign w2997 = w2994 & w2996;
assign w2998 = w2986 & w2997;
assign w2999 = w2964 & w2998;
assign w3000 = w1006 & w2999;
assign w3001 = w2937 & w3000;
assign v898 = ~(w2937 | w3000);
assign w3002 = v898;
assign v899 = ~(w221 | w299);
assign w3003 = v899;
assign w3004 = w2465 & w3003;
assign w3005 = w1109 & w1955;
assign w3006 = w3004 & w3005;
assign v900 = ~(w168 | w742);
assign w3007 = v900;
assign v901 = ~(w451 | w484);
assign w3008 = v901;
assign v902 = ~(w409 | w427);
assign w3009 = v902;
assign w3010 = w3008 & w3009;
assign w3011 = w3007 & w3010;
assign w3012 = w3006 & w3011;
assign v903 = ~(w550 | w630);
assign w3013 = v903;
assign v904 = ~(w151 | w238);
assign w3014 = v904;
assign v905 = ~(w370 | w525);
assign w3015 = v905;
assign w3016 = w3014 & w3015;
assign w3017 = w3013 & w3016;
assign w3018 = w1417 & w3017;
assign w3019 = w3012 & w3018;
assign w3020 = ~w530 & w1613;
assign w3021 = w1503 & w3020;
assign v906 = ~(w244 | w378);
assign w3022 = v906;
assign w3023 = w3021 & w3022;
assign w3024 = w3019 & w3023;
assign w3025 = ~w53 & w726;
assign w3026 = w1321 & w3025;
assign w3027 = w279 & w3026;
assign w3028 = w2687 & w3027;
assign w3029 = w3024 & w3028;
assign w3030 = w290 & w549;
assign w3031 = w2736 & w3030;
assign v907 = ~(w715 | w989);
assign w3032 = v907;
assign w3033 = w1647 & w3032;
assign w3034 = w1693 & w3033;
assign w3035 = w1258 & w3034;
assign w3036 = w3031 & w3035;
assign v908 = ~(w128 | w180);
assign w3037 = v908;
assign w3038 = ~w158 & w3037;
assign v909 = ~(w37 | w248);
assign w3039 = v909;
assign w3040 = w3038 & w3039;
assign w3041 = w1000 & w28152;
assign w3042 = w3040 & w3041;
assign v910 = ~(w232 | w593);
assign w3043 = v910;
assign v911 = ~(w234 | w308);
assign w3044 = v911;
assign v912 = ~(w194 | w692);
assign w3045 = v912;
assign w3046 = w3044 & w3045;
assign w3047 = w3043 & w3046;
assign v913 = ~(w195 | w639);
assign w3048 = v913;
assign w3049 = w3046 & w28153;
assign w3050 = w3042 & w3049;
assign v914 = ~(w177 | w247);
assign w3051 = v914;
assign w3052 = ~w291 & w1868;
assign w3053 = w3051 & w3052;
assign v915 = ~(w120 | w343);
assign w3054 = v915;
assign w3055 = ~w753 & w3054;
assign w3056 = w2182 & w3055;
assign w3057 = w3053 & w3056;
assign w3058 = ~w78 & w1442;
assign w3059 = w1106 & w3058;
assign v916 = ~(w90 | w642);
assign w3060 = v916;
assign v917 = ~(w144 | w595);
assign w3061 = v917;
assign w3062 = w3060 & w3061;
assign w3063 = w3059 & w3062;
assign w3064 = w3057 & w3063;
assign w3065 = w3050 & w3064;
assign w3066 = w2293 & w3065;
assign w3067 = w3036 & w3066;
assign w3068 = w3029 & w3067;
assign w3069 = w3000 & w3068;
assign v918 = ~(w3000 | w3068);
assign w3070 = v918;
assign v919 = ~(w123 | w259);
assign w3071 = v919;
assign w3072 = w265 & w3071;
assign w3073 = w625 & w3072;
assign w3074 = ~w286 & w3073;
assign v920 = ~(w165 | w731);
assign w3075 = v920;
assign v921 = ~(w220 | w454);
assign w3076 = v921;
assign w3077 = w3075 & w3076;
assign w3078 = w2863 & w3077;
assign w3079 = w1492 & w28154;
assign w3080 = w3074 & w3079;
assign w3081 = w1359 & w1822;
assign w3082 = w667 & w1099;
assign v922 = ~(w100 | w463);
assign w3083 = v922;
assign w3084 = w1228 & w3083;
assign w3085 = w3082 & w3084;
assign v923 = ~(w384 | w1134);
assign w3086 = v923;
assign w3087 = w2508 & w3086;
assign v924 = ~(w176 | w438);
assign w3088 = v924;
assign w3089 = w3087 & w3088;
assign w3090 = w3085 & w3089;
assign v925 = ~(w329 | w652);
assign w3091 = v925;
assign w3092 = ~w200 & w3091;
assign w3093 = w3092 & w28155;
assign w3094 = w3090 & w3093;
assign w3095 = w3081 & w3094;
assign w3096 = ~w493 & w1636;
assign w3097 = ~w558 & w3096;
assign w3098 = w1406 & w3097;
assign w3099 = ~w462 & w1840;
assign w3100 = ~w241 & w2052;
assign w3101 = w3099 & w3100;
assign w3102 = w225 & w1200;
assign w3103 = w2661 & w3102;
assign w3104 = w3101 & w3103;
assign v926 = ~(w281 | w387);
assign w3105 = v926;
assign w3106 = w1475 & w3105;
assign v927 = ~(w531 | w886);
assign w3107 = v927;
assign w3108 = w3106 & w3107;
assign w3109 = w3104 & w3108;
assign w3110 = w3098 & w3109;
assign w3111 = w3095 & w3110;
assign w3112 = w3080 & w3111;
assign v928 = ~(w359 | w548);
assign w3113 = v928;
assign w3114 = ~w469 & w3113;
assign v929 = ~(w892 | w978);
assign w3115 = v929;
assign w3116 = w2889 & w3115;
assign w3117 = w3114 & w3116;
assign w3118 = w115 & w3117;
assign v930 = ~(w479 | w673);
assign w3119 = v930;
assign w3120 = w597 & w3119;
assign w3121 = w304 & ~w1207;
assign w3122 = w3120 & w3121;
assign w3123 = w3065 & w28156;
assign w3124 = w3112 & w3123;
assign v931 = ~(w3068 | w3124);
assign w3125 = v931;
assign w3126 = w3068 & w3124;
assign v932 = ~(w3125 | w3126);
assign w3127 = v932;
assign v933 = ~(w244 | w437);
assign w3128 = v933;
assign w3129 = w2835 & w3128;
assign v934 = ~(w112 | w192);
assign w3130 = v934;
assign w3131 = w3129 & w3130;
assign w3132 = w3058 & w3131;
assign v935 = ~(w191 | w469);
assign w3133 = v935;
assign v936 = ~(w248 | w292);
assign w3134 = v936;
assign v937 = ~(w70 | w414);
assign w3135 = v937;
assign w3136 = ~w150 & w3135;
assign w3137 = w3134 & w3136;
assign w3138 = w3133 & w3137;
assign w3139 = w3132 & w3138;
assign v938 = ~(w263 | w331);
assign w3140 = v938;
assign w3141 = ~w82 & w594;
assign w3142 = w3140 & w3141;
assign w3143 = w553 & w1330;
assign w3144 = w188 & w3143;
assign w3145 = w3142 & w3144;
assign w3146 = ~w541 & w3145;
assign w3147 = w3139 & w3146;
assign w3148 = w2087 & w3147;
assign v939 = ~(w128 | w613);
assign w3149 = v939;
assign w3150 = w1238 & w3149;
assign w3151 = w573 & w3150;
assign v940 = ~(w37 | w384);
assign w3152 = v940;
assign v941 = ~(w103 | w488);
assign w3153 = v941;
assign w3154 = w3152 & w3153;
assign w3155 = ~w99 & w3154;
assign w3156 = w3151 & w3155;
assign w3157 = w1109 & w3156;
assign v942 = ~(w134 | w317);
assign w3158 = v942;
assign w3159 = w2299 & w3158;
assign w3160 = w3157 & w3159;
assign w3161 = w1704 & w3160;
assign w3162 = w3148 & w3161;
assign w3163 = w3124 & w3162;
assign w3164 = ~w21 & w2444;
assign w3165 = w2369 & w3164;
assign v943 = ~(w220 | w656);
assign w3166 = v943;
assign w3167 = ~w640 & w3166;
assign w3168 = w3165 & w3167;
assign v944 = ~(w82 | w329);
assign w3169 = v944;
assign w3170 = w1799 & w3169;
assign w3171 = w1043 & w3170;
assign w3172 = w1682 & w3071;
assign w3173 = w3171 & w3172;
assign w3174 = w3168 & w3173;
assign w3175 = ~w945 & w3086;
assign w3176 = w3086 & w27994;
assign w3177 = ~w271 & w3176;
assign w3178 = w2276 & w3177;
assign w3179 = w3174 & w3178;
assign w3180 = w551 & w31154;
assign w3181 = w284 & w1593;
assign w3182 = w3181 & w31155;
assign v945 = ~(w216 | w605);
assign w3183 = v945;
assign w3184 = ~w428 & w3183;
assign v946 = ~(w248 | w874);
assign w3185 = v946;
assign w3186 = ~w287 & w3185;
assign w3187 = w174 & w3186;
assign w3188 = w3184 & w3187;
assign v947 = ~(w209 | w430);
assign w3189 = v947;
assign w3190 = ~w112 & w3189;
assign w3191 = w3187 & w31156;
assign w3192 = w3182 & w3191;
assign w3193 = w3179 & w3192;
assign v948 = ~(w425 | w441);
assign w3194 = v948;
assign w3195 = w2689 & w3194;
assign v949 = ~(w503 | w666);
assign w3196 = v949;
assign v950 = ~(w176 | w372);
assign w3197 = v950;
assign w3198 = w3196 & w3197;
assign w3199 = w3195 & w3198;
assign v951 = ~(w533 | w674);
assign w3200 = v951;
assign w3201 = w1418 & w28473;
assign w3202 = ~w37 & w3201;
assign w3203 = w109 & w1048;
assign w3204 = ~w1032 & w3203;
assign v952 = ~(w150 | w877);
assign w3205 = v952;
assign w3206 = w615 & w3205;
assign w3207 = w3204 & w3206;
assign w3208 = w3207 & w28474;
assign w3209 = w3199 & w3208;
assign w3210 = w748 & w3209;
assign w3211 = w3193 & w3210;
assign w3212 = ~w463 & w2970;
assign w3213 = w76 & w3013;
assign v953 = ~(w141 | w398);
assign w3214 = v953;
assign w3215 = w2768 & w3214;
assign w3216 = w859 & w1131;
assign v954 = ~(w493 | w692);
assign w3217 = v954;
assign v955 = ~(w263 | w812);
assign w3218 = v955;
assign w3219 = w3217 & w3218;
assign w3220 = w3216 & w3219;
assign w3221 = w3215 & w3220;
assign w3222 = w3213 & w3221;
assign w3223 = w740 & w1878;
assign w3224 = w2078 & w3223;
assign w3225 = w2243 & w3224;
assign w3226 = w1342 & w3225;
assign w3227 = w3222 & w3226;
assign w3228 = w3212 & w3227;
assign v956 = ~(w316 | w451);
assign w3229 = v956;
assign w3230 = ~w298 & w3229;
assign v957 = ~(w160 | w454);
assign w3231 = v957;
assign v958 = ~(w93 | w742);
assign w3232 = v958;
assign w3233 = w3231 & w3232;
assign w3234 = w3230 & w3233;
assign v959 = ~(w245 | w420);
assign w3235 = v959;
assign w3236 = w2015 & w3235;
assign w3237 = w490 & ~w624;
assign w3238 = w3236 & w3237;
assign w3239 = w2740 & w3238;
assign w3240 = w3234 & w3239;
assign v960 = ~(w151 | w291);
assign w3241 = v960;
assign w3242 = w2076 & w3241;
assign w3243 = w1853 & w3242;
assign w3244 = w676 & w3243;
assign w3245 = w3240 & w3244;
assign w3246 = w3179 & w3245;
assign w3247 = w416 & w1065;
assign w3248 = ~w56 & w2606;
assign v961 = ~(w183 | w387);
assign w3249 = v961;
assign w3250 = ~w128 & w3249;
assign w3251 = w3248 & w3250;
assign w3252 = ~w531 & w1118;
assign w3253 = w3251 & w3252;
assign w3254 = w3247 & w3253;
assign v962 = ~(w127 | w437);
assign w3255 = v962;
assign w3256 = w233 & w3255;
assign w3257 = ~w685 & w3256;
assign w3258 = ~w192 & w3257;
assign w3259 = w1003 & w3258;
assign w3260 = w3254 & w3259;
assign w3261 = w3246 & w3260;
assign w3262 = w3228 & w3261;
assign w3263 = w3162 & w3262;
assign v963 = ~(w3211 | w3263);
assign w3264 = v963;
assign w3265 = w57 & w213;
assign w3266 = ~w27 & w2427;
assign v964 = ~(w474 | w530);
assign w3267 = v964;
assign v965 = ~(w272 | w481);
assign w3268 = v965;
assign w3269 = w3267 & w3268;
assign w3270 = w3266 & w3269;
assign v966 = ~(w484 | w692);
assign w3271 = v966;
assign w3272 = w366 & w3271;
assign w3273 = w196 & w3272;
assign w3274 = w3270 & w3273;
assign w3275 = w3265 & w3274;
assign w3276 = ~w388 & w2452;
assign v967 = ~(w264 | w753);
assign w3277 = v967;
assign w3278 = w2849 & w3277;
assign w3279 = w2749 & w3189;
assign w3280 = w3166 & w3279;
assign w3281 = w3278 & w3280;
assign w3282 = w3276 & w3281;
assign w3283 = w3275 & w3282;
assign w3284 = w869 & w3283;
assign v968 = ~(w522 | w624);
assign w3285 = v968;
assign w3286 = w3133 & w3285;
assign w3287 = w2134 & w3286;
assign w3288 = ~w373 & w894;
assign w3289 = w2196 & w3288;
assign w3290 = w3287 & w3289;
assign w3291 = ~w581 & w1535;
assign w3292 = w1050 & w3291;
assign v969 = ~(w42 | w892);
assign w3293 = v969;
assign w3294 = w3292 & w3293;
assign w3295 = w3290 & w3294;
assign w3296 = w1371 & w3030;
assign w3297 = w3295 & w3296;
assign w3298 = ~w749 & w1041;
assign w3299 = w358 & w3298;
assign v970 = ~(w312 | w384);
assign w3300 = v970;
assign v971 = ~(w337 | w595);
assign w3301 = v971;
assign w3302 = w2478 & w3301;
assign w3303 = w3300 & w3302;
assign v972 = ~(w588 | w999);
assign w3304 = v972;
assign w3305 = ~w731 & w3304;
assign w3306 = w2733 & w3305;
assign w3307 = w3303 & w3306;
assign w3308 = w3299 & w3307;
assign w3309 = ~w418 & w1010;
assign w3310 = w3308 & w3309;
assign w3311 = w3297 & w3310;
assign v973 = ~(w559 | w605);
assign w3312 = v973;
assign w3313 = w638 & w3312;
assign w3314 = w580 & w600;
assign w3315 = w1144 & w3314;
assign w3316 = w3313 & w3315;
assign v974 = ~(w65 | w431);
assign w3317 = v974;
assign v975 = ~(w135 | w258);
assign w3318 = v975;
assign w3319 = w3317 & w3318;
assign v976 = ~(w420 | w564);
assign w3320 = v976;
assign w3321 = ~w150 & w3320;
assign w3322 = w3319 & w3321;
assign v977 = ~(w224 | w711);
assign w3323 = v977;
assign w3324 = w1457 & w3323;
assign w3325 = ~w326 & w1600;
assign w3326 = ~w422 & w1536;
assign w3327 = w3325 & w3326;
assign w3328 = w3324 & w3327;
assign w3329 = w3322 & w3328;
assign w3330 = w3316 & w3329;
assign w3331 = w3311 & w3330;
assign w3332 = w3284 & w3331;
assign v978 = ~(w3162 | w3262);
assign w3333 = v978;
assign w3334 = ~w3332 & w3333;
assign v979 = ~(w3264 | w3334);
assign w3335 = v979;
assign v980 = ~(w3124 | w3162);
assign w3336 = v980;
assign v981 = ~(w3163 | w3336);
assign w3337 = v981;
assign w3338 = w3335 & w3337;
assign w3339 = (~w3163 & ~w3335) | (~w3163 & w27995) | (~w3335 & w27995);
assign w3340 = w3127 & w3339;
assign w3341 = (w3339 & w28275) | (w3339 & w28276) | (w28275 & w28276);
assign w3342 = (w3341 & w28690) | (w3341 & w28691) | (w28690 & w28691);
assign w3343 = (~w3341 & w28956) | (~w3341 & w28957) | (w28956 & w28957);
assign w3344 = (w3341 & w29461) | (w3341 & w29462) | (w29461 & w29462);
assign w3345 = w2814 & ~w3344;
assign w3346 = (w3341 & w29828) | (w3341 & w29829) | (w29828 & w29829);
assign w3347 = w2727 & w3346;
assign w3348 = (~w2725 & ~w3346) | (~w2725 & w29830) | (~w3346 & w29830);
assign w3349 = w2596 & w2669;
assign v982 = ~(w2670 | w3349);
assign w3350 = v982;
assign w3351 = (w3346 & w29995) | (w3346 & w29996) | (w29995 & w29996);
assign w3352 = (~w3346 & w30140) | (~w3346 & w30141) | (w30140 & w30141);
assign w3353 = w2568 & w2596;
assign v983 = ~(w2597 | w3353);
assign w3354 = v983;
assign w3355 = (w3346 & w30306) | (w3346 & w30307) | (w30306 & w30307);
assign w3356 = (~w3346 & w30474) | (~w3346 & w30475) | (w30474 & w30475);
assign w3357 = w2492 & w2568;
assign v984 = ~(w2569 | w3357);
assign w3358 = v984;
assign w3359 = (w3346 & w30583) | (w3346 & w30584) | (w30583 & w30584);
assign v985 = ~(w2569 | w3359);
assign w3360 = v985;
assign w3361 = w2424 & w2492;
assign v986 = ~(w2493 | w3361);
assign w3362 = v986;
assign w3363 = (w3346 & w30996) | (w3346 & w30997) | (w30996 & w30997);
assign v987 = ~(w2493 | w3363);
assign w3364 = v987;
assign w3365 = w2339 & w2424;
assign v988 = ~(w2425 | w3365);
assign w3366 = v988;
assign w3367 = (w3366 & w3363) | (w3366 & w31157) | (w3363 & w31157);
assign w3368 = (~w3363 & w31254) | (~w3363 & w31255) | (w31254 & w31255);
assign w3369 = w2290 & w2339;
assign v989 = ~(w2340 | w3369);
assign w3370 = v989;
assign w3371 = ~w3368 & w3370;
assign v990 = ~(w2340 | w3371);
assign w3372 = v990;
assign w3373 = w2202 & w2290;
assign v991 = ~(w2291 | w3373);
assign w3374 = v991;
assign w3375 = ~w3372 & w3374;
assign v992 = ~(w2291 | w3375);
assign w3376 = v992;
assign w3377 = w2089 & w2202;
assign v993 = ~(w2203 | w3377);
assign w3378 = v993;
assign w3379 = ~w3376 & w3378;
assign v994 = ~(w2203 | w3379);
assign w3380 = v994;
assign w3381 = ~w2091 & w3380;
assign v995 = ~(w2090 | w3381);
assign w3382 = v995;
assign w3383 = w2041 & w3382;
assign v996 = ~(w2039 | w3383);
assign w3384 = v996;
assign v997 = ~(w1944 | w3384);
assign w3385 = v997;
assign v998 = ~(w1943 | w3385);
assign w3386 = v998;
assign w3387 = w1863 & ~w3386;
assign v999 = ~(w1861 | w3387);
assign w3388 = v999;
assign w3389 = w1798 & ~w3388;
assign v1000 = ~(w1796 | w3389);
assign w3390 = v1000;
assign v1001 = ~(w1676 | w3390);
assign w3391 = v1001;
assign v1002 = ~(w1675 | w3391);
assign w3392 = v1002;
assign v1003 = ~(w1611 | w3392);
assign w3393 = v1003;
assign v1004 = ~(w1610 | w3393);
assign w3394 = v1004;
assign w3395 = w1499 & ~w3394;
assign w3396 = ~w1499 & w3394;
assign v1005 = ~(w3395 | w3396);
assign w3397 = v1005;
assign w3398 = w928 & w3397;
assign w3399 = pi31 & w18;
assign w3400 = ~w1609 & w3399;
assign v1006 = ~(pi31 | w18);
assign w3401 = v1006;
assign v1007 = ~(w927 | w3401);
assign w3402 = v1007;
assign w3403 = ~w1496 & w3402;
assign v1008 = ~(w3400 | w3403);
assign w3404 = v1008;
assign v1009 = ~(w29 | w45);
assign w3405 = v1009;
assign v1010 = ~(pi31 | w3405);
assign w3406 = v1010;
assign w3407 = ~w1387 & w3406;
assign w3408 = w3404 & ~w3407;
assign w3409 = ~w3398 & w3408;
assign w3410 = w1279 & ~w3409;
assign w3411 = ~w1279 & w3409;
assign v1011 = ~(w3410 | w3411);
assign w3412 = v1011;
assign v1012 = ~(pi20 | w1274);
assign w3413 = v1012;
assign v1013 = ~(w1275 | w3413);
assign w3414 = v1013;
assign w3415 = w358 & w1157;
assign w3416 = ~w488 & w3415;
assign v1014 = ~(w88 | w331);
assign w3417 = v1014;
assign w3418 = w1302 & w3417;
assign w3419 = w3416 & w3418;
assign w3420 = w121 & w3419;
assign w3421 = ~w404 & w1415;
assign v1015 = ~(w100 | w165);
assign w3422 = v1015;
assign w3423 = w1462 & w3422;
assign w3424 = w3421 & w3423;
assign w3425 = w46 & w72;
assign w3426 = ~w989 & w1560;
assign w3427 = ~w3425 & w3426;
assign w3428 = w3424 & w3427;
assign w3429 = w3420 & w3428;
assign w3430 = ~w414 & w2245;
assign w3431 = ~w613 & w3430;
assign w3432 = w450 & w3231;
assign w3433 = ~w593 & w3432;
assign v1016 = ~(w107 | w191);
assign w3434 = v1016;
assign w3435 = ~w405 & w3434;
assign w3436 = ~w680 & w3435;
assign w3437 = w3433 & w3436;
assign v1017 = ~(w77 | w353);
assign w3438 = v1017;
assign w3439 = ~w177 & w3438;
assign w3440 = w1905 & w3439;
assign w3441 = w3437 & w3440;
assign w3442 = w3431 & w3441;
assign w3443 = w3429 & w3442;
assign w3444 = w419 & w3443;
assign w3445 = ~w308 & w1048;
assign w3446 = ~w74 & w3445;
assign v1018 = ~(w278 | w422);
assign w3447 = v1018;
assign w3448 = ~w112 & w3447;
assign w3449 = w3446 & w3448;
assign v1019 = ~(w224 | w466);
assign w3450 = v1019;
assign w3451 = ~w253 & w3450;
assign w3452 = w1842 & w3451;
assign w3453 = w1603 & w2188;
assign w3454 = w565 & w3453;
assign w3455 = w3452 & w3454;
assign w3456 = w3449 & w3455;
assign v1020 = ~(w475 | w584);
assign w3457 = v1020;
assign v1021 = ~(w624 | w888);
assign w3458 = v1021;
assign w3459 = w1754 & w3458;
assign v1022 = ~(w312 | w1032);
assign w3460 = v1022;
assign w3461 = ~w245 & w3460;
assign w3462 = w3459 & w3461;
assign w3463 = w3457 & w3462;
assign v1023 = ~(w99 | w108);
assign w3464 = v1023;
assign v1024 = ~(w78 | w337);
assign w3465 = v1024;
assign w3466 = w3464 & w3465;
assign v1025 = ~(w90 | w812);
assign w3467 = v1025;
assign w3468 = w1722 & w3467;
assign w3469 = w3466 & w3468;
assign w3470 = w2319 & w3469;
assign w3471 = w3463 & w3470;
assign w3472 = w3456 & w3471;
assign v1026 = ~(w82 | w479);
assign w3473 = v1026;
assign w3474 = ~w731 & w3473;
assign v1027 = ~(w220 | w550);
assign w3475 = v1027;
assign v1028 = ~(w469 | w758);
assign w3476 = v1028;
assign w3477 = w3475 & w3476;
assign w3478 = w3474 & w3477;
assign w3479 = w2010 & w2866;
assign w3480 = w3478 & w3479;
assign w3481 = w3472 & w3480;
assign w3482 = w1041 & w2602;
assign w3483 = w1813 & w3482;
assign w3484 = w1540 & w3483;
assign w3485 = w1256 & w3484;
assign w3486 = w3481 & w3485;
assign w3487 = w3444 & w3486;
assign w3488 = ~w1153 & w3487;
assign w3489 = w1153 & ~w3487;
assign v1029 = ~(w3488 | w3489);
assign w3490 = v1029;
assign w3491 = ~w1675 & w3391;
assign v1030 = ~(w1675 | w1676);
assign w3492 = v1030;
assign w3493 = w3390 & ~w3492;
assign v1031 = ~(w3491 | w3493);
assign w3494 = v1031;
assign w3495 = w928 & w3494;
assign w3496 = ~w1795 & w3399;
assign w3497 = ~w1609 & w3406;
assign v1032 = ~(w3496 | w3497);
assign w3498 = v1032;
assign w3499 = ~w1674 & w3402;
assign w3500 = w3498 & ~w3499;
assign w3501 = ~w3495 & w3500;
assign w3502 = w3490 & w3501;
assign v1033 = ~(w3488 | w3502);
assign w3503 = v1033;
assign w3504 = ~w3414 & w3503;
assign w3505 = w3414 & ~w3503;
assign v1034 = ~(w3504 | w3505);
assign w3506 = v1034;
assign v1035 = ~(w1610 | w1611);
assign w3507 = v1035;
assign w3508 = w3392 & w3507;
assign v1036 = ~(w3392 | w3507);
assign w3509 = v1036;
assign v1037 = ~(w3508 | w3509);
assign w3510 = v1037;
assign w3511 = w928 & ~w3510;
assign w3512 = ~w1609 & w3402;
assign w3513 = ~w1496 & w3406;
assign v1038 = ~(w3512 | w3513);
assign w3514 = v1038;
assign w3515 = ~w1674 & w3399;
assign w3516 = w3514 & ~w3515;
assign w3517 = ~w3511 & w3516;
assign w3518 = w3506 & ~w3517;
assign v1039 = ~(w3504 | w3518);
assign w3519 = v1039;
assign w3520 = w3412 & ~w3519;
assign w3521 = ~w3412 & w3519;
assign v1040 = ~(w3520 | w3521);
assign w3522 = v1040;
assign v1041 = ~(pi26 | pi27);
assign w3523 = v1041;
assign w3524 = pi26 & pi27;
assign v1042 = ~(w3523 | w3524);
assign w3525 = v1042;
assign v1043 = ~(pi28 | pi29);
assign w3526 = v1043;
assign w3527 = pi28 & pi29;
assign v1044 = ~(w3526 | w3527);
assign w3528 = v1044;
assign w3529 = w3525 & w3528;
assign v1045 = ~(w169 | w173);
assign w3530 = v1045;
assign v1046 = ~(w286 | w997);
assign w3531 = v1046;
assign w3532 = ~w110 & w3531;
assign w3533 = w3530 & w3532;
assign w3534 = w222 & w3533;
assign w3535 = w185 & w366;
assign w3536 = w2707 & w3535;
assign w3537 = w3534 & w3536;
assign w3538 = ~w312 & w2630;
assign w3539 = ~w448 & w565;
assign w3540 = w3538 & w3539;
assign w3541 = ~w642 & w3540;
assign w3542 = w2643 & w3541;
assign w3543 = w3537 & w3542;
assign v1047 = ~(w125 | w609);
assign w3544 = v1047;
assign v1048 = ~(w165 | w697);
assign w3545 = v1048;
assign w3546 = w101 & w3545;
assign w3547 = w3544 & w3546;
assign v1049 = ~(w378 | w420);
assign w3548 = v1049;
assign w3549 = w382 & w3548;
assign w3550 = w2988 & w3549;
assign w3551 = w3547 & w3550;
assign v1050 = ~(w215 | w874);
assign w3552 = v1050;
assign w3553 = ~w309 & w452;
assign w3554 = w3552 & w3553;
assign w3555 = w2887 & w3554;
assign w3556 = w3551 & w3555;
assign v1051 = ~(w633 | w749);
assign w3557 = v1051;
assign v1052 = ~(w194 | w463);
assign w3558 = v1052;
assign w3559 = w3557 & w3558;
assign w3560 = ~w639 & w3559;
assign w3561 = w834 & w3560;
assign w3562 = w3556 & w3561;
assign w3563 = ~w643 & w2625;
assign v1053 = ~(w65 | w108);
assign w3564 = v1053;
assign w3565 = w3563 & w3564;
assign w3566 = w3562 & w3565;
assign w3567 = w3543 & w3566;
assign v1054 = ~(w224 | w252);
assign w3568 = v1054;
assign v1055 = ~(w167 | w886);
assign w3569 = v1055;
assign v1056 = ~(w324 | w418);
assign w3570 = v1056;
assign w3571 = ~w260 & w1409;
assign w3572 = w3570 & w3571;
assign v1057 = ~(w298 | w457);
assign w3573 = v1057;
assign w3574 = ~w123 & w3573;
assign w3575 = w3572 & w3574;
assign w3576 = w2156 & w2507;
assign v1058 = ~(w103 | w191);
assign w3577 = v1058;
assign w3578 = ~w271 & w3577;
assign w3579 = w3576 & w3578;
assign v1059 = ~(w390 | w465);
assign w3580 = v1059;
assign w3581 = w1186 & w3580;
assign w3582 = w3579 & w3581;
assign w3583 = w3575 & w3582;
assign w3584 = w3569 & w3583;
assign w3585 = w3568 & w3584;
assign w3586 = w1461 & w3585;
assign w3587 = w3567 & w3586;
assign w3588 = ~w53 & w970;
assign v1060 = ~(w214 | w877);
assign w3589 = v1060;
assign v1061 = ~(w584 | w656);
assign w3590 = v1061;
assign w3591 = w3589 & w3590;
assign w3592 = w1786 & w3591;
assign w3593 = w3588 & w3592;
assign w3594 = w1093 & w2381;
assign w3595 = w419 & w3594;
assign v1062 = ~(w235 | w430);
assign w3596 = v1062;
assign w3597 = w1574 & w3596;
assign v1063 = ~(w263 | w338);
assign w3598 = v1063;
assign v1064 = ~(w183 | w253);
assign w3599 = v1064;
assign w3600 = w3598 & w3599;
assign w3601 = w3597 & w3600;
assign w3602 = w3595 & w3601;
assign w3603 = ~w331 & w2349;
assign w3604 = w1888 & w3603;
assign w3605 = w1632 & w3604;
assign w3606 = w3602 & w3605;
assign w3607 = w1602 & w1717;
assign w3608 = ~w685 & w2788;
assign w3609 = ~w388 & w3608;
assign w3610 = w3607 & w3609;
assign w3611 = w3606 & w3610;
assign w3612 = w3593 & w3611;
assign w3613 = ~w195 & w979;
assign w3614 = w1226 & w3613;
assign v1065 = ~(w640 | w749);
assign w3615 = v1065;
assign w3616 = w1345 & w3615;
assign w3617 = w990 & w3616;
assign w3618 = w3614 & w3617;
assign w3619 = w455 & w3618;
assign v1066 = ~(w260 | w613);
assign w3620 = v1066;
assign w3621 = w3196 & w3620;
assign w3622 = w3619 & w3621;
assign w3623 = w1462 & w2704;
assign v1067 = ~(w56 | w244);
assign w3624 = v1067;
assign w3625 = w3623 & w3624;
assign v1068 = ~(w63 | w144);
assign w3626 = v1068;
assign w3627 = w318 & w2142;
assign w3628 = w3626 & w3627;
assign w3629 = w3625 & w3628;
assign w3630 = w1623 & w3629;
assign w3631 = w3622 & w3630;
assign v1069 = ~(w180 | w223);
assign w3632 = v1069;
assign w3633 = w1056 & w3632;
assign w3634 = ~w711 & w3633;
assign w3635 = ~w99 & w2681;
assign v1070 = ~(w128 | w633);
assign w3636 = v1070;
assign w3637 = ~w337 & w3636;
assign w3638 = w3635 & w3637;
assign w3639 = w3634 & w3638;
assign w3640 = ~w145 & w1935;
assign w3641 = w442 & w3640;
assign w3642 = w3639 & w3641;
assign w3643 = w3631 & w3642;
assign v1071 = ~(w177 | w642);
assign w3644 = v1071;
assign w3645 = w2728 & w3644;
assign w3646 = ~w373 & w1162;
assign w3647 = w3645 & w3646;
assign w3648 = w3446 & w3647;
assign w3649 = w1596 & w2341;
assign v1072 = ~(w162 | w997);
assign w3650 = v1072;
assign v1073 = ~(w150 | w312);
assign w3651 = v1073;
assign w3652 = w3650 & w3651;
assign w3653 = w217 & w3652;
assign v1074 = ~(w343 | w378);
assign w3654 = v1074;
assign w3655 = ~w462 & w3654;
assign w3656 = w1287 & w3655;
assign w3657 = w3653 & w3656;
assign v1075 = ~(w282 | w463);
assign w3658 = v1075;
assign v1076 = ~(w208 | w680);
assign w3659 = v1076;
assign w3660 = w3658 & w3659;
assign w3661 = w1921 & w3660;
assign w3662 = w3657 & w3661;
assign w3663 = w3649 & w3662;
assign w3664 = w3648 & w3663;
assign w3665 = w3643 & w3664;
assign w3666 = w3612 & w3665;
assign v1077 = ~(w3587 | w3666);
assign w3667 = v1077;
assign w3668 = w3587 & w3666;
assign v1078 = ~(w3667 | w3668);
assign w3669 = v1078;
assign w3670 = w1387 & w3666;
assign v1079 = ~(w1387 | w3666);
assign w3671 = v1079;
assign v1080 = ~(w1497 | w3395);
assign w3672 = v1080;
assign w3673 = ~w3671 & w3672;
assign v1081 = ~(w3670 | w3673);
assign w3674 = v1081;
assign w3675 = w3669 & w3674;
assign v1082 = ~(w3667 | w3675);
assign w3676 = v1082;
assign v1083 = ~(w151 | w168);
assign w3677 = v1083;
assign w3678 = ~w390 & w3677;
assign v1084 = ~(w27 | w125);
assign w3679 = v1084;
assign w3680 = w3545 & w3679;
assign w3681 = w2405 & w3680;
assign w3682 = w3678 & w3681;
assign w3683 = w306 & w3682;
assign w3684 = w959 & ~w997;
assign w3685 = w2033 & w3684;
assign v1085 = ~(w169 | w541);
assign w3686 = v1085;
assign w3687 = w2478 & w3686;
assign w3688 = w3685 & w3687;
assign w3689 = ~w88 & w2043;
assign w3690 = w1853 & w3689;
assign v1086 = ~(w278 | w311);
assign w3691 = v1086;
assign w3692 = w1462 & w3691;
assign w3693 = w761 & w3692;
assign w3694 = w3690 & w3693;
assign w3695 = w3688 & w3694;
assign w3696 = w3683 & w3695;
assign v1087 = ~(w65 | w220);
assign w3697 = v1087;
assign w3698 = w3696 & w3697;
assign v1088 = ~(w287 | w566);
assign w3699 = v1088;
assign w3700 = w1893 & w3699;
assign v1089 = ~(w202 | w281);
assign w3701 = v1089;
assign w3702 = w1475 & w3701;
assign w3703 = w375 & w3702;
assign w3704 = w3700 & w3703;
assign w3705 = w707 & w3658;
assign w3706 = w1409 & w1536;
assign w3707 = w3705 & w3706;
assign w3708 = w1080 & w3707;
assign w3709 = w1722 & w1884;
assign w3710 = w2078 & w3709;
assign w3711 = w3708 & w3710;
assign w3712 = w3704 & w3711;
assign w3713 = w2268 & w2749;
assign w3714 = ~w742 & w3713;
assign v1090 = ~(w462 | w978);
assign w3715 = v1090;
assign w3716 = w2239 & w3715;
assign w3717 = w3439 & w3716;
assign w3718 = w3714 & w3717;
assign w3719 = w1141 & w3718;
assign w3720 = w3712 & w3719;
assign w3721 = w3698 & w3720;
assign v1091 = ~(w418 | w488);
assign w3722 = v1091;
assign v1092 = ~(w120 | w252);
assign w3723 = v1092;
assign v1093 = ~(w454 | w1207);
assign w3724 = v1093;
assign w3725 = w1398 & w3724;
assign w3726 = w3723 & w3725;
assign w3727 = w57 & w2650;
assign w3728 = w1864 & w3727;
assign w3729 = w3726 & w3728;
assign v1094 = ~(w822 | w999);
assign w3730 = v1094;
assign w3731 = w785 & w3730;
assign w3732 = w3729 & w3731;
assign v1095 = ~(w215 | w224);
assign w3733 = v1095;
assign w3734 = w1255 & w3733;
assign v1096 = ~(w216 | w564);
assign w3735 = v1096;
assign w3736 = w2955 & w3735;
assign v1097 = ~(w379 | w422);
assign w3737 = v1097;
assign v1098 = ~(w266 | w343);
assign w3738 = v1098;
assign w3739 = w3737 & w3738;
assign w3740 = w3736 & w3739;
assign v1099 = ~(w405 | w674);
assign w3741 = v1099;
assign w3742 = ~w531 & w3741;
assign w3743 = w3038 & w3742;
assign w3744 = w3740 & w3743;
assign w3745 = ~w451 & w1177;
assign v1100 = ~(w90 | w588);
assign w3746 = v1100;
assign w3747 = w3745 & w3746;
assign w3748 = w3744 & w3747;
assign w3749 = w3734 & w3748;
assign w3750 = w3732 & w3749;
assign w3751 = w3722 & w3750;
assign w3752 = w3721 & w3751;
assign w3753 = w3587 & w3752;
assign v1101 = ~(w3587 | w3752);
assign w3754 = v1101;
assign v1102 = ~(w3753 | w3754);
assign w3755 = v1102;
assign w3756 = w3676 & ~w3755;
assign w3757 = ~w3676 & w3755;
assign v1103 = ~(w3756 | w3757);
assign w3758 = v1103;
assign w3759 = w3529 & w3758;
assign w3760 = w3525 & ~w3528;
assign w3761 = ~w3752 & w3760;
assign v1104 = ~(w19 | w40);
assign w3762 = v1104;
assign w3763 = ~w3525 & w3762;
assign w3764 = ~w3587 & w3763;
assign v1105 = ~(w3761 | w3764);
assign w3765 = v1105;
assign w3766 = ~w3525 & w3528;
assign w3767 = ~w3762 & w3766;
assign w3768 = ~w3666 & w3767;
assign w3769 = w3765 & ~w3768;
assign w3770 = ~w3759 & w3769;
assign w3771 = ~pi29 & w3770;
assign w3772 = pi29 & ~w3770;
assign v1106 = ~(w3771 | w3772);
assign w3773 = v1106;
assign w3774 = w3522 & w3773;
assign v1107 = ~(w3520 | w3774);
assign w3775 = v1107;
assign v1108 = ~(w1277 | w3410);
assign w3776 = v1108;
assign w3777 = ~w652 & w3015;
assign w3778 = ~w531 & w3777;
assign w3779 = w3058 & w3778;
assign v1109 = ~(w159 | w466);
assign w3780 = v1109;
assign w3781 = ~w999 & w3780;
assign w3782 = ~w978 & w3781;
assign w3783 = w3779 & w3782;
assign v1110 = ~(w74 | w302);
assign w3784 = v1110;
assign w3785 = ~w88 & w768;
assign w3786 = w3784 & w3785;
assign w3787 = ~w359 & w1552;
assign w3788 = w2661 & w3787;
assign w3789 = w3786 & w3788;
assign w3790 = ~w742 & w3789;
assign w3791 = w3783 & w3790;
assign w3792 = ~w158 & w3577;
assign w3793 = w1619 & w3792;
assign w3794 = w2253 & w2532;
assign w3795 = w3793 & w3794;
assign w3796 = ~w558 & w3475;
assign w3797 = w2729 & w3796;
assign w3798 = w3609 & w3797;
assign w3799 = w3795 & w3798;
assign w3800 = w801 & w3799;
assign w3801 = w2100 & w3599;
assign w3802 = ~w405 & w3801;
assign v1111 = ~(w180 | w711);
assign w3803 = v1111;
assign w3804 = ~w400 & w3803;
assign v1112 = ~(w168 | w307);
assign w3805 = v1112;
assign w3806 = w3804 & w3805;
assign w3807 = w3802 & w3806;
assign v1113 = ~(w324 | w329);
assign w3808 = v1113;
assign w3809 = w2527 & w3808;
assign v1114 = ~(w200 | w378);
assign w3810 = v1114;
assign w3811 = w3809 & w3810;
assign w3812 = w3807 & w3811;
assign w3813 = ~w192 & w990;
assign w3814 = ~w223 & w3813;
assign w3815 = w3199 & w3814;
assign w3816 = w34 & ~w1563;
assign w3817 = w1239 & ~w3816;
assign v1115 = ~(w160 | w892);
assign w3818 = v1115;
assign w3819 = w889 & w3818;
assign w3820 = ~w282 & w3819;
assign w3821 = w3817 & w3820;
assign w3822 = w3815 & w3821;
assign w3823 = w3812 & w3822;
assign w3824 = w3800 & w3823;
assign w3825 = ~w715 & w1888;
assign w3826 = w2374 & w3825;
assign w3827 = ~w522 & w2003;
assign w3828 = ~w559 & w3827;
assign w3829 = w3826 & w3828;
assign w3830 = w489 & w3829;
assign w3831 = w2167 & w3830;
assign w3832 = w3824 & w3831;
assign w3833 = w3791 & w3832;
assign w3834 = w1055 & ~w3833;
assign w3835 = ~w1055 & w3833;
assign v1116 = ~(w3834 | w3835);
assign w3836 = v1116;
assign w3837 = w3776 & w3836;
assign v1117 = ~(w3776 | w3836);
assign w3838 = v1117;
assign v1118 = ~(w3837 | w3838);
assign w3839 = v1118;
assign v1119 = ~(w3670 | w3671);
assign w3840 = v1119;
assign w3841 = w3672 & ~w3840;
assign w3842 = ~w3672 & w3840;
assign v1120 = ~(w3841 | w3842);
assign w3843 = v1120;
assign w3844 = w928 & w3843;
assign w3845 = w3406 & ~w3666;
assign w3846 = ~w1387 & w3402;
assign v1121 = ~(w3845 | w3846);
assign w3847 = v1121;
assign w3848 = ~w1496 & w3399;
assign w3849 = w3847 & ~w3848;
assign w3850 = ~w3844 & w3849;
assign v1122 = ~(w3839 | w3850);
assign w3851 = v1122;
assign w3852 = w3839 & w3850;
assign v1123 = ~(w3851 | w3852);
assign w3853 = v1123;
assign w3854 = ~w3775 & w3853;
assign w3855 = w3775 & ~w3853;
assign v1124 = ~(w3854 | w3855);
assign w3856 = v1124;
assign w3857 = ~w3587 & w3767;
assign v1125 = ~(w112 | w238);
assign w3858 = v1125;
assign w3859 = w1834 & w3858;
assign w3860 = w587 & w3859;
assign v1126 = ~(w437 | w475);
assign w3861 = v1126;
assign w3862 = w1226 & w3861;
assign w3863 = w2283 & w3140;
assign w3864 = w3862 & w3863;
assign v1127 = ~(w874 | w945);
assign w3865 = v1127;
assign w3866 = w698 & w2229;
assign w3867 = w1512 & w2268;
assign w3868 = w3866 & w3867;
assign w3869 = w3865 & w3868;
assign w3870 = w3864 & w3869;
assign w3871 = ~w168 & w1722;
assign w3872 = w783 & w3871;
assign v1128 = ~(w223 | w609);
assign w3873 = v1128;
assign w3874 = w3872 & w3873;
assign w3875 = w3870 & w3874;
assign w3876 = w403 & w3875;
assign w3877 = w3860 & w3876;
assign v1129 = ~(w173 | w324);
assign w3878 = v1129;
assign w3879 = w1161 & w3878;
assign w3880 = ~w531 & w3879;
assign w3881 = w1813 & w3880;
assign w3882 = ~w73 & w1057;
assign v1130 = ~(w742 | w1032);
assign w3883 = v1130;
assign w3884 = w2235 & w3883;
assign w3885 = w3882 & w3884;
assign v1131 = ~(w184 | w474);
assign w3886 = v1131;
assign v1132 = ~(w140 | w505);
assign w3887 = v1132;
assign w3888 = ~w93 & w3887;
assign w3889 = ~w177 & w3888;
assign w3890 = w3886 & w3889;
assign w3891 = w3885 & w3890;
assign w3892 = ~w125 & w2546;
assign w3893 = w3122 & w3892;
assign w3894 = w3891 & w3893;
assign w3895 = w3881 & w3894;
assign w3896 = ~w390 & w1559;
assign w3897 = w1028 & w1853;
assign w3898 = w3896 & w3897;
assign w3899 = ~w588 & w3730;
assign w3900 = w3898 & w3899;
assign w3901 = w798 & w3900;
assign v1133 = ~(w186 | w212);
assign w3902 = v1133;
assign w3903 = ~w447 & w3902;
assign v1134 = ~(w280 | w370);
assign w3904 = v1134;
assign w3905 = w993 & w3904;
assign w3906 = w3903 & w3905;
assign w3907 = w1980 & w3906;
assign w3908 = w415 & w607;
assign w3909 = ~w548 & w3271;
assign w3910 = w3908 & w3909;
assign v1135 = ~(w388 | w530);
assign w3911 = v1135;
assign v1136 = ~(w31 | w812);
assign w3912 = v1136;
assign w3913 = w3911 & w3912;
assign w3914 = w3910 & w3913;
assign w3915 = w204 & ~w264;
assign w3916 = w3914 & w3915;
assign w3917 = w3907 & w3916;
assign w3918 = w3901 & w3917;
assign w3919 = w3895 & w3918;
assign w3920 = w3877 & w3919;
assign v1137 = ~(w3752 | w3920);
assign w3921 = v1137;
assign w3922 = w3752 & w3920;
assign v1138 = ~(w3921 | w3922);
assign w3923 = v1138;
assign v1139 = ~(w3676 | w3753);
assign w3924 = v1139;
assign v1140 = ~(w3754 | w3924);
assign w3925 = v1140;
assign v1141 = ~(w3923 | w3925);
assign w3926 = v1141;
assign w3927 = w3923 & w3925;
assign v1142 = ~(w3926 | w3927);
assign w3928 = v1142;
assign w3929 = w3529 & ~w3928;
assign w3930 = ~w3752 & w3763;
assign w3931 = w3760 & ~w3920;
assign v1143 = ~(w3930 | w3931);
assign w3932 = v1143;
assign w3933 = ~w3929 & w3932;
assign w3934 = ~w3857 & w3933;
assign w3935 = pi29 & w3934;
assign v1144 = ~(pi29 | w3934);
assign w3936 = v1144;
assign v1145 = ~(w3935 | w3936);
assign w3937 = v1145;
assign w3938 = w3856 & ~w3937;
assign w3939 = ~w3856 & w3937;
assign v1146 = ~(w3938 | w3939);
assign w3940 = v1146;
assign w3941 = w615 & w2636;
assign w3942 = w2918 & w3941;
assign w3943 = w859 & w3942;
assign v1147 = ~(w143 | w247);
assign w3944 = v1147;
assign w3945 = ~w409 & w3944;
assign w3946 = ~w184 & w3945;
assign v1148 = ~(w307 | w581);
assign w3947 = v1148;
assign w3948 = ~w132 & w3947;
assign w3949 = ~w463 & w3948;
assign w3950 = w3946 & w3949;
assign w3951 = w967 & w3697;
assign v1149 = ~(w469 | w1032);
assign w3952 = v1149;
assign w3953 = w1132 & w3952;
assign w3954 = w3951 & w3953;
assign w3955 = w596 & w3954;
assign w3956 = w3950 & w3955;
assign w3957 = w1559 & w3119;
assign w3958 = w1326 & w3957;
assign w3959 = w3956 & w3958;
assign w3960 = w366 & w2545;
assign w3961 = w3959 & w3960;
assign w3962 = ~w311 & w1378;
assign w3963 = ~w299 & w3962;
assign w3964 = w3714 & w3963;
assign v1150 = ~(w312 | w405);
assign w3965 = v1150;
assign w3966 = w657 & w3965;
assign w3967 = ~w541 & w3966;
assign w3968 = w1331 & w2768;
assign w3969 = w3967 & w3968;
assign w3970 = w3251 & w3969;
assign w3971 = ~w685 & w3970;
assign w3972 = w3964 & w3971;
assign w3973 = w3961 & w3972;
assign w3974 = ~w37 & w1447;
assign w3975 = w2052 & w3974;
assign w3976 = w1613 & w1888;
assign w3977 = ~w224 & w3976;
assign w3978 = w3975 & w3977;
assign w3979 = w3914 & w3978;
assign w3980 = w3973 & w3979;
assign w3981 = w3943 & w3980;
assign v1151 = ~(w298 | w639);
assign w3982 = v1151;
assign w3983 = w2069 & w3982;
assign v1152 = ~(w191 | w674);
assign w3984 = v1152;
assign w3985 = ~w82 & w3984;
assign w3986 = w3983 & w3985;
assign w3987 = w1771 & w3986;
assign w3988 = ~w281 & w3987;
assign w3989 = ~w88 & w397;
assign w3990 = w375 & w2107;
assign w3991 = w3989 & w3990;
assign v1153 = ~(w234 | w739);
assign w3992 = v1153;
assign w3993 = ~w168 & w3887;
assign w3994 = w3992 & w3993;
assign w3995 = w1911 & w3994;
assign w3996 = w3991 & w3995;
assign w3997 = w3988 & w3996;
assign w3998 = ~w248 & w3285;
assign w3999 = ~w338 & w3998;
assign v1154 = ~(w119 | w241);
assign w4000 = v1154;
assign w4001 = w3735 & w4000;
assign w4002 = w1130 & w4001;
assign w4003 = w3999 & w4002;
assign v1155 = ~(w385 | w420);
assign w4004 = v1155;
assign w4005 = w240 & w4004;
assign w4006 = w3730 & w4005;
assign w4007 = w4003 & w4006;
assign w4008 = w3997 & w4007;
assign w4009 = ~w70 & w561;
assign v1156 = ~(w21 | w337);
assign w4010 = v1156;
assign w4011 = w1238 & w4010;
assign w4012 = w426 & w4011;
assign w4013 = w4009 & w4012;
assign w4014 = ~w258 & w4013;
assign w4015 = ~w277 & w4014;
assign w4016 = w4008 & w4015;
assign v1157 = ~(w192 | w640);
assign w4017 = v1157;
assign w4018 = w3087 & w4017;
assign v1158 = ~(w232 | w456);
assign w4019 = v1158;
assign w4020 = ~w287 & w4019;
assign v1159 = ~(w99 | w278);
assign w4021 = v1159;
assign w4022 = w4020 & w4021;
assign w4023 = w4018 & w4022;
assign w4024 = pi25 & pi26;
assign v1160 = ~(pi25 | pi26);
assign w4025 = v1160;
assign v1161 = ~(w4024 | w4025);
assign w4026 = v1161;
assign v1162 = ~(w38 | w47);
assign w4027 = v1162;
assign w4028 = ~w61 & w4027;
assign w4029 = w122 & ~w4028;
assign w4030 = w4026 & w4029;
assign v1163 = ~(w187 | w4030);
assign w4031 = v1163;
assign w4032 = w4023 & w4031;
assign w4033 = ~w353 & w4032;
assign w4034 = w4016 & w4033;
assign w4035 = w3981 & w4034;
assign w4036 = ~w99 & w1561;
assign v1164 = ~(w277 | w685);
assign w4037 = v1164;
assign w4038 = w1647 & w4037;
assign w4039 = ~w753 & w4038;
assign w4040 = w4036 & w4039;
assign v1165 = ~(w162 | w731);
assign w4041 = v1165;
assign w4042 = w1228 & w3570;
assign w4043 = w4041 & w4042;
assign v1166 = ~(w90 | w711);
assign w4044 = v1166;
assign w4045 = ~w286 & w4044;
assign v1167 = ~(w317 | w466);
assign w4046 = v1167;
assign w4047 = w4045 & w4046;
assign w4048 = w4043 & w4047;
assign w4049 = w4040 & w4048;
assign w4050 = ~w173 & w3943;
assign w4051 = w1761 & w2334;
assign v1168 = ~(w209 | w548);
assign w4052 = v1168;
assign w4053 = ~w997 & w2982;
assign w4054 = w4052 & w4053;
assign v1169 = ~(w232 | w353);
assign w4055 = v1169;
assign w4056 = w965 & w4055;
assign w4057 = w4054 & w4056;
assign w4058 = w4051 & w4057;
assign w4059 = w3568 & w4058;
assign w4060 = w4050 & w4059;
assign w4061 = w2897 & w4060;
assign w4062 = w1188 & w1350;
assign w4063 = ~w195 & w4062;
assign w4064 = w573 & w2138;
assign v1170 = ~(w499 | w888);
assign w4065 = v1170;
assign w4066 = w1414 & w4065;
assign w4067 = w4064 & w4066;
assign w4068 = w1878 & w4067;
assign w4069 = w4063 & w4068;
assign v1171 = ~(w73 | w112);
assign w4070 = v1171;
assign w4071 = ~w95 & w4070;
assign w4072 = ~w245 & w4071;
assign w4073 = ~w331 & w4072;
assign w4074 = w4069 & w4073;
assign w4075 = ~w699 & w3544;
assign w4076 = w330 & w4075;
assign w4077 = w1586 & w4076;
assign w4078 = w4074 & w4077;
assign w4079 = w4061 & w4078;
assign w4080 = ~w172 & w4079;
assign w4081 = w4049 & w4080;
assign w4082 = ~w214 & w4081;
assign w4083 = w4035 & w4082;
assign v1172 = ~(w4035 | w4082);
assign w4084 = v1172;
assign v1173 = ~(w4083 | w4084);
assign w4085 = v1173;
assign w4086 = w1022 & w3902;
assign w4087 = w2092 & w4086;
assign w4088 = w2494 & w3013;
assign w4089 = ~w431 & w4088;
assign w4090 = w4087 & w4089;
assign w4091 = ~w145 & w3229;
assign w4092 = w210 & w2517;
assign w4093 = w565 & w1042;
assign w4094 = w4092 & w4093;
assign w4095 = w4091 & w4094;
assign w4096 = w4090 & w4095;
assign v1174 = ~(w141 | w292);
assign w4097 = v1174;
assign v1175 = ~(w93 | w169);
assign w4098 = v1175;
assign w4099 = ~w241 & w4098;
assign w4100 = w4097 & w4099;
assign w4101 = w4096 & w4100;
assign w4102 = w1161 & w1864;
assign v1176 = ~(w215 | w223);
assign w4103 = v1176;
assign w4104 = w4102 & w4103;
assign w4105 = ~w272 & w2885;
assign w4106 = w4104 & w4105;
assign w4107 = w1538 & w4106;
assign w4108 = w504 & w2677;
assign w4109 = w2429 & w4108;
assign w4110 = w1225 & w4109;
assign w4111 = w4107 & w4110;
assign w4112 = w3988 & w4111;
assign w4113 = w4101 & w4112;
assign w4114 = w2347 & w4045;
assign w4115 = ~w886 & w1118;
assign w4116 = w3999 & w4115;
assign w4117 = w4114 & w4116;
assign v1177 = ~(w98 | w329);
assign w4118 = v1177;
assign w4119 = ~w753 & w4118;
assign w4120 = w3304 & w4119;
assign v1178 = ~(w531 | w877);
assign w4121 = v1178;
assign w4122 = ~w127 & w4121;
assign w4123 = ~w697 & w4122;
assign w4124 = w4120 & w4123;
assign w4125 = w1535 & w1722;
assign w4126 = w467 & w1888;
assign w4127 = w4125 & w4126;
assign w4128 = w1063 & w3548;
assign w4129 = w740 & w4128;
assign w4130 = w4127 & w4129;
assign w4131 = w4124 & w4130;
assign w4132 = w4117 & w4131;
assign w4133 = w3996 & w4132;
assign w4134 = w4113 & w4133;
assign v1179 = ~(w4035 | w4134);
assign w4135 = v1179;
assign v1180 = ~(w3920 | w4134);
assign w4136 = v1180;
assign w4137 = w3920 & w4134;
assign v1181 = ~(w4136 | w4137);
assign w4138 = v1181;
assign w4139 = ~w3921 & w3925;
assign v1182 = ~(w3922 | w4139);
assign w4140 = v1182;
assign w4141 = w4138 & w4140;
assign v1183 = ~(w4136 | w4141);
assign w4142 = v1183;
assign w4143 = w4035 & w4134;
assign v1184 = ~(w4135 | w4143);
assign w4144 = v1184;
assign w4145 = ~w4142 & w4144;
assign v1185 = ~(w4135 | w4145);
assign w4146 = v1185;
assign w4147 = w4085 & w4146;
assign v1186 = ~(w4085 | w4146);
assign w4148 = v1186;
assign v1187 = ~(w4147 | w4148);
assign w4149 = v1187;
assign v1188 = ~(pi23 | pi24);
assign w4150 = v1188;
assign w4151 = pi23 & pi24;
assign v1189 = ~(w4150 | w4151);
assign w4152 = v1189;
assign w4153 = w4026 & w4152;
assign w4154 = ~w4149 & w4153;
assign w4155 = ~w4026 & w4152;
assign w4156 = ~w4082 & w4155;
assign v1190 = ~(w2873 | w4134);
assign w4157 = v1190;
assign w4158 = w4027 & ~w4152;
assign w4159 = ~w4035 & w4158;
assign v1191 = ~(w4157 | w4159);
assign w4160 = v1191;
assign w4161 = ~w4156 & w4160;
assign w4162 = ~w4154 & w4161;
assign w4163 = pi26 & ~w4162;
assign w4164 = ~pi26 & w4162;
assign v1192 = ~(w4163 | w4164);
assign w4165 = v1192;
assign w4166 = w3940 & w4165;
assign v1193 = ~(w3938 | w4166);
assign w4167 = v1193;
assign v1194 = ~(w4083 | w4147);
assign w4168 = v1194;
assign w4169 = ~w316 & w4098;
assign w4170 = w1074 & w2239;
assign w4171 = w4169 & w4170;
assign w4172 = ~w201 & w1613;
assign w4173 = w3129 & w4172;
assign w4174 = w4171 & w4173;
assign v1195 = ~(w199 | w308);
assign w4175 = v1195;
assign w4176 = w3054 & w4175;
assign w4177 = w1718 & w4176;
assign w4178 = w1066 & w2465;
assign w4179 = w4177 & w4178;
assign w4180 = w4174 & w4179;
assign v1196 = ~(w100 | w187);
assign w4181 = v1196;
assign w4182 = w1424 & w4181;
assign w4183 = w1888 & w2282;
assign w4184 = ~w758 & w4183;
assign w4185 = w4182 & w4184;
assign w4186 = w4180 & w4185;
assign w4187 = ~w267 & w4186;
assign v1197 = ~(w214 | w4030);
assign w4188 = v1197;
assign w4189 = w4187 & w4188;
assign w4190 = w4081 & w4189;
assign w4191 = w4049 & w4189;
assign v1198 = ~(w4082 | w4191);
assign w4192 = v1198;
assign v1199 = ~(w4190 | w4192);
assign w4193 = v1199;
assign w4194 = w4168 & w4193;
assign v1200 = ~(w4168 | w4193);
assign w4195 = v1200;
assign v1201 = ~(w4194 | w4195);
assign w4196 = v1201;
assign w4197 = w4153 & w4196;
assign w4198 = ~w4082 & w4158;
assign w4199 = w4155 & ~w4191;
assign v1202 = ~(w2873 | w4035);
assign w4200 = v1202;
assign v1203 = ~(w4199 | w4200);
assign w4201 = v1203;
assign w4202 = ~w4198 & w4201;
assign w4203 = ~w4197 & w4202;
assign w4204 = pi26 & ~w4203;
assign w4205 = ~pi26 & w4203;
assign v1204 = ~(w4204 | w4205);
assign w4206 = v1204;
assign w4207 = ~w4167 & w4206;
assign v1205 = ~(w3851 | w3854);
assign w4208 = v1205;
assign v1206 = ~(w3834 | w3837);
assign w4209 = v1206;
assign v1207 = ~(w74 | w447);
assign w4210 = v1207;
assign w4211 = ~w812 & w4210;
assign w4212 = ~w167 & w4211;
assign v1208 = ~(w231 | w999);
assign w4213 = v1208;
assign w4214 = ~w505 & w4213;
assign v1209 = ~(w110 | w317);
assign w4215 = v1209;
assign w4216 = w3285 & w4215;
assign w4217 = w4214 & w4216;
assign v1210 = ~(w493 | w593);
assign w4218 = v1210;
assign w4219 = w1772 & w4218;
assign w4220 = w2517 & w3214;
assign w4221 = w4219 & w4220;
assign w4222 = w4217 & w4221;
assign w4223 = w4212 & w4222;
assign w4224 = w1741 & w2108;
assign v1211 = ~(w98 | w201);
assign w4225 = v1211;
assign w4226 = w1587 & w4225;
assign w4227 = w4224 & w4226;
assign w4228 = w2707 & w4227;
assign w4229 = w4223 & w4228;
assign v1212 = ~(w437 | w466);
assign w4230 = v1212;
assign w4231 = w1066 & w4230;
assign w4232 = ~w409 & w4231;
assign w4233 = w1374 & w4232;
assign w4234 = w1483 & w2134;
assign w4235 = w440 & w1682;
assign w4236 = w4234 & w4235;
assign w4237 = w547 & w4236;
assign w4238 = w4233 & w4237;
assign w4239 = w213 & w2010;
assign v1213 = ~(w216 | w870);
assign w4240 = v1213;
assign w4241 = w3944 & w4240;
assign w4242 = w4239 & w4241;
assign w4243 = w2348 & w4242;
assign w4244 = ~w51 & w4243;
assign w4245 = ~w278 & w1840;
assign v1214 = ~(w271 | w749);
assign w4246 = v1214;
assign w4247 = w236 & w4246;
assign w4248 = w4245 & w4247;
assign w4249 = w1073 & w4248;
assign w4250 = w4244 & w4249;
assign w4251 = w4238 & w4250;
assign w4252 = w4229 & w4251;
assign w4253 = ~w177 & w1242;
assign v1215 = ~(w581 | w692);
assign w4254 = v1215;
assign w4255 = w818 & w4254;
assign w4256 = w4253 & w4255;
assign v1216 = ~(w499 | w633);
assign w4257 = v1216;
assign w4258 = ~w194 & w4257;
assign w4259 = w4256 & w4258;
assign w4260 = w1154 & w2758;
assign w4261 = w1707 & w4260;
assign w4262 = w335 & w534;
assign w4263 = w2233 & w4262;
assign w4264 = ~w405 & w4263;
assign w4265 = w4261 & w4264;
assign w4266 = w4259 & w4265;
assign w4267 = w2849 & w3858;
assign w4268 = w1358 & w4267;
assign v1217 = ~(w462 | w609);
assign w4269 = v1217;
assign w4270 = w412 & w1437;
assign w4271 = w4269 & w4270;
assign w4272 = w4268 & w4271;
assign w4273 = w315 & w4272;
assign v1218 = ~(w331 | w630);
assign w4274 = v1218;
assign v1219 = ~(w90 | w288);
assign w4275 = v1219;
assign w4276 = w4274 & w4275;
assign v1220 = ~(w150 | w874);
assign w4277 = v1220;
assign w4278 = w121 & w4277;
assign w4279 = w4276 & w4278;
assign w4280 = w4273 & w4279;
assign w4281 = w1948 & w4280;
assign w4282 = w4266 & w4281;
assign w4283 = w4252 & w4282;
assign w4284 = w3833 & w4283;
assign v1221 = ~(w3833 | w4283);
assign w4285 = v1221;
assign v1222 = ~(w4284 | w4285);
assign w4286 = v1222;
assign w4287 = pi23 & w4286;
assign v1223 = ~(pi23 | w4286);
assign w4288 = v1223;
assign v1224 = ~(w4287 | w4288);
assign w4289 = v1224;
assign v1225 = ~(w3669 | w3674);
assign w4290 = v1225;
assign v1226 = ~(w3675 | w4290);
assign w4291 = v1226;
assign w4292 = w928 & w4291;
assign w4293 = ~w1387 & w3399;
assign w4294 = w3406 & ~w3587;
assign v1227 = ~(w4293 | w4294);
assign w4295 = v1227;
assign w4296 = w3402 & ~w3666;
assign w4297 = w4295 & ~w4296;
assign w4298 = ~w4292 & w4297;
assign v1228 = ~(w4289 | w4298);
assign w4299 = v1228;
assign w4300 = w4289 & w4298;
assign v1229 = ~(w4299 | w4300);
assign w4301 = v1229;
assign w4302 = w4209 & w4301;
assign v1230 = ~(w4209 | w4301);
assign w4303 = v1230;
assign v1231 = ~(w4302 | w4303);
assign w4304 = v1231;
assign w4305 = ~w4208 & w4304;
assign w4306 = w4208 & ~w4304;
assign v1232 = ~(w4305 | w4306);
assign w4307 = v1232;
assign v1233 = ~(w4138 | w4140);
assign w4308 = v1233;
assign v1234 = ~(w4141 | w4308);
assign w4309 = v1234;
assign w4310 = w3529 & w4309;
assign w4311 = w3763 & ~w3920;
assign w4312 = ~w3752 & w3767;
assign w4313 = w3760 & ~w4134;
assign v1235 = ~(w4312 | w4313);
assign w4314 = v1235;
assign w4315 = ~w4311 & w4314;
assign w4316 = ~w4310 & w4315;
assign w4317 = pi29 & ~w4316;
assign w4318 = ~pi29 & w4316;
assign v1236 = ~(w4317 | w4318);
assign w4319 = v1236;
assign w4320 = w4307 & w4319;
assign v1237 = ~(w4307 | w4319);
assign w4321 = v1237;
assign v1238 = ~(w4320 | w4321);
assign w4322 = v1238;
assign w4323 = w4167 & ~w4206;
assign v1239 = ~(w4207 | w4323);
assign w4324 = v1239;
assign w4325 = w4322 & w4324;
assign v1240 = ~(w4207 | w4325);
assign w4326 = v1240;
assign v1241 = ~(w4305 | w4320);
assign w4327 = v1241;
assign w4328 = w625 & w1202;
assign w4329 = w615 & w4010;
assign w4330 = w4328 & w4329;
assign w4331 = w2955 & w4330;
assign w4332 = w3271 & w4331;
assign w4333 = w1109 & w4332;
assign w4334 = w2337 & w4333;
assign v1242 = ~(w107 | w172);
assign w4335 = v1242;
assign w4336 = ~w870 & w4335;
assign w4337 = ~w438 & w4336;
assign w4338 = w837 & w4337;
assign v1243 = ~(w99 | w252);
assign w4339 = v1243;
assign v1244 = ~(w123 | w727);
assign w4340 = v1244;
assign w4341 = ~w208 & w4340;
assign v1245 = ~(w184 | w248);
assign w4342 = v1245;
assign w4343 = w4341 & w4342;
assign w4344 = w4339 & w4343;
assign w4345 = w4338 & w4344;
assign w4346 = ~w274 & w3691;
assign v1246 = ~(w168 | w425);
assign w4347 = v1246;
assign w4348 = w79 & w4347;
assign w4349 = w4346 & w4348;
assign w4350 = w2541 & w2598;
assign w4351 = w4349 & w4350;
assign v1247 = ~(w221 | w280);
assign w4352 = v1247;
assign w4353 = w4351 & w4352;
assign w4354 = w4345 & w4353;
assign w4355 = ~w497 & w752;
assign w4356 = w1396 & w1423;
assign w4357 = w4355 & w4356;
assign w4358 = w2370 & w4357;
assign w4359 = w4214 & w4358;
assign w4360 = w4354 & w4359;
assign v1248 = ~(w93 | w548);
assign w4361 = v1248;
assign v1249 = ~(w144 | w656);
assign w4362 = v1249;
assign w4363 = w1435 & w4362;
assign w4364 = w2830 & w4363;
assign w4365 = w4361 & w4364;
assign v1250 = ~(w111 | w422);
assign w4366 = v1250;
assign w4367 = ~w1134 & w4366;
assign w4368 = w1409 & w1414;
assign w4369 = ~w209 & w4368;
assign w4370 = w4367 & w4369;
assign v1251 = ~(w307 | w374);
assign w4371 = v1251;
assign w4372 = ~w245 & w4371;
assign w4373 = ~w300 & w4372;
assign w4374 = w4370 & w4373;
assign w4375 = w4365 & w4374;
assign w4376 = w765 & ~w892;
assign w4377 = w2462 & w2533;
assign w4378 = w4376 & w4377;
assign w4379 = ~w303 & w3632;
assign w4380 = w1587 & w4379;
assign w4381 = w4378 & w4380;
assign w4382 = w3312 & w4381;
assign w4383 = w4375 & w4382;
assign w4384 = w4360 & w4383;
assign w4385 = w4334 & w4384;
assign v1252 = ~(w4284 | w4287);
assign w4386 = v1252;
assign w4387 = w4385 & w4386;
assign v1253 = ~(w4385 | w4386);
assign w4388 = v1253;
assign v1254 = ~(w4387 | w4388);
assign w4389 = v1254;
assign w4390 = w928 & w3758;
assign w4391 = w3399 & ~w3666;
assign w4392 = w3402 & ~w3587;
assign v1255 = ~(w4391 | w4392);
assign w4393 = v1255;
assign w4394 = w3406 & ~w3752;
assign w4395 = w4393 & ~w4394;
assign w4396 = ~w4390 & w4395;
assign w4397 = w4389 & ~w4396;
assign w4398 = ~w4389 & w4396;
assign v1256 = ~(w4397 | w4398);
assign w4399 = v1256;
assign v1257 = ~(w4299 | w4302);
assign w4400 = v1257;
assign w4401 = w4399 & ~w4400;
assign w4402 = ~w4399 & w4400;
assign v1258 = ~(w4401 | w4402);
assign w4403 = v1258;
assign w4404 = w4142 & ~w4144;
assign v1259 = ~(w4145 | w4404);
assign w4405 = v1259;
assign w4406 = w3529 & w4405;
assign w4407 = w3760 & ~w4035;
assign w4408 = w3767 & ~w3920;
assign w4409 = w3763 & ~w4134;
assign v1260 = ~(w4408 | w4409);
assign w4410 = v1260;
assign w4411 = ~w4407 & w4410;
assign w4412 = ~w4406 & w4411;
assign w4413 = pi29 & ~w4412;
assign w4414 = ~pi29 & w4412;
assign v1261 = ~(w4413 | w4414);
assign w4415 = v1261;
assign w4416 = w4403 & w4415;
assign v1262 = ~(w4403 | w4415);
assign w4417 = v1262;
assign v1263 = ~(w4416 | w4417);
assign w4418 = v1263;
assign w4419 = ~w4327 & w4418;
assign w4420 = w4327 & ~w4418;
assign v1264 = ~(w4419 | w4420);
assign w4421 = v1264;
assign w4422 = w4082 & ~w4168;
assign v1265 = ~(w4191 | w4422);
assign w4423 = v1265;
assign w4424 = w4191 & ~w4194;
assign v1266 = ~(w4423 | w4424);
assign w4425 = v1266;
assign w4426 = w4153 & w4425;
assign v1267 = ~(w2873 | w4082);
assign w4427 = v1267;
assign w4428 = w4158 & ~w4191;
assign v1268 = ~(w4427 | w4428);
assign w4429 = v1268;
assign w4430 = ~w4426 & w4429;
assign w4431 = ~pi26 & w4430;
assign w4432 = pi26 & ~w4430;
assign v1269 = ~(w4431 | w4432);
assign w4433 = v1269;
assign w4434 = w4421 & w4433;
assign v1270 = ~(w4421 | w4433);
assign w4435 = v1270;
assign v1271 = ~(w4434 | w4435);
assign w4436 = v1271;
assign w4437 = ~w4326 & w4436;
assign w4438 = ~w3506 & w3517;
assign v1272 = ~(w3518 | w4438);
assign w4439 = v1272;
assign w4440 = ~w1387 & w3767;
assign w4441 = w3529 & w4291;
assign w4442 = ~w3666 & w3763;
assign w4443 = ~w3587 & w3760;
assign v1273 = ~(w4442 | w4443);
assign w4444 = v1273;
assign w4445 = ~w4441 & w4444;
assign w4446 = ~w4440 & w4445;
assign w4447 = pi29 & w4446;
assign v1274 = ~(pi29 | w4446);
assign w4448 = v1274;
assign v1275 = ~(w4447 | w4448);
assign w4449 = v1275;
assign w4450 = w4439 & ~w4449;
assign w4451 = ~w420 & w2852;
assign w4452 = ~w945 & w4451;
assign w4453 = w1349 & w4452;
assign w4454 = w2932 & w4453;
assign w4455 = w3110 & w4454;
assign v1276 = ~(w253 | w469);
assign w4456 = v1276;
assign w4457 = ~w201 & w894;
assign w4458 = w4456 & w4457;
assign w4459 = w2076 & w2350;
assign w4460 = w1581 & w4459;
assign w4461 = w4458 & w4460;
assign w4462 = ~w251 & w339;
assign w4463 = w1786 & w4462;
assign w4464 = w129 & w4463;
assign w4465 = w4461 & w4464;
assign w4466 = w4096 & w4465;
assign w4467 = w1295 & w4466;
assign w4468 = w3696 & w4467;
assign w4469 = w4455 & w4468;
assign w4470 = w1642 & w2244;
assign w4471 = ~w448 & w4470;
assign w4472 = w1800 & w4471;
assign w4473 = ~w739 & w2526;
assign w4474 = ~w692 & w4473;
assign w4475 = ~w82 & w174;
assign w4476 = w121 & w1934;
assign w4477 = w4475 & w4476;
assign w4478 = w4474 & w4477;
assign w4479 = w4472 & w4478;
assign w4480 = w1916 & w2043;
assign w4481 = w1884 & w4480;
assign w4482 = w852 & w2350;
assign w4483 = w1681 & w4482;
assign w4484 = w4481 & w4483;
assign v1277 = ~(w132 | w281);
assign w4485 = v1277;
assign w4486 = w254 & w4485;
assign v1278 = ~(w78 | w1108);
assign w4487 = v1278;
assign v1279 = ~(w169 | w877);
assign w4488 = v1279;
assign w4489 = w4487 & w4488;
assign w4490 = w4486 & w4489;
assign v1280 = ~(w245 | w469);
assign w4491 = v1280;
assign w4492 = w3014 & w3733;
assign w4493 = w4491 & w4492;
assign w4494 = w4490 & w4493;
assign w4495 = w4484 & w4494;
assign w4496 = ~w629 & w1165;
assign w4497 = w1058 & w4496;
assign w4498 = w1870 & w3460;
assign w4499 = w4497 & w4498;
assign w4500 = w2116 & w4499;
assign w4501 = w4495 & w4500;
assign w4502 = w2393 & w3714;
assign v1281 = ~(w49 | w187);
assign w4503 = v1281;
assign v1282 = ~(w93 | w209);
assign w4504 = v1282;
assign w4505 = w4503 & w4504;
assign w4506 = w2316 & w4505;
assign w4507 = w4502 & w4506;
assign w4508 = w4501 & w4507;
assign w4509 = w4479 & w4508;
assign w4510 = w3643 & w4509;
assign w4511 = w4469 & w4510;
assign v1283 = ~(w4469 | w4510);
assign w4512 = v1283;
assign v1284 = ~(w4511 | w4512);
assign w4513 = v1284;
assign w4514 = pi17 & w4513;
assign v1285 = ~(w4511 | w4514);
assign w4515 = v1285;
assign w4516 = w1153 & w4515;
assign v1286 = ~(w1153 | w4515);
assign w4517 = v1286;
assign v1287 = ~(w4516 | w4517);
assign w4518 = v1287;
assign w4519 = ~w1798 & w3388;
assign v1288 = ~(w3389 | w4519);
assign w4520 = v1288;
assign w4521 = w928 & w4520;
assign w4522 = ~w1674 & w3406;
assign w4523 = ~w1860 & w3399;
assign v1289 = ~(w4522 | w4523);
assign w4524 = v1289;
assign w4525 = ~w1795 & w3402;
assign w4526 = w4524 & ~w4525;
assign w4527 = ~w4521 & w4526;
assign w4528 = w4518 & ~w4527;
assign v1290 = ~(w4516 | w4528);
assign w4529 = v1290;
assign v1291 = ~(w3490 | w3501);
assign w4530 = v1291;
assign v1292 = ~(w3502 | w4530);
assign w4531 = v1292;
assign v1293 = ~(w4529 | w4531);
assign w4532 = v1293;
assign w4533 = ~w4518 & w4527;
assign v1294 = ~(w4528 | w4533);
assign w4534 = v1294;
assign v1295 = ~(pi17 | w4513);
assign w4535 = v1295;
assign v1296 = ~(w4514 | w4535);
assign w4536 = v1296;
assign w4537 = ~w1863 & w3386;
assign v1297 = ~(w3387 | w4537);
assign w4538 = v1297;
assign w4539 = w928 & w4538;
assign w4540 = ~w1795 & w3406;
assign w4541 = ~w1860 & w3402;
assign v1298 = ~(w4540 | w4541);
assign w4542 = v1298;
assign w4543 = ~w1942 & w3399;
assign w4544 = w4542 & ~w4543;
assign w4545 = ~w4539 & w4544;
assign v1299 = ~(w4536 | w4545);
assign w4546 = v1299;
assign w4547 = w1729 & w2712;
assign w4548 = ~w141 & w667;
assign w4549 = ~w563 & w4548;
assign w4550 = ~w183 & w3304;
assign w4551 = ~w437 & w1442;
assign w4552 = w4550 & w4551;
assign w4553 = w4549 & w4552;
assign v1300 = ~(w282 | w291);
assign w4554 = v1300;
assign v1301 = ~(w68 | w238);
assign w4555 = v1301;
assign w4556 = w838 & w4555;
assign w4557 = w4554 & w4556;
assign w4558 = w4041 & w4557;
assign w4559 = w4553 & w4558;
assign w4560 = w4547 & w4559;
assign v1302 = ~(w77 | w605);
assign w4561 = v1302;
assign w4562 = w3194 & w4561;
assign w4563 = w625 & w3569;
assign w4564 = ~w989 & w3175;
assign w4565 = w4563 & w4564;
assign w4566 = w4562 & w4565;
assign w4567 = w4560 & w4566;
assign v1303 = ~(w221 | w899);
assign w4568 = v1303;
assign w4569 = ~w639 & w4568;
assign w4570 = ~w234 & w1396;
assign v1304 = ~(w123 | w463);
assign w4571 = v1304;
assign w4572 = w4570 & w4571;
assign w4573 = w4569 & w4572;
assign w4574 = w1092 & w4573;
assign v1305 = ~(w251 | w274);
assign w4575 = v1305;
assign w4576 = w1840 & w4575;
assign w4577 = w900 & w4576;
assign v1306 = ~(w231 | w481);
assign w4578 = v1306;
assign w4579 = w2766 & w4578;
assign w4580 = w4577 & w4579;
assign w4581 = w4574 & w4580;
assign w4582 = w969 & w1110;
assign w4583 = w2909 & w4582;
assign w4584 = w4581 & w4583;
assign w4585 = w1026 & w2974;
assign w4586 = w1562 & w4585;
assign w4587 = w117 & w4586;
assign v1307 = ~(w272 | w457);
assign w4588 = v1307;
assign w4589 = w943 & w4588;
assign w4590 = w2877 & w3220;
assign w4591 = w4589 & w4590;
assign w4592 = w4587 & w4591;
assign w4593 = w4584 & w4592;
assign w4594 = w4567 & w4593;
assign w4595 = ~w4469 & w4594;
assign v1308 = ~(w183 | w337);
assign w4596 = v1308;
assign w4597 = w156 & w4596;
assign w4598 = w665 & ~w1032;
assign w4599 = w3177 & w4598;
assign w4600 = ~w522 & w2256;
assign w4601 = w2486 & w4600;
assign v1309 = ~(w302 | w630);
assign w4602 = v1309;
assign w4603 = w4569 & w4602;
assign w4604 = w4601 & w4603;
assign w4605 = w1218 & w2181;
assign w4606 = w1889 & w3647;
assign w4607 = w4605 & w4606;
assign w4608 = w4604 & w4607;
assign w4609 = w4599 & w4608;
assign v1310 = ~(w212 | w385);
assign w4610 = v1310;
assign w4611 = ~w680 & w4610;
assign w4612 = w984 & w4611;
assign w4613 = w2078 & w3568;
assign w4614 = w4612 & w4613;
assign w4615 = ~w404 & w3304;
assign w4616 = w1068 & w4615;
assign w4617 = w4614 & w4616;
assign w4618 = w4609 & w4617;
assign v1311 = ~(w209 | w390);
assign w4619 = v1311;
assign w4620 = w760 & w2749;
assign w4621 = ~w168 & w174;
assign v1312 = ~(w405 | w548);
assign w4622 = v1312;
assign w4623 = w4621 & w4622;
assign w4624 = w4620 & w4623;
assign v1313 = ~(w21 | w742);
assign w4625 = v1313;
assign w4626 = w2272 & w4625;
assign w4627 = w4624 & w4626;
assign w4628 = w473 & w4627;
assign w4629 = w4619 & w4628;
assign w4630 = w4618 & w4629;
assign w4631 = w4597 & w4630;
assign w4632 = ~w398 & w2709;
assign w4633 = w1168 & w4632;
assign w4634 = w2398 & w3267;
assign v1314 = ~(w119 | w479);
assign w4635 = v1314;
assign w4636 = w2929 & w4635;
assign w4637 = w4634 & w4636;
assign w4638 = w4505 & w4637;
assign w4639 = w4633 & w4638;
assign w4640 = w1127 & w3589;
assign v1315 = ~(w441 | w1134);
assign w4641 = v1315;
assign w4642 = w2117 & w4641;
assign w4643 = w4640 & w4642;
assign w4644 = w3744 & w4643;
assign v1316 = ~(w127 | w303);
assign w4645 = v1316;
assign w4646 = w4253 & w4645;
assign w4647 = ~w27 & w4646;
assign w4648 = w4549 & w4647;
assign w4649 = w4644 & w4648;
assign w4650 = w4639 & w4649;
assign v1317 = ~(w499 | w624);
assign w4651 = v1317;
assign w4652 = w1650 & w4651;
assign w4653 = w810 & w4652;
assign w4654 = ~w77 & w4653;
assign v1318 = ~(w258 | w374);
assign w4655 = v1318;
assign w4656 = w1877 & w4655;
assign w4657 = w3048 & w4656;
assign w4658 = w1031 & w3706;
assign w4659 = w4657 & w4658;
assign w4660 = w4654 & w4659;
assign w4661 = w965 & w2156;
assign w4662 = w1612 & w4661;
assign v1319 = ~(w267 | w541);
assign w4663 = v1319;
assign w4664 = ~w291 & w4663;
assign w4665 = w1781 & w4664;
assign w4666 = w4662 & w4665;
assign w4667 = w996 & w2912;
assign w4668 = w4666 & w4667;
assign w4669 = ~w469 & w1041;
assign w4670 = w1020 & w4669;
assign w4671 = w4218 & w4670;
assign w4672 = w3469 & w4671;
assign w4673 = w4668 & w4672;
assign w4674 = w389 & ~w870;
assign w4675 = w2553 & w4674;
assign v1320 = ~(w111 | w414);
assign w4676 = v1320;
assign w4677 = ~w384 & w4676;
assign v1321 = ~(w298 | w369);
assign w4678 = v1321;
assign w4679 = ~w259 & w4678;
assign w4680 = w4677 & w4679;
assign w4681 = w1975 & w4680;
assign w4682 = w4675 & w4681;
assign w4683 = w1767 & w2193;
assign w4684 = w2440 & w2708;
assign v1322 = ~(w224 | w692);
assign w4685 = v1322;
assign w4686 = w1118 & w4685;
assign w4687 = w4684 & w4686;
assign w4688 = w4683 & w4687;
assign w4689 = w4682 & w4688;
assign w4690 = w4673 & w4689;
assign w4691 = w4660 & w4690;
assign w4692 = w4650 & w4691;
assign w4693 = w4631 & w4692;
assign v1323 = ~(w4631 | w4692);
assign w4694 = v1323;
assign v1324 = ~(w4693 | w4694);
assign w4695 = v1324;
assign w4696 = pi14 & w4695;
assign v1325 = ~(w4693 | w4696);
assign w4697 = v1325;
assign w4698 = w4594 & w4697;
assign v1326 = ~(w4594 | w4697);
assign w4699 = v1326;
assign v1327 = ~(w4698 | w4699);
assign w4700 = v1327;
assign v1328 = ~(w2041 | w3382);
assign w4701 = v1328;
assign v1329 = ~(w3383 | w4701);
assign w4702 = v1329;
assign w4703 = w928 & w4702;
assign w4704 = ~w2038 & w3402;
assign w4705 = ~w2089 & w3399;
assign v1330 = ~(w4704 | w4705);
assign w4706 = v1330;
assign w4707 = ~w1942 & w3406;
assign w4708 = w4706 & ~w4707;
assign w4709 = ~w4703 & w4708;
assign w4710 = w4700 & ~w4709;
assign v1331 = ~(w4698 | w4710);
assign w4711 = v1331;
assign w4712 = w4469 & ~w4594;
assign v1332 = ~(w4595 | w4712);
assign w4713 = v1332;
assign w4714 = w4711 & w4713;
assign v1333 = ~(w4595 | w4714);
assign w4715 = v1333;
assign w4716 = w4536 & w4545;
assign v1334 = ~(w4546 | w4716);
assign w4717 = v1334;
assign w4718 = w4715 & w4717;
assign v1335 = ~(w4546 | w4718);
assign w4719 = v1335;
assign w4720 = w4534 & ~w4719;
assign w4721 = ~w4534 & w4719;
assign v1336 = ~(w4720 | w4721);
assign w4722 = v1336;
assign w4723 = w3397 & w3529;
assign w4724 = ~w1496 & w3763;
assign w4725 = ~w1387 & w3760;
assign v1337 = ~(w4724 | w4725);
assign w4726 = v1337;
assign w4727 = ~w1609 & w3767;
assign w4728 = w4726 & ~w4727;
assign w4729 = ~w4723 & w4728;
assign w4730 = ~pi29 & w4729;
assign w4731 = pi29 & ~w4729;
assign v1338 = ~(w4730 | w4731);
assign w4732 = v1338;
assign w4733 = w4722 & w4732;
assign v1339 = ~(w4720 | w4733);
assign w4734 = v1339;
assign w4735 = w4529 & w4531;
assign v1340 = ~(w4532 | w4735);
assign w4736 = v1340;
assign w4737 = ~w4734 & w4736;
assign v1341 = ~(w4532 | w4737);
assign w4738 = v1341;
assign w4739 = ~w4439 & w4449;
assign v1342 = ~(w4450 | w4739);
assign w4740 = v1342;
assign w4741 = ~w4738 & w4740;
assign v1343 = ~(w4450 | w4741);
assign w4742 = v1343;
assign v1344 = ~(w3522 | w3773);
assign w4743 = v1344;
assign v1345 = ~(w3774 | w4743);
assign w4744 = v1345;
assign w4745 = ~w4742 & w4744;
assign w4746 = w4742 & ~w4744;
assign v1346 = ~(w4745 | w4746);
assign w4747 = v1346;
assign w4748 = w4153 & w4405;
assign w4749 = ~w4035 & w4155;
assign w4750 = ~w4134 & w4158;
assign v1347 = ~(w4749 | w4750);
assign w4751 = v1347;
assign v1348 = ~(w2873 | w3920);
assign w4752 = v1348;
assign w4753 = w4751 & ~w4752;
assign w4754 = ~w4748 & w4753;
assign w4755 = ~pi26 & w4754;
assign w4756 = pi26 & ~w4754;
assign v1349 = ~(w4755 | w4756);
assign w4757 = v1349;
assign w4758 = w4747 & w4757;
assign v1350 = ~(w4745 | w4758);
assign w4759 = v1350;
assign v1351 = ~(pi22 | pi23);
assign w4760 = v1351;
assign w4761 = pi22 & pi23;
assign v1352 = ~(w4760 | w4761);
assign w4762 = v1352;
assign w4763 = w11 & w4762;
assign w4764 = w10 & w4762;
assign w4765 = ~w4422 & w4764;
assign v1353 = ~(w4763 | w4765);
assign w4766 = v1353;
assign v1354 = ~(w4191 | w4766);
assign w4767 = v1354;
assign w4768 = ~pi23 & w4767;
assign w4769 = pi23 & ~w4767;
assign v1355 = ~(w4768 | w4769);
assign w4770 = v1355;
assign v1356 = ~(w4759 | w4770);
assign w4771 = v1356;
assign v1357 = ~(w3940 | w4165);
assign w4772 = v1357;
assign v1358 = ~(w4166 | w4772);
assign w4773 = v1358;
assign w4774 = w4759 & w4770;
assign v1359 = ~(w4771 | w4774);
assign w4775 = v1359;
assign w4776 = w4773 & w4775;
assign v1360 = ~(w4771 | w4776);
assign w4777 = v1360;
assign v1361 = ~(w4322 | w4324);
assign w4778 = v1361;
assign v1362 = ~(w4325 | w4778);
assign w4779 = v1362;
assign w4780 = ~w4777 & w4779;
assign w4781 = w4777 & ~w4779;
assign v1363 = ~(w4780 | w4781);
assign w4782 = v1363;
assign v1364 = ~(w4773 | w4775);
assign w4783 = v1364;
assign v1365 = ~(w4776 | w4783);
assign w4784 = v1365;
assign w4785 = w4738 & ~w4740;
assign v1366 = ~(w4741 | w4785);
assign w4786 = v1366;
assign w4787 = w4153 & w4309;
assign w4788 = ~w3920 & w4158;
assign v1367 = ~(w2873 | w3752);
assign w4789 = v1367;
assign w4790 = ~w4134 & w4155;
assign v1368 = ~(w4789 | w4790);
assign w4791 = v1368;
assign w4792 = ~w4788 & w4791;
assign w4793 = ~w4787 & w4792;
assign w4794 = pi26 & ~w4793;
assign w4795 = ~pi26 & w4793;
assign v1369 = ~(w4794 | w4795);
assign w4796 = v1369;
assign w4797 = w4786 & w4796;
assign w4798 = w4734 & ~w4736;
assign v1370 = ~(w4737 | w4798);
assign w4799 = v1370;
assign w4800 = w3529 & w3843;
assign w4801 = ~w3666 & w3760;
assign w4802 = ~w1496 & w3767;
assign w4803 = ~w1387 & w3763;
assign v1371 = ~(w4802 | w4803);
assign w4804 = v1371;
assign w4805 = ~w4801 & w4804;
assign w4806 = ~w4800 & w4805;
assign w4807 = pi29 & ~w4806;
assign w4808 = ~pi29 & w4806;
assign v1372 = ~(w4807 | w4808);
assign w4809 = v1372;
assign w4810 = w4799 & w4809;
assign v1373 = ~(w4799 | w4809);
assign w4811 = v1373;
assign v1374 = ~(w4810 | w4811);
assign w4812 = v1374;
assign w4813 = ~w3928 & w4153;
assign w4814 = ~w3920 & w4155;
assign w4815 = ~w3752 & w4158;
assign v1375 = ~(w4814 | w4815);
assign w4816 = v1375;
assign v1376 = ~(w2873 | w3587);
assign w4817 = v1376;
assign w4818 = w4816 & ~w4817;
assign w4819 = ~w4813 & w4818;
assign w4820 = ~pi26 & w4819;
assign w4821 = pi26 & ~w4819;
assign v1377 = ~(w4820 | w4821);
assign w4822 = v1377;
assign w4823 = w4812 & w4822;
assign v1378 = ~(w4810 | w4823);
assign w4824 = v1378;
assign v1379 = ~(w4786 | w4796);
assign w4825 = v1379;
assign v1380 = ~(w4797 | w4825);
assign w4826 = v1380;
assign w4827 = ~w4824 & w4826;
assign v1381 = ~(w4797 | w4827);
assign w4828 = v1381;
assign v1382 = ~(w4747 | w4757);
assign w4829 = v1382;
assign v1383 = ~(w4758 | w4829);
assign w4830 = v1383;
assign w4831 = ~w4828 & w4830;
assign w4832 = w4828 & ~w4830;
assign v1384 = ~(w4831 | w4832);
assign w4833 = v1384;
assign w4834 = w4425 & w4764;
assign w4835 = ~w4082 & w4763;
assign w4836 = w7 & ~w10;
assign w4837 = ~w4191 & w4836;
assign v1385 = ~(w4835 | w4837);
assign w4838 = v1385;
assign w4839 = ~w4834 & w4838;
assign w4840 = ~pi23 & w4839;
assign w4841 = pi23 & ~w4839;
assign v1386 = ~(w4840 | w4841);
assign w4842 = v1386;
assign w4843 = w4833 & w4842;
assign v1387 = ~(w4831 | w4843);
assign w4844 = v1387;
assign w4845 = w4784 & ~w4844;
assign w4846 = ~w4784 & w4844;
assign v1388 = ~(w4812 | w4822);
assign w4847 = v1388;
assign v1389 = ~(w4823 | w4847);
assign w4848 = v1389;
assign v1390 = ~(w4711 | w4713);
assign w4849 = v1390;
assign v1391 = ~(w4714 | w4849);
assign w4850 = v1391;
assign v1392 = ~(w1943 | w1944);
assign w4851 = v1392;
assign w4852 = w3384 & ~w4851;
assign w4853 = ~w3384 & w4851;
assign v1393 = ~(w4852 | w4853);
assign w4854 = v1393;
assign w4855 = w928 & w4854;
assign w4856 = ~w1860 & w3406;
assign w4857 = ~w2038 & w3399;
assign v1394 = ~(w4856 | w4857);
assign w4858 = v1394;
assign w4859 = ~w1942 & w3402;
assign w4860 = w4858 & ~w4859;
assign w4861 = ~w4855 & w4860;
assign v1395 = ~(w4850 | w4861);
assign w4862 = v1395;
assign w4863 = w4850 & w4861;
assign v1396 = ~(w4862 | w4863);
assign w4864 = v1396;
assign w4865 = w3494 & w3529;
assign w4866 = ~w1609 & w3760;
assign w4867 = ~w1674 & w3763;
assign v1397 = ~(w4866 | w4867);
assign w4868 = v1397;
assign w4869 = ~w1795 & w3767;
assign w4870 = w4868 & ~w4869;
assign w4871 = ~w4865 & w4870;
assign w4872 = ~pi29 & w4871;
assign w4873 = pi29 & ~w4871;
assign v1398 = ~(w4872 | w4873);
assign w4874 = v1398;
assign w4875 = w4864 & w4874;
assign v1399 = ~(w4862 | w4875);
assign w4876 = v1399;
assign v1400 = ~(w4715 | w4717);
assign w4877 = v1400;
assign v1401 = ~(w4718 | w4877);
assign w4878 = v1401;
assign w4879 = ~w4876 & w4878;
assign w4880 = w4876 & ~w4878;
assign v1402 = ~(w4879 | w4880);
assign w4881 = v1402;
assign w4882 = ~w3510 & w3529;
assign w4883 = ~w1496 & w3760;
assign w4884 = ~w1609 & w3763;
assign v1403 = ~(w4883 | w4884);
assign w4885 = v1403;
assign w4886 = ~w1674 & w3767;
assign w4887 = w4885 & ~w4886;
assign w4888 = ~w4882 & w4887;
assign w4889 = ~pi29 & w4888;
assign w4890 = pi29 & ~w4888;
assign v1404 = ~(w4889 | w4890);
assign w4891 = v1404;
assign w4892 = w4881 & w4891;
assign v1405 = ~(w4879 | w4892);
assign w4893 = v1405;
assign v1406 = ~(w4722 | w4732);
assign w4894 = v1406;
assign v1407 = ~(w4733 | w4894);
assign w4895 = v1407;
assign w4896 = ~w4893 & w4895;
assign w4897 = w4893 & ~w4895;
assign v1408 = ~(w4896 | w4897);
assign w4898 = v1408;
assign w4899 = w3758 & w4153;
assign w4900 = ~w3752 & w4155;
assign v1409 = ~(w2873 | w3666);
assign w4901 = v1409;
assign w4902 = ~w3587 & w4158;
assign v1410 = ~(w4901 | w4902);
assign w4903 = v1410;
assign w4904 = ~w4900 & w4903;
assign w4905 = ~w4899 & w4904;
assign w4906 = pi26 & ~w4905;
assign w4907 = ~pi26 & w4905;
assign v1411 = ~(w4906 | w4907);
assign w4908 = v1411;
assign w4909 = w4898 & w4908;
assign v1412 = ~(w4896 | w4909);
assign w4910 = v1412;
assign w4911 = w4848 & ~w4910;
assign w4912 = ~w4149 & w4764;
assign w4913 = w10 & ~w4762;
assign w4914 = ~w4082 & w4913;
assign w4915 = ~w4134 & w4763;
assign w4916 = ~w4035 & w4836;
assign v1413 = ~(w4915 | w4916);
assign w4917 = v1413;
assign w4918 = ~w4914 & w4917;
assign w4919 = ~w4912 & w4918;
assign w4920 = pi23 & ~w4919;
assign w4921 = ~pi23 & w4919;
assign v1414 = ~(w4920 | w4921);
assign w4922 = v1414;
assign w4923 = ~w4848 & w4910;
assign v1415 = ~(w4911 | w4923);
assign w4924 = v1415;
assign w4925 = w4922 & w4924;
assign v1416 = ~(w4911 | w4925);
assign w4926 = v1416;
assign w4927 = w4196 & w4764;
assign w4928 = ~w4082 & w4836;
assign w4929 = ~w4191 & w4913;
assign w4930 = ~w4035 & w4763;
assign v1417 = ~(w4929 | w4930);
assign w4931 = v1417;
assign w4932 = ~w4928 & w4931;
assign w4933 = ~w4927 & w4932;
assign w4934 = pi23 & ~w4933;
assign w4935 = ~pi23 & w4933;
assign v1418 = ~(w4934 | w4935);
assign w4936 = v1418;
assign w4937 = ~w4926 & w4936;
assign w4938 = w4824 & ~w4826;
assign v1419 = ~(w4827 | w4938);
assign w4939 = v1419;
assign w4940 = w4926 & ~w4936;
assign v1420 = ~(w4937 | w4940);
assign w4941 = v1420;
assign w4942 = w4939 & w4941;
assign v1421 = ~(w4937 | w4942);
assign w4943 = v1421;
assign v1422 = ~(w4833 | w4842);
assign w4944 = v1422;
assign v1423 = ~(w4843 | w4944);
assign w4945 = v1423;
assign w4946 = ~w4943 & w4945;
assign v1424 = ~(w4939 | w4941);
assign w4947 = v1424;
assign v1425 = ~(w4942 | w4947);
assign w4948 = v1425;
assign v1426 = ~(w4898 | w4908);
assign w4949 = v1426;
assign v1427 = ~(w4909 | w4949);
assign w4950 = v1427;
assign v1428 = ~(w4881 | w4891);
assign w4951 = v1428;
assign v1429 = ~(w4892 | w4951);
assign w4952 = v1429;
assign w4953 = ~w3587 & w4155;
assign w4954 = w4153 & w4291;
assign w4955 = ~w3666 & w4158;
assign v1430 = ~(w1387 | w2873);
assign w4956 = v1430;
assign v1431 = ~(w4955 | w4956);
assign w4957 = v1431;
assign w4958 = ~w4954 & w4957;
assign w4959 = ~w4953 & w4958;
assign w4960 = pi26 & w4959;
assign v1432 = ~(pi26 | w4959);
assign w4961 = v1432;
assign v1433 = ~(w4960 | w4961);
assign w4962 = v1433;
assign w4963 = w4952 & ~w4962;
assign w4964 = ~w4700 & w4709;
assign v1434 = ~(w4710 | w4964);
assign w4965 = v1434;
assign v1435 = ~(pi14 | w4695);
assign w4966 = v1435;
assign v1436 = ~(w4696 | w4966);
assign w4967 = v1436;
assign w4968 = ~w381 & w2955;
assign w4969 = ~w187 & w4968;
assign w4970 = ~w98 & w1490;
assign w4971 = w1330 & w4970;
assign w4972 = w4456 & w4971;
assign w4973 = w4969 & w4972;
assign v1437 = ~(w272 | w630);
assign w4974 = v1437;
assign w4975 = w3624 & w4974;
assign w4976 = w3475 & w4975;
assign w4977 = w1814 & w2043;
assign v1438 = ~(w162 | w398);
assign w4978 = v1438;
assign w4979 = w4977 & w4978;
assign w4980 = w4976 & w4979;
assign w4981 = w386 & w626;
assign v1439 = ~(w53 | w699);
assign w4982 = v1439;
assign w4983 = w4981 & w4982;
assign w4984 = w1428 & w4983;
assign w4985 = w4980 & w4984;
assign w4986 = w4973 & w4985;
assign v1440 = ~(w286 | w559);
assign w4987 = v1440;
assign w4988 = w506 & w4987;
assign v1441 = ~(w131 | w140);
assign w4989 = v1441;
assign w4990 = w1470 & w4989;
assign w4991 = ~w674 & w4990;
assign w4992 = w4988 & w4991;
assign v1442 = ~(w127 | w311);
assign w4993 = v1442;
assign w4994 = ~w99 & w4993;
assign w4995 = ~w308 & w4994;
assign w4996 = w1129 & w1281;
assign w4997 = w4995 & w4996;
assign w4998 = w4992 & w4997;
assign w4999 = w171 & w2824;
assign v1443 = ~(w82 | w231);
assign w5000 = v1443;
assign v1444 = ~(w183 | w447);
assign w5001 = v1444;
assign w5002 = w5000 & w5001;
assign w5003 = w4999 & w5002;
assign w5004 = w2465 & w4010;
assign w5005 = ~w264 & w5004;
assign w5006 = w1799 & w4371;
assign v1445 = ~(w202 | w888);
assign w5007 = v1445;
assign w5008 = w5006 & w5007;
assign w5009 = w5005 & w5008;
assign w5010 = w5003 & w5009;
assign w5011 = w4998 & w5010;
assign v1446 = ~(w184 | w640);
assign w5012 = v1446;
assign w5013 = w178 & w5012;
assign w5014 = w2820 & w5013;
assign w5015 = w483 & w2381;
assign w5016 = w5014 & w5015;
assign w5017 = w5011 & w5016;
assign w5018 = w2626 & w2728;
assign w5019 = ~w300 & w1679;
assign w5020 = ~w172 & w1008;
assign w5021 = w1033 & w5020;
assign w5022 = w5019 & w5021;
assign w5023 = w1263 & w5022;
assign w5024 = w5018 & w5023;
assign w5025 = w436 & w2642;
assign w5026 = w5024 & w5025;
assign w5027 = w5017 & w5026;
assign w5028 = w4986 & w5027;
assign w5029 = ~w4631 & w5028;
assign w5030 = w4631 & ~w5028;
assign v1447 = ~(w5029 | w5030);
assign w5031 = v1447;
assign w5032 = w3376 & ~w3378;
assign v1448 = ~(w3379 | w5032);
assign w5033 = v1448;
assign w5034 = w928 & w5033;
assign w5035 = ~w2202 & w3402;
assign w5036 = ~w2089 & w3406;
assign v1449 = ~(w5035 | w5036);
assign w5037 = v1449;
assign w5038 = ~w2290 & w3399;
assign w5039 = w5037 & ~w5038;
assign w5040 = ~w5034 & w5039;
assign w5041 = w5031 & w5040;
assign v1450 = ~(w5029 | w5041);
assign w5042 = v1450;
assign w5043 = ~w4967 & w5042;
assign w5044 = w4967 & ~w5042;
assign v1451 = ~(w5043 | w5044);
assign w5045 = v1451;
assign v1452 = ~(w2090 | w2091);
assign w5046 = v1452;
assign w5047 = w3380 & ~w5046;
assign w5048 = ~w3380 & w5046;
assign v1453 = ~(w5047 | w5048);
assign w5049 = v1453;
assign w5050 = w928 & w5049;
assign w5051 = ~w2202 & w3399;
assign w5052 = ~w2089 & w3402;
assign v1454 = ~(w5051 | w5052);
assign w5053 = v1454;
assign w5054 = ~w2038 & w3406;
assign w5055 = w5053 & ~w5054;
assign w5056 = ~w5050 & w5055;
assign w5057 = w5045 & ~w5056;
assign v1455 = ~(w5043 | w5057);
assign w5058 = v1455;
assign w5059 = w4965 & ~w5058;
assign w5060 = ~w4965 & w5058;
assign v1456 = ~(w5059 | w5060);
assign w5061 = v1456;
assign w5062 = w3529 & w4520;
assign w5063 = ~w1795 & w3763;
assign w5064 = ~w1674 & w3760;
assign w5065 = ~w1860 & w3767;
assign v1457 = ~(w5064 | w5065);
assign w5066 = v1457;
assign w5067 = ~w5063 & w5066;
assign w5068 = ~w5062 & w5067;
assign w5069 = pi29 & ~w5068;
assign w5070 = ~pi29 & w5068;
assign v1458 = ~(w5069 | w5070);
assign w5071 = v1458;
assign w5072 = w5061 & w5071;
assign v1459 = ~(w5059 | w5072);
assign w5073 = v1459;
assign v1460 = ~(w4864 | w4874);
assign w5074 = v1460;
assign v1461 = ~(w4875 | w5074);
assign w5075 = v1461;
assign w5076 = ~w5073 & w5075;
assign w5077 = w3843 & w4153;
assign v1462 = ~(w1496 | w2873);
assign w5078 = v1462;
assign w5079 = ~w3666 & w4155;
assign w5080 = ~w1387 & w4158;
assign v1463 = ~(w5079 | w5080);
assign w5081 = v1463;
assign w5082 = ~w5078 & w5081;
assign w5083 = ~w5077 & w5082;
assign w5084 = pi26 & ~w5083;
assign w5085 = ~pi26 & w5083;
assign v1464 = ~(w5084 | w5085);
assign w5086 = v1464;
assign w5087 = w5073 & ~w5075;
assign v1465 = ~(w5076 | w5087);
assign w5088 = v1465;
assign w5089 = w5086 & w5088;
assign v1466 = ~(w5076 | w5089);
assign w5090 = v1466;
assign w5091 = ~w4952 & w4962;
assign v1467 = ~(w4963 | w5091);
assign w5092 = v1467;
assign w5093 = ~w5090 & w5092;
assign v1468 = ~(w4963 | w5093);
assign w5094 = v1468;
assign w5095 = w4950 & ~w5094;
assign w5096 = ~w4950 & w5094;
assign v1469 = ~(w5095 | w5096);
assign w5097 = v1469;
assign w5098 = w4405 & w4764;
assign w5099 = ~w4035 & w4913;
assign w5100 = ~w4134 & w4836;
assign v1470 = ~(w5099 | w5100);
assign w5101 = v1470;
assign w5102 = ~w3920 & w4763;
assign w5103 = w5101 & ~w5102;
assign w5104 = ~w5098 & w5103;
assign w5105 = pi23 & w5104;
assign v1471 = ~(pi23 | w5104);
assign w5106 = v1471;
assign v1472 = ~(w5105 | w5106);
assign w5107 = v1472;
assign w5108 = w5097 & ~w5107;
assign v1473 = ~(w5095 | w5108);
assign w5109 = v1473;
assign v1474 = ~(pi19 | pi20);
assign w5110 = v1474;
assign w5111 = pi19 & pi20;
assign v1475 = ~(w5110 | w5111);
assign w5112 = v1475;
assign w5113 = w916 & w5112;
assign w5114 = w912 & w5112;
assign w5115 = ~w4422 & w5114;
assign v1476 = ~(w5113 | w5115);
assign w5116 = v1476;
assign v1477 = ~(w4191 | w5116);
assign w5117 = v1477;
assign w5118 = ~pi20 & w5117;
assign w5119 = pi20 & ~w5117;
assign v1478 = ~(w5118 | w5119);
assign w5120 = v1478;
assign v1479 = ~(w5109 | w5120);
assign w5121 = v1479;
assign v1480 = ~(w4922 | w4924);
assign w5122 = v1480;
assign v1481 = ~(w4925 | w5122);
assign w5123 = v1481;
assign w5124 = w5109 & w5120;
assign v1482 = ~(w5121 | w5124);
assign w5125 = v1482;
assign w5126 = w5123 & w5125;
assign v1483 = ~(w5121 | w5126);
assign w5127 = v1483;
assign w5128 = w4948 & ~w5127;
assign w5129 = ~w4948 & w5127;
assign v1484 = ~(w5128 | w5129);
assign w5130 = v1484;
assign v1485 = ~(w5123 | w5125);
assign w5131 = v1485;
assign v1486 = ~(w5126 | w5131);
assign w5132 = v1486;
assign w5133 = ~w5097 & w5107;
assign v1487 = ~(w5108 | w5133);
assign w5134 = v1487;
assign w5135 = w5090 & ~w5092;
assign v1488 = ~(w5093 | w5135);
assign w5136 = v1488;
assign w5137 = w4309 & w4764;
assign w5138 = ~w3920 & w4836;
assign w5139 = ~w3752 & w4763;
assign w5140 = ~w4134 & w4913;
assign v1489 = ~(w5139 | w5140);
assign w5141 = v1489;
assign w5142 = ~w5138 & w5141;
assign w5143 = ~w5137 & w5142;
assign w5144 = pi23 & ~w5143;
assign w5145 = ~pi23 & w5143;
assign v1490 = ~(w5144 | w5145);
assign w5146 = v1490;
assign w5147 = w5136 & w5146;
assign v1491 = ~(w5086 | w5088);
assign w5148 = v1491;
assign v1492 = ~(w5089 | w5148);
assign w5149 = v1492;
assign w5150 = ~w5045 & w5056;
assign v1493 = ~(w5057 | w5150);
assign w5151 = v1493;
assign w5152 = w3529 & w4538;
assign w5153 = ~w1860 & w3763;
assign w5154 = ~w1942 & w3767;
assign v1494 = ~(w5153 | w5154);
assign w5155 = v1494;
assign w5156 = ~w1795 & w3760;
assign w5157 = w5155 & ~w5156;
assign w5158 = ~w5152 & w5157;
assign w5159 = ~pi29 & w5158;
assign w5160 = pi29 & ~w5158;
assign v1495 = ~(w5159 | w5160);
assign w5161 = v1495;
assign w5162 = w5151 & w5161;
assign v1496 = ~(w37 | w474);
assign w5163 = v1496;
assign w5164 = w698 & w5163;
assign w5165 = ~w200 & w2672;
assign w5166 = ~w438 & w5165;
assign w5167 = w5164 & w5166;
assign w5168 = w964 & w2157;
assign v1497 = ~(w112 | w300);
assign w5169 = v1497;
assign v1498 = ~(w258 | w1207);
assign w5170 = v1498;
assign w5171 = ~w145 & w5170;
assign w5172 = w5169 & w5171;
assign w5173 = w5168 & w5172;
assign v1499 = ~(w135 | w558);
assign w5174 = v1499;
assign v1500 = ~(w195 | w223);
assign w5175 = v1500;
assign w5176 = w3580 & w5175;
assign w5177 = w5174 & w5176;
assign w5178 = w2561 & w3992;
assign w5179 = w5177 & w5178;
assign w5180 = w5173 & w5179;
assign w5181 = w5167 & w5180;
assign w5182 = w2404 & w4571;
assign w5183 = w1186 & w5182;
assign w5184 = w5181 & w5183;
assign w5185 = w210 & w4678;
assign w5186 = ~w235 & w3723;
assign w5187 = ~w248 & w752;
assign w5188 = w5186 & w5187;
assign w5189 = w5185 & w5188;
assign w5190 = w366 & w2960;
assign w5191 = w789 & w4097;
assign w5192 = w5190 & w5191;
assign w5193 = w4181 & w5192;
assign w5194 = w5189 & w5193;
assign w5195 = w4624 & w5194;
assign v1501 = ~(w176 | w379);
assign w5196 = v1501;
assign w5197 = ~w191 & w5196;
assign w5198 = ~w1134 & w1681;
assign w5199 = w5197 & w5198;
assign w5200 = ~w629 & w5199;
assign w5201 = w5195 & w5200;
assign v1502 = ~(w167 | w533);
assign w5202 = v1502;
assign w5203 = ~w566 & w5202;
assign w5204 = w285 & w5203;
assign w5205 = w1377 & w5204;
assign w5206 = w5201 & w5205;
assign w5207 = w5184 & w5206;
assign w5208 = w1033 & w3102;
assign v1503 = ~(w201 | w559);
assign w5209 = v1503;
assign w5210 = ~w143 & w5209;
assign w5211 = w5208 & w5210;
assign w5212 = ~w168 & w2022;
assign w5213 = ~w564 & w5212;
assign w5214 = w716 & w5213;
assign w5215 = w5211 & w5214;
assign v1504 = ~(w317 | w488);
assign w5216 = v1504;
assign w5217 = w1414 & w5216;
assign v1505 = ~(w169 | w438);
assign w5218 = v1505;
assign w5219 = w5217 & w5218;
assign w5220 = w1659 & w5219;
assign w5221 = w1934 & w2505;
assign v1506 = ~(w398 | w503);
assign w5222 = v1506;
assign w5223 = w681 & w823;
assign w5224 = w5222 & w5223;
assign w5225 = w5221 & w5224;
assign w5226 = ~w108 & w440;
assign w5227 = w846 & w5226;
assign v1507 = ~(w374 | w692);
assign w5228 = v1507;
assign w5229 = w5227 & w5228;
assign w5230 = w5225 & w5229;
assign w5231 = w5220 & w5230;
assign w5232 = w5215 & w5231;
assign w5233 = w1905 & w1952;
assign w5234 = w52 & w1780;
assign w5235 = w1829 & w5234;
assign w5236 = w5233 & w5235;
assign v1508 = ~(w68 | w727);
assign w5237 = v1508;
assign w5238 = w1682 & w5237;
assign w5239 = w382 & w2835;
assign w5240 = w5238 & w5239;
assign w5241 = w5236 & w5240;
assign w5242 = w3799 & w5241;
assign v1509 = ~(w37 | w456);
assign w5243 = v1509;
assign w5244 = ~w258 & w5243;
assign w5245 = ~w652 & w5244;
assign w5246 = w313 & w5245;
assign w5247 = w1102 & w5246;
assign w5248 = w5194 & w5247;
assign w5249 = w818 & w2854;
assign w5250 = w5248 & w5249;
assign w5251 = w5242 & w5250;
assign w5252 = w5232 & w5251;
assign w5253 = w5207 & w5252;
assign v1510 = ~(w5207 | w5252);
assign w5254 = v1510;
assign v1511 = ~(w5253 | w5254);
assign w5255 = v1511;
assign w5256 = pi11 & w5255;
assign v1512 = ~(w5253 | w5256);
assign w5257 = v1512;
assign w5258 = w4631 & w5257;
assign v1513 = ~(w4631 | w5257);
assign w5259 = v1513;
assign v1514 = ~(w5258 | w5259);
assign w5260 = v1514;
assign w5261 = w3372 & ~w3374;
assign v1515 = ~(w3375 | w5261);
assign w5262 = v1515;
assign w5263 = w928 & w5262;
assign w5264 = ~w2202 & w3406;
assign w5265 = ~w2339 & w3399;
assign v1516 = ~(w5264 | w5265);
assign w5266 = v1516;
assign w5267 = ~w2290 & w3402;
assign w5268 = w5266 & ~w5267;
assign w5269 = ~w5263 & w5268;
assign w5270 = w5260 & ~w5269;
assign v1517 = ~(w5258 | w5270);
assign w5271 = v1517;
assign v1518 = ~(w5031 | w5040);
assign w5272 = v1518;
assign v1519 = ~(w5041 | w5272);
assign w5273 = v1519;
assign v1520 = ~(w5271 | w5273);
assign w5274 = v1520;
assign w5275 = ~w5260 & w5269;
assign v1521 = ~(w5270 | w5275);
assign w5276 = v1521;
assign v1522 = ~(pi11 | w5255);
assign w5277 = v1522;
assign v1523 = ~(w5256 | w5277);
assign w5278 = v1523;
assign w5279 = w3368 & ~w3370;
assign v1524 = ~(w3371 | w5279);
assign w5280 = v1524;
assign w5281 = w928 & w5280;
assign w5282 = ~w2424 & w3399;
assign w5283 = ~w2339 & w3402;
assign v1525 = ~(w5282 | w5283);
assign w5284 = v1525;
assign w5285 = ~w2290 & w3406;
assign w5286 = w5284 & ~w5285;
assign w5287 = ~w5281 & w5286;
assign v1526 = ~(w5278 | w5287);
assign w5288 = v1526;
assign w5289 = ~w125 & w2319;
assign w5290 = ~w245 & w5289;
assign w5291 = ~w384 & w2156;
assign w5292 = ~w739 & w5291;
assign w5293 = w5290 & w5292;
assign w5294 = w3821 & w5293;
assign w5295 = w2422 & w5294;
assign w5296 = w1980 & w2076;
assign w5297 = ~w541 & w5296;
assign w5298 = ~w369 & w5297;
assign v1527 = ~(w258 | w281);
assign w5299 = v1527;
assign w5300 = w5298 & w5299;
assign w5301 = w3009 & w3071;
assign w5302 = w703 & w2661;
assign w5303 = w5163 & w5302;
assign w5304 = w5301 & w5303;
assign w5305 = w2378 & w5304;
assign w5306 = w5300 & w5305;
assign w5307 = w954 & w1751;
assign w5308 = w5306 & w5307;
assign w5309 = w5295 & w5308;
assign w5310 = ~w5207 & w5309;
assign v1528 = ~(w99 | w666);
assign w5311 = v1528;
assign w5312 = ~w369 & w5311;
assign w5313 = w4588 & w5312;
assign w5314 = w2870 & w5313;
assign w5315 = ~w241 & w5314;
assign w5316 = w1001 & w1915;
assign w5317 = w2315 & w5316;
assign w5318 = w5315 & w5317;
assign w5319 = ~w550 & w1632;
assign v1529 = ~(w31 | w53);
assign w5320 = v1529;
assign w5321 = w5319 & w5320;
assign w5322 = w967 & w3904;
assign w5323 = w5321 & w5322;
assign v1530 = ~(w522 | w731);
assign w5324 = v1530;
assign w5325 = w3818 & w5324;
assign w5326 = w4119 & w5325;
assign v1531 = ~(w131 | w564);
assign w5327 = v1531;
assign w5328 = ~w685 & w5327;
assign w5329 = ~w639 & w5328;
assign w5330 = w5326 & w5329;
assign w5331 = ~w173 & w468;
assign w5332 = ~w299 & w5331;
assign w5333 = w5330 & w5332;
assign w5334 = w5323 & w5333;
assign w5335 = w5318 & w5334;
assign v1532 = ~(w42 | w1032);
assign w5336 = v1532;
assign w5337 = ~w438 & w5336;
assign w5338 = w2768 & w4676;
assign w5339 = w283 & w5338;
assign w5340 = w5337 & w5339;
assign v1533 = ~(w381 | w1134);
assign w5341 = v1533;
assign w5342 = w5226 & w5341;
assign w5343 = w5340 & w5342;
assign v1534 = ~(w95 | w989);
assign w5344 = v1534;
assign w5345 = w583 & w5344;
assign w5346 = w5343 & w5345;
assign w5347 = w5335 & w5346;
assign w5348 = ~w484 & w4654;
assign w5349 = w3076 & w3241;
assign w5350 = w1007 & w1154;
assign w5351 = w5349 & w5350;
assign v1535 = ~(w172 | w874);
assign w5352 = v1535;
assign w5353 = w1666 & w2849;
assign w5354 = w5352 & w5353;
assign w5355 = w5351 & w5354;
assign w5356 = ~w70 & w358;
assign v1536 = ~(w56 | w877);
assign w5357 = v1536;
assign w5358 = w1414 & w5357;
assign w5359 = w1088 & w5358;
assign w5360 = w5356 & w5359;
assign w5361 = w5355 & w5360;
assign w5362 = w5348 & w5361;
assign v1537 = ~(w110 | w656);
assign w5363 = v1537;
assign v1538 = ~(w343 | w505);
assign w5364 = v1538;
assign w5365 = w5363 & w5364;
assign w5366 = ~w822 & w4978;
assign w5367 = w3060 & w5366;
assign w5368 = ~w420 & w5367;
assign v1539 = ~(w251 | w379);
assign w5369 = v1539;
assign w5370 = w2560 & w5369;
assign w5371 = w5368 & w5370;
assign w5372 = w700 & w1371;
assign w5373 = w1989 & w5372;
assign w5374 = ~w338 & w1945;
assign w5375 = ~w287 & w2282;
assign w5376 = w5374 & w5375;
assign w5377 = w5373 & w5376;
assign w5378 = w5243 & w5377;
assign w5379 = w5371 & w5378;
assign w5380 = w5365 & w5379;
assign w5381 = w5362 & w5380;
assign w5382 = w5347 & w5381;
assign w5383 = w1093 & w2138;
assign w5384 = w1398 & w3271;
assign w5385 = w1423 & w5384;
assign w5386 = w5383 & w5385;
assign w5387 = ~w214 & w3184;
assign v1540 = ~(w135 | w680);
assign w5388 = v1540;
assign w5389 = w5387 & w5388;
assign w5390 = w5386 & w5389;
assign w5391 = ~w95 & w4655;
assign w5392 = w3427 & w5391;
assign w5393 = w5390 & w5392;
assign w5394 = ~w298 & w1813;
assign w5395 = w707 & w1632;
assign w5396 = w5175 & w5395;
assign w5397 = w3416 & w5396;
assign w5398 = w5394 & w5397;
assign v1541 = ~(w98 | w202);
assign w5399 = v1541;
assign w5400 = w318 & w5399;
assign v1542 = ~(w31 | w184);
assign w5401 = v1542;
assign w5402 = w5237 & w5401;
assign w5403 = w5400 & w5402;
assign w5404 = w1028 & w2912;
assign w5405 = w3061 & w5404;
assign w5406 = w5403 & w5405;
assign v1543 = ~(w125 | w1207);
assign w5407 = v1543;
assign w5408 = w2363 & w5407;
assign w5409 = w1066 & w5408;
assign w5410 = ~w566 & w1239;
assign w5411 = w1200 & w5410;
assign w5412 = w5409 & w5411;
assign w5413 = w5406 & w5412;
assign w5414 = w1853 & w4993;
assign v1544 = ~(w120 | w404);
assign w5415 = v1544;
assign w5416 = w580 & w5415;
assign w5417 = w5414 & w5416;
assign w5418 = w3128 & w5417;
assign w5419 = w5413 & w5418;
assign w5420 = w5398 & w5419;
assign w5421 = ~w300 & w657;
assign w5422 = ~w630 & w5421;
assign v1545 = ~(w271 | w287);
assign w5423 = v1545;
assign w5424 = w1020 & w5423;
assign w5425 = w4503 & w5424;
assign w5426 = w5422 & w5425;
assign w5427 = w348 & w2401;
assign v1546 = ~(w65 | w238);
assign w5428 = v1546;
assign w5429 = ~w209 & w5428;
assign w5430 = w3686 & w5429;
assign v1547 = ~(w70 | w215);
assign w5431 = v1547;
assign w5432 = w304 & w1647;
assign w5433 = w5431 & w5432;
assign w5434 = w5430 & w5433;
assign w5435 = w5427 & w5434;
assign w5436 = w5426 & w5435;
assign w5437 = w3472 & w5436;
assign w5438 = w5420 & w5437;
assign w5439 = w5393 & w5438;
assign w5440 = w5382 & w5439;
assign v1548 = ~(w5382 | w5439);
assign w5441 = v1548;
assign v1549 = ~(w5440 | w5441);
assign w5442 = v1549;
assign w5443 = pi08 & w5442;
assign v1550 = ~(w5440 | w5443);
assign w5444 = v1550;
assign w5445 = w5207 & w5444;
assign v1551 = ~(w5207 | w5444);
assign w5446 = v1551;
assign v1552 = ~(w5445 | w5446);
assign w5447 = v1552;
assign w5448 = w3360 & ~w3362;
assign v1553 = ~(w3363 | w5448);
assign w5449 = v1553;
assign w5450 = w928 & w5449;
assign w5451 = ~w2568 & w3399;
assign w5452 = ~w2492 & w3402;
assign v1554 = ~(w5451 | w5452);
assign w5453 = v1554;
assign w5454 = ~w2424 & w3406;
assign w5455 = w5453 & ~w5454;
assign w5456 = ~w5450 & w5455;
assign w5457 = w5447 & ~w5456;
assign v1555 = ~(w5445 | w5457);
assign w5458 = v1555;
assign w5459 = w5207 & ~w5309;
assign v1556 = ~(w5310 | w5459);
assign w5460 = v1556;
assign w5461 = w5458 & w5460;
assign v1557 = ~(w5310 | w5461);
assign w5462 = v1557;
assign w5463 = w5278 & w5287;
assign v1558 = ~(w5288 | w5463);
assign w5464 = v1558;
assign w5465 = w5462 & w5464;
assign v1559 = ~(w5288 | w5465);
assign w5466 = v1559;
assign w5467 = w5276 & ~w5466;
assign w5468 = ~w5276 & w5466;
assign v1560 = ~(w5467 | w5468);
assign w5469 = v1560;
assign w5470 = w3529 & w4702;
assign w5471 = ~w2089 & w3767;
assign w5472 = ~w1942 & w3760;
assign w5473 = ~w2038 & w3763;
assign v1561 = ~(w5472 | w5473);
assign w5474 = v1561;
assign w5475 = ~w5471 & w5474;
assign w5476 = ~w5470 & w5475;
assign w5477 = pi29 & ~w5476;
assign w5478 = ~pi29 & w5476;
assign v1562 = ~(w5477 | w5478);
assign w5479 = v1562;
assign w5480 = w5469 & w5479;
assign v1563 = ~(w5467 | w5480);
assign w5481 = v1563;
assign w5482 = w5271 & w5273;
assign v1564 = ~(w5274 | w5482);
assign w5483 = v1564;
assign w5484 = ~w5481 & w5483;
assign v1565 = ~(w5274 | w5484);
assign w5485 = v1565;
assign v1566 = ~(w5151 | w5161);
assign w5486 = v1566;
assign v1567 = ~(w5162 | w5486);
assign w5487 = v1567;
assign w5488 = ~w5485 & w5487;
assign v1568 = ~(w5162 | w5488);
assign w5489 = v1568;
assign v1569 = ~(w5061 | w5071);
assign w5490 = v1569;
assign v1570 = ~(w5072 | w5490);
assign w5491 = v1570;
assign w5492 = ~w5489 & w5491;
assign w5493 = w5489 & ~w5491;
assign v1571 = ~(w5492 | w5493);
assign w5494 = v1571;
assign w5495 = w3397 & w4153;
assign w5496 = ~w1387 & w4155;
assign w5497 = ~w1496 & w4158;
assign v1572 = ~(w1609 | w2873);
assign w5498 = v1572;
assign v1573 = ~(w5497 | w5498);
assign w5499 = v1573;
assign w5500 = ~w5496 & w5499;
assign w5501 = ~w5495 & w5500;
assign w5502 = pi26 & ~w5501;
assign w5503 = ~pi26 & w5501;
assign v1574 = ~(w5502 | w5503);
assign w5504 = v1574;
assign w5505 = w5494 & w5504;
assign v1575 = ~(w5492 | w5505);
assign w5506 = v1575;
assign w5507 = w5149 & ~w5506;
assign w5508 = ~w5149 & w5506;
assign v1576 = ~(w5507 | w5508);
assign w5509 = v1576;
assign w5510 = ~w3928 & w4764;
assign w5511 = ~w3587 & w4763;
assign w5512 = ~w3752 & w4836;
assign v1577 = ~(w5511 | w5512);
assign w5513 = v1577;
assign w5514 = ~w3920 & w4913;
assign w5515 = w5513 & ~w5514;
assign w5516 = ~w5510 & w5515;
assign w5517 = pi23 & w5516;
assign v1578 = ~(pi23 | w5516);
assign w5518 = v1578;
assign v1579 = ~(w5517 | w5518);
assign w5519 = v1579;
assign w5520 = w5509 & ~w5519;
assign v1580 = ~(w5507 | w5520);
assign w5521 = v1580;
assign v1581 = ~(w5136 | w5146);
assign w5522 = v1581;
assign v1582 = ~(w5147 | w5522);
assign w5523 = v1582;
assign w5524 = ~w5521 & w5523;
assign v1583 = ~(w5147 | w5524);
assign w5525 = v1583;
assign w5526 = w5134 & ~w5525;
assign w5527 = ~w5134 & w5525;
assign v1584 = ~(w5526 | w5527);
assign w5528 = v1584;
assign w5529 = w4425 & w5114;
assign w5530 = ~w4082 & w5113;
assign w5531 = ~w912 & w915;
assign w5532 = ~w4191 & w5531;
assign v1585 = ~(w5530 | w5532);
assign w5533 = v1585;
assign w5534 = ~w5529 & w5533;
assign w5535 = pi20 & ~w5534;
assign w5536 = ~pi20 & w5534;
assign v1586 = ~(w5535 | w5536);
assign w5537 = v1586;
assign w5538 = w5528 & w5537;
assign v1587 = ~(w5526 | w5538);
assign w5539 = v1587;
assign w5540 = ~w5132 & w5539;
assign w5541 = w5132 & ~w5539;
assign v1588 = ~(w5528 | w5537);
assign w5542 = v1588;
assign v1589 = ~(w5538 | w5542);
assign w5543 = v1589;
assign w5544 = ~w5509 & w5519;
assign v1590 = ~(w5520 | w5544);
assign w5545 = v1590;
assign v1591 = ~(w5494 | w5504);
assign w5546 = v1591;
assign v1592 = ~(w5505 | w5546);
assign w5547 = v1592;
assign w5548 = w5485 & ~w5487;
assign v1593 = ~(w5488 | w5548);
assign w5549 = v1593;
assign w5550 = ~w3510 & w4153;
assign w5551 = ~w1496 & w4155;
assign w5552 = ~w1609 & w4158;
assign v1594 = ~(w1674 | w2873);
assign w5553 = v1594;
assign v1595 = ~(w5552 | w5553);
assign w5554 = v1595;
assign w5555 = ~w5551 & w5554;
assign w5556 = ~w5550 & w5555;
assign w5557 = pi26 & ~w5556;
assign w5558 = ~pi26 & w5556;
assign v1596 = ~(w5557 | w5558);
assign w5559 = v1596;
assign w5560 = w5549 & w5559;
assign w5561 = w5481 & ~w5483;
assign v1597 = ~(w5484 | w5561);
assign w5562 = v1597;
assign w5563 = w3529 & w4854;
assign w5564 = ~w1860 & w3760;
assign w5565 = ~w2038 & w3767;
assign w5566 = ~w1942 & w3763;
assign v1598 = ~(w5565 | w5566);
assign w5567 = v1598;
assign w5568 = ~w5564 & w5567;
assign w5569 = ~w5563 & w5568;
assign w5570 = pi29 & ~w5569;
assign w5571 = ~pi29 & w5569;
assign v1599 = ~(w5570 | w5571);
assign w5572 = v1599;
assign w5573 = w5562 & w5572;
assign v1600 = ~(w5562 | w5572);
assign w5574 = v1600;
assign v1601 = ~(w5573 | w5574);
assign w5575 = v1601;
assign v1602 = ~(w1795 | w2873);
assign w5576 = v1602;
assign w5577 = w3494 & w4153;
assign w5578 = ~w1609 & w4155;
assign w5579 = ~w1674 & w4158;
assign v1603 = ~(w5578 | w5579);
assign w5580 = v1603;
assign w5581 = ~w5577 & w5580;
assign w5582 = ~w5576 & w5581;
assign w5583 = pi26 & w5582;
assign v1604 = ~(pi26 | w5582);
assign w5584 = v1604;
assign v1605 = ~(w5583 | w5584);
assign w5585 = v1605;
assign w5586 = w5575 & ~w5585;
assign v1606 = ~(w5573 | w5586);
assign w5587 = v1606;
assign v1607 = ~(w5549 | w5559);
assign w5588 = v1607;
assign v1608 = ~(w5560 | w5588);
assign w5589 = v1608;
assign w5590 = ~w5587 & w5589;
assign v1609 = ~(w5560 | w5590);
assign w5591 = v1609;
assign w5592 = w5547 & ~w5591;
assign w5593 = ~w5547 & w5591;
assign v1610 = ~(w5592 | w5593);
assign w5594 = v1610;
assign w5595 = w3758 & w4764;
assign w5596 = ~w3587 & w4836;
assign w5597 = ~w3666 & w4763;
assign w5598 = ~w3752 & w4913;
assign v1611 = ~(w5597 | w5598);
assign w5599 = v1611;
assign w5600 = ~w5596 & w5599;
assign w5601 = ~w5595 & w5600;
assign w5602 = pi23 & ~w5601;
assign w5603 = ~pi23 & w5601;
assign v1612 = ~(w5602 | w5603);
assign w5604 = v1612;
assign w5605 = w5594 & w5604;
assign v1613 = ~(w5592 | w5605);
assign w5606 = v1613;
assign w5607 = w5545 & ~w5606;
assign w5608 = ~w5545 & w5606;
assign v1614 = ~(w5607 | w5608);
assign w5609 = v1614;
assign w5610 = w912 & ~w5112;
assign w5611 = ~w4082 & w5610;
assign w5612 = ~w4149 & w5114;
assign w5613 = ~w4134 & w5113;
assign w5614 = ~w4035 & w5531;
assign v1615 = ~(w5613 | w5614);
assign w5615 = v1615;
assign w5616 = ~w5612 & w5615;
assign w5617 = ~w5611 & w5616;
assign w5618 = pi20 & w5617;
assign v1616 = ~(pi20 | w5617);
assign w5619 = v1616;
assign v1617 = ~(w5618 | w5619);
assign w5620 = v1617;
assign w5621 = w5609 & ~w5620;
assign v1618 = ~(w5607 | w5621);
assign w5622 = v1618;
assign w5623 = w4196 & w5114;
assign w5624 = ~w4082 & w5531;
assign w5625 = ~w4191 & w5610;
assign w5626 = ~w4035 & w5113;
assign v1619 = ~(w5625 | w5626);
assign w5627 = v1619;
assign w5628 = ~w5624 & w5627;
assign w5629 = ~w5623 & w5628;
assign w5630 = pi20 & ~w5629;
assign w5631 = ~pi20 & w5629;
assign v1620 = ~(w5630 | w5631);
assign w5632 = v1620;
assign w5633 = ~w5622 & w5632;
assign w5634 = w5521 & ~w5523;
assign v1621 = ~(w5524 | w5634);
assign w5635 = v1621;
assign w5636 = w5622 & ~w5632;
assign v1622 = ~(w5633 | w5636);
assign w5637 = v1622;
assign w5638 = w5635 & w5637;
assign v1623 = ~(w5633 | w5638);
assign w5639 = v1623;
assign w5640 = w5543 & ~w5639;
assign w5641 = ~w5543 & w5639;
assign v1624 = ~(w5640 | w5641);
assign w5642 = v1624;
assign v1625 = ~(w5594 | w5604);
assign w5643 = v1625;
assign v1626 = ~(w5605 | w5643);
assign w5644 = v1626;
assign w5645 = w5587 & ~w5589;
assign v1627 = ~(w5590 | w5645);
assign w5646 = v1627;
assign w5647 = w4291 & w4764;
assign w5648 = ~w3587 & w4913;
assign w5649 = ~w3666 & w4836;
assign v1628 = ~(w5648 | w5649);
assign w5650 = v1628;
assign w5651 = ~w1387 & w4763;
assign w5652 = w5650 & ~w5651;
assign w5653 = ~w5647 & w5652;
assign w5654 = ~pi23 & w5653;
assign w5655 = pi23 & ~w5653;
assign v1629 = ~(w5654 | w5655);
assign w5656 = v1629;
assign w5657 = w5646 & w5656;
assign v1630 = ~(w5646 | w5656);
assign w5658 = v1630;
assign v1631 = ~(w5657 | w5658);
assign w5659 = v1631;
assign w5660 = ~w5575 & w5585;
assign v1632 = ~(w5586 | w5660);
assign w5661 = v1632;
assign v1633 = ~(w5458 | w5460);
assign w5662 = v1633;
assign v1634 = ~(w5461 | w5662);
assign w5663 = v1634;
assign w5664 = w3364 & ~w3366;
assign v1635 = ~(w3367 | w5664);
assign w5665 = v1635;
assign w5666 = w928 & w5665;
assign w5667 = ~w2492 & w3399;
assign w5668 = ~w2424 & w3402;
assign v1636 = ~(w5667 | w5668);
assign w5669 = v1636;
assign w5670 = ~w2339 & w3406;
assign w5671 = w5669 & ~w5670;
assign w5672 = ~w5666 & w5671;
assign v1637 = ~(w5663 | w5672);
assign w5673 = v1637;
assign w5674 = w5663 & w5672;
assign v1638 = ~(w5673 | w5674);
assign w5675 = v1638;
assign w5676 = w3529 & w5033;
assign w5677 = ~w2290 & w3767;
assign w5678 = ~w2089 & w3760;
assign w5679 = ~w2202 & w3763;
assign v1639 = ~(w5678 | w5679);
assign w5680 = v1639;
assign w5681 = ~w5677 & w5680;
assign w5682 = ~w5676 & w5681;
assign w5683 = pi29 & ~w5682;
assign w5684 = ~pi29 & w5682;
assign v1640 = ~(w5683 | w5684);
assign w5685 = v1640;
assign w5686 = w5675 & w5685;
assign v1641 = ~(w5673 | w5686);
assign w5687 = v1641;
assign v1642 = ~(w5462 | w5464);
assign w5688 = v1642;
assign v1643 = ~(w5465 | w5688);
assign w5689 = v1643;
assign w5690 = ~w5687 & w5689;
assign w5691 = w5687 & ~w5689;
assign v1644 = ~(w5690 | w5691);
assign w5692 = v1644;
assign w5693 = ~w2202 & w3767;
assign w5694 = w3529 & w5049;
assign w5695 = ~w2089 & w3763;
assign w5696 = ~w2038 & w3760;
assign v1645 = ~(w5695 | w5696);
assign w5697 = v1645;
assign w5698 = ~w5694 & w5697;
assign w5699 = ~w5693 & w5698;
assign w5700 = pi29 & w5699;
assign v1646 = ~(pi29 | w5699);
assign w5701 = v1646;
assign v1647 = ~(w5700 | w5701);
assign w5702 = v1647;
assign w5703 = w5692 & ~w5702;
assign v1648 = ~(w5690 | w5703);
assign w5704 = v1648;
assign v1649 = ~(w5469 | w5479);
assign w5705 = v1649;
assign v1650 = ~(w5480 | w5705);
assign w5706 = v1650;
assign w5707 = ~w5704 & w5706;
assign w5708 = w5704 & ~w5706;
assign v1651 = ~(w5707 | w5708);
assign w5709 = v1651;
assign w5710 = w4153 & w4520;
assign w5711 = ~w1795 & w4158;
assign w5712 = ~w1674 & w4155;
assign v1652 = ~(w5711 | w5712);
assign w5713 = v1652;
assign v1653 = ~(w1860 | w2873);
assign w5714 = v1653;
assign w5715 = w5713 & ~w5714;
assign w5716 = ~w5710 & w5715;
assign w5717 = ~pi26 & w5716;
assign w5718 = pi26 & ~w5716;
assign v1654 = ~(w5717 | w5718);
assign w5719 = v1654;
assign w5720 = w5709 & w5719;
assign v1655 = ~(w5707 | w5720);
assign w5721 = v1655;
assign w5722 = w5661 & ~w5721;
assign w5723 = ~w5661 & w5721;
assign v1656 = ~(w5722 | w5723);
assign w5724 = v1656;
assign w5725 = w3843 & w4764;
assign w5726 = ~w1387 & w4836;
assign w5727 = ~w1496 & w4763;
assign v1657 = ~(w5726 | w5727);
assign w5728 = v1657;
assign w5729 = ~w3666 & w4913;
assign w5730 = w5728 & ~w5729;
assign w5731 = ~w5725 & w5730;
assign w5732 = ~pi23 & w5731;
assign w5733 = pi23 & ~w5731;
assign v1658 = ~(w5732 | w5733);
assign w5734 = v1658;
assign w5735 = w5724 & w5734;
assign v1659 = ~(w5722 | w5735);
assign w5736 = v1659;
assign w5737 = w5659 & ~w5736;
assign v1660 = ~(w5657 | w5737);
assign w5738 = v1660;
assign w5739 = w5644 & ~w5738;
assign w5740 = ~w5644 & w5738;
assign v1661 = ~(w5739 | w5740);
assign w5741 = v1661;
assign w5742 = w4405 & w5114;
assign w5743 = ~w4035 & w5610;
assign w5744 = ~w4134 & w5531;
assign v1662 = ~(w5743 | w5744);
assign w5745 = v1662;
assign w5746 = ~w3920 & w5113;
assign w5747 = w5745 & ~w5746;
assign w5748 = ~w5742 & w5747;
assign w5749 = ~pi20 & w5748;
assign w5750 = pi20 & ~w5748;
assign v1663 = ~(w5749 | w5750);
assign w5751 = v1663;
assign w5752 = w5741 & w5751;
assign v1664 = ~(w5739 | w5752);
assign w5753 = v1664;
assign v1665 = ~(pi14 | pi15);
assign w5754 = v1665;
assign w5755 = pi14 & pi15;
assign v1666 = ~(w5754 | w5755);
assign w5756 = v1666;
assign v1667 = ~(pi15 | pi16);
assign w5757 = v1667;
assign w5758 = pi15 & pi16;
assign v1668 = ~(w5757 | w5758);
assign w5759 = v1668;
assign v1669 = ~(w5756 | w5759);
assign w5760 = v1669;
assign v1670 = ~(pi16 | pi17);
assign w5761 = v1670;
assign w5762 = pi16 & pi17;
assign v1671 = ~(w5761 | w5762);
assign w5763 = v1671;
assign w5764 = w5760 & w5763;
assign w5765 = w5756 & w5763;
assign w5766 = ~w4422 & w5765;
assign v1672 = ~(w5764 | w5766);
assign w5767 = v1672;
assign v1673 = ~(w4191 | w5767);
assign w5768 = v1673;
assign w5769 = ~pi17 & w5768;
assign w5770 = pi17 & ~w5768;
assign v1674 = ~(w5769 | w5770);
assign w5771 = v1674;
assign v1675 = ~(w5753 | w5771);
assign w5772 = v1675;
assign w5773 = ~w5609 & w5620;
assign v1676 = ~(w5621 | w5773);
assign w5774 = v1676;
assign w5775 = w5753 & w5771;
assign v1677 = ~(w5772 | w5775);
assign w5776 = v1677;
assign w5777 = w5774 & w5776;
assign v1678 = ~(w5772 | w5777);
assign w5778 = v1678;
assign v1679 = ~(w5635 | w5637);
assign w5779 = v1679;
assign v1680 = ~(w5638 | w5779);
assign w5780 = v1680;
assign w5781 = ~w5778 & w5780;
assign w5782 = w5778 & ~w5780;
assign v1681 = ~(w5781 | w5782);
assign w5783 = v1681;
assign v1682 = ~(w5774 | w5776);
assign w5784 = v1682;
assign v1683 = ~(w5777 | w5784);
assign w5785 = v1683;
assign v1684 = ~(w5741 | w5751);
assign w5786 = v1684;
assign v1685 = ~(w5752 | w5786);
assign w5787 = v1685;
assign w5788 = ~w5659 & w5736;
assign v1686 = ~(w5737 | w5788);
assign w5789 = v1686;
assign w5790 = w4309 & w5114;
assign w5791 = ~w3920 & w5531;
assign w5792 = ~w3752 & w5113;
assign w5793 = ~w4134 & w5610;
assign v1687 = ~(w5792 | w5793);
assign w5794 = v1687;
assign w5795 = ~w5791 & w5794;
assign w5796 = ~w5790 & w5795;
assign w5797 = pi20 & ~w5796;
assign w5798 = ~pi20 & w5796;
assign v1688 = ~(w5797 | w5798);
assign w5799 = v1688;
assign w5800 = w5789 & w5799;
assign v1689 = ~(w5724 | w5734);
assign w5801 = v1689;
assign v1690 = ~(w5735 | w5801);
assign w5802 = v1690;
assign v1691 = ~(w5709 | w5719);
assign w5803 = v1691;
assign v1692 = ~(w5720 | w5803);
assign w5804 = v1692;
assign w5805 = ~w5692 & w5702;
assign v1693 = ~(w5703 | w5805);
assign w5806 = v1693;
assign w5807 = w4153 & w4538;
assign w5808 = ~w1795 & w4155;
assign w5809 = ~w1860 & w4158;
assign v1694 = ~(w5808 | w5809);
assign w5810 = v1694;
assign v1695 = ~(w1942 | w2873);
assign w5811 = v1695;
assign w5812 = w5810 & ~w5811;
assign w5813 = ~w5807 & w5812;
assign w5814 = pi26 & w5813;
assign v1696 = ~(pi26 | w5813);
assign w5815 = v1696;
assign v1697 = ~(w5814 | w5815);
assign w5816 = v1697;
assign w5817 = w5806 & ~w5816;
assign w5818 = ~w5447 & w5456;
assign v1698 = ~(w5457 | w5818);
assign w5819 = v1698;
assign v1699 = ~(pi08 | w5442);
assign w5820 = v1699;
assign v1700 = ~(w5443 | w5820);
assign w5821 = v1700;
assign w5822 = w4555 & w5417;
assign w5823 = w5340 & w5822;
assign w5824 = w1654 & w1688;
assign w5825 = w5823 & w5824;
assign w5826 = w96 & ~w427;
assign w5827 = ~w692 & w5826;
assign w5828 = w3778 & w5827;
assign w5829 = w219 & w2363;
assign w5830 = w5828 & w5829;
assign w5831 = ~w674 & w2207;
assign w5832 = w3559 & w4118;
assign w5833 = ~w184 & w476;
assign w5834 = w5832 & w5833;
assign w5835 = w5831 & w5834;
assign w5836 = w5830 & w5835;
assign v1701 = ~(w70 | w727);
assign w5837 = v1701;
assign w5838 = ~w499 & w5837;
assign w5839 = w419 & w1031;
assign w5840 = w1546 & w5839;
assign w5841 = w5838 & w5840;
assign w5842 = w1821 & w3865;
assign v1702 = ~(w267 | w550);
assign w5843 = v1702;
assign w5844 = w5842 & w5843;
assign w5845 = w5841 & w5844;
assign w5846 = w5836 & w5845;
assign w5847 = w1248 & w5846;
assign w5848 = w5825 & w5847;
assign w5849 = ~w5382 & w5848;
assign w5850 = ~w639 & w3650;
assign w5851 = w554 & w5850;
assign v1703 = ~(w302 | w989);
assign w5852 = v1703;
assign w5853 = w2301 & w5852;
assign w5854 = w5851 & w5853;
assign w5855 = w2547 & w5854;
assign w5856 = w1339 & w1935;
assign w5857 = w4982 & w5856;
assign w5858 = w5855 & w5857;
assign w5859 = w1624 & w5858;
assign w5860 = w1048 & w1312;
assign v1704 = ~(w74 | w98);
assign w5861 = v1704;
assign w5862 = ~w338 & w5861;
assign w5863 = ~w410 & w5862;
assign v1705 = ~(w110 | w112);
assign w5864 = v1705;
assign w5865 = w1535 & w5864;
assign w5866 = w5863 & w5865;
assign w5867 = w5860 & w5866;
assign w5868 = w5859 & w5867;
assign w5869 = w4360 & w4650;
assign w5870 = w5868 & w5869;
assign v1706 = ~(pi02 | w5870);
assign w5871 = v1706;
assign w5872 = pi02 & w5870;
assign v1707 = ~(w5871 | w5872);
assign w5873 = v1707;
assign w5874 = ~pi05 & w5873;
assign v1708 = ~(w5871 | w5874);
assign w5875 = v1708;
assign w5876 = w5382 & ~w5875;
assign w5877 = ~w5382 & w5875;
assign v1709 = ~(w5876 | w5877);
assign w5878 = v1709;
assign w5879 = w3348 & ~w3350;
assign v1710 = ~(w3351 | w5879);
assign w5880 = v1710;
assign w5881 = w928 & w5880;
assign w5882 = ~w2724 & w3399;
assign w5883 = ~w2596 & w3406;
assign v1711 = ~(w5882 | w5883);
assign w5884 = v1711;
assign w5885 = ~w2669 & w3402;
assign w5886 = w5884 & ~w5885;
assign w5887 = ~w5881 & w5886;
assign w5888 = w5878 & ~w5887;
assign v1712 = ~(w5876 | w5888);
assign w5889 = v1712;
assign w5890 = w5382 & ~w5848;
assign v1713 = ~(w5849 | w5890);
assign w5891 = v1713;
assign w5892 = w5889 & w5891;
assign v1714 = ~(w5849 | w5892);
assign w5893 = v1714;
assign w5894 = ~w5821 & w5893;
assign w5895 = w5821 & ~w5893;
assign v1715 = ~(w5894 | w5895);
assign w5896 = v1715;
assign w5897 = w3356 & ~w3358;
assign v1716 = ~(w3359 | w5897);
assign w5898 = v1716;
assign w5899 = w928 & w5898;
assign w5900 = ~w2568 & w3402;
assign w5901 = ~w2492 & w3406;
assign v1717 = ~(w5900 | w5901);
assign w5902 = v1717;
assign w5903 = ~w2596 & w3399;
assign w5904 = w5902 & ~w5903;
assign w5905 = ~w5899 & w5904;
assign w5906 = w5896 & ~w5905;
assign v1718 = ~(w5894 | w5906);
assign w5907 = v1718;
assign w5908 = w5819 & ~w5907;
assign w5909 = ~w5819 & w5907;
assign v1719 = ~(w5908 | w5909);
assign w5910 = v1719;
assign w5911 = w3529 & w5262;
assign w5912 = ~w2202 & w3760;
assign w5913 = ~w2339 & w3767;
assign w5914 = ~w2290 & w3763;
assign v1720 = ~(w5913 | w5914);
assign w5915 = v1720;
assign w5916 = ~w5912 & w5915;
assign w5917 = ~w5911 & w5916;
assign w5918 = pi29 & ~w5917;
assign w5919 = ~pi29 & w5917;
assign v1721 = ~(w5918 | w5919);
assign w5920 = v1721;
assign w5921 = w5910 & w5920;
assign v1722 = ~(w5908 | w5921);
assign w5922 = v1722;
assign v1723 = ~(w5675 | w5685);
assign w5923 = v1723;
assign v1724 = ~(w5686 | w5923);
assign w5924 = v1724;
assign w5925 = ~w5922 & w5924;
assign w5926 = w5922 & ~w5924;
assign v1725 = ~(w5925 | w5926);
assign w5927 = v1725;
assign v1726 = ~(w2038 | w2873);
assign w5928 = v1726;
assign w5929 = w4153 & w4854;
assign w5930 = ~w1942 & w4158;
assign w5931 = ~w1860 & w4155;
assign v1727 = ~(w5930 | w5931);
assign w5932 = v1727;
assign w5933 = ~w5929 & w5932;
assign w5934 = ~w5928 & w5933;
assign w5935 = pi26 & w5934;
assign v1728 = ~(pi26 | w5934);
assign w5936 = v1728;
assign v1729 = ~(w5935 | w5936);
assign w5937 = v1729;
assign w5938 = w5927 & ~w5937;
assign v1730 = ~(w5925 | w5938);
assign w5939 = v1730;
assign w5940 = ~w5806 & w5816;
assign v1731 = ~(w5817 | w5940);
assign w5941 = v1731;
assign w5942 = ~w5939 & w5941;
assign v1732 = ~(w5817 | w5942);
assign w5943 = v1732;
assign w5944 = w5804 & ~w5943;
assign w5945 = ~w5804 & w5943;
assign v1733 = ~(w5944 | w5945);
assign w5946 = v1733;
assign w5947 = w3397 & w4764;
assign w5948 = ~w1387 & w4913;
assign w5949 = ~w1609 & w4763;
assign w5950 = ~w1496 & w4836;
assign v1734 = ~(w5949 | w5950);
assign w5951 = v1734;
assign w5952 = ~w5948 & w5951;
assign w5953 = ~w5947 & w5952;
assign w5954 = pi23 & ~w5953;
assign w5955 = ~pi23 & w5953;
assign v1735 = ~(w5954 | w5955);
assign w5956 = v1735;
assign w5957 = w5946 & w5956;
assign v1736 = ~(w5944 | w5957);
assign w5958 = v1736;
assign w5959 = w5802 & ~w5958;
assign w5960 = ~w5802 & w5958;
assign v1737 = ~(w5959 | w5960);
assign w5961 = v1737;
assign w5962 = ~w3928 & w5114;
assign w5963 = ~w3920 & w5610;
assign w5964 = ~w3752 & w5531;
assign v1738 = ~(w5963 | w5964);
assign w5965 = v1738;
assign w5966 = ~w3587 & w5113;
assign w5967 = w5965 & ~w5966;
assign w5968 = ~w5962 & w5967;
assign w5969 = pi20 & ~w5968;
assign w5970 = ~pi20 & w5968;
assign v1739 = ~(w5969 | w5970);
assign w5971 = v1739;
assign w5972 = w5961 & w5971;
assign v1740 = ~(w5959 | w5972);
assign w5973 = v1740;
assign v1741 = ~(w5789 | w5799);
assign w5974 = v1741;
assign v1742 = ~(w5800 | w5974);
assign w5975 = v1742;
assign w5976 = ~w5973 & w5975;
assign v1743 = ~(w5800 | w5976);
assign w5977 = v1743;
assign w5978 = w5787 & ~w5977;
assign w5979 = ~w5787 & w5977;
assign v1744 = ~(w5978 | w5979);
assign w5980 = v1744;
assign w5981 = w4425 & w5765;
assign w5982 = ~w4082 & w5764;
assign w5983 = ~w5756 & w5759;
assign w5984 = ~w4191 & w5983;
assign v1745 = ~(w5982 | w5984);
assign w5985 = v1745;
assign w5986 = ~w5981 & w5985;
assign w5987 = pi17 & ~w5986;
assign w5988 = ~pi17 & w5986;
assign v1746 = ~(w5987 | w5988);
assign w5989 = v1746;
assign w5990 = w5980 & w5989;
assign v1747 = ~(w5978 | w5990);
assign w5991 = v1747;
assign w5992 = ~w5785 & w5991;
assign w5993 = w5785 & ~w5991;
assign v1748 = ~(w5980 | w5989);
assign w5994 = v1748;
assign v1749 = ~(w5990 | w5994);
assign w5995 = v1749;
assign v1750 = ~(w5961 | w5971);
assign w5996 = v1750;
assign v1751 = ~(w5972 | w5996);
assign w5997 = v1751;
assign v1752 = ~(w5946 | w5956);
assign w5998 = v1752;
assign v1753 = ~(w5957 | w5998);
assign w5999 = v1753;
assign w6000 = w5939 & ~w5941;
assign v1754 = ~(w5942 | w6000);
assign w6001 = v1754;
assign w6002 = ~w3510 & w4764;
assign w6003 = ~w1496 & w4913;
assign w6004 = ~w1609 & w4836;
assign v1755 = ~(w6003 | w6004);
assign w6005 = v1755;
assign w6006 = ~w1674 & w4763;
assign w6007 = w6005 & ~w6006;
assign w6008 = ~w6002 & w6007;
assign w6009 = ~pi23 & w6008;
assign w6010 = pi23 & ~w6008;
assign v1756 = ~(w6009 | w6010);
assign w6011 = v1756;
assign w6012 = w6001 & w6011;
assign w6013 = ~w5927 & w5937;
assign v1757 = ~(w5938 | w6013);
assign w6014 = v1757;
assign w6015 = ~w5896 & w5905;
assign v1758 = ~(w5906 | w6015);
assign w6016 = v1758;
assign w6017 = ~w2290 & w3760;
assign w6018 = w3529 & w5280;
assign w6019 = ~w2339 & w3763;
assign w6020 = ~w2424 & w3767;
assign v1759 = ~(w6019 | w6020);
assign w6021 = v1759;
assign w6022 = ~w6018 & w6021;
assign w6023 = ~w6017 & w6022;
assign w6024 = pi29 & w6023;
assign v1760 = ~(pi29 | w6023);
assign w6025 = v1760;
assign v1761 = ~(w6024 | w6025);
assign w6026 = v1761;
assign w6027 = w6016 & ~w6026;
assign v1762 = ~(w5889 | w5891);
assign w6028 = v1762;
assign v1763 = ~(w5892 | w6028);
assign w6029 = v1763;
assign w6030 = w3352 & ~w3354;
assign v1764 = ~(w3355 | w6030);
assign w6031 = v1764;
assign w6032 = w928 & w6031;
assign w6033 = ~w2568 & w3406;
assign w6034 = ~w2596 & w3402;
assign v1765 = ~(w6033 | w6034);
assign w6035 = v1765;
assign w6036 = ~w2669 & w3399;
assign w6037 = w6035 & ~w6036;
assign w6038 = ~w6032 & w6037;
assign v1766 = ~(w6029 | w6038);
assign w6039 = v1766;
assign w6040 = ~w5878 & w5887;
assign v1767 = ~(w5888 | w6040);
assign w6041 = v1767;
assign w6042 = pi05 & ~w5873;
assign v1768 = ~(w5874 | w6042);
assign w6043 = v1768;
assign v1769 = ~(w892 | w1207);
assign w6044 = v1769;
assign w6045 = ~w208 & w1988;
assign w6046 = w6044 & w6045;
assign w6047 = w502 & w6046;
assign v1770 = ~(w245 | w635);
assign w6048 = v1770;
assign w6049 = ~w200 & w6048;
assign w6050 = w3231 & w6049;
assign w6051 = w829 & w3598;
assign w6052 = w6050 & w6051;
assign w6053 = w4371 & w6052;
assign w6054 = w1921 & w4596;
assign w6055 = w6053 & w6054;
assign w6056 = w6047 & w6055;
assign w6057 = w5213 & w5292;
assign w6058 = w3065 & w6057;
assign w6059 = w589 & ~w699;
assign w6060 = w3556 & w6059;
assign w6061 = w2796 & w6060;
assign w6062 = w6058 & w6061;
assign w6063 = w6056 & w6062;
assign w6064 = pi02 & ~w6063;
assign w6065 = ~pi02 & w6063;
assign v1771 = ~(w6064 | w6065);
assign w6066 = v1771;
assign w6067 = w1374 & w1458;
assign w6068 = w589 & w3475;
assign w6069 = w1142 & w6068;
assign w6070 = w6067 & w6069;
assign w6071 = w1482 & w4382;
assign v1772 = ~(w184 | w563);
assign w6072 = v1772;
assign w6073 = w2299 & w6072;
assign w6074 = w1340 & w2995;
assign w6075 = ~w410 & w6074;
assign w6076 = w138 & w6075;
assign w6077 = w6073 & w6076;
assign w6078 = ~w232 & w1613;
assign w6079 = w3453 & w6078;
assign w6080 = ~w98 & w6079;
assign w6081 = w6077 & w6080;
assign w6082 = w6071 & w6081;
assign w6083 = w748 & w6082;
assign w6084 = w6070 & w6083;
assign w6085 = pi02 & ~w6084;
assign w6086 = ~pi02 & w6084;
assign w6087 = w1921 & w5290;
assign w6088 = w1580 & w6087;
assign v1773 = ~(w253 | w454);
assign w6089 = v1773;
assign w6090 = ~w63 & w6089;
assign w6091 = ~w251 & w2498;
assign w6092 = w1878 & w6091;
assign w6093 = w6090 & w6092;
assign w6094 = w693 & w2349;
assign w6095 = w3691 & w6094;
assign w6096 = ~w134 & w6095;
assign w6097 = w6093 & w6096;
assign w6098 = w6088 & w6097;
assign w6099 = w5368 & w6098;
assign w6100 = w1490 & w6099;
assign v1774 = ~(w21 | w493);
assign w6101 = v1774;
assign w6102 = w336 & w6101;
assign v1775 = ~(w231 | w1134);
assign w6103 = v1775;
assign w6104 = w4371 & w6103;
assign w6105 = w6102 & w6104;
assign w6106 = w2877 & w6105;
assign v1776 = ~(w281 | w370);
assign w6107 = v1776;
assign w6108 = ~w390 & w6107;
assign v1777 = ~(w605 | w978);
assign w6109 = v1777;
assign w6110 = ~w73 & w6109;
assign w6111 = w6108 & w6110;
assign w6112 = w133 & w6111;
assign w6113 = w6106 & w6112;
assign w6114 = w3308 & w6113;
assign v1778 = ~(w119 | w263);
assign w6115 = v1778;
assign w6116 = w3043 & w6115;
assign v1779 = ~(w65 | w140);
assign w6117 = v1779;
assign w6118 = w2348 & w6117;
assign w6119 = w1902 & w6118;
assign w6120 = w6116 & w6119;
assign w6121 = w3267 & w4974;
assign w6122 = w6120 & w6121;
assign w6123 = w6114 & w6122;
assign w6124 = w3323 & w6123;
assign w6125 = w2154 & w6124;
assign w6126 = w6100 & w6125;
assign w6127 = pi02 & ~w6126;
assign w6128 = ~pi02 & w6126;
assign w6129 = (~w3341 & w29463) | (~w3341 & w29464) | (w29463 & w29464);
assign v1780 = ~(w3342 | w6129);
assign w6130 = v1780;
assign w6131 = w928 & w6130;
assign w6132 = ~w3000 & w3399;
assign w6133 = ~w2846 & w3406;
assign w6134 = ~w2937 & w3402;
assign v1781 = ~(w6133 | w6134);
assign w6135 = v1781;
assign w6136 = ~w6132 & w6135;
assign w6137 = ~w6131 & w6136;
assign v1782 = ~(w6128 | w6137);
assign w6138 = v1782;
assign v1783 = ~(w6127 | w6138);
assign w6139 = v1783;
assign v1784 = ~(w6086 | w6139);
assign w6140 = v1784;
assign v1785 = ~(w6085 | w6140);
assign w6141 = v1785;
assign w6142 = w6066 & ~w6141;
assign v1786 = ~(w6064 | w6142);
assign w6143 = v1786;
assign w6144 = w6043 & ~w6143;
assign w6145 = ~w6043 & w6143;
assign v1787 = ~(w6144 | w6145);
assign w6146 = v1787;
assign v1788 = ~(w2727 | w3346);
assign w6147 = v1788;
assign v1789 = ~(w3347 | w6147);
assign w6148 = v1789;
assign w6149 = w928 & w6148;
assign w6150 = ~w2724 & w3402;
assign w6151 = ~w2811 & w3399;
assign v1790 = ~(w6150 | w6151);
assign w6152 = v1790;
assign w6153 = ~w2669 & w3406;
assign w6154 = w6152 & ~w6153;
assign w6155 = ~w6149 & w6154;
assign w6156 = w6146 & ~w6155;
assign v1791 = ~(w6144 | w6156);
assign w6157 = v1791;
assign w6158 = w6041 & ~w6157;
assign w6159 = ~w6041 & w6157;
assign v1792 = ~(w6158 | w6159);
assign w6160 = v1792;
assign w6161 = w3529 & w5449;
assign w6162 = ~w2568 & w3767;
assign w6163 = ~w2492 & w3763;
assign w6164 = ~w2424 & w3760;
assign v1793 = ~(w6163 | w6164);
assign w6165 = v1793;
assign w6166 = ~w6162 & w6165;
assign w6167 = ~w6161 & w6166;
assign w6168 = pi29 & ~w6167;
assign w6169 = ~pi29 & w6167;
assign v1794 = ~(w6168 | w6169);
assign w6170 = v1794;
assign w6171 = w6160 & w6170;
assign v1795 = ~(w6158 | w6171);
assign w6172 = v1795;
assign w6173 = w6029 & w6038;
assign v1796 = ~(w6039 | w6173);
assign w6174 = v1796;
assign w6175 = ~w6172 & w6174;
assign v1797 = ~(w6039 | w6175);
assign w6176 = v1797;
assign w6177 = ~w6016 & w6026;
assign v1798 = ~(w6027 | w6177);
assign w6178 = v1798;
assign w6179 = ~w6176 & w6178;
assign v1799 = ~(w6027 | w6179);
assign w6180 = v1799;
assign v1800 = ~(w5910 | w5920);
assign w6181 = v1800;
assign v1801 = ~(w5921 | w6181);
assign w6182 = v1801;
assign w6183 = ~w6180 & w6182;
assign w6184 = w6180 & ~w6182;
assign v1802 = ~(w6183 | w6184);
assign w6185 = v1802;
assign w6186 = w4153 & w4702;
assign v1803 = ~(w2089 | w2873);
assign w6187 = v1803;
assign w6188 = ~w1942 & w4155;
assign w6189 = ~w2038 & w4158;
assign v1804 = ~(w6188 | w6189);
assign w6190 = v1804;
assign w6191 = ~w6187 & w6190;
assign w6192 = ~w6186 & w6191;
assign w6193 = pi26 & ~w6192;
assign w6194 = ~pi26 & w6192;
assign v1805 = ~(w6193 | w6194);
assign w6195 = v1805;
assign w6196 = w6185 & w6195;
assign v1806 = ~(w6183 | w6196);
assign w6197 = v1806;
assign w6198 = w6014 & ~w6197;
assign w6199 = ~w6014 & w6197;
assign v1807 = ~(w6198 | w6199);
assign w6200 = v1807;
assign w6201 = ~w1795 & w4763;
assign w6202 = w3494 & w4764;
assign w6203 = ~w1609 & w4913;
assign w6204 = ~w1674 & w4836;
assign v1808 = ~(w6203 | w6204);
assign w6205 = v1808;
assign w6206 = ~w6202 & w6205;
assign w6207 = ~w6201 & w6206;
assign w6208 = pi23 & w6207;
assign v1809 = ~(pi23 | w6207);
assign w6209 = v1809;
assign v1810 = ~(w6208 | w6209);
assign w6210 = v1810;
assign w6211 = w6200 & ~w6210;
assign v1811 = ~(w6198 | w6211);
assign w6212 = v1811;
assign v1812 = ~(w6001 | w6011);
assign w6213 = v1812;
assign v1813 = ~(w6012 | w6213);
assign w6214 = v1813;
assign w6215 = ~w6212 & w6214;
assign v1814 = ~(w6012 | w6215);
assign w6216 = v1814;
assign w6217 = w5999 & ~w6216;
assign w6218 = ~w5999 & w6216;
assign v1815 = ~(w6217 | w6218);
assign w6219 = v1815;
assign w6220 = w3758 & w5114;
assign w6221 = ~w3752 & w5610;
assign w6222 = ~w3587 & w5531;
assign v1816 = ~(w6221 | w6222);
assign w6223 = v1816;
assign w6224 = ~w3666 & w5113;
assign w6225 = w6223 & ~w6224;
assign w6226 = ~w6220 & w6225;
assign w6227 = ~pi20 & w6226;
assign w6228 = pi20 & ~w6226;
assign v1817 = ~(w6227 | w6228);
assign w6229 = v1817;
assign w6230 = w6219 & w6229;
assign v1818 = ~(w6217 | w6230);
assign w6231 = v1818;
assign w6232 = w5997 & ~w6231;
assign w6233 = ~w5997 & w6231;
assign v1819 = ~(w6232 | w6233);
assign w6234 = v1819;
assign w6235 = ~w4149 & w5765;
assign w6236 = w5756 & ~w5763;
assign w6237 = ~w4082 & w6236;
assign w6238 = ~w4134 & w5764;
assign w6239 = ~w4035 & w5983;
assign v1820 = ~(w6238 | w6239);
assign w6240 = v1820;
assign w6241 = ~w6237 & w6240;
assign w6242 = ~w6235 & w6241;
assign w6243 = pi17 & ~w6242;
assign w6244 = ~pi17 & w6242;
assign v1821 = ~(w6243 | w6244);
assign w6245 = v1821;
assign w6246 = w6234 & w6245;
assign v1822 = ~(w6232 | w6246);
assign w6247 = v1822;
assign w6248 = w4196 & w5765;
assign w6249 = ~w4082 & w5983;
assign w6250 = ~w4191 & w6236;
assign w6251 = ~w4035 & w5764;
assign v1823 = ~(w6250 | w6251);
assign w6252 = v1823;
assign w6253 = ~w6249 & w6252;
assign w6254 = ~w6248 & w6253;
assign w6255 = pi17 & ~w6254;
assign w6256 = ~pi17 & w6254;
assign v1824 = ~(w6255 | w6256);
assign w6257 = v1824;
assign w6258 = ~w6247 & w6257;
assign w6259 = w5973 & ~w5975;
assign v1825 = ~(w5976 | w6259);
assign w6260 = v1825;
assign w6261 = w6247 & ~w6257;
assign v1826 = ~(w6258 | w6261);
assign w6262 = v1826;
assign w6263 = w6260 & w6262;
assign v1827 = ~(w6258 | w6263);
assign w6264 = v1827;
assign w6265 = w5995 & ~w6264;
assign v1828 = ~(w6219 | w6229);
assign w6266 = v1828;
assign v1829 = ~(w6230 | w6266);
assign w6267 = v1829;
assign w6268 = w6212 & ~w6214;
assign v1830 = ~(w6215 | w6268);
assign w6269 = v1830;
assign w6270 = w4291 & w5114;
assign w6271 = ~w3587 & w5610;
assign w6272 = ~w3666 & w5531;
assign v1831 = ~(w6271 | w6272);
assign w6273 = v1831;
assign w6274 = ~w1387 & w5113;
assign w6275 = w6273 & ~w6274;
assign w6276 = ~w6270 & w6275;
assign w6277 = ~pi20 & w6276;
assign w6278 = pi20 & ~w6276;
assign v1832 = ~(w6277 | w6278);
assign w6279 = v1832;
assign w6280 = w6269 & w6279;
assign w6281 = ~w6200 & w6210;
assign v1833 = ~(w6211 | w6281);
assign w6282 = v1833;
assign v1834 = ~(w6185 | w6195);
assign w6283 = v1834;
assign v1835 = ~(w6196 | w6283);
assign w6284 = v1835;
assign w6285 = w6176 & ~w6178;
assign v1836 = ~(w6179 | w6285);
assign w6286 = v1836;
assign w6287 = w4153 & w5049;
assign v1837 = ~(w2202 | w2873);
assign w6288 = v1837;
assign w6289 = ~w2089 & w4158;
assign w6290 = ~w2038 & w4155;
assign v1838 = ~(w6289 | w6290);
assign w6291 = v1838;
assign w6292 = ~w6288 & w6291;
assign w6293 = ~w6287 & w6292;
assign w6294 = pi26 & ~w6293;
assign w6295 = ~pi26 & w6293;
assign v1839 = ~(w6294 | w6295);
assign w6296 = v1839;
assign w6297 = w6286 & w6296;
assign w6298 = w6172 & ~w6174;
assign v1840 = ~(w6175 | w6298);
assign w6299 = v1840;
assign w6300 = w3529 & w5665;
assign w6301 = ~w2492 & w3767;
assign w6302 = ~w2424 & w3763;
assign w6303 = ~w2339 & w3760;
assign v1841 = ~(w6302 | w6303);
assign w6304 = v1841;
assign w6305 = ~w6301 & w6304;
assign w6306 = ~w6300 & w6305;
assign w6307 = pi29 & ~w6306;
assign w6308 = ~pi29 & w6306;
assign v1842 = ~(w6307 | w6308);
assign w6309 = v1842;
assign w6310 = w6299 & w6309;
assign v1843 = ~(w6299 | w6309);
assign w6311 = v1843;
assign v1844 = ~(w6310 | w6311);
assign w6312 = v1844;
assign v1845 = ~(w2290 | w2873);
assign w6313 = v1845;
assign w6314 = w4153 & w5033;
assign w6315 = ~w2089 & w4155;
assign w6316 = ~w2202 & w4158;
assign v1846 = ~(w6315 | w6316);
assign w6317 = v1846;
assign w6318 = ~w6314 & w6317;
assign w6319 = ~w6313 & w6318;
assign w6320 = pi26 & w6319;
assign v1847 = ~(pi26 | w6319);
assign w6321 = v1847;
assign v1848 = ~(w6320 | w6321);
assign w6322 = v1848;
assign w6323 = w6312 & ~w6322;
assign v1849 = ~(w6310 | w6323);
assign w6324 = v1849;
assign v1850 = ~(w6286 | w6296);
assign w6325 = v1850;
assign v1851 = ~(w6297 | w6325);
assign w6326 = v1851;
assign w6327 = ~w6324 & w6326;
assign v1852 = ~(w6297 | w6327);
assign w6328 = v1852;
assign w6329 = w6284 & ~w6328;
assign w6330 = ~w6284 & w6328;
assign v1853 = ~(w6329 | w6330);
assign w6331 = v1853;
assign w6332 = w4520 & w4764;
assign w6333 = ~w1795 & w4836;
assign w6334 = ~w1860 & w4763;
assign w6335 = ~w1674 & w4913;
assign v1854 = ~(w6334 | w6335);
assign w6336 = v1854;
assign w6337 = ~w6333 & w6336;
assign w6338 = ~w6332 & w6337;
assign w6339 = pi23 & ~w6338;
assign w6340 = ~pi23 & w6338;
assign v1855 = ~(w6339 | w6340);
assign w6341 = v1855;
assign w6342 = w6331 & w6341;
assign v1856 = ~(w6329 | w6342);
assign w6343 = v1856;
assign w6344 = w6282 & ~w6343;
assign w6345 = ~w6282 & w6343;
assign v1857 = ~(w6344 | w6345);
assign w6346 = v1857;
assign w6347 = w3843 & w5114;
assign w6348 = ~w1387 & w5531;
assign w6349 = ~w1496 & w5113;
assign v1858 = ~(w6348 | w6349);
assign w6350 = v1858;
assign w6351 = ~w3666 & w5610;
assign w6352 = w6350 & ~w6351;
assign w6353 = ~w6347 & w6352;
assign w6354 = ~pi20 & w6353;
assign w6355 = pi20 & ~w6353;
assign v1859 = ~(w6354 | w6355);
assign w6356 = v1859;
assign w6357 = w6346 & w6356;
assign v1860 = ~(w6344 | w6357);
assign w6358 = v1860;
assign v1861 = ~(w6269 | w6279);
assign w6359 = v1861;
assign v1862 = ~(w6280 | w6359);
assign w6360 = v1862;
assign w6361 = ~w6358 & w6360;
assign v1863 = ~(w6280 | w6361);
assign w6362 = v1863;
assign w6363 = w6267 & ~w6362;
assign w6364 = ~w6267 & w6362;
assign v1864 = ~(w6363 | w6364);
assign w6365 = v1864;
assign w6366 = w4405 & w5765;
assign w6367 = ~w4035 & w6236;
assign w6368 = ~w4134 & w5983;
assign v1865 = ~(w6367 | w6368);
assign w6369 = v1865;
assign w6370 = ~w3920 & w5764;
assign w6371 = w6369 & ~w6370;
assign w6372 = ~w6366 & w6371;
assign w6373 = pi17 & w6372;
assign v1866 = ~(pi17 | w6372);
assign w6374 = v1866;
assign v1867 = ~(w6373 | w6374);
assign w6375 = v1867;
assign w6376 = w6365 & ~w6375;
assign v1868 = ~(w6363 | w6376);
assign w6377 = v1868;
assign w6378 = ~pi13 & pi14;
assign w6379 = pi13 & ~pi14;
assign v1869 = ~(w6378 | w6379);
assign w6380 = v1869;
assign v1870 = ~(pi11 | pi12);
assign w6381 = v1870;
assign w6382 = pi11 & pi12;
assign v1871 = ~(w6381 | w6382);
assign w6383 = v1871;
assign v1872 = ~(pi12 | pi13);
assign w6384 = v1872;
assign w6385 = pi12 & pi13;
assign v1873 = ~(w6384 | w6385);
assign w6386 = v1873;
assign v1874 = ~(w6383 | w6386);
assign w6387 = v1874;
assign w6388 = ~w6380 & w6387;
assign w6389 = ~w6380 & w6383;
assign w6390 = ~w4422 & w6389;
assign v1875 = ~(w6388 | w6390);
assign w6391 = v1875;
assign v1876 = ~(w4191 | w6391);
assign w6392 = v1876;
assign w6393 = ~pi14 & w6392;
assign w6394 = pi14 & ~w6392;
assign v1877 = ~(w6393 | w6394);
assign w6395 = v1877;
assign v1878 = ~(w6377 | w6395);
assign w6396 = v1878;
assign v1879 = ~(w6234 | w6245);
assign w6397 = v1879;
assign v1880 = ~(w6246 | w6397);
assign w6398 = v1880;
assign w6399 = w6377 & w6395;
assign v1881 = ~(w6396 | w6399);
assign w6400 = v1881;
assign w6401 = w6398 & w6400;
assign v1882 = ~(w6396 | w6401);
assign w6402 = v1882;
assign v1883 = ~(w6260 | w6262);
assign w6403 = v1883;
assign v1884 = ~(w6263 | w6403);
assign w6404 = v1884;
assign w6405 = ~w6402 & w6404;
assign w6406 = w6402 & ~w6404;
assign v1885 = ~(w6405 | w6406);
assign w6407 = v1885;
assign v1886 = ~(w6398 | w6400);
assign w6408 = v1886;
assign v1887 = ~(w6401 | w6408);
assign w6409 = v1887;
assign w6410 = w6358 & ~w6360;
assign v1888 = ~(w6361 | w6410);
assign w6411 = v1888;
assign w6412 = w4309 & w5765;
assign w6413 = ~w3920 & w5983;
assign w6414 = ~w3752 & w5764;
assign w6415 = ~w4134 & w6236;
assign v1889 = ~(w6414 | w6415);
assign w6416 = v1889;
assign w6417 = ~w6413 & w6416;
assign w6418 = ~w6412 & w6417;
assign w6419 = pi17 & ~w6418;
assign w6420 = ~pi17 & w6418;
assign v1890 = ~(w6419 | w6420);
assign w6421 = v1890;
assign w6422 = w6411 & w6421;
assign v1891 = ~(w6346 | w6356);
assign w6423 = v1891;
assign v1892 = ~(w6357 | w6423);
assign w6424 = v1892;
assign v1893 = ~(w6331 | w6341);
assign w6425 = v1893;
assign v1894 = ~(w6342 | w6425);
assign w6426 = v1894;
assign w6427 = w6324 & ~w6326;
assign v1895 = ~(w6327 | w6427);
assign w6428 = v1895;
assign w6429 = w4538 & w4764;
assign w6430 = ~w1795 & w4913;
assign w6431 = ~w1942 & w4763;
assign w6432 = ~w1860 & w4836;
assign v1896 = ~(w6431 | w6432);
assign w6433 = v1896;
assign w6434 = ~w6430 & w6433;
assign w6435 = ~w6429 & w6434;
assign w6436 = pi23 & ~w6435;
assign w6437 = ~pi23 & w6435;
assign v1897 = ~(w6436 | w6437);
assign w6438 = v1897;
assign w6439 = w6428 & w6438;
assign w6440 = ~w6312 & w6322;
assign v1898 = ~(w6323 | w6440);
assign w6441 = v1898;
assign w6442 = ~w6146 & w6155;
assign v1899 = ~(w6156 | w6442);
assign w6443 = v1899;
assign w6444 = ~w6066 & w6141;
assign v1900 = ~(w6142 | w6444);
assign w6445 = v1900;
assign w6446 = ~w2814 & w3344;
assign v1901 = ~(w3345 | w6446);
assign w6447 = v1901;
assign w6448 = w928 & ~w6447;
assign w6449 = ~w2811 & w3402;
assign w6450 = ~w2724 & w3406;
assign v1902 = ~(w6449 | w6450);
assign w6451 = v1902;
assign w6452 = ~w2846 & w3399;
assign w6453 = w6451 & ~w6452;
assign w6454 = ~w6448 & w6453;
assign w6455 = w6445 & ~w6454;
assign v1903 = ~(w2847 | w2848);
assign w6456 = v1903;
assign w6457 = w3343 & ~w6456;
assign w6458 = ~w3343 & w6456;
assign v1904 = ~(w6457 | w6458);
assign w6459 = v1904;
assign w6460 = w928 & w6459;
assign w6461 = ~w2937 & w3399;
assign w6462 = ~w2811 & w3406;
assign v1905 = ~(w6461 | w6462);
assign w6463 = v1905;
assign w6464 = ~w2846 & w3402;
assign w6465 = w6463 & ~w6464;
assign w6466 = ~w6460 & w6465;
assign v1906 = ~(w6085 | w6086);
assign w6467 = v1906;
assign w6468 = w6139 & ~w6467;
assign w6469 = ~w6139 & w6467;
assign v1907 = ~(w6468 | w6469);
assign w6470 = v1907;
assign w6471 = ~w6466 & w6470;
assign w6472 = w1814 & w2107;
assign w6473 = w2296 & w6472;
assign w6474 = w148 & w6473;
assign w6475 = ~w158 & w1165;
assign w6476 = w717 & w6475;
assign w6477 = w1189 & w6072;
assign v1908 = ~(w51 | w387);
assign w6478 = v1908;
assign w6479 = ~w298 & w6478;
assign w6480 = w6477 & w6479;
assign w6481 = w1379 & w6480;
assign w6482 = w6476 & w6481;
assign w6483 = w2551 & w6482;
assign w6484 = w6474 & w6483;
assign w6485 = ~w160 & w5363;
assign w6486 = w1301 & w6485;
assign w6487 = ~w456 & w1340;
assign w6488 = w4341 & w6487;
assign w6489 = w240 & w2188;
assign w6490 = w6488 & w6489;
assign w6491 = w6486 & w6490;
assign w6492 = w4673 & w6491;
assign w6493 = w6484 & w6492;
assign v1909 = ~(w186 | w274);
assign w6494 = v1909;
assign w6495 = w3650 & w6494;
assign w6496 = w1641 & w6495;
assign w6497 = w2452 & w3149;
assign w6498 = w562 & w6497;
assign w6499 = w6496 & w6498;
assign w6500 = w4639 & w6499;
assign w6501 = w6493 & w6500;
assign v1910 = ~(w3001 | w3002);
assign w6502 = v1910;
assign w6503 = ~w3341 & w6502;
assign w6504 = w3341 & ~w6502;
assign v1911 = ~(w6503 | w6504);
assign w6505 = v1911;
assign w6506 = w928 & ~w6505;
assign w6507 = ~w2937 & w3406;
assign w6508 = ~w3000 & w3402;
assign w6509 = ~w3068 & w3399;
assign v1912 = ~(w6508 | w6509);
assign w6510 = v1912;
assign w6511 = ~w6507 & w6510;
assign w6512 = ~w6506 & w6511;
assign v1913 = ~(w6501 | w6512);
assign w6513 = v1913;
assign w6514 = w852 & w2082;
assign w6515 = w2398 & w6514;
assign w6516 = w361 & w6515;
assign v1914 = ~(w216 | w311);
assign w6517 = v1914;
assign w6518 = w6516 & w6517;
assign w6519 = w5215 & w6518;
assign v1915 = ~(w151 | w999);
assign w6520 = v1915;
assign v1916 = ~(w184 | w584);
assign w6521 = v1916;
assign w6522 = w1991 & w6521;
assign w6523 = w1603 & w6522;
assign w6524 = w6520 & w6523;
assign w6525 = w1284 & w6524;
assign w6526 = w2465 & w3620;
assign w6527 = w339 & w2443;
assign w6528 = w3706 & w6527;
assign w6529 = w6526 & w6528;
assign w6530 = w883 & w6529;
assign w6531 = w6525 & w6530;
assign w6532 = w6519 & w6531;
assign w6533 = w2009 & w5171;
assign v1917 = ~(w451 | w699);
assign w6534 = v1917;
assign w6535 = w2540 & w6534;
assign w6536 = w1903 & w2214;
assign w6537 = w6535 & w6536;
assign w6538 = w4490 & w6537;
assign w6539 = ~w277 & w1287;
assign w6540 = w4578 & w6539;
assign v1918 = ~(w49 | w211);
assign w6541 = v1918;
assign w6542 = ~w463 & w6541;
assign w6543 = w6540 & w6542;
assign w6544 = w6538 & w6543;
assign w6545 = w6533 & w6544;
assign w6546 = w1403 & w6545;
assign w6547 = w6532 & w6546;
assign v1919 = ~(w3069 | w3070);
assign w6548 = v1919;
assign w6549 = (~w3339 & w28476) | (~w3339 & w28477) | (w28476 & w28477);
assign w6550 = (w3339 & w28478) | (w3339 & w28479) | (w28478 & w28479);
assign v1920 = ~(w6549 | w6550);
assign w6551 = v1920;
assign w6552 = w928 & ~w6551;
assign w6553 = ~w3068 & w3402;
assign w6554 = ~w3000 & w3406;
assign w6555 = ~w3124 & w3399;
assign v1921 = ~(w6554 | w6555);
assign w6556 = v1921;
assign w6557 = ~w6553 & w6556;
assign w6558 = ~w6552 & w6557;
assign v1922 = ~(w6547 | w6558);
assign w6559 = v1922;
assign w6560 = w1073 & w2738;
assign v1923 = ~(w410 | w499);
assign w6561 = v1923;
assign w6562 = ~w431 & w1465;
assign w6563 = w6561 & w6562;
assign w6564 = ~w200 & w1423;
assign w6565 = w6563 & w6564;
assign w6566 = w6560 & w6565;
assign w6567 = w3885 & w6566;
assign w6568 = ~w428 & w984;
assign w6569 = w5369 & w6568;
assign w6570 = w2959 & w6569;
assign w6571 = w6567 & w6570;
assign w6572 = w5335 & w6571;
assign v1924 = ~(w78 | w497);
assign w6573 = v1924;
assign w6574 = w2411 & w6573;
assign w6575 = w1536 & w3083;
assign w6576 = w6574 & w6575;
assign w6577 = w1110 & w6576;
assign w6578 = w2207 & w5297;
assign w6579 = w6577 & w6578;
assign w6580 = w2517 & w3158;
assign w6581 = ~w224 & w6580;
assign w6582 = ~w68 & w6581;
assign w6583 = ~w448 & w1722;
assign w6584 = w2380 & w6583;
assign w6585 = ~w172 & w580;
assign w6586 = w3008 & w6585;
assign w6587 = w6584 & w6586;
assign w6588 = w6582 & w6587;
assign w6589 = w6579 & w6588;
assign v1925 = ~(w286 | w488);
assign w6590 = v1925;
assign w6591 = w554 & ~w588;
assign w6592 = w6590 & w6591;
assign v1926 = ~(w258 | w307);
assign w6593 = v1926;
assign w6594 = ~w282 & w6593;
assign w6595 = ~w145 & w6594;
assign w6596 = w6592 & w6595;
assign w6597 = w6589 & w6596;
assign w6598 = w2095 & w6597;
assign w6599 = w6572 & w6598;
assign v1927 = ~(w3163 | w3335);
assign w6600 = v1927;
assign v1928 = ~(w3127 | w3336);
assign w6601 = v1928;
assign w6602 = ~w6600 & w6601;
assign v1929 = ~(w3340 | w6602);
assign w6603 = v1929;
assign w6604 = ~w3068 & w3406;
assign w6605 = ~w3162 & w3399;
assign w6606 = ~w3124 & w3402;
assign v1930 = ~(w6605 | w6606);
assign w6607 = v1930;
assign w6608 = ~w6604 & w6607;
assign w6609 = (w6603 & w31256) | (w6603 & w31257) | (w31256 & w31257);
assign w6610 = ~w238 & w375;
assign v1931 = ~(w212 | w441);
assign w6611 = v1931;
assign w6612 = w3474 & w6611;
assign w6613 = w6610 & w6612;
assign w6614 = w222 & w1660;
assign w6615 = w762 & w2319;
assign w6616 = w6614 & w6615;
assign w6617 = w1485 & w6616;
assign w6618 = w6613 & w6617;
assign w6619 = w133 & w783;
assign w6620 = w2369 & w6619;
assign v1932 = ~(w215 | w418);
assign w6621 = v1932;
assign w6622 = w2024 & w6621;
assign w6623 = w1754 & w6622;
assign w6624 = w6620 & w6623;
assign v1933 = ~(w108 | w997);
assign w6625 = v1933;
assign w6626 = w1613 & w6625;
assign w6627 = ~w53 & w2476;
assign w6628 = w6626 & w6627;
assign w6629 = w901 & w990;
assign w6630 = w6628 & w6629;
assign w6631 = w6624 & w6630;
assign w6632 = ~w125 & w965;
assign w6633 = w439 & w2952;
assign w6634 = w6632 & w6633;
assign w6635 = w650 & w6634;
assign w6636 = w4212 & w6635;
assign w6637 = w6631 & w6636;
assign w6638 = w6618 & w6637;
assign w6639 = w2883 & w6638;
assign v1934 = ~(w3335 | w3337);
assign w6640 = v1934;
assign v1935 = ~(w3338 | w6640);
assign w6641 = v1935;
assign w6642 = ~w3124 & w3406;
assign w6643 = ~w3211 & w3399;
assign w6644 = ~w3162 & w3402;
assign v1936 = ~(w6643 | w6644);
assign w6645 = v1936;
assign w6646 = (~w6641 & w31159) | (~w6641 & w31160) | (w31159 & w31160);
assign w6647 = w893 & w1542;
assign w6648 = ~w870 & w6647;
assign w6649 = w823 & w6648;
assign w6650 = ~w331 & w3813;
assign w6651 = ~w221 & w6650;
assign w6652 = w1287 & w3805;
assign w6653 = w6651 & w6652;
assign w6654 = ~w639 & w6561;
assign w6655 = w6653 & w6654;
assign w6656 = w6649 & w6655;
assign v1937 = ~(w267 | w899);
assign w6657 = v1937;
assign v1938 = ~(w241 | w298);
assign w6658 = v1938;
assign w6659 = w6657 & w6658;
assign w6660 = ~w388 & w6659;
assign v1939 = ~(w150 | w558);
assign w6661 = v1939;
assign w6662 = ~w165 & w6661;
assign w6663 = w1475 & w6662;
assign w6664 = w6660 & w6663;
assign w6665 = w1177 & w1738;
assign w6666 = w1811 & w6665;
assign w6667 = w1360 & w6666;
assign w6668 = w6664 & w6667;
assign w6669 = w2808 & w6668;
assign w6670 = w4229 & w4501;
assign w6671 = w6669 & w6670;
assign w6672 = w6656 & w6671;
assign w6673 = ~w3262 & w3332;
assign w6674 = w3211 & ~w6673;
assign w6675 = ~w3211 & w6673;
assign v1940 = ~(w6674 | w6675);
assign w6676 = v1940;
assign w6677 = (w3399 & ~w3331) | (w3399 & w31161) | (~w3331 & w31161);
assign w6678 = (w3406 & ~w3210) | (w3406 & w31000) | (~w3210 & w31000);
assign w6679 = (w3402 & ~w3261) | (w3402 & w31001) | (~w3261 & w31001);
assign v1941 = ~(w6678 | w6679);
assign w6680 = v1941;
assign w6681 = (~w6676 & w30787) | (~w6676 & w30788) | (w30787 & w30788);
assign w6682 = (w6676 & w31002) | (w6676 & w31003) | (w31002 & w31003);
assign w6683 = ~w530 & w3557;
assign w6684 = ~w1134 & w6683;
assign w6685 = w2434 & w6684;
assign w6686 = ~w888 & w2797;
assign w6687 = w1087 & w3060;
assign w6688 = w998 & w6687;
assign w6689 = w6686 & w6688;
assign w6690 = w6685 & w6689;
assign v1942 = ~(w337 | w753);
assign w6691 = v1942;
assign w6692 = w3658 & w6691;
assign v1943 = ~(w331 | w666);
assign w6693 = v1943;
assign w6694 = w1042 & w6693;
assign w6695 = w6692 & w6694;
assign w6696 = w210 & w2413;
assign w6697 = w6695 & w6696;
assign v1944 = ~(w176 | w211);
assign w6698 = v1944;
assign w6699 = w1689 & w6698;
assign w6700 = w990 & w6699;
assign v1945 = ~(w239 | w680);
assign w6701 = v1945;
assign v1946 = ~(w78 | w370);
assign w6702 = v1946;
assign w6703 = w6701 & w6702;
assign w6704 = w6700 & w6703;
assign w6705 = w6697 & w6704;
assign w6706 = w6690 & w6705;
assign w6707 = ~w697 & w1214;
assign w6708 = w2924 & w6707;
assign w6709 = w2061 & w6708;
assign v1947 = ~(w278 | w316);
assign w6710 = v1947;
assign v1948 = ~(w31 | w329);
assign w6711 = v1948;
assign w6712 = w6710 & w6711;
assign w6713 = w6709 & w6712;
assign w6714 = ~w457 & w960;
assign v1949 = ~(w70 | w288);
assign w6715 = v1949;
assign w6716 = w1475 & w6715;
assign w6717 = w6714 & w6716;
assign w6718 = ~w201 & w1840;
assign w6719 = ~w183 & w6718;
assign w6720 = w6717 & w6719;
assign w6721 = w2396 & w6720;
assign w6722 = w6713 & w6721;
assign v1950 = ~(w388 | w484);
assign w6723 = v1950;
assign w6724 = w3202 & w6723;
assign w6725 = w3188 & w6724;
assign w6726 = w6722 & w6725;
assign w6727 = w2227 & w6726;
assign w6728 = w6706 & w6727;
assign w6729 = (w6676 & w31258) | (w6676 & w31259) | (w31258 & w31259);
assign w6730 = (~w6676 & w31260) | (~w6676 & w31261) | (w31260 & w31261);
assign v1951 = ~(w6729 | w6730);
assign w6731 = v1951;
assign v1952 = ~(w3263 | w3333);
assign w6732 = v1952;
assign w6733 = w6674 & ~w6732;
assign w6734 = ~w6674 & w6732;
assign v1953 = ~(w6733 | w6734);
assign w6735 = v1953;
assign w6736 = ~w3162 & w3406;
assign w6737 = ~w3262 & w3399;
assign w6738 = ~w3211 & w3402;
assign v1954 = ~(w6737 | w6738);
assign w6739 = v1954;
assign w6740 = (~w6735 & w31162) | (~w6735 & w31163) | (w31162 & w31163);
assign w6741 = w6731 & ~w6740;
assign w6742 = (~w6729 & ~w6731) | (~w6729 & w31164) | (~w6731 & w31164);
assign w6743 = (w6641 & w31165) | (w6641 & w31166) | (w31165 & w31166);
assign v1955 = ~(w6646 | w6743);
assign w6744 = v1955;
assign w6745 = ~w6742 & w6744;
assign v1956 = ~(w6646 | w6745);
assign w6746 = v1956;
assign w6747 = (~w6603 & w31262) | (~w6603 & w31263) | (w31262 & w31263);
assign v1957 = ~(w6609 | w6747);
assign w6748 = v1957;
assign w6749 = ~w6746 & w6748;
assign w6750 = (~w6609 & w6746) | (~w6609 & w31264) | (w6746 & w31264);
assign w6751 = w6547 & w6558;
assign v1958 = ~(w6559 | w6751);
assign w6752 = v1958;
assign w6753 = ~w6750 & w6752;
assign v1959 = ~(w6559 | w6753);
assign w6754 = v1959;
assign w6755 = w6501 & w6512;
assign v1960 = ~(w6513 | w6755);
assign w6756 = v1960;
assign w6757 = ~w6754 & w6756;
assign v1961 = ~(w6513 | w6757);
assign w6758 = v1961;
assign v1962 = ~(w6127 | w6128);
assign w6759 = v1962;
assign w6760 = w6137 & w6759;
assign v1963 = ~(w6137 | w6759);
assign w6761 = v1963;
assign v1964 = ~(w6760 | w6761);
assign w6762 = v1964;
assign v1965 = ~(w6758 | w6762);
assign w6763 = v1965;
assign w6764 = w6758 & w6762;
assign v1966 = ~(w6763 | w6764);
assign w6765 = v1966;
assign w6766 = w3529 & w6148;
assign w6767 = ~w2811 & w3767;
assign w6768 = ~w2724 & w3763;
assign v1967 = ~(w6767 | w6768);
assign w6769 = v1967;
assign w6770 = ~w2669 & w3760;
assign w6771 = w6769 & ~w6770;
assign w6772 = ~w6766 & w6771;
assign w6773 = pi29 & w6772;
assign v1968 = ~(pi29 | w6772);
assign w6774 = v1968;
assign v1969 = ~(w6773 | w6774);
assign w6775 = v1969;
assign w6776 = w6765 & ~w6775;
assign v1970 = ~(w6763 | w6776);
assign w6777 = v1970;
assign w6778 = w6466 & ~w6470;
assign v1971 = ~(w6471 | w6778);
assign w6779 = v1971;
assign w6780 = ~w6777 & w6779;
assign v1972 = ~(w6471 | w6780);
assign w6781 = v1972;
assign w6782 = ~w6445 & w6454;
assign v1973 = ~(w6455 | w6782);
assign w6783 = v1973;
assign w6784 = ~w6781 & w6783;
assign v1974 = ~(w6455 | w6784);
assign w6785 = v1974;
assign w6786 = w6443 & ~w6785;
assign w6787 = ~w6443 & w6785;
assign v1975 = ~(w6786 | w6787);
assign w6788 = v1975;
assign w6789 = w3529 & w5898;
assign w6790 = ~w2568 & w3763;
assign w6791 = ~w2596 & w3767;
assign w6792 = ~w2492 & w3760;
assign v1976 = ~(w6791 | w6792);
assign w6793 = v1976;
assign w6794 = ~w6790 & w6793;
assign w6795 = ~w6789 & w6794;
assign w6796 = pi29 & ~w6795;
assign w6797 = ~pi29 & w6795;
assign v1977 = ~(w6796 | w6797);
assign w6798 = v1977;
assign w6799 = w6788 & w6798;
assign v1978 = ~(w6786 | w6799);
assign w6800 = v1978;
assign v1979 = ~(w6160 | w6170);
assign w6801 = v1979;
assign v1980 = ~(w6171 | w6801);
assign w6802 = v1980;
assign w6803 = ~w6800 & w6802;
assign w6804 = w6800 & ~w6802;
assign v1981 = ~(w6803 | w6804);
assign w6805 = v1981;
assign w6806 = w4153 & w5262;
assign w6807 = ~w2202 & w4155;
assign v1982 = ~(w2339 | w2873);
assign w6808 = v1982;
assign w6809 = ~w2290 & w4158;
assign v1983 = ~(w6808 | w6809);
assign w6810 = v1983;
assign w6811 = ~w6807 & w6810;
assign w6812 = ~w6806 & w6811;
assign w6813 = pi26 & ~w6812;
assign w6814 = ~pi26 & w6812;
assign v1984 = ~(w6813 | w6814);
assign w6815 = v1984;
assign w6816 = w6805 & w6815;
assign v1985 = ~(w6803 | w6816);
assign w6817 = v1985;
assign w6818 = w6441 & ~w6817;
assign w6819 = ~w6441 & w6817;
assign v1986 = ~(w6818 | w6819);
assign w6820 = v1986;
assign w6821 = w4764 & w4854;
assign w6822 = ~w1860 & w4913;
assign w6823 = ~w2038 & w4763;
assign w6824 = ~w1942 & w4836;
assign v1987 = ~(w6823 | w6824);
assign w6825 = v1987;
assign w6826 = ~w6822 & w6825;
assign w6827 = ~w6821 & w6826;
assign w6828 = pi23 & ~w6827;
assign w6829 = ~pi23 & w6827;
assign v1988 = ~(w6828 | w6829);
assign w6830 = v1988;
assign w6831 = w6820 & w6830;
assign v1989 = ~(w6818 | w6831);
assign w6832 = v1989;
assign v1990 = ~(w6428 | w6438);
assign w6833 = v1990;
assign v1991 = ~(w6439 | w6833);
assign w6834 = v1991;
assign w6835 = ~w6832 & w6834;
assign v1992 = ~(w6439 | w6835);
assign w6836 = v1992;
assign w6837 = w6426 & ~w6836;
assign w6838 = ~w6426 & w6836;
assign v1993 = ~(w6837 | w6838);
assign w6839 = v1993;
assign w6840 = w3397 & w5114;
assign w6841 = ~w1496 & w5531;
assign w6842 = ~w1609 & w5113;
assign w6843 = ~w1387 & w5610;
assign v1994 = ~(w6842 | w6843);
assign w6844 = v1994;
assign w6845 = ~w6841 & w6844;
assign w6846 = ~w6840 & w6845;
assign w6847 = pi20 & ~w6846;
assign w6848 = ~pi20 & w6846;
assign v1995 = ~(w6847 | w6848);
assign w6849 = v1995;
assign w6850 = w6839 & w6849;
assign v1996 = ~(w6837 | w6850);
assign w6851 = v1996;
assign w6852 = w6424 & ~w6851;
assign w6853 = ~w6424 & w6851;
assign v1997 = ~(w6852 | w6853);
assign w6854 = v1997;
assign w6855 = ~w3928 & w5765;
assign w6856 = ~w3752 & w5983;
assign w6857 = ~w3587 & w5764;
assign v1998 = ~(w6856 | w6857);
assign w6858 = v1998;
assign w6859 = ~w3920 & w6236;
assign w6860 = w6858 & ~w6859;
assign w6861 = ~w6855 & w6860;
assign w6862 = ~pi17 & w6861;
assign w6863 = pi17 & ~w6861;
assign v1999 = ~(w6862 | w6863);
assign w6864 = v1999;
assign w6865 = w6854 & w6864;
assign v2000 = ~(w6852 | w6865);
assign w6866 = v2000;
assign v2001 = ~(w6411 | w6421);
assign w6867 = v2001;
assign v2002 = ~(w6422 | w6867);
assign w6868 = v2002;
assign w6869 = ~w6866 & w6868;
assign v2003 = ~(w6422 | w6869);
assign w6870 = v2003;
assign w6871 = ~w6383 & w6386;
assign w6872 = ~w4191 & w6871;
assign w6873 = w4425 & w6389;
assign w6874 = ~w4082 & w6388;
assign v2004 = ~(w6873 | w6874);
assign w6875 = v2004;
assign w6876 = ~w6872 & w6875;
assign w6877 = pi14 & w6876;
assign v2005 = ~(pi14 | w6876);
assign w6878 = v2005;
assign v2006 = ~(w6877 | w6878);
assign w6879 = v2006;
assign v2007 = ~(w6870 | w6879);
assign w6880 = v2007;
assign w6881 = ~w6365 & w6375;
assign v2008 = ~(w6376 | w6881);
assign w6882 = v2008;
assign w6883 = w6870 & w6879;
assign v2009 = ~(w6880 | w6883);
assign w6884 = v2009;
assign w6885 = w6882 & w6884;
assign v2010 = ~(w6880 | w6885);
assign w6886 = v2010;
assign w6887 = ~w6409 & w6886;
assign v2011 = ~(w6854 | w6864);
assign w6888 = v2011;
assign v2012 = ~(w6865 | w6888);
assign w6889 = v2012;
assign v2013 = ~(w6839 | w6849);
assign w6890 = v2013;
assign v2014 = ~(w6850 | w6890);
assign w6891 = v2014;
assign w6892 = w6832 & ~w6834;
assign v2015 = ~(w6835 | w6892);
assign w6893 = v2015;
assign w6894 = ~w3510 & w5114;
assign w6895 = ~w1609 & w5531;
assign w6896 = ~w1674 & w5113;
assign w6897 = ~w1496 & w5610;
assign v2016 = ~(w6896 | w6897);
assign w6898 = v2016;
assign w6899 = ~w6895 & w6898;
assign w6900 = ~w6894 & w6899;
assign w6901 = pi20 & ~w6900;
assign w6902 = ~pi20 & w6900;
assign v2017 = ~(w6901 | w6902);
assign w6903 = v2017;
assign w6904 = w6893 & w6903;
assign v2018 = ~(w6820 | w6830);
assign w6905 = v2018;
assign v2019 = ~(w6831 | w6905);
assign w6906 = v2019;
assign v2020 = ~(w6805 | w6815);
assign w6907 = v2020;
assign v2021 = ~(w6816 | w6907);
assign w6908 = v2021;
assign v2022 = ~(w6788 | w6798);
assign w6909 = v2022;
assign v2023 = ~(w6799 | w6909);
assign w6910 = v2023;
assign w6911 = w4153 & w5280;
assign w6912 = ~w2290 & w4155;
assign w6913 = ~w2339 & w4158;
assign v2024 = ~(w2424 | w2873);
assign w6914 = v2024;
assign v2025 = ~(w6913 | w6914);
assign w6915 = v2025;
assign w6916 = ~w6912 & w6915;
assign w6917 = ~w6911 & w6916;
assign w6918 = pi26 & ~w6917;
assign w6919 = ~pi26 & w6917;
assign v2026 = ~(w6918 | w6919);
assign w6920 = v2026;
assign w6921 = w6910 & w6920;
assign w6922 = w6781 & ~w6783;
assign v2027 = ~(w6784 | w6922);
assign w6923 = v2027;
assign w6924 = w3529 & w6031;
assign w6925 = ~w2568 & w3760;
assign w6926 = ~w2596 & w3763;
assign w6927 = ~w2669 & w3767;
assign v2028 = ~(w6926 | w6927);
assign w6928 = v2028;
assign w6929 = ~w6925 & w6928;
assign w6930 = ~w6924 & w6929;
assign w6931 = pi29 & ~w6930;
assign w6932 = ~pi29 & w6930;
assign v2029 = ~(w6931 | w6932);
assign w6933 = v2029;
assign w6934 = w6923 & w6933;
assign w6935 = w4153 & w5665;
assign v2030 = ~(w2492 | w2873);
assign w6936 = v2030;
assign w6937 = ~w2424 & w4158;
assign w6938 = ~w2339 & w4155;
assign v2031 = ~(w6937 | w6938);
assign w6939 = v2031;
assign w6940 = ~w6936 & w6939;
assign w6941 = ~w6935 & w6940;
assign w6942 = pi26 & ~w6941;
assign w6943 = ~pi26 & w6941;
assign v2032 = ~(w6942 | w6943);
assign w6944 = v2032;
assign v2033 = ~(w6923 | w6933);
assign w6945 = v2033;
assign v2034 = ~(w6934 | w6945);
assign w6946 = v2034;
assign w6947 = w6944 & w6946;
assign v2035 = ~(w6934 | w6947);
assign w6948 = v2035;
assign v2036 = ~(w6910 | w6920);
assign w6949 = v2036;
assign v2037 = ~(w6921 | w6949);
assign w6950 = v2037;
assign w6951 = ~w6948 & w6950;
assign v2038 = ~(w6921 | w6951);
assign w6952 = v2038;
assign w6953 = w6908 & ~w6952;
assign w6954 = ~w6908 & w6952;
assign v2039 = ~(w6953 | w6954);
assign w6955 = v2039;
assign w6956 = w4702 & w4764;
assign w6957 = ~w2089 & w4763;
assign w6958 = ~w1942 & w4913;
assign w6959 = ~w2038 & w4836;
assign v2040 = ~(w6958 | w6959);
assign w6960 = v2040;
assign w6961 = ~w6957 & w6960;
assign w6962 = ~w6956 & w6961;
assign w6963 = pi23 & ~w6962;
assign w6964 = ~pi23 & w6962;
assign v2041 = ~(w6963 | w6964);
assign w6965 = v2041;
assign w6966 = w6955 & w6965;
assign v2042 = ~(w6953 | w6966);
assign w6967 = v2042;
assign w6968 = w6906 & ~w6967;
assign w6969 = ~w6906 & w6967;
assign v2043 = ~(w6968 | w6969);
assign w6970 = v2043;
assign w6971 = w3494 & w5114;
assign w6972 = ~w1609 & w5610;
assign w6973 = ~w1674 & w5531;
assign v2044 = ~(w6972 | w6973);
assign w6974 = v2044;
assign w6975 = ~w1795 & w5113;
assign w6976 = w6974 & ~w6975;
assign w6977 = ~w6971 & w6976;
assign w6978 = pi20 & ~w6977;
assign w6979 = ~pi20 & w6977;
assign v2045 = ~(w6978 | w6979);
assign w6980 = v2045;
assign w6981 = w6970 & w6980;
assign v2046 = ~(w6968 | w6981);
assign w6982 = v2046;
assign v2047 = ~(w6893 | w6903);
assign w6983 = v2047;
assign v2048 = ~(w6904 | w6983);
assign w6984 = v2048;
assign w6985 = ~w6982 & w6984;
assign v2049 = ~(w6904 | w6985);
assign w6986 = v2049;
assign w6987 = w6891 & ~w6986;
assign w6988 = ~w6891 & w6986;
assign v2050 = ~(w6987 | w6988);
assign w6989 = v2050;
assign w6990 = w3758 & w5765;
assign w6991 = ~w3587 & w5983;
assign w6992 = ~w3666 & w5764;
assign v2051 = ~(w6991 | w6992);
assign w6993 = v2051;
assign w6994 = ~w3752 & w6236;
assign w6995 = w6993 & ~w6994;
assign w6996 = ~w6990 & w6995;
assign w6997 = pi17 & w6996;
assign v2052 = ~(pi17 | w6996);
assign w6998 = v2052;
assign v2053 = ~(w6997 | w6998);
assign w6999 = v2053;
assign w7000 = w6989 & ~w6999;
assign v2054 = ~(w6987 | w7000);
assign w7001 = v2054;
assign w7002 = w6889 & ~w7001;
assign w7003 = ~w4149 & w6389;
assign w7004 = w6380 & w6383;
assign w7005 = ~w4082 & w7004;
assign w7006 = ~w4134 & w6388;
assign w7007 = ~w4035 & w6871;
assign v2055 = ~(w7006 | w7007);
assign w7008 = v2055;
assign w7009 = ~w7005 & w7008;
assign w7010 = ~w7003 & w7009;
assign w7011 = pi14 & ~w7010;
assign w7012 = ~pi14 & w7010;
assign v2056 = ~(w7011 | w7012);
assign w7013 = v2056;
assign w7014 = ~w6889 & w7001;
assign v2057 = ~(w7002 | w7014);
assign w7015 = v2057;
assign w7016 = w7013 & w7015;
assign v2058 = ~(w7002 | w7016);
assign w7017 = v2058;
assign w7018 = w4196 & w6389;
assign w7019 = ~w4082 & w6871;
assign w7020 = ~w4191 & w7004;
assign w7021 = ~w4035 & w6388;
assign v2059 = ~(w7020 | w7021);
assign w7022 = v2059;
assign w7023 = ~w7019 & w7022;
assign w7024 = ~w7018 & w7023;
assign w7025 = pi14 & ~w7024;
assign w7026 = ~pi14 & w7024;
assign v2060 = ~(w7025 | w7026);
assign w7027 = v2060;
assign w7028 = ~w7017 & w7027;
assign w7029 = w6866 & ~w6868;
assign v2061 = ~(w6869 | w7029);
assign w7030 = v2061;
assign w7031 = w7017 & ~w7027;
assign v2062 = ~(w7028 | w7031);
assign w7032 = v2062;
assign w7033 = w7030 & w7032;
assign v2063 = ~(w7028 | w7033);
assign w7034 = v2063;
assign v2064 = ~(w6882 | w6884);
assign w7035 = v2064;
assign v2065 = ~(w6885 | w7035);
assign w7036 = v2065;
assign w7037 = ~w7034 & w7036;
assign w7038 = ~w6989 & w6999;
assign v2066 = ~(w7000 | w7038);
assign w7039 = v2066;
assign w7040 = w6982 & ~w6984;
assign v2067 = ~(w6985 | w7040);
assign w7041 = v2067;
assign w7042 = w4291 & w5765;
assign w7043 = ~w3587 & w6236;
assign w7044 = ~w3666 & w5983;
assign v2068 = ~(w7043 | w7044);
assign w7045 = v2068;
assign w7046 = ~w1387 & w5764;
assign w7047 = w7045 & ~w7046;
assign w7048 = ~w7042 & w7047;
assign w7049 = ~pi17 & w7048;
assign w7050 = pi17 & ~w7048;
assign v2069 = ~(w7049 | w7050);
assign w7051 = v2069;
assign w7052 = w7041 & w7051;
assign v2070 = ~(w7041 | w7051);
assign w7053 = v2070;
assign v2071 = ~(w7052 | w7053);
assign w7054 = v2071;
assign v2072 = ~(w6970 | w6980);
assign w7055 = v2072;
assign v2073 = ~(w6981 | w7055);
assign w7056 = v2073;
assign v2074 = ~(w6955 | w6965);
assign w7057 = v2074;
assign v2075 = ~(w6966 | w7057);
assign w7058 = v2075;
assign w7059 = w6948 & ~w6950;
assign v2076 = ~(w6951 | w7059);
assign w7060 = v2076;
assign w7061 = w4764 & w5049;
assign w7062 = ~w2202 & w4763;
assign w7063 = ~w2038 & w4913;
assign w7064 = ~w2089 & w4836;
assign v2077 = ~(w7063 | w7064);
assign w7065 = v2077;
assign w7066 = ~w7062 & w7065;
assign w7067 = ~w7061 & w7066;
assign w7068 = pi23 & ~w7067;
assign w7069 = ~pi23 & w7067;
assign v2078 = ~(w7068 | w7069);
assign w7070 = v2078;
assign w7071 = w7060 & w7070;
assign v2079 = ~(w6944 | w6946);
assign w7072 = v2079;
assign v2080 = ~(w6947 | w7072);
assign w7073 = v2080;
assign w7074 = w6777 & ~w6779;
assign v2081 = ~(w6780 | w7074);
assign w7075 = v2081;
assign w7076 = w3529 & w5880;
assign w7077 = ~w2669 & w3763;
assign w7078 = ~w2596 & w3760;
assign v2082 = ~(w7077 | w7078);
assign w7079 = v2082;
assign w7080 = ~w2724 & w3767;
assign w7081 = w7079 & ~w7080;
assign w7082 = ~w7076 & w7081;
assign w7083 = ~pi29 & w7082;
assign w7084 = pi29 & ~w7082;
assign v2083 = ~(w7083 | w7084);
assign w7085 = v2083;
assign w7086 = w7075 & w7085;
assign v2084 = ~(w7075 | w7085);
assign w7087 = v2084;
assign v2085 = ~(w7086 | w7087);
assign w7088 = v2085;
assign v2086 = ~(w2568 | w2873);
assign w7089 = v2086;
assign w7090 = w4153 & w5449;
assign w7091 = ~w2492 & w4158;
assign w7092 = ~w2424 & w4155;
assign v2087 = ~(w7091 | w7092);
assign w7093 = v2087;
assign w7094 = ~w7090 & w7093;
assign w7095 = ~w7089 & w7094;
assign w7096 = pi26 & w7095;
assign v2088 = ~(pi26 | w7095);
assign w7097 = v2088;
assign v2089 = ~(w7096 | w7097);
assign w7098 = v2089;
assign w7099 = w7088 & ~w7098;
assign v2090 = ~(w7086 | w7099);
assign w7100 = v2090;
assign w7101 = w7073 & ~w7100;
assign w7102 = ~w7073 & w7100;
assign v2091 = ~(w7101 | w7102);
assign w7103 = v2091;
assign w7104 = w4764 & w5033;
assign w7105 = ~w2202 & w4836;
assign w7106 = ~w2089 & w4913;
assign w7107 = ~w2290 & w4763;
assign v2092 = ~(w7106 | w7107);
assign w7108 = v2092;
assign w7109 = ~w7105 & w7108;
assign w7110 = ~w7104 & w7109;
assign w7111 = pi23 & ~w7110;
assign w7112 = ~pi23 & w7110;
assign v2093 = ~(w7111 | w7112);
assign w7113 = v2093;
assign w7114 = w7103 & w7113;
assign v2094 = ~(w7101 | w7114);
assign w7115 = v2094;
assign v2095 = ~(w7060 | w7070);
assign w7116 = v2095;
assign v2096 = ~(w7071 | w7116);
assign w7117 = v2096;
assign w7118 = ~w7115 & w7117;
assign v2097 = ~(w7071 | w7118);
assign w7119 = v2097;
assign w7120 = w7058 & ~w7119;
assign w7121 = ~w7058 & w7119;
assign v2098 = ~(w7120 | w7121);
assign w7122 = v2098;
assign w7123 = w4520 & w5114;
assign w7124 = ~w1795 & w5531;
assign w7125 = ~w1674 & w5610;
assign w7126 = ~w1860 & w5113;
assign v2099 = ~(w7125 | w7126);
assign w7127 = v2099;
assign w7128 = ~w7124 & w7127;
assign w7129 = ~w7123 & w7128;
assign w7130 = pi20 & ~w7129;
assign w7131 = ~pi20 & w7129;
assign v2100 = ~(w7130 | w7131);
assign w7132 = v2100;
assign w7133 = w7122 & w7132;
assign v2101 = ~(w7120 | w7133);
assign w7134 = v2101;
assign w7135 = w7056 & ~w7134;
assign w7136 = ~w7056 & w7134;
assign v2102 = ~(w7135 | w7136);
assign w7137 = v2102;
assign w7138 = w3843 & w5765;
assign w7139 = ~w1387 & w5983;
assign w7140 = ~w1496 & w5764;
assign v2103 = ~(w7139 | w7140);
assign w7141 = v2103;
assign w7142 = ~w3666 & w6236;
assign w7143 = w7141 & ~w7142;
assign w7144 = ~w7138 & w7143;
assign w7145 = ~pi17 & w7144;
assign w7146 = pi17 & ~w7144;
assign v2104 = ~(w7145 | w7146);
assign w7147 = v2104;
assign w7148 = w7137 & w7147;
assign v2105 = ~(w7135 | w7148);
assign w7149 = v2105;
assign w7150 = w7054 & ~w7149;
assign v2106 = ~(w7052 | w7150);
assign w7151 = v2106;
assign w7152 = w7039 & ~w7151;
assign w7153 = ~w7039 & w7151;
assign v2107 = ~(w7152 | w7153);
assign w7154 = v2107;
assign w7155 = w4405 & w6389;
assign w7156 = ~w4035 & w7004;
assign w7157 = ~w3920 & w6388;
assign w7158 = ~w4134 & w6871;
assign v2108 = ~(w7157 | w7158);
assign w7159 = v2108;
assign w7160 = ~w7156 & w7159;
assign w7161 = ~w7155 & w7160;
assign w7162 = pi14 & ~w7161;
assign w7163 = ~pi14 & w7161;
assign v2109 = ~(w7162 | w7163);
assign w7164 = v2109;
assign w7165 = w7154 & w7164;
assign v2110 = ~(w7152 | w7165);
assign w7166 = v2110;
assign w7167 = pi10 & ~pi11;
assign w7168 = ~pi10 & pi11;
assign v2111 = ~(w7167 | w7168);
assign w7169 = v2111;
assign v2112 = ~(pi08 | pi09);
assign w7170 = v2112;
assign w7171 = pi08 & pi09;
assign v2113 = ~(w7170 | w7171);
assign w7172 = v2113;
assign v2114 = ~(pi09 | pi10);
assign w7173 = v2114;
assign w7174 = pi09 & pi10;
assign v2115 = ~(w7173 | w7174);
assign w7175 = v2115;
assign v2116 = ~(w7172 | w7175);
assign w7176 = v2116;
assign w7177 = ~w7169 & w7176;
assign w7178 = ~w7169 & w7172;
assign w7179 = ~w4422 & w7178;
assign v2117 = ~(w7177 | w7179);
assign w7180 = v2117;
assign v2118 = ~(w4191 | w7180);
assign w7181 = v2118;
assign w7182 = ~pi11 & w7181;
assign w7183 = pi11 & ~w7181;
assign v2119 = ~(w7182 | w7183);
assign w7184 = v2119;
assign v2120 = ~(w7166 | w7184);
assign w7185 = v2120;
assign v2121 = ~(w7013 | w7015);
assign w7186 = v2121;
assign v2122 = ~(w7016 | w7186);
assign w7187 = v2122;
assign w7188 = w7166 & w7184;
assign v2123 = ~(w7185 | w7188);
assign w7189 = v2123;
assign w7190 = w7187 & w7189;
assign v2124 = ~(w7185 | w7190);
assign w7191 = v2124;
assign v2125 = ~(w7030 | w7032);
assign w7192 = v2125;
assign v2126 = ~(w7033 | w7192);
assign w7193 = v2126;
assign w7194 = ~w7191 & w7193;
assign w7195 = w7191 & ~w7193;
assign v2127 = ~(w7194 | w7195);
assign w7196 = v2127;
assign v2128 = ~(w7187 | w7189);
assign w7197 = v2128;
assign v2129 = ~(w7190 | w7197);
assign w7198 = v2129;
assign w7199 = ~w7054 & w7149;
assign v2130 = ~(w7150 | w7199);
assign w7200 = v2130;
assign w7201 = w4309 & w6389;
assign w7202 = ~w3920 & w6871;
assign w7203 = ~w3752 & w6388;
assign w7204 = ~w4134 & w7004;
assign v2131 = ~(w7203 | w7204);
assign w7205 = v2131;
assign w7206 = ~w7202 & w7205;
assign w7207 = ~w7201 & w7206;
assign w7208 = pi14 & ~w7207;
assign w7209 = ~pi14 & w7207;
assign v2132 = ~(w7208 | w7209);
assign w7210 = v2132;
assign w7211 = w7200 & w7210;
assign v2133 = ~(w7137 | w7147);
assign w7212 = v2133;
assign v2134 = ~(w7148 | w7212);
assign w7213 = v2134;
assign v2135 = ~(w7122 | w7132);
assign w7214 = v2135;
assign v2136 = ~(w7133 | w7214);
assign w7215 = v2136;
assign w7216 = w7115 & ~w7117;
assign v2137 = ~(w7118 | w7216);
assign w7217 = v2137;
assign w7218 = w4538 & w5114;
assign w7219 = ~w1795 & w5610;
assign w7220 = ~w1860 & w5531;
assign w7221 = ~w1942 & w5113;
assign v2138 = ~(w7220 | w7221);
assign w7222 = v2138;
assign w7223 = ~w7219 & w7222;
assign w7224 = ~w7218 & w7223;
assign w7225 = pi20 & ~w7224;
assign w7226 = ~pi20 & w7224;
assign v2139 = ~(w7225 | w7226);
assign w7227 = v2139;
assign w7228 = w7217 & w7227;
assign v2140 = ~(w7103 | w7113);
assign w7229 = v2140;
assign v2141 = ~(w7114 | w7229);
assign w7230 = v2141;
assign w7231 = ~w7088 & w7098;
assign v2142 = ~(w7099 | w7231);
assign w7232 = v2142;
assign w7233 = w6754 & ~w6756;
assign v2143 = ~(w6757 | w7233);
assign w7234 = v2143;
assign w7235 = w3529 & ~w6447;
assign w7236 = ~w2846 & w3767;
assign w7237 = ~w2811 & w3763;
assign w7238 = ~w2724 & w3760;
assign v2144 = ~(w7237 | w7238);
assign w7239 = v2144;
assign w7240 = ~w7236 & w7239;
assign w7241 = ~w7235 & w7240;
assign w7242 = pi29 & ~w7241;
assign w7243 = ~pi29 & w7241;
assign v2145 = ~(w7242 | w7243);
assign w7244 = v2145;
assign w7245 = w7234 & w7244;
assign w7246 = w6750 & ~w6752;
assign v2146 = ~(w6753 | w7246);
assign w7247 = v2146;
assign w7248 = ~w2937 & w3767;
assign w7249 = w3529 & w6459;
assign w7250 = ~w2846 & w3763;
assign w7251 = ~w2811 & w3760;
assign v2147 = ~(w7250 | w7251);
assign w7252 = v2147;
assign w7253 = ~w7249 & w7252;
assign w7254 = ~w7248 & w7253;
assign w7255 = ~pi29 & w7254;
assign w7256 = pi29 & ~w7254;
assign v2148 = ~(w7255 | w7256);
assign w7257 = v2148;
assign w7258 = w7247 & w7257;
assign w7259 = w6746 & ~w6748;
assign v2149 = ~(w6749 | w7259);
assign w7260 = v2149;
assign w7261 = w3529 & w6130;
assign w7262 = ~w2846 & w3760;
assign w7263 = ~w3000 & w3767;
assign w7264 = ~w2937 & w3763;
assign v2150 = ~(w7263 | w7264);
assign w7265 = v2150;
assign w7266 = ~w7262 & w7265;
assign w7267 = ~w7261 & w7266;
assign w7268 = ~pi29 & w7267;
assign w7269 = pi29 & ~w7267;
assign v2151 = ~(w7268 | w7269);
assign w7270 = v2151;
assign w7271 = w7260 & w7270;
assign w7272 = w6742 & ~w6744;
assign v2152 = ~(w6745 | w7272);
assign w7273 = v2152;
assign w7274 = w3529 & ~w6505;
assign w7275 = ~w3000 & w3763;
assign w7276 = ~w2937 & w3760;
assign v2153 = ~(w7275 | w7276);
assign w7277 = v2153;
assign w7278 = ~w3068 & w3767;
assign w7279 = w7277 & ~w7278;
assign w7280 = ~w7274 & w7279;
assign v2154 = ~(pi29 | w7280);
assign w7281 = v2154;
assign w7282 = pi29 & w7280;
assign v2155 = ~(w7281 | w7282);
assign w7283 = v2155;
assign w7284 = w7273 & ~w7283;
assign w7285 = ~w6731 & w6740;
assign v2156 = ~(w6741 | w7285);
assign w7286 = v2156;
assign w7287 = ~w3068 & w3763;
assign w7288 = ~w3124 & w3767;
assign w7289 = ~w3000 & w3760;
assign v2157 = ~(w7288 | w7289);
assign w7290 = v2157;
assign w7291 = ~w7287 & w7290;
assign w7292 = (w7291 & w6551) | (w7291 & w31167) | (w6551 & w31167);
assign w7293 = ~pi29 & w7292;
assign w7294 = pi29 & ~w7292;
assign v2158 = ~(w7293 | w7294);
assign w7295 = v2158;
assign w7296 = w7286 & w7295;
assign w7297 = w6672 & w6681;
assign v2159 = ~(w6682 | w7297);
assign w7298 = v2159;
assign w7299 = ~w3124 & w3763;
assign w7300 = ~w3068 & w3760;
assign v2160 = ~(w7299 | w7300);
assign w7301 = v2160;
assign w7302 = ~w3162 & w3767;
assign w7303 = w7301 & ~w7302;
assign w7304 = (w6603 & w31005) | (w6603 & w31006) | (w31005 & w31006);
assign w7305 = (~w6603 & w31007) | (~w6603 & w31008) | (w31007 & w31008);
assign v2161 = ~(w7304 | w7305);
assign w7306 = v2161;
assign w7307 = w7298 & ~w7306;
assign w7308 = w3262 & ~w3332;
assign v2162 = ~(w6673 | w7308);
assign w7309 = v2162;
assign w7310 = w928 & ~w7309;
assign w7311 = ~w3332 & w3402;
assign w7312 = ~w3262 & w3406;
assign v2163 = ~(w7311 | w7312);
assign w7313 = v2163;
assign w7314 = ~w7310 & w7313;
assign w7315 = ~w3211 & w3767;
assign w7316 = ~w3124 & w3760;
assign v2164 = ~(w7315 | w7316);
assign w7317 = v2164;
assign w7318 = ~w3162 & w3763;
assign w7319 = w7317 & ~w7318;
assign w7320 = (~w6641 & w30790) | (~w6641 & w30791) | (w30790 & w30791);
assign w7321 = (w6641 & w30792) | (w6641 & w30793) | (w30792 & w30793);
assign v2165 = ~(w7320 | w7321);
assign w7322 = v2165;
assign v2166 = ~(w7314 | w7322);
assign w7323 = v2166;
assign v2167 = ~(w3332 | w3405);
assign w7324 = v2167;
assign w7325 = ~w3332 & w3525;
assign w7326 = w3529 & ~w7309;
assign w7327 = (w3760 & ~w3261) | (w3760 & w30794) | (~w3261 & w30794);
assign w7328 = (w3763 & ~w3331) | (w3763 & w30795) | (~w3331 & w30795);
assign v2168 = ~(w7327 | w7328);
assign w7329 = v2168;
assign w7330 = ~w7326 & w7329;
assign w7331 = ~w7326 & w30796;
assign w7332 = ~w3262 & w3763;
assign w7333 = (w3767 & ~w3331) | (w3767 & w31009) | (~w3331 & w31009);
assign w7334 = (w3760 & ~w3210) | (w3760 & w31010) | (~w3210 & w31010);
assign v2169 = ~(w7333 | w7334);
assign w7335 = v2169;
assign w7336 = (~w6676 & w30797) | (~w6676 & w30798) | (w30797 & w30798);
assign w7337 = w7331 & w7336;
assign w7338 = w7324 & w7337;
assign v2170 = ~(w7324 | w7337);
assign w7339 = v2170;
assign v2171 = ~(w7338 | w7339);
assign w7340 = v2171;
assign w7341 = ~w3162 & w3760;
assign w7342 = (w3767 & ~w3261) | (w3767 & w31168) | (~w3261 & w31168);
assign w7343 = (w3763 & ~w3210) | (w3763 & w31169) | (~w3210 & w31169);
assign v2172 = ~(w7342 | w7343);
assign w7344 = v2172;
assign w7345 = ~w7341 & w7344;
assign w7346 = (w6735 & w31011) | (w6735 & w31012) | (w31011 & w31012);
assign w7347 = (~w6735 & w31013) | (~w6735 & w31014) | (w31013 & w31014);
assign v2173 = ~(w7346 | w7347);
assign w7348 = v2173;
assign w7349 = w7340 & w7348;
assign w7350 = (~w7338 & ~w7340) | (~w7338 & w31015) | (~w7340 & w31015);
assign w7351 = w7314 & w7322;
assign v2174 = ~(w7323 | w7351);
assign w7352 = v2174;
assign w7353 = ~w7350 & w7352;
assign w7354 = (~w7323 & ~w7352) | (~w7323 & w31016) | (~w7352 & w31016);
assign w7355 = ~w7298 & w7306;
assign v2175 = ~(w7307 | w7355);
assign w7356 = v2175;
assign w7357 = ~w7354 & w7356;
assign v2176 = ~(w7307 | w7357);
assign w7358 = v2176;
assign v2177 = ~(w7286 | w7295);
assign w7359 = v2177;
assign v2178 = ~(w7296 | w7359);
assign w7360 = v2178;
assign w7361 = ~w7358 & w7360;
assign w7362 = (~w7296 & w7358) | (~w7296 & w31170) | (w7358 & w31170);
assign w7363 = ~w7273 & w7283;
assign v2179 = ~(w7284 | w7363);
assign w7364 = v2179;
assign w7365 = ~w7362 & w7364;
assign v2180 = ~(w7284 | w7365);
assign w7366 = v2180;
assign v2181 = ~(w7260 | w7270);
assign w7367 = v2181;
assign v2182 = ~(w7271 | w7367);
assign w7368 = v2182;
assign w7369 = ~w7366 & w7368;
assign v2183 = ~(w7271 | w7369);
assign w7370 = v2183;
assign v2184 = ~(w7247 | w7257);
assign w7371 = v2184;
assign v2185 = ~(w7258 | w7371);
assign w7372 = v2185;
assign w7373 = ~w7370 & w7372;
assign v2186 = ~(w7258 | w7373);
assign w7374 = v2186;
assign v2187 = ~(w7234 | w7244);
assign w7375 = v2187;
assign v2188 = ~(w7245 | w7375);
assign w7376 = v2188;
assign w7377 = ~w7374 & w7376;
assign v2189 = ~(w7245 | w7377);
assign w7378 = v2189;
assign w7379 = ~w6765 & w6775;
assign v2190 = ~(w6776 | w7379);
assign w7380 = v2190;
assign w7381 = ~w7378 & w7380;
assign w7382 = w7378 & ~w7380;
assign v2191 = ~(w7381 | w7382);
assign w7383 = v2191;
assign w7384 = w4153 & w5898;
assign w7385 = ~w2568 & w4158;
assign v2192 = ~(w2596 | w2873);
assign w7386 = v2192;
assign w7387 = ~w2492 & w4155;
assign v2193 = ~(w7386 | w7387);
assign w7388 = v2193;
assign w7389 = ~w7385 & w7388;
assign w7390 = ~w7384 & w7389;
assign w7391 = pi26 & ~w7390;
assign w7392 = ~pi26 & w7390;
assign v2194 = ~(w7391 | w7392);
assign w7393 = v2194;
assign w7394 = w7383 & w7393;
assign v2195 = ~(w7381 | w7394);
assign w7395 = v2195;
assign w7396 = w7232 & ~w7395;
assign w7397 = w4764 & w5262;
assign w7398 = ~w2202 & w4913;
assign w7399 = ~w2339 & w4763;
assign w7400 = ~w2290 & w4836;
assign v2196 = ~(w7399 | w7400);
assign w7401 = v2196;
assign w7402 = ~w7398 & w7401;
assign w7403 = ~w7397 & w7402;
assign w7404 = pi23 & ~w7403;
assign w7405 = ~pi23 & w7403;
assign v2197 = ~(w7404 | w7405);
assign w7406 = v2197;
assign w7407 = ~w7232 & w7395;
assign v2198 = ~(w7396 | w7407);
assign w7408 = v2198;
assign w7409 = w7406 & w7408;
assign v2199 = ~(w7396 | w7409);
assign w7410 = v2199;
assign w7411 = w7230 & ~w7410;
assign w7412 = ~w7230 & w7410;
assign v2200 = ~(w7411 | w7412);
assign w7413 = v2200;
assign w7414 = w4854 & w5114;
assign w7415 = ~w1860 & w5610;
assign w7416 = ~w2038 & w5113;
assign w7417 = ~w1942 & w5531;
assign v2201 = ~(w7416 | w7417);
assign w7418 = v2201;
assign w7419 = ~w7415 & w7418;
assign w7420 = ~w7414 & w7419;
assign w7421 = pi20 & ~w7420;
assign w7422 = ~pi20 & w7420;
assign v2202 = ~(w7421 | w7422);
assign w7423 = v2202;
assign w7424 = w7413 & w7423;
assign v2203 = ~(w7411 | w7424);
assign w7425 = v2203;
assign v2204 = ~(w7217 | w7227);
assign w7426 = v2204;
assign v2205 = ~(w7228 | w7426);
assign w7427 = v2205;
assign w7428 = ~w7425 & w7427;
assign v2206 = ~(w7228 | w7428);
assign w7429 = v2206;
assign w7430 = w7215 & ~w7429;
assign w7431 = ~w7215 & w7429;
assign v2207 = ~(w7430 | w7431);
assign w7432 = v2207;
assign w7433 = ~w1387 & w6236;
assign w7434 = w3397 & w5765;
assign w7435 = ~w1496 & w5983;
assign w7436 = ~w1609 & w5764;
assign v2208 = ~(w7435 | w7436);
assign w7437 = v2208;
assign w7438 = ~w7434 & w7437;
assign w7439 = ~w7433 & w7438;
assign w7440 = pi17 & w7439;
assign v2209 = ~(pi17 | w7439);
assign w7441 = v2209;
assign v2210 = ~(w7440 | w7441);
assign w7442 = v2210;
assign w7443 = w7432 & ~w7442;
assign v2211 = ~(w7430 | w7443);
assign w7444 = v2211;
assign w7445 = w7213 & ~w7444;
assign w7446 = ~w7213 & w7444;
assign v2212 = ~(w7445 | w7446);
assign w7447 = v2212;
assign w7448 = ~w3928 & w6389;
assign w7449 = ~w3752 & w6871;
assign w7450 = ~w3587 & w6388;
assign w7451 = ~w3920 & w7004;
assign v2213 = ~(w7450 | w7451);
assign w7452 = v2213;
assign w7453 = ~w7449 & w7452;
assign w7454 = ~w7448 & w7453;
assign w7455 = pi14 & ~w7454;
assign w7456 = ~pi14 & w7454;
assign v2214 = ~(w7455 | w7456);
assign w7457 = v2214;
assign w7458 = w7447 & w7457;
assign v2215 = ~(w7445 | w7458);
assign w7459 = v2215;
assign v2216 = ~(w7200 | w7210);
assign w7460 = v2216;
assign v2217 = ~(w7211 | w7460);
assign w7461 = v2217;
assign w7462 = ~w7459 & w7461;
assign v2218 = ~(w7211 | w7462);
assign w7463 = v2218;
assign w7464 = w4425 & w7178;
assign w7465 = ~w4082 & w7177;
assign w7466 = ~w7172 & w7175;
assign w7467 = ~w4191 & w7466;
assign v2219 = ~(w7465 | w7467);
assign w7468 = v2219;
assign w7469 = ~w7464 & w7468;
assign w7470 = pi11 & ~w7469;
assign w7471 = ~pi11 & w7469;
assign v2220 = ~(w7470 | w7471);
assign w7472 = v2220;
assign w7473 = ~w7463 & w7472;
assign v2221 = ~(w7154 | w7164);
assign w7474 = v2221;
assign v2222 = ~(w7165 | w7474);
assign w7475 = v2222;
assign w7476 = w7463 & ~w7472;
assign v2223 = ~(w7473 | w7476);
assign w7477 = v2223;
assign w7478 = w7475 & w7477;
assign v2224 = ~(w7473 | w7478);
assign w7479 = v2224;
assign w7480 = w7198 & ~w7479;
assign w7481 = ~w7198 & w7479;
assign v2225 = ~(w7447 | w7457);
assign w7482 = v2225;
assign v2226 = ~(w7458 | w7482);
assign w7483 = v2226;
assign w7484 = ~w7432 & w7442;
assign v2227 = ~(w7443 | w7484);
assign w7485 = v2227;
assign w7486 = w7425 & ~w7427;
assign v2228 = ~(w7428 | w7486);
assign w7487 = v2228;
assign w7488 = ~w3510 & w5765;
assign w7489 = ~w1496 & w6236;
assign w7490 = ~w1609 & w5983;
assign v2229 = ~(w7489 | w7490);
assign w7491 = v2229;
assign w7492 = ~w1674 & w5764;
assign w7493 = w7491 & ~w7492;
assign w7494 = ~w7488 & w7493;
assign w7495 = ~pi17 & w7494;
assign w7496 = pi17 & ~w7494;
assign v2230 = ~(w7495 | w7496);
assign w7497 = v2230;
assign w7498 = w7487 & w7497;
assign v2231 = ~(w7413 | w7423);
assign w7499 = v2231;
assign v2232 = ~(w7424 | w7499);
assign w7500 = v2232;
assign v2233 = ~(w7406 | w7408);
assign w7501 = v2233;
assign v2234 = ~(w7409 | w7501);
assign w7502 = v2234;
assign w7503 = w7374 & ~w7376;
assign v2235 = ~(w7377 | w7503);
assign w7504 = v2235;
assign w7505 = w4153 & w6031;
assign w7506 = ~w2568 & w4155;
assign w7507 = ~w2596 & w4158;
assign v2236 = ~(w7506 | w7507);
assign w7508 = v2236;
assign v2237 = ~(w2669 | w2873);
assign w7509 = v2237;
assign w7510 = w7508 & ~w7509;
assign w7511 = ~w7505 & w7510;
assign w7512 = ~pi26 & w7511;
assign w7513 = pi26 & ~w7511;
assign v2238 = ~(w7512 | w7513);
assign w7514 = v2238;
assign w7515 = w7504 & w7514;
assign w7516 = w7370 & ~w7372;
assign v2239 = ~(w7373 | w7516);
assign w7517 = v2239;
assign w7518 = w4153 & w5880;
assign w7519 = ~w2669 & w4158;
assign w7520 = ~w2596 & w4155;
assign v2240 = ~(w2724 | w2873);
assign w7521 = v2240;
assign v2241 = ~(w7520 | w7521);
assign w7522 = v2241;
assign w7523 = ~w7519 & w7522;
assign w7524 = ~w7518 & w7523;
assign w7525 = pi26 & ~w7524;
assign w7526 = ~pi26 & w7524;
assign v2242 = ~(w7525 | w7526);
assign w7527 = v2242;
assign w7528 = w7517 & w7527;
assign w7529 = w7366 & ~w7368;
assign v2243 = ~(w7369 | w7529);
assign w7530 = v2243;
assign w7531 = ~w2669 & w4155;
assign w7532 = w4153 & w6148;
assign v2244 = ~(w2811 | w2873);
assign w7533 = v2244;
assign w7534 = ~w2724 & w4158;
assign v2245 = ~(w7533 | w7534);
assign w7535 = v2245;
assign w7536 = ~w7532 & w7535;
assign w7537 = ~w7531 & w7536;
assign w7538 = pi26 & w7537;
assign v2246 = ~(pi26 | w7537);
assign w7539 = v2246;
assign v2247 = ~(w7538 | w7539);
assign w7540 = v2247;
assign w7541 = w7530 & ~w7540;
assign w7542 = w7362 & ~w7364;
assign v2248 = ~(w7365 | w7542);
assign w7543 = v2248;
assign w7544 = w4153 & ~w6447;
assign w7545 = ~w2724 & w4155;
assign w7546 = ~w2811 & w4158;
assign v2249 = ~(w7545 | w7546);
assign w7547 = v2249;
assign v2250 = ~(w2846 | w2873);
assign w7548 = v2250;
assign w7549 = w7547 & ~w7548;
assign w7550 = ~w7544 & w7549;
assign w7551 = ~pi26 & w7550;
assign w7552 = pi26 & ~w7550;
assign v2251 = ~(w7551 | w7552);
assign w7553 = v2251;
assign w7554 = w7543 & w7553;
assign w7555 = w7358 & ~w7360;
assign v2252 = ~(w7361 | w7555);
assign w7556 = v2252;
assign w7557 = w4153 & w6459;
assign v2253 = ~(w2873 | w2937);
assign w7558 = v2253;
assign w7559 = ~w2811 & w4155;
assign w7560 = ~w2846 & w4158;
assign v2254 = ~(w7559 | w7560);
assign w7561 = v2254;
assign w7562 = ~w7558 & w7561;
assign w7563 = ~w7557 & w7562;
assign w7564 = pi26 & ~w7563;
assign w7565 = ~pi26 & w7563;
assign v2255 = ~(w7564 | w7565);
assign w7566 = v2255;
assign w7567 = w7556 & w7566;
assign w7568 = w7354 & ~w7356;
assign v2256 = ~(w7357 | w7568);
assign w7569 = v2256;
assign w7570 = w4153 & w6130;
assign w7571 = ~w2846 & w4155;
assign v2257 = ~(w2873 | w3000);
assign w7572 = v2257;
assign w7573 = ~w2937 & w4158;
assign v2258 = ~(w7572 | w7573);
assign w7574 = v2258;
assign w7575 = ~w7571 & w7574;
assign w7576 = ~w7570 & w7575;
assign w7577 = ~pi26 & w7576;
assign w7578 = pi26 & ~w7576;
assign v2259 = ~(w7577 | w7578);
assign w7579 = v2259;
assign w7580 = w7569 & w7579;
assign w7581 = w7350 & ~w7352;
assign v2260 = ~(w7353 | w7581);
assign w7582 = v2260;
assign w7583 = ~w3000 & w4158;
assign w7584 = ~w2937 & w4155;
assign v2261 = ~(w7583 | w7584);
assign w7585 = v2261;
assign v2262 = ~(w2873 | w3068);
assign w7586 = v2262;
assign w7587 = w7585 & ~w7586;
assign w7588 = (w7587 & w6505) | (w7587 & w31017) | (w6505 & w31017);
assign w7589 = pi26 & w7588;
assign v2263 = ~(pi26 | w7588);
assign w7590 = v2263;
assign v2264 = ~(w7589 | w7590);
assign w7591 = v2264;
assign w7592 = w7582 & ~w7591;
assign v2265 = ~(w7340 | w7348);
assign w7593 = v2265;
assign v2266 = ~(w7349 | w7593);
assign w7594 = v2266;
assign w7595 = ~w3000 & w4155;
assign w7596 = ~w3068 & w4158;
assign v2267 = ~(w7595 | w7596);
assign w7597 = v2267;
assign v2268 = ~(w2873 | w3124);
assign w7598 = v2268;
assign w7599 = w7597 & ~w7598;
assign w7600 = (w6551 & w31018) | (w6551 & w31019) | (w31018 & w31019);
assign w7601 = (~w6551 & w31020) | (~w6551 & w31021) | (w31020 & w31021);
assign v2269 = ~(w7600 | w7601);
assign w7602 = v2269;
assign w7603 = w7594 & ~w7602;
assign w7604 = ~w3124 & w4158;
assign w7605 = ~w3068 & w4155;
assign v2270 = ~(w7604 | w7605);
assign w7606 = v2270;
assign v2271 = ~(w2873 | w3162);
assign w7607 = v2271;
assign w7608 = w7606 & ~w7607;
assign w7609 = (w6603 & w30589) | (w6603 & w30590) | (w30589 & w30590);
assign w7610 = (~w6603 & w30591) | (~w6603 & w30592) | (w30591 & w30592);
assign v2272 = ~(w7609 | w7610);
assign w7611 = v2272;
assign w7612 = pi29 & ~w7331;
assign w7613 = ~w7336 & w7612;
assign w7614 = w7336 & ~w7612;
assign v2273 = ~(w7613 | w7614);
assign w7615 = v2273;
assign w7616 = ~w7611 & w7615;
assign w7617 = pi29 & w7325;
assign v2274 = ~(w7330 | w7617);
assign w7618 = v2274;
assign w7619 = w7330 & w7617;
assign v2275 = ~(w7618 | w7619);
assign w7620 = v2275;
assign w7621 = ~w3124 & w4155;
assign v2276 = ~(w2873 | w3211);
assign w7622 = v2276;
assign w7623 = ~w3162 & w4158;
assign v2277 = ~(w7622 | w7623);
assign w7624 = v2277;
assign w7625 = ~w7621 & w7624;
assign w7626 = (~w6641 & w30477) | (~w6641 & w30478) | (w30477 & w30478);
assign w7627 = (w6641 & w30479) | (w6641 & w30480) | (w30479 & w30480);
assign v2278 = ~(w7626 | w7627);
assign w7628 = v2278;
assign v2279 = ~(w7620 | w7628);
assign w7629 = v2279;
assign w7630 = ~w3332 & w4152;
assign w7631 = w4153 & ~w7309;
assign w7632 = (w4158 & ~w3331) | (w4158 & w30481) | (~w3331 & w30481);
assign w7633 = (w4155 & ~w3261) | (w4155 & w30482) | (~w3261 & w30482);
assign v2280 = ~(w7632 | w7633);
assign w7634 = v2280;
assign w7635 = ~w7631 & w7634;
assign w7636 = ~w7631 & w30483;
assign w7637 = ~w3262 & w4158;
assign w7638 = (~w2873 & ~w3331) | (~w2873 & w30593) | (~w3331 & w30593);
assign w7639 = (w4155 & ~w3210) | (w4155 & w30594) | (~w3210 & w30594);
assign v2281 = ~(w7638 | w7639);
assign w7640 = v2281;
assign w7641 = (~w6676 & w30484) | (~w6676 & w30485) | (w30484 & w30485);
assign w7642 = w7636 & w7641;
assign w7643 = w7325 & w7642;
assign v2282 = ~(w7325 | w7642);
assign w7644 = v2282;
assign v2283 = ~(w7643 | w7644);
assign w7645 = v2283;
assign w7646 = (w4158 & ~w3210) | (w4158 & w30800) | (~w3210 & w30800);
assign w7647 = ~w3162 & w4155;
assign v2284 = ~(w7646 | w7647);
assign w7648 = v2284;
assign v2285 = ~(w2873 | w3262);
assign w7649 = v2285;
assign w7650 = (~w6735 & w30595) | (~w6735 & w30596) | (w30595 & w30596);
assign w7651 = (w6735 & w30597) | (w6735 & w30598) | (w30597 & w30598);
assign v2286 = ~(w7650 | w7651);
assign w7652 = v2286;
assign w7653 = w7645 & ~w7652;
assign w7654 = (~w7643 & ~w7645) | (~w7643 & w30599) | (~w7645 & w30599);
assign w7655 = w7620 & w7628;
assign v2287 = ~(w7629 | w7655);
assign w7656 = v2287;
assign w7657 = ~w7654 & w7656;
assign w7658 = (~w7629 & ~w7656) | (~w7629 & w30600) | (~w7656 & w30600);
assign w7659 = w7611 & ~w7615;
assign v2288 = ~(w7616 | w7659);
assign w7660 = v2288;
assign w7661 = ~w7658 & w7660;
assign v2289 = ~(w7616 | w7661);
assign w7662 = v2289;
assign w7663 = ~w7594 & w7602;
assign v2290 = ~(w7603 | w7663);
assign w7664 = v2290;
assign w7665 = ~w7662 & w7664;
assign w7666 = (~w7603 & w7662) | (~w7603 & w30801) | (w7662 & w30801);
assign w7667 = ~w7582 & w7591;
assign v2291 = ~(w7592 | w7667);
assign w7668 = v2291;
assign w7669 = ~w7666 & w7668;
assign v2292 = ~(w7592 | w7669);
assign w7670 = v2292;
assign v2293 = ~(w7569 | w7579);
assign w7671 = v2293;
assign v2294 = ~(w7580 | w7671);
assign w7672 = v2294;
assign w7673 = ~w7670 & w7672;
assign w7674 = (~w7580 & w7670) | (~w7580 & w31022) | (w7670 & w31022);
assign v2295 = ~(w7556 | w7566);
assign w7675 = v2295;
assign v2296 = ~(w7567 | w7675);
assign w7676 = v2296;
assign w7677 = ~w7674 & w7676;
assign v2297 = ~(w7567 | w7677);
assign w7678 = v2297;
assign v2298 = ~(w7543 | w7553);
assign w7679 = v2298;
assign v2299 = ~(w7554 | w7679);
assign w7680 = v2299;
assign w7681 = ~w7678 & w7680;
assign w7682 = (~w7554 & w7678) | (~w7554 & w31171) | (w7678 & w31171);
assign w7683 = ~w7530 & w7540;
assign v2300 = ~(w7541 | w7683);
assign w7684 = v2300;
assign w7685 = ~w7682 & w7684;
assign v2301 = ~(w7541 | w7685);
assign w7686 = v2301;
assign v2302 = ~(w7517 | w7527);
assign w7687 = v2302;
assign v2303 = ~(w7528 | w7687);
assign w7688 = v2303;
assign w7689 = ~w7686 & w7688;
assign v2304 = ~(w7528 | w7689);
assign w7690 = v2304;
assign v2305 = ~(w7504 | w7514);
assign w7691 = v2305;
assign v2306 = ~(w7515 | w7691);
assign w7692 = v2306;
assign w7693 = ~w7690 & w7692;
assign v2307 = ~(w7515 | w7693);
assign w7694 = v2307;
assign v2308 = ~(w7383 | w7393);
assign w7695 = v2308;
assign v2309 = ~(w7394 | w7695);
assign w7696 = v2309;
assign w7697 = ~w7694 & w7696;
assign w7698 = w7694 & ~w7696;
assign v2310 = ~(w7697 | w7698);
assign w7699 = v2310;
assign w7700 = w4764 & w5280;
assign w7701 = ~w2290 & w4913;
assign w7702 = ~w2339 & w4836;
assign w7703 = ~w2424 & w4763;
assign v2311 = ~(w7702 | w7703);
assign w7704 = v2311;
assign w7705 = ~w7701 & w7704;
assign w7706 = ~w7700 & w7705;
assign w7707 = pi23 & ~w7706;
assign w7708 = ~pi23 & w7706;
assign v2312 = ~(w7707 | w7708);
assign w7709 = v2312;
assign w7710 = w7699 & w7709;
assign v2313 = ~(w7697 | w7710);
assign w7711 = v2313;
assign w7712 = w7502 & ~w7711;
assign w7713 = ~w7502 & w7711;
assign v2314 = ~(w7712 | w7713);
assign w7714 = v2314;
assign w7715 = w4702 & w5114;
assign w7716 = ~w2089 & w5113;
assign w7717 = ~w2038 & w5531;
assign v2315 = ~(w7716 | w7717);
assign w7718 = v2315;
assign w7719 = ~w1942 & w5610;
assign w7720 = w7718 & ~w7719;
assign w7721 = ~w7715 & w7720;
assign w7722 = ~pi20 & w7721;
assign w7723 = pi20 & ~w7721;
assign v2316 = ~(w7722 | w7723);
assign w7724 = v2316;
assign w7725 = w7714 & w7724;
assign v2317 = ~(w7712 | w7725);
assign w7726 = v2317;
assign w7727 = w7500 & ~w7726;
assign w7728 = ~w7500 & w7726;
assign v2318 = ~(w7727 | w7728);
assign w7729 = v2318;
assign w7730 = w3494 & w5765;
assign w7731 = ~w1609 & w6236;
assign w7732 = ~w1674 & w5983;
assign v2319 = ~(w7731 | w7732);
assign w7733 = v2319;
assign w7734 = ~w1795 & w5764;
assign w7735 = w7733 & ~w7734;
assign w7736 = ~w7730 & w7735;
assign w7737 = ~pi17 & w7736;
assign w7738 = pi17 & ~w7736;
assign v2320 = ~(w7737 | w7738);
assign w7739 = v2320;
assign w7740 = w7729 & w7739;
assign v2321 = ~(w7727 | w7740);
assign w7741 = v2321;
assign v2322 = ~(w7487 | w7497);
assign w7742 = v2322;
assign v2323 = ~(w7498 | w7742);
assign w7743 = v2323;
assign w7744 = ~w7741 & w7743;
assign v2324 = ~(w7498 | w7744);
assign w7745 = v2324;
assign w7746 = w7485 & ~w7745;
assign w7747 = ~w7485 & w7745;
assign v2325 = ~(w7746 | w7747);
assign w7748 = v2325;
assign w7749 = w3758 & w6389;
assign w7750 = ~w3752 & w7004;
assign w7751 = ~w3587 & w6871;
assign v2326 = ~(w7750 | w7751);
assign w7752 = v2326;
assign w7753 = ~w3666 & w6388;
assign w7754 = w7752 & ~w7753;
assign w7755 = ~w7749 & w7754;
assign w7756 = pi14 & ~w7755;
assign w7757 = ~pi14 & w7755;
assign v2327 = ~(w7756 | w7757);
assign w7758 = v2327;
assign w7759 = w7748 & w7758;
assign v2328 = ~(w7746 | w7759);
assign w7760 = v2328;
assign w7761 = w7483 & ~w7760;
assign w7762 = ~w7483 & w7760;
assign v2329 = ~(w7761 | w7762);
assign w7763 = v2329;
assign w7764 = ~w4149 & w7178;
assign w7765 = w7169 & w7172;
assign w7766 = ~w4082 & w7765;
assign w7767 = ~w4134 & w7177;
assign w7768 = ~w4035 & w7466;
assign v2330 = ~(w7767 | w7768);
assign w7769 = v2330;
assign w7770 = ~w7766 & w7769;
assign w7771 = ~w7764 & w7770;
assign w7772 = pi11 & ~w7771;
assign w7773 = ~pi11 & w7771;
assign v2331 = ~(w7772 | w7773);
assign w7774 = v2331;
assign w7775 = w7763 & w7774;
assign v2332 = ~(w7761 | w7775);
assign w7776 = v2332;
assign w7777 = w4196 & w7178;
assign w7778 = ~w4082 & w7466;
assign w7779 = ~w4191 & w7765;
assign w7780 = ~w4035 & w7177;
assign v2333 = ~(w7779 | w7780);
assign w7781 = v2333;
assign w7782 = ~w7778 & w7781;
assign w7783 = ~w7777 & w7782;
assign w7784 = pi11 & ~w7783;
assign w7785 = ~pi11 & w7783;
assign v2334 = ~(w7784 | w7785);
assign w7786 = v2334;
assign w7787 = ~w7776 & w7786;
assign w7788 = w7459 & ~w7461;
assign v2335 = ~(w7462 | w7788);
assign w7789 = v2335;
assign w7790 = w7776 & ~w7786;
assign v2336 = ~(w7787 | w7790);
assign w7791 = v2336;
assign w7792 = w7789 & w7791;
assign v2337 = ~(w7787 | w7792);
assign w7793 = v2337;
assign v2338 = ~(w7475 | w7477);
assign w7794 = v2338;
assign v2339 = ~(w7478 | w7794);
assign w7795 = v2339;
assign w7796 = ~w7793 & w7795;
assign w7797 = w7793 & ~w7795;
assign v2340 = ~(w7796 | w7797);
assign w7798 = v2340;
assign v2341 = ~(w7789 | w7791);
assign w7799 = v2341;
assign v2342 = ~(w7792 | w7799);
assign w7800 = v2342;
assign v2343 = ~(w7748 | w7758);
assign w7801 = v2343;
assign v2344 = ~(w7759 | w7801);
assign w7802 = v2344;
assign w7803 = w7741 & ~w7743;
assign v2345 = ~(w7744 | w7803);
assign w7804 = v2345;
assign w7805 = w4291 & w6389;
assign w7806 = ~w3587 & w7004;
assign w7807 = ~w3666 & w6871;
assign w7808 = ~w1387 & w6388;
assign v2346 = ~(w7807 | w7808);
assign w7809 = v2346;
assign w7810 = ~w7806 & w7809;
assign w7811 = ~w7805 & w7810;
assign w7812 = pi14 & ~w7811;
assign w7813 = ~pi14 & w7811;
assign v2347 = ~(w7812 | w7813);
assign w7814 = v2347;
assign w7815 = w7804 & w7814;
assign v2348 = ~(w7729 | w7739);
assign w7816 = v2348;
assign v2349 = ~(w7740 | w7816);
assign w7817 = v2349;
assign v2350 = ~(w7714 | w7724);
assign w7818 = v2350;
assign v2351 = ~(w7725 | w7818);
assign w7819 = v2351;
assign w7820 = w7690 & ~w7692;
assign v2352 = ~(w7693 | w7820);
assign w7821 = v2352;
assign w7822 = w4764 & w5665;
assign w7823 = ~w2492 & w4763;
assign w7824 = ~w2424 & w4836;
assign w7825 = ~w2339 & w4913;
assign v2353 = ~(w7824 | w7825);
assign w7826 = v2353;
assign w7827 = ~w7823 & w7826;
assign w7828 = ~w7822 & w7827;
assign w7829 = pi23 & ~w7828;
assign w7830 = ~pi23 & w7828;
assign v2354 = ~(w7829 | w7830);
assign w7831 = v2354;
assign w7832 = w7821 & w7831;
assign w7833 = w7686 & ~w7688;
assign v2355 = ~(w7689 | w7833);
assign w7834 = v2355;
assign w7835 = ~w2568 & w4763;
assign w7836 = w4764 & w5449;
assign w7837 = ~w2492 & w4836;
assign w7838 = ~w2424 & w4913;
assign v2356 = ~(w7837 | w7838);
assign w7839 = v2356;
assign w7840 = ~w7836 & w7839;
assign w7841 = ~w7835 & w7840;
assign w7842 = pi23 & w7841;
assign v2357 = ~(pi23 | w7841);
assign w7843 = v2357;
assign v2358 = ~(w7842 | w7843);
assign w7844 = v2358;
assign w7845 = w7834 & ~w7844;
assign w7846 = w7682 & ~w7684;
assign v2359 = ~(w7685 | w7846);
assign w7847 = v2359;
assign w7848 = w4764 & w5898;
assign w7849 = ~w2568 & w4836;
assign w7850 = ~w2596 & w4763;
assign w7851 = ~w2492 & w4913;
assign v2360 = ~(w7850 | w7851);
assign w7852 = v2360;
assign w7853 = ~w7849 & w7852;
assign w7854 = ~w7848 & w7853;
assign w7855 = pi23 & ~w7854;
assign w7856 = ~pi23 & w7854;
assign v2361 = ~(w7855 | w7856);
assign w7857 = v2361;
assign w7858 = w7847 & w7857;
assign w7859 = w7678 & ~w7680;
assign v2362 = ~(w7681 | w7859);
assign w7860 = v2362;
assign w7861 = w4764 & w6031;
assign w7862 = ~w2568 & w4913;
assign w7863 = ~w2596 & w4836;
assign w7864 = ~w2669 & w4763;
assign v2363 = ~(w7863 | w7864);
assign w7865 = v2363;
assign w7866 = ~w7862 & w7865;
assign w7867 = ~w7861 & w7866;
assign w7868 = pi23 & ~w7867;
assign w7869 = ~pi23 & w7867;
assign v2364 = ~(w7868 | w7869);
assign w7870 = v2364;
assign w7871 = w7860 & w7870;
assign w7872 = w7674 & ~w7676;
assign v2365 = ~(w7677 | w7872);
assign w7873 = v2365;
assign w7874 = w4764 & w5880;
assign w7875 = ~w2669 & w4836;
assign w7876 = ~w2724 & w4763;
assign v2366 = ~(w7875 | w7876);
assign w7877 = v2366;
assign w7878 = ~w2596 & w4913;
assign w7879 = w7877 & ~w7878;
assign w7880 = ~w7874 & w7879;
assign w7881 = pi23 & ~w7880;
assign w7882 = ~pi23 & w7880;
assign v2367 = ~(w7881 | w7882);
assign w7883 = v2367;
assign w7884 = w7873 & w7883;
assign w7885 = w7670 & ~w7672;
assign v2368 = ~(w7673 | w7885);
assign w7886 = v2368;
assign w7887 = w4764 & w6148;
assign w7888 = ~w2669 & w4913;
assign w7889 = ~w2724 & w4836;
assign v2369 = ~(w7888 | w7889);
assign w7890 = v2369;
assign w7891 = ~w2811 & w4763;
assign w7892 = w7890 & ~w7891;
assign w7893 = ~w7887 & w7892;
assign w7894 = pi23 & w7893;
assign v2370 = ~(pi23 | w7893);
assign w7895 = v2370;
assign v2371 = ~(w7894 | w7895);
assign w7896 = v2371;
assign w7897 = w7886 & ~w7896;
assign w7898 = w7666 & ~w7668;
assign v2372 = ~(w7669 | w7898);
assign w7899 = v2372;
assign w7900 = ~w2846 & w4763;
assign w7901 = w4764 & ~w6447;
assign w7902 = ~w2811 & w4836;
assign w7903 = ~w2724 & w4913;
assign v2373 = ~(w7902 | w7903);
assign w7904 = v2373;
assign w7905 = ~w7901 & w7904;
assign w7906 = ~w7900 & w7905;
assign w7907 = pi23 & w7906;
assign v2374 = ~(pi23 | w7906);
assign w7908 = v2374;
assign v2375 = ~(w7907 | w7908);
assign w7909 = v2375;
assign w7910 = w7899 & ~w7909;
assign w7911 = w7662 & ~w7664;
assign v2376 = ~(w7665 | w7911);
assign w7912 = v2376;
assign w7913 = w4764 & w6459;
assign w7914 = ~w2937 & w4763;
assign w7915 = ~w2846 & w4836;
assign v2377 = ~(w7914 | w7915);
assign w7916 = v2377;
assign w7917 = ~w2811 & w4913;
assign w7918 = w7916 & ~w7917;
assign w7919 = ~w7913 & w7918;
assign w7920 = ~pi23 & w7919;
assign w7921 = pi23 & ~w7919;
assign v2378 = ~(w7920 | w7921);
assign w7922 = v2378;
assign w7923 = w7912 & w7922;
assign w7924 = w7658 & ~w7660;
assign v2379 = ~(w7661 | w7924);
assign w7925 = v2379;
assign w7926 = w4764 & w6130;
assign w7927 = ~w2846 & w4913;
assign w7928 = ~w2937 & w4836;
assign v2380 = ~(w7927 | w7928);
assign w7929 = v2380;
assign w7930 = ~w3000 & w4763;
assign w7931 = w7929 & ~w7930;
assign w7932 = ~w7926 & w7931;
assign v2381 = ~(pi23 | w7932);
assign w7933 = v2381;
assign w7934 = pi23 & w7932;
assign v2382 = ~(w7933 | w7934);
assign w7935 = v2382;
assign w7936 = w7925 & ~w7935;
assign w7937 = w7654 & ~w7656;
assign v2383 = ~(w7657 | w7937);
assign w7938 = v2383;
assign w7939 = ~w3000 & w4836;
assign w7940 = ~w2937 & w4913;
assign v2384 = ~(w7939 | w7940);
assign w7941 = v2384;
assign w7942 = ~w3068 & w4763;
assign w7943 = w7941 & ~w7942;
assign w7944 = (w7943 & w6505) | (w7943 & w30601) | (w6505 & w30601);
assign w7945 = pi23 & w7944;
assign v2385 = ~(pi23 | w7944);
assign w7946 = v2385;
assign v2386 = ~(w7945 | w7946);
assign w7947 = v2386;
assign w7948 = w7938 & ~w7947;
assign w7949 = ~w7645 & w7652;
assign v2387 = ~(w7653 | w7949);
assign w7950 = v2387;
assign w7951 = ~w3000 & w4913;
assign w7952 = ~w3068 & w4836;
assign v2388 = ~(w7951 | w7952);
assign w7953 = v2388;
assign w7954 = ~w3124 & w4763;
assign w7955 = w7953 & ~w7954;
assign w7956 = (w6551 & w30602) | (w6551 & w30603) | (w30602 & w30603);
assign w7957 = (~w6551 & w30604) | (~w6551 & w30605) | (w30604 & w30605);
assign v2389 = ~(w7956 | w7957);
assign w7958 = v2389;
assign w7959 = w7950 & ~w7958;
assign w7960 = ~w3124 & w4836;
assign w7961 = ~w3068 & w4913;
assign v2390 = ~(w7960 | w7961);
assign w7962 = v2390;
assign w7963 = ~w3162 & w4763;
assign w7964 = w7962 & ~w7963;
assign w7965 = (w6603 & w30311) | (w6603 & w30312) | (w30311 & w30312);
assign w7966 = (~w6603 & w30313) | (~w6603 & w30314) | (w30313 & w30314);
assign v2391 = ~(w7965 | w7966);
assign w7967 = v2391;
assign w7968 = pi26 & ~w7636;
assign w7969 = ~w7641 & w7968;
assign w7970 = w7641 & ~w7968;
assign v2392 = ~(w7969 | w7970);
assign w7971 = v2392;
assign w7972 = ~w7967 & w7971;
assign w7973 = pi26 & w7630;
assign v2393 = ~(w7635 | w7973);
assign w7974 = v2393;
assign w7975 = w7635 & w7973;
assign v2394 = ~(w7974 | w7975);
assign w7976 = v2394;
assign w7977 = ~w3162 & w4836;
assign w7978 = ~w3211 & w4763;
assign v2395 = ~(w7977 | w7978);
assign w7979 = v2395;
assign w7980 = ~w3124 & w4913;
assign w7981 = w7979 & ~w7980;
assign w7982 = (~w6641 & w30143) | (~w6641 & w30144) | (w30143 & w30144);
assign w7983 = (w6641 & w30145) | (w6641 & w30146) | (w30145 & w30146);
assign v2396 = ~(w7982 | w7983);
assign w7984 = v2396;
assign v2397 = ~(w7976 | w7984);
assign w7985 = v2397;
assign w7986 = w10 & ~w3332;
assign w7987 = w4764 & ~w7309;
assign w7988 = (w4913 & ~w3261) | (w4913 & w30147) | (~w3261 & w30147);
assign w7989 = (w4836 & ~w3331) | (w4836 & w30148) | (~w3331 & w30148);
assign v2398 = ~(w7988 | w7989);
assign w7990 = v2398;
assign w7991 = ~w7987 & w7990;
assign w7992 = ~w7987 & w30149;
assign w7993 = ~w3211 & w4913;
assign w7994 = (w4836 & ~w3261) | (w4836 & w30315) | (~w3261 & w30315);
assign w7995 = (w4763 & ~w3331) | (w4763 & w30316) | (~w3331 & w30316);
assign v2399 = ~(w7994 | w7995);
assign w7996 = v2399;
assign w7997 = (~w6676 & w30150) | (~w6676 & w30151) | (w30150 & w30151);
assign w7998 = w7992 & w7997;
assign w7999 = w7630 & w7998;
assign v2400 = ~(w7630 | w7998);
assign w8000 = v2400;
assign v2401 = ~(w7999 | w8000);
assign w8001 = v2401;
assign w8002 = (w4836 & ~w3210) | (w4836 & w30487) | (~w3210 & w30487);
assign w8003 = (w4763 & ~w3261) | (w4763 & w30488) | (~w3261 & w30488);
assign v2402 = ~(w8002 | w8003);
assign w8004 = v2402;
assign w8005 = ~w3162 & w4913;
assign w8006 = w8004 & ~w8005;
assign w8007 = (~w6735 & w30317) | (~w6735 & w30318) | (w30317 & w30318);
assign w8008 = (w6735 & w30319) | (w6735 & w30320) | (w30319 & w30320);
assign v2403 = ~(w8007 | w8008);
assign w8009 = v2403;
assign w8010 = w8001 & ~w8009;
assign w8011 = (~w7999 & ~w8001) | (~w7999 & w30321) | (~w8001 & w30321);
assign w8012 = w7976 & w7984;
assign v2404 = ~(w7985 | w8012);
assign w8013 = v2404;
assign w8014 = ~w8011 & w8013;
assign w8015 = (~w7985 & ~w8013) | (~w7985 & w30322) | (~w8013 & w30322);
assign w8016 = w7967 & ~w7971;
assign v2405 = ~(w7972 | w8016);
assign w8017 = v2405;
assign w8018 = ~w8015 & w8017;
assign v2406 = ~(w7972 | w8018);
assign w8019 = v2406;
assign w8020 = ~w7950 & w7958;
assign v2407 = ~(w7959 | w8020);
assign w8021 = v2407;
assign w8022 = ~w8019 & w8021;
assign w8023 = (~w7959 & w8019) | (~w7959 & w30489) | (w8019 & w30489);
assign w8024 = ~w7938 & w7947;
assign v2408 = ~(w7948 | w8024);
assign w8025 = v2408;
assign w8026 = ~w8023 & w8025;
assign v2409 = ~(w7948 | w8026);
assign w8027 = v2409;
assign w8028 = ~w7925 & w7935;
assign v2410 = ~(w7936 | w8028);
assign w8029 = v2410;
assign w8030 = ~w8027 & w8029;
assign w8031 = (~w7936 & w8027) | (~w7936 & w30606) | (w8027 & w30606);
assign v2411 = ~(w7912 | w7922);
assign w8032 = v2411;
assign v2412 = ~(w7923 | w8032);
assign w8033 = v2412;
assign w8034 = ~w8031 & w8033;
assign v2413 = ~(w7923 | w8034);
assign w8035 = v2413;
assign w8036 = ~w7899 & w7909;
assign v2414 = ~(w7910 | w8036);
assign w8037 = v2414;
assign w8038 = ~w8035 & w8037;
assign w8039 = (~w7910 & w8035) | (~w7910 & w30802) | (w8035 & w30802);
assign w8040 = ~w7886 & w7896;
assign v2415 = ~(w7897 | w8040);
assign w8041 = v2415;
assign w8042 = ~w8039 & w8041;
assign v2416 = ~(w7897 | w8042);
assign w8043 = v2416;
assign v2417 = ~(w7873 | w7883);
assign w8044 = v2417;
assign v2418 = ~(w7884 | w8044);
assign w8045 = v2418;
assign w8046 = ~w8043 & w8045;
assign w8047 = (~w7884 & w8043) | (~w7884 & w31023) | (w8043 & w31023);
assign v2419 = ~(w7860 | w7870);
assign w8048 = v2419;
assign v2420 = ~(w7871 | w8048);
assign w8049 = v2420;
assign w8050 = ~w8047 & w8049;
assign v2421 = ~(w7871 | w8050);
assign w8051 = v2421;
assign v2422 = ~(w7847 | w7857);
assign w8052 = v2422;
assign v2423 = ~(w7858 | w8052);
assign w8053 = v2423;
assign w8054 = ~w8051 & w8053;
assign w8055 = (~w7858 & w8051) | (~w7858 & w31172) | (w8051 & w31172);
assign w8056 = ~w7834 & w7844;
assign v2424 = ~(w7845 | w8056);
assign w8057 = v2424;
assign w8058 = ~w8055 & w8057;
assign v2425 = ~(w7845 | w8058);
assign w8059 = v2425;
assign v2426 = ~(w7821 | w7831);
assign w8060 = v2426;
assign v2427 = ~(w7832 | w8060);
assign w8061 = v2427;
assign w8062 = ~w8059 & w8061;
assign v2428 = ~(w7832 | w8062);
assign w8063 = v2428;
assign v2429 = ~(w7699 | w7709);
assign w8064 = v2429;
assign v2430 = ~(w7710 | w8064);
assign w8065 = v2430;
assign w8066 = ~w8063 & w8065;
assign w8067 = w8063 & ~w8065;
assign v2431 = ~(w8066 | w8067);
assign w8068 = v2431;
assign w8069 = ~w2202 & w5113;
assign w8070 = w5049 & w5114;
assign w8071 = ~w2089 & w5531;
assign w8072 = ~w2038 & w5610;
assign v2432 = ~(w8071 | w8072);
assign w8073 = v2432;
assign w8074 = ~w8070 & w8073;
assign w8075 = ~w8069 & w8074;
assign w8076 = pi20 & w8075;
assign v2433 = ~(pi20 | w8075);
assign w8077 = v2433;
assign v2434 = ~(w8076 | w8077);
assign w8078 = v2434;
assign w8079 = w8068 & ~w8078;
assign v2435 = ~(w8066 | w8079);
assign w8080 = v2435;
assign w8081 = w7819 & ~w8080;
assign w8082 = ~w7819 & w8080;
assign v2436 = ~(w8081 | w8082);
assign w8083 = v2436;
assign w8084 = w4520 & w5765;
assign w8085 = ~w1795 & w5983;
assign w8086 = ~w1674 & w6236;
assign w8087 = ~w1860 & w5764;
assign v2437 = ~(w8086 | w8087);
assign w8088 = v2437;
assign w8089 = ~w8085 & w8088;
assign w8090 = ~w8084 & w8089;
assign w8091 = pi17 & ~w8090;
assign w8092 = ~pi17 & w8090;
assign v2438 = ~(w8091 | w8092);
assign w8093 = v2438;
assign w8094 = w8083 & w8093;
assign v2439 = ~(w8081 | w8094);
assign w8095 = v2439;
assign w8096 = w7817 & ~w8095;
assign w8097 = ~w7817 & w8095;
assign v2440 = ~(w8096 | w8097);
assign w8098 = v2440;
assign w8099 = w3843 & w6389;
assign w8100 = ~w1387 & w6871;
assign w8101 = ~w3666 & w7004;
assign w8102 = ~w1496 & w6388;
assign v2441 = ~(w8101 | w8102);
assign w8103 = v2441;
assign w8104 = ~w8100 & w8103;
assign w8105 = ~w8099 & w8104;
assign w8106 = pi14 & ~w8105;
assign w8107 = ~pi14 & w8105;
assign v2442 = ~(w8106 | w8107);
assign w8108 = v2442;
assign w8109 = w8098 & w8108;
assign v2443 = ~(w8096 | w8109);
assign w8110 = v2443;
assign v2444 = ~(w7804 | w7814);
assign w8111 = v2444;
assign v2445 = ~(w7815 | w8111);
assign w8112 = v2445;
assign w8113 = ~w8110 & w8112;
assign v2446 = ~(w7815 | w8113);
assign w8114 = v2446;
assign w8115 = w7802 & ~w8114;
assign w8116 = ~w7802 & w8114;
assign v2447 = ~(w8115 | w8116);
assign w8117 = v2447;
assign w8118 = w4405 & w7178;
assign w8119 = ~w4035 & w7765;
assign w8120 = ~w3920 & w7177;
assign w8121 = ~w4134 & w7466;
assign v2448 = ~(w8120 | w8121);
assign w8122 = v2448;
assign w8123 = ~w8119 & w8122;
assign w8124 = ~w8118 & w8123;
assign w8125 = pi11 & ~w8124;
assign w8126 = ~pi11 & w8124;
assign v2449 = ~(w8125 | w8126);
assign w8127 = v2449;
assign w8128 = w8117 & w8127;
assign v2450 = ~(w8115 | w8128);
assign w8129 = v2450;
assign w8130 = ~pi07 & pi08;
assign w8131 = pi07 & ~pi08;
assign v2451 = ~(w8130 | w8131);
assign w8132 = v2451;
assign v2452 = ~(pi06 | pi07);
assign w8133 = v2452;
assign w8134 = pi06 & pi07;
assign v2453 = ~(w8133 | w8134);
assign w8135 = v2453;
assign v2454 = ~(pi05 | pi06);
assign w8136 = v2454;
assign w8137 = pi05 & pi06;
assign v2455 = ~(w8136 | w8137);
assign w8138 = v2455;
assign v2456 = ~(w8135 | w8138);
assign w8139 = v2456;
assign w8140 = ~w8132 & w8139;
assign w8141 = ~w8132 & w8138;
assign w8142 = ~w4422 & w8141;
assign v2457 = ~(w8140 | w8142);
assign w8143 = v2457;
assign v2458 = ~(w4191 | w8143);
assign w8144 = v2458;
assign w8145 = ~pi08 & w8144;
assign w8146 = pi08 & ~w8144;
assign v2459 = ~(w8145 | w8146);
assign w8147 = v2459;
assign v2460 = ~(w8129 | w8147);
assign w8148 = v2460;
assign v2461 = ~(w7763 | w7774);
assign w8149 = v2461;
assign v2462 = ~(w7775 | w8149);
assign w8150 = v2462;
assign w8151 = w8129 & w8147;
assign v2463 = ~(w8148 | w8151);
assign w8152 = v2463;
assign w8153 = w8150 & w8152;
assign v2464 = ~(w8148 | w8153);
assign w8154 = v2464;
assign w8155 = w7800 & ~w8154;
assign w8156 = ~w7800 & w8154;
assign v2465 = ~(w8155 | w8156);
assign w8157 = v2465;
assign v2466 = ~(w8150 | w8152);
assign w8158 = v2466;
assign v2467 = ~(w8153 | w8158);
assign w8159 = v2467;
assign v2468 = ~(w8098 | w8108);
assign w8160 = v2468;
assign v2469 = ~(w8109 | w8160);
assign w8161 = v2469;
assign v2470 = ~(w8083 | w8093);
assign w8162 = v2470;
assign v2471 = ~(w8094 | w8162);
assign w8163 = v2471;
assign w8164 = w8059 & ~w8061;
assign v2472 = ~(w8062 | w8164);
assign w8165 = v2472;
assign w8166 = w5033 & w5114;
assign w8167 = ~w2202 & w5531;
assign w8168 = ~w2089 & w5610;
assign v2473 = ~(w8167 | w8168);
assign w8169 = v2473;
assign w8170 = ~w2290 & w5113;
assign w8171 = w8169 & ~w8170;
assign w8172 = ~w8166 & w8171;
assign w8173 = ~pi20 & w8172;
assign w8174 = pi20 & ~w8172;
assign v2474 = ~(w8173 | w8174);
assign w8175 = v2474;
assign w8176 = w8165 & w8175;
assign w8177 = w8055 & ~w8057;
assign v2475 = ~(w8058 | w8177);
assign w8178 = v2475;
assign w8179 = w5114 & w5262;
assign w8180 = ~w2202 & w5610;
assign w8181 = ~w2339 & w5113;
assign w8182 = ~w2290 & w5531;
assign v2476 = ~(w8181 | w8182);
assign w8183 = v2476;
assign w8184 = ~w8180 & w8183;
assign w8185 = ~w8179 & w8184;
assign w8186 = pi20 & ~w8185;
assign w8187 = ~pi20 & w8185;
assign v2477 = ~(w8186 | w8187);
assign w8188 = v2477;
assign w8189 = w8178 & w8188;
assign w8190 = w8051 & ~w8053;
assign v2478 = ~(w8054 | w8190);
assign w8191 = v2478;
assign w8192 = ~w2290 & w5610;
assign w8193 = w5114 & w5280;
assign w8194 = ~w2339 & w5531;
assign w8195 = ~w2424 & w5113;
assign v2479 = ~(w8194 | w8195);
assign w8196 = v2479;
assign w8197 = ~w8193 & w8196;
assign w8198 = ~w8192 & w8197;
assign w8199 = pi20 & w8198;
assign v2480 = ~(pi20 | w8198);
assign w8200 = v2480;
assign v2481 = ~(w8199 | w8200);
assign w8201 = v2481;
assign w8202 = w8191 & ~w8201;
assign w8203 = w8047 & ~w8049;
assign v2482 = ~(w8050 | w8203);
assign w8204 = v2482;
assign w8205 = ~w2492 & w5113;
assign w8206 = w5114 & w5665;
assign w8207 = ~w2424 & w5531;
assign w8208 = ~w2339 & w5610;
assign v2483 = ~(w8207 | w8208);
assign w8209 = v2483;
assign w8210 = ~w8206 & w8209;
assign w8211 = ~w8205 & w8210;
assign w8212 = pi20 & w8211;
assign v2484 = ~(pi20 | w8211);
assign w8213 = v2484;
assign v2485 = ~(w8212 | w8213);
assign w8214 = v2485;
assign w8215 = w8204 & ~w8214;
assign w8216 = w8043 & ~w8045;
assign v2486 = ~(w8046 | w8216);
assign w8217 = v2486;
assign w8218 = w5114 & w5449;
assign w8219 = ~w2424 & w5610;
assign w8220 = ~w2492 & w5531;
assign w8221 = ~w2568 & w5113;
assign v2487 = ~(w8220 | w8221);
assign w8222 = v2487;
assign w8223 = ~w8219 & w8222;
assign w8224 = ~w8218 & w8223;
assign w8225 = pi20 & ~w8224;
assign w8226 = ~pi20 & w8224;
assign v2488 = ~(w8225 | w8226);
assign w8227 = v2488;
assign w8228 = w8217 & w8227;
assign w8229 = w8039 & ~w8041;
assign v2489 = ~(w8042 | w8229);
assign w8230 = v2489;
assign w8231 = w5114 & w5898;
assign w8232 = ~w2568 & w5531;
assign w8233 = ~w2596 & w5113;
assign w8234 = ~w2492 & w5610;
assign v2490 = ~(w8233 | w8234);
assign w8235 = v2490;
assign w8236 = ~w8232 & w8235;
assign w8237 = ~w8231 & w8236;
assign w8238 = pi20 & ~w8237;
assign w8239 = ~pi20 & w8237;
assign v2491 = ~(w8238 | w8239);
assign w8240 = v2491;
assign w8241 = w8230 & w8240;
assign w8242 = w8035 & ~w8037;
assign v2492 = ~(w8038 | w8242);
assign w8243 = v2492;
assign w8244 = w5114 & w6031;
assign w8245 = ~w2568 & w5610;
assign w8246 = ~w2596 & w5531;
assign v2493 = ~(w8245 | w8246);
assign w8247 = v2493;
assign w8248 = ~w2669 & w5113;
assign w8249 = w8247 & ~w8248;
assign w8250 = ~w8244 & w8249;
assign w8251 = ~pi20 & w8250;
assign w8252 = pi20 & ~w8250;
assign v2494 = ~(w8251 | w8252);
assign w8253 = v2494;
assign w8254 = w8243 & w8253;
assign w8255 = w8031 & ~w8033;
assign v2495 = ~(w8034 | w8255);
assign w8256 = v2495;
assign w8257 = w5114 & w5880;
assign w8258 = ~w2669 & w5531;
assign w8259 = ~w2724 & w5113;
assign w8260 = ~w2596 & w5610;
assign v2496 = ~(w8259 | w8260);
assign w8261 = v2496;
assign w8262 = ~w8258 & w8261;
assign w8263 = ~w8257 & w8262;
assign w8264 = pi20 & ~w8263;
assign w8265 = ~pi20 & w8263;
assign v2497 = ~(w8264 | w8265);
assign w8266 = v2497;
assign w8267 = w8256 & w8266;
assign w8268 = w8027 & ~w8029;
assign v2498 = ~(w8030 | w8268);
assign w8269 = v2498;
assign w8270 = w5114 & w6148;
assign w8271 = ~w2724 & w5531;
assign w8272 = ~w2669 & w5610;
assign w8273 = ~w2811 & w5113;
assign v2499 = ~(w8272 | w8273);
assign w8274 = v2499;
assign w8275 = ~w8271 & w8274;
assign w8276 = ~w8270 & w8275;
assign w8277 = pi20 & ~w8276;
assign w8278 = ~pi20 & w8276;
assign v2500 = ~(w8277 | w8278);
assign w8279 = v2500;
assign w8280 = w8269 & w8279;
assign w8281 = w8023 & ~w8025;
assign v2501 = ~(w8026 | w8281);
assign w8282 = v2501;
assign w8283 = w5114 & ~w6447;
assign w8284 = ~w2846 & w5113;
assign w8285 = ~w2811 & w5531;
assign w8286 = ~w2724 & w5610;
assign v2502 = ~(w8285 | w8286);
assign w8287 = v2502;
assign w8288 = ~w8284 & w8287;
assign w8289 = ~w8283 & w8288;
assign w8290 = pi20 & ~w8289;
assign w8291 = ~pi20 & w8289;
assign v2503 = ~(w8290 | w8291);
assign w8292 = v2503;
assign w8293 = w8282 & w8292;
assign w8294 = w8019 & ~w8021;
assign v2504 = ~(w8022 | w8294);
assign w8295 = v2504;
assign w8296 = w5114 & w6459;
assign w8297 = ~w2811 & w5610;
assign w8298 = ~w2846 & w5531;
assign w8299 = ~w2937 & w5113;
assign v2505 = ~(w8298 | w8299);
assign w8300 = v2505;
assign w8301 = ~w8297 & w8300;
assign w8302 = ~w8296 & w8301;
assign w8303 = pi20 & ~w8302;
assign w8304 = ~pi20 & w8302;
assign v2506 = ~(w8303 | w8304);
assign w8305 = v2506;
assign w8306 = w8295 & w8305;
assign w8307 = w8015 & ~w8017;
assign v2507 = ~(w8018 | w8307);
assign w8308 = v2507;
assign w8309 = w5114 & w6130;
assign w8310 = ~w2846 & w5610;
assign w8311 = ~w2937 & w5531;
assign v2508 = ~(w8310 | w8311);
assign w8312 = v2508;
assign w8313 = ~w3000 & w5113;
assign w8314 = w8312 & ~w8313;
assign w8315 = ~w8309 & w8314;
assign w8316 = pi20 & w8315;
assign v2509 = ~(pi20 | w8315);
assign w8317 = v2509;
assign v2510 = ~(w8316 | w8317);
assign w8318 = v2510;
assign w8319 = w8308 & ~w8318;
assign w8320 = w8011 & ~w8013;
assign v2511 = ~(w8014 | w8320);
assign w8321 = v2511;
assign w8322 = ~w3000 & w5531;
assign w8323 = ~w2937 & w5610;
assign v2512 = ~(w8322 | w8323);
assign w8324 = v2512;
assign w8325 = ~w3068 & w5113;
assign w8326 = w8324 & ~w8325;
assign w8327 = (w8326 & w6505) | (w8326 & w30323) | (w6505 & w30323);
assign w8328 = pi20 & w8327;
assign v2513 = ~(pi20 | w8327);
assign w8329 = v2513;
assign v2514 = ~(w8328 | w8329);
assign w8330 = v2514;
assign w8331 = w8321 & ~w8330;
assign w8332 = ~w8001 & w8009;
assign v2515 = ~(w8010 | w8332);
assign w8333 = v2515;
assign w8334 = ~w3068 & w5531;
assign w8335 = ~w3124 & w5113;
assign w8336 = ~w3000 & w5610;
assign v2516 = ~(w8335 | w8336);
assign w8337 = v2516;
assign w8338 = ~w8334 & w8337;
assign w8339 = (w6551 & w30324) | (w6551 & w30325) | (w30324 & w30325);
assign w8340 = (~w6551 & w30326) | (~w6551 & w30327) | (w30326 & w30327);
assign v2517 = ~(w8339 | w8340);
assign w8341 = v2517;
assign w8342 = w8333 & w8341;
assign w8343 = ~w3124 & w5531;
assign w8344 = ~w3068 & w5610;
assign v2518 = ~(w8343 | w8344);
assign w8345 = v2518;
assign w8346 = ~w3162 & w5113;
assign w8347 = w8345 & ~w8346;
assign w8348 = (~w6603 & w30000) | (~w6603 & w30001) | (w30000 & w30001);
assign w8349 = (w6603 & w30002) | (w6603 & w30003) | (w30002 & w30003);
assign v2519 = ~(w8348 | w8349);
assign w8350 = v2519;
assign w8351 = pi23 & ~w7992;
assign w8352 = ~w7997 & w8351;
assign w8353 = w7997 & ~w8351;
assign v2520 = ~(w8352 | w8353);
assign w8354 = v2520;
assign w8355 = ~w8350 & w8354;
assign w8356 = pi23 & w7986;
assign v2521 = ~(w7991 | w8356);
assign w8357 = v2521;
assign w8358 = w7991 & w8356;
assign v2522 = ~(w8357 | w8358);
assign w8359 = v2522;
assign w8360 = ~w3162 & w5531;
assign w8361 = ~w3124 & w5610;
assign v2523 = ~(w8360 | w8361);
assign w8362 = v2523;
assign w8363 = ~w3211 & w5113;
assign w8364 = w8362 & ~w8363;
assign w8365 = (w6641 & w29832) | (w6641 & w29833) | (w29832 & w29833);
assign w8366 = (~w6641 & w29834) | (~w6641 & w29835) | (w29834 & w29835);
assign v2524 = ~(w8365 | w8366);
assign w8367 = v2524;
assign v2525 = ~(w8359 | w8367);
assign w8368 = v2525;
assign w8369 = ~w3262 & w5531;
assign w8370 = (w5610 & ~w3210) | (w5610 & w30004) | (~w3210 & w30004);
assign w8371 = (w5113 & ~w3331) | (w5113 & w30005) | (~w3331 & w30005);
assign v2526 = ~(w8370 | w8371);
assign w8372 = v2526;
assign w8373 = (~w6676 & w29836) | (~w6676 & w29837) | (w29836 & w29837);
assign w8374 = w912 & ~w3332;
assign w8375 = (w29838 & ~w3331) | (w29838 & w30006) | (~w3331 & w30006);
assign w8376 = w5114 & ~w7309;
assign w8377 = (w5531 & ~w3331) | (w5531 & w29839) | (~w3331 & w29839);
assign w8378 = (w5610 & ~w3261) | (w5610 & w29840) | (~w3261 & w29840);
assign v2527 = ~(w8377 | w8378);
assign w8379 = v2527;
assign w8380 = ~w8376 & w8379;
assign w8381 = ~w8376 & w29645;
assign w8382 = ~w8376 & w29841;
assign w8383 = w8373 & w8382;
assign w8384 = w7986 & w8383;
assign v2528 = ~(w7986 | w8383);
assign w8385 = v2528;
assign v2529 = ~(w8384 | w8385);
assign w8386 = v2529;
assign w8387 = ~w3162 & w5610;
assign w8388 = (w5113 & ~w3261) | (w5113 & w30153) | (~w3261 & w30153);
assign w8389 = (w5531 & ~w3210) | (w5531 & w30154) | (~w3210 & w30154);
assign v2530 = ~(w8388 | w8389);
assign w8390 = v2530;
assign w8391 = ~w8387 & w8390;
assign w8392 = (w6735 & w30007) | (w6735 & w30008) | (w30007 & w30008);
assign w8393 = (~w6735 & w30009) | (~w6735 & w30010) | (w30009 & w30010);
assign v2531 = ~(w8392 | w8393);
assign w8394 = v2531;
assign w8395 = w8386 & w8394;
assign w8396 = (~w8384 & ~w8386) | (~w8384 & w30011) | (~w8386 & w30011);
assign w8397 = w8359 & w8367;
assign v2532 = ~(w8368 | w8397);
assign w8398 = v2532;
assign w8399 = ~w8396 & w8398;
assign w8400 = (~w8368 & ~w8398) | (~w8368 & w30012) | (~w8398 & w30012);
assign w8401 = w8350 & ~w8354;
assign v2533 = ~(w8355 | w8401);
assign w8402 = v2533;
assign w8403 = ~w8400 & w8402;
assign v2534 = ~(w8355 | w8403);
assign w8404 = v2534;
assign v2535 = ~(w8333 | w8341);
assign w8405 = v2535;
assign v2536 = ~(w8342 | w8405);
assign w8406 = v2536;
assign w8407 = ~w8404 & w8406;
assign w8408 = (~w8342 & w8404) | (~w8342 & w30155) | (w8404 & w30155);
assign w8409 = ~w8321 & w8330;
assign v2537 = ~(w8331 | w8409);
assign w8410 = v2537;
assign w8411 = ~w8408 & w8410;
assign v2538 = ~(w8331 | w8411);
assign w8412 = v2538;
assign w8413 = ~w8308 & w8318;
assign v2539 = ~(w8319 | w8413);
assign w8414 = v2539;
assign w8415 = ~w8412 & w8414;
assign w8416 = (~w8319 & w8412) | (~w8319 & w30328) | (w8412 & w30328);
assign v2540 = ~(w8295 | w8305);
assign w8417 = v2540;
assign v2541 = ~(w8306 | w8417);
assign w8418 = v2541;
assign w8419 = ~w8416 & w8418;
assign v2542 = ~(w8306 | w8419);
assign w8420 = v2542;
assign v2543 = ~(w8282 | w8292);
assign w8421 = v2543;
assign v2544 = ~(w8293 | w8421);
assign w8422 = v2544;
assign w8423 = ~w8420 & w8422;
assign w8424 = (~w8293 & w8420) | (~w8293 & w30490) | (w8420 & w30490);
assign v2545 = ~(w8269 | w8279);
assign w8425 = v2545;
assign v2546 = ~(w8280 | w8425);
assign w8426 = v2546;
assign w8427 = ~w8424 & w8426;
assign v2547 = ~(w8280 | w8427);
assign w8428 = v2547;
assign v2548 = ~(w8256 | w8266);
assign w8429 = v2548;
assign v2549 = ~(w8267 | w8429);
assign w8430 = v2549;
assign w8431 = ~w8428 & w8430;
assign w8432 = (~w8267 & w8428) | (~w8267 & w30607) | (w8428 & w30607);
assign v2550 = ~(w8243 | w8253);
assign w8433 = v2550;
assign v2551 = ~(w8254 | w8433);
assign w8434 = v2551;
assign w8435 = ~w8432 & w8434;
assign v2552 = ~(w8254 | w8435);
assign w8436 = v2552;
assign v2553 = ~(w8230 | w8240);
assign w8437 = v2553;
assign v2554 = ~(w8241 | w8437);
assign w8438 = v2554;
assign w8439 = ~w8436 & w8438;
assign w8440 = (~w8241 & w8436) | (~w8241 & w30803) | (w8436 & w30803);
assign v2555 = ~(w8217 | w8227);
assign w8441 = v2555;
assign v2556 = ~(w8228 | w8441);
assign w8442 = v2556;
assign w8443 = ~w8440 & w8442;
assign v2557 = ~(w8228 | w8443);
assign w8444 = v2557;
assign w8445 = ~w8204 & w8214;
assign v2558 = ~(w8215 | w8445);
assign w8446 = v2558;
assign w8447 = ~w8444 & w8446;
assign w8448 = (~w8215 & w8444) | (~w8215 & w31024) | (w8444 & w31024);
assign w8449 = ~w8191 & w8201;
assign v2559 = ~(w8202 | w8449);
assign w8450 = v2559;
assign w8451 = ~w8448 & w8450;
assign v2560 = ~(w8202 | w8451);
assign w8452 = v2560;
assign v2561 = ~(w8178 | w8188);
assign w8453 = v2561;
assign v2562 = ~(w8189 | w8453);
assign w8454 = v2562;
assign w8455 = ~w8452 & w8454;
assign w8456 = (~w8189 & w8452) | (~w8189 & w31173) | (w8452 & w31173);
assign v2563 = ~(w8165 | w8175);
assign w8457 = v2563;
assign v2564 = ~(w8176 | w8457);
assign w8458 = v2564;
assign w8459 = ~w8456 & w8458;
assign v2565 = ~(w8176 | w8459);
assign w8460 = v2565;
assign w8461 = ~w8068 & w8078;
assign v2566 = ~(w8079 | w8461);
assign w8462 = v2566;
assign w8463 = w8460 & ~w8462;
assign w8464 = ~w8460 & w8462;
assign w8465 = w4538 & w5765;
assign w8466 = ~w1860 & w5983;
assign w8467 = ~w1942 & w5764;
assign v2567 = ~(w8466 | w8467);
assign w8468 = v2567;
assign w8469 = ~w1795 & w6236;
assign w8470 = w8468 & ~w8469;
assign w8471 = ~w8465 & w8470;
assign w8472 = pi17 & ~w8471;
assign w8473 = ~pi17 & w8471;
assign v2568 = ~(w8472 | w8473);
assign w8474 = v2568;
assign v2569 = ~(w8464 | w8474);
assign w8475 = v2569;
assign v2570 = ~(w8463 | w8475);
assign w8476 = v2570;
assign w8477 = w8163 & w8476;
assign v2571 = ~(w8163 | w8476);
assign w8478 = v2571;
assign v2572 = ~(w8477 | w8478);
assign w8479 = v2572;
assign w8480 = w3397 & w6389;
assign w8481 = ~w1387 & w7004;
assign w8482 = ~w1496 & w6871;
assign v2573 = ~(w8481 | w8482);
assign w8483 = v2573;
assign w8484 = ~w1609 & w6388;
assign w8485 = w8483 & ~w8484;
assign w8486 = ~w8480 & w8485;
assign w8487 = pi14 & ~w8486;
assign w8488 = ~pi14 & w8486;
assign v2574 = ~(w8487 | w8488);
assign w8489 = v2574;
assign w8490 = w8479 & w8489;
assign v2575 = ~(w8477 | w8490);
assign w8491 = v2575;
assign w8492 = w8161 & ~w8491;
assign w8493 = ~w8161 & w8491;
assign v2576 = ~(w8492 | w8493);
assign w8494 = v2576;
assign w8495 = ~w3928 & w7178;
assign w8496 = ~w3752 & w7466;
assign w8497 = ~w3587 & w7177;
assign w8498 = ~w3920 & w7765;
assign v2577 = ~(w8497 | w8498);
assign w8499 = v2577;
assign w8500 = ~w8496 & w8499;
assign w8501 = ~w8495 & w8500;
assign w8502 = pi11 & ~w8501;
assign w8503 = ~pi11 & w8501;
assign v2578 = ~(w8502 | w8503);
assign w8504 = v2578;
assign w8505 = w8494 & w8504;
assign v2579 = ~(w8492 | w8505);
assign w8506 = v2579;
assign w8507 = w4309 & w7178;
assign w8508 = ~w3920 & w7466;
assign w8509 = ~w3752 & w7177;
assign w8510 = ~w4134 & w7765;
assign v2580 = ~(w8509 | w8510);
assign w8511 = v2580;
assign w8512 = ~w8508 & w8511;
assign w8513 = ~w8507 & w8512;
assign w8514 = pi11 & ~w8513;
assign w8515 = ~pi11 & w8513;
assign v2581 = ~(w8514 | w8515);
assign w8516 = v2581;
assign w8517 = ~w8506 & w8516;
assign w8518 = w8110 & ~w8112;
assign v2582 = ~(w8113 | w8518);
assign w8519 = v2582;
assign w8520 = w8506 & ~w8516;
assign v2583 = ~(w8517 | w8520);
assign w8521 = v2583;
assign w8522 = w8519 & w8521;
assign v2584 = ~(w8517 | w8522);
assign w8523 = v2584;
assign w8524 = w4425 & w8141;
assign w8525 = ~w4082 & w8140;
assign w8526 = w8135 & ~w8138;
assign w8527 = ~w4191 & w8526;
assign v2585 = ~(w8525 | w8527);
assign w8528 = v2585;
assign w8529 = ~w8524 & w8528;
assign w8530 = ~pi08 & w8529;
assign w8531 = pi08 & ~w8529;
assign v2586 = ~(w8530 | w8531);
assign w8532 = v2586;
assign w8533 = ~w8523 & w8532;
assign v2587 = ~(w8117 | w8127);
assign w8534 = v2587;
assign v2588 = ~(w8128 | w8534);
assign w8535 = v2588;
assign w8536 = w8523 & ~w8532;
assign v2589 = ~(w8533 | w8536);
assign w8537 = v2589;
assign w8538 = w8535 & w8537;
assign v2590 = ~(w8533 | w8538);
assign w8539 = v2590;
assign w8540 = w8159 & ~w8539;
assign w8541 = ~w8159 & w8539;
assign v2591 = ~(w8494 | w8504);
assign w8542 = v2591;
assign v2592 = ~(w8505 | w8542);
assign w8543 = v2592;
assign v2593 = ~(w8479 | w8489);
assign w8544 = v2593;
assign v2594 = ~(w8490 | w8544);
assign w8545 = v2594;
assign w8546 = ~w3510 & w6389;
assign w8547 = ~w1609 & w6871;
assign w8548 = ~w1496 & w7004;
assign v2595 = ~(w8547 | w8548);
assign w8549 = v2595;
assign w8550 = ~w1674 & w6388;
assign w8551 = w8549 & ~w8550;
assign w8552 = ~w8546 & w8551;
assign w8553 = ~pi14 & w8552;
assign w8554 = pi14 & ~w8552;
assign v2596 = ~(w8553 | w8554);
assign w8555 = v2596;
assign v2597 = ~(w8463 | w8464);
assign w8556 = v2597;
assign w8557 = ~w8474 & w8556;
assign w8558 = w8474 & ~w8556;
assign v2598 = ~(w8557 | w8558);
assign w8559 = v2598;
assign w8560 = w8555 & ~w8559;
assign w8561 = ~w8555 & w8559;
assign v2599 = ~(w8560 | w8561);
assign w8562 = v2599;
assign w8563 = w4854 & w5765;
assign w8564 = ~w1860 & w6236;
assign w8565 = ~w2038 & w5764;
assign w8566 = ~w1942 & w5983;
assign v2600 = ~(w8565 | w8566);
assign w8567 = v2600;
assign w8568 = ~w8564 & w8567;
assign w8569 = ~w8563 & w8568;
assign w8570 = pi17 & ~w8569;
assign w8571 = ~pi17 & w8569;
assign v2601 = ~(w8570 | w8571);
assign w8572 = v2601;
assign w8573 = w8456 & ~w8458;
assign v2602 = ~(w8459 | w8573);
assign w8574 = v2602;
assign v2603 = ~(w8572 | w8574);
assign w8575 = v2603;
assign w8576 = w8572 & w8574;
assign w8577 = w8452 & ~w8454;
assign v2604 = ~(w8455 | w8577);
assign w8578 = v2604;
assign w8579 = w4702 & w5765;
assign w8580 = ~w2089 & w5764;
assign w8581 = ~w2038 & w5983;
assign v2605 = ~(w8580 | w8581);
assign w8582 = v2605;
assign w8583 = ~w1942 & w6236;
assign w8584 = w8582 & ~w8583;
assign w8585 = ~w8579 & w8584;
assign w8586 = ~pi17 & w8585;
assign w8587 = pi17 & ~w8585;
assign v2606 = ~(w8586 | w8587);
assign w8588 = v2606;
assign w8589 = w8578 & w8588;
assign v2607 = ~(w8578 | w8588);
assign w8590 = v2607;
assign w8591 = w8448 & ~w8450;
assign v2608 = ~(w8451 | w8591);
assign w8592 = v2608;
assign w8593 = w5049 & w5765;
assign w8594 = ~w2202 & w5764;
assign w8595 = ~w2089 & w5983;
assign w8596 = ~w2038 & w6236;
assign v2609 = ~(w8595 | w8596);
assign w8597 = v2609;
assign w8598 = ~w8594 & w8597;
assign w8599 = ~w8593 & w8598;
assign w8600 = pi17 & ~w8599;
assign w8601 = ~pi17 & w8599;
assign v2610 = ~(w8600 | w8601);
assign w8602 = v2610;
assign v2611 = ~(w8592 | w8602);
assign w8603 = v2611;
assign w8604 = w8592 & w8602;
assign w8605 = w8444 & ~w8446;
assign v2612 = ~(w8447 | w8605);
assign w8606 = v2612;
assign w8607 = w5033 & w5765;
assign w8608 = ~w2290 & w5764;
assign w8609 = ~w2089 & w6236;
assign w8610 = ~w2202 & w5983;
assign v2613 = ~(w8609 | w8610);
assign w8611 = v2613;
assign w8612 = ~w8608 & w8611;
assign w8613 = ~w8607 & w8612;
assign w8614 = pi17 & ~w8613;
assign w8615 = ~pi17 & w8613;
assign v2614 = ~(w8614 | w8615);
assign w8616 = v2614;
assign w8617 = w8606 & w8616;
assign w8618 = w5262 & w5765;
assign w8619 = ~w2202 & w6236;
assign w8620 = ~w2339 & w5764;
assign w8621 = ~w2290 & w5983;
assign v2615 = ~(w8620 | w8621);
assign w8622 = v2615;
assign w8623 = ~w8619 & w8622;
assign w8624 = ~w8618 & w8623;
assign w8625 = pi17 & ~w8624;
assign w8626 = ~pi17 & w8624;
assign v2616 = ~(w8625 | w8626);
assign w8627 = v2616;
assign w8628 = w8440 & ~w8442;
assign v2617 = ~(w8443 | w8628);
assign w8629 = v2617;
assign w8630 = w8627 & w8629;
assign w8631 = w8436 & ~w8438;
assign v2618 = ~(w8439 | w8631);
assign w8632 = v2618;
assign w8633 = w5280 & w5765;
assign w8634 = ~w2290 & w6236;
assign w8635 = ~w2339 & w5983;
assign w8636 = ~w2424 & w5764;
assign v2619 = ~(w8635 | w8636);
assign w8637 = v2619;
assign w8638 = ~w8634 & w8637;
assign w8639 = ~w8633 & w8638;
assign w8640 = pi17 & ~w8639;
assign w8641 = ~pi17 & w8639;
assign v2620 = ~(w8640 | w8641);
assign w8642 = v2620;
assign w8643 = w8632 & w8642;
assign w8644 = w8432 & ~w8434;
assign v2621 = ~(w8435 | w8644);
assign w8645 = v2621;
assign w8646 = ~w2492 & w5764;
assign w8647 = w5665 & w5765;
assign w8648 = ~w2424 & w5983;
assign w8649 = ~w2339 & w6236;
assign v2622 = ~(w8648 | w8649);
assign w8650 = v2622;
assign w8651 = ~w8647 & w8650;
assign w8652 = ~w8646 & w8651;
assign w8653 = pi17 & w8652;
assign v2623 = ~(pi17 | w8652);
assign w8654 = v2623;
assign v2624 = ~(w8653 | w8654);
assign w8655 = v2624;
assign w8656 = w8645 & ~w8655;
assign w8657 = w8428 & ~w8430;
assign v2625 = ~(w8431 | w8657);
assign w8658 = v2625;
assign w8659 = w5449 & w5765;
assign w8660 = ~w2424 & w6236;
assign w8661 = ~w2492 & w5983;
assign w8662 = ~w2568 & w5764;
assign v2626 = ~(w8661 | w8662);
assign w8663 = v2626;
assign w8664 = ~w8660 & w8663;
assign w8665 = ~w8659 & w8664;
assign w8666 = pi17 & ~w8665;
assign w8667 = ~pi17 & w8665;
assign v2627 = ~(w8666 | w8667);
assign w8668 = v2627;
assign w8669 = w8658 & w8668;
assign w8670 = w8424 & ~w8426;
assign v2628 = ~(w8427 | w8670);
assign w8671 = v2628;
assign w8672 = w5765 & w5898;
assign w8673 = ~w2568 & w5983;
assign w8674 = ~w2596 & w5764;
assign w8675 = ~w2492 & w6236;
assign v2629 = ~(w8674 | w8675);
assign w8676 = v2629;
assign w8677 = ~w8673 & w8676;
assign w8678 = ~w8672 & w8677;
assign w8679 = pi17 & ~w8678;
assign w8680 = ~pi17 & w8678;
assign v2630 = ~(w8679 | w8680);
assign w8681 = v2630;
assign w8682 = w8671 & w8681;
assign w8683 = w8420 & ~w8422;
assign v2631 = ~(w8423 | w8683);
assign w8684 = v2631;
assign w8685 = w5765 & w6031;
assign w8686 = ~w2669 & w5764;
assign w8687 = ~w2596 & w5983;
assign w8688 = ~w2568 & w6236;
assign v2632 = ~(w8687 | w8688);
assign w8689 = v2632;
assign w8690 = ~w8686 & w8689;
assign w8691 = ~w8685 & w8690;
assign w8692 = pi17 & ~w8691;
assign w8693 = ~pi17 & w8691;
assign v2633 = ~(w8692 | w8693);
assign w8694 = v2633;
assign w8695 = w8684 & w8694;
assign v2634 = ~(w8684 | w8694);
assign w8696 = v2634;
assign v2635 = ~(w8695 | w8696);
assign w8697 = v2635;
assign w8698 = w8416 & ~w8418;
assign v2636 = ~(w8419 | w8698);
assign w8699 = v2636;
assign w8700 = w5765 & w5880;
assign w8701 = ~w2669 & w5983;
assign w8702 = ~w2724 & w5764;
assign w8703 = ~w2596 & w6236;
assign v2637 = ~(w8702 | w8703);
assign w8704 = v2637;
assign w8705 = ~w8701 & w8704;
assign w8706 = ~w8700 & w8705;
assign w8707 = pi17 & ~w8706;
assign w8708 = ~pi17 & w8706;
assign v2638 = ~(w8707 | w8708);
assign w8709 = v2638;
assign w8710 = w8699 & w8709;
assign w8711 = w8412 & ~w8414;
assign v2639 = ~(w8415 | w8711);
assign w8712 = v2639;
assign w8713 = w5765 & w6148;
assign w8714 = ~w2811 & w5764;
assign w8715 = ~w2724 & w5983;
assign v2640 = ~(w8714 | w8715);
assign w8716 = v2640;
assign w8717 = ~w2669 & w6236;
assign w8718 = w8716 & ~w8717;
assign w8719 = ~w8713 & w8718;
assign w8720 = pi17 & w8719;
assign v2641 = ~(pi17 | w8719);
assign w8721 = v2641;
assign v2642 = ~(w8720 | w8721);
assign w8722 = v2642;
assign w8723 = w8712 & ~w8722;
assign w8724 = w8408 & ~w8410;
assign v2643 = ~(w8411 | w8724);
assign w8725 = v2643;
assign w8726 = ~w2846 & w5764;
assign w8727 = w5765 & ~w6447;
assign w8728 = ~w2811 & w5983;
assign w8729 = ~w2724 & w6236;
assign v2644 = ~(w8728 | w8729);
assign w8730 = v2644;
assign w8731 = ~w8727 & w8730;
assign w8732 = ~w8726 & w8731;
assign w8733 = pi17 & w8732;
assign v2645 = ~(pi17 | w8732);
assign w8734 = v2645;
assign v2646 = ~(w8733 | w8734);
assign w8735 = v2646;
assign w8736 = w8725 & ~w8735;
assign w8737 = w8404 & ~w8406;
assign v2647 = ~(w8407 | w8737);
assign w8738 = v2647;
assign w8739 = ~w2937 & w5764;
assign w8740 = w5765 & w6459;
assign w8741 = ~w2811 & w6236;
assign w8742 = ~w2846 & w5983;
assign v2648 = ~(w8741 | w8742);
assign w8743 = v2648;
assign w8744 = ~w8740 & w8743;
assign w8745 = ~w8739 & w8744;
assign w8746 = pi17 & w8745;
assign v2649 = ~(pi17 | w8745);
assign w8747 = v2649;
assign v2650 = ~(w8746 | w8747);
assign w8748 = v2650;
assign w8749 = w8738 & ~w8748;
assign w8750 = w8400 & ~w8402;
assign v2651 = ~(w8403 | w8750);
assign w8751 = v2651;
assign w8752 = w5765 & w6130;
assign w8753 = ~w2846 & w6236;
assign w8754 = ~w2937 & w5983;
assign v2652 = ~(w8753 | w8754);
assign w8755 = v2652;
assign w8756 = ~w3000 & w5764;
assign w8757 = w8755 & ~w8756;
assign w8758 = ~w8752 & w8757;
assign w8759 = pi17 & w8758;
assign v2653 = ~(pi17 | w8758);
assign w8760 = v2653;
assign v2654 = ~(w8759 | w8760);
assign w8761 = v2654;
assign w8762 = w8751 & ~w8761;
assign w8763 = w8396 & ~w8398;
assign v2655 = ~(w8399 | w8763);
assign w8764 = v2655;
assign w8765 = ~w3000 & w5983;
assign w8766 = ~w2937 & w6236;
assign v2656 = ~(w8765 | w8766);
assign w8767 = v2656;
assign w8768 = ~w3068 & w5764;
assign w8769 = w8767 & ~w8768;
assign w8770 = (w8769 & w6505) | (w8769 & w30013) | (w6505 & w30013);
assign w8771 = pi17 & w8770;
assign v2657 = ~(pi17 | w8770);
assign w8772 = v2657;
assign v2658 = ~(w8771 | w8772);
assign w8773 = v2658;
assign w8774 = w8764 & ~w8773;
assign v2659 = ~(w8386 | w8394);
assign w8775 = v2659;
assign v2660 = ~(w8395 | w8775);
assign w8776 = v2660;
assign w8777 = ~w3124 & w5764;
assign w8778 = ~w3068 & w5983;
assign v2661 = ~(w8777 | w8778);
assign w8779 = v2661;
assign w8780 = ~w3000 & w6236;
assign w8781 = w8779 & ~w8780;
assign w8782 = (w6551 & w30014) | (w6551 & w30015) | (w30014 & w30015);
assign w8783 = (~w6551 & w30016) | (~w6551 & w30017) | (w30016 & w30017);
assign v2662 = ~(w8782 | w8783);
assign w8784 = v2662;
assign w8785 = w8776 & ~w8784;
assign w8786 = ~w3124 & w5983;
assign w8787 = ~w3068 & w6236;
assign v2663 = ~(w8786 | w8787);
assign w8788 = v2663;
assign w8789 = ~w3162 & w5764;
assign w8790 = w8788 & ~w8789;
assign w8791 = (w6603 & w29646) | (w6603 & w29647) | (w29646 & w29647);
assign w8792 = (~w6603 & w29648) | (~w6603 & w29649) | (w29648 & w29649);
assign v2664 = ~(w8791 | w8792);
assign w8793 = v2664;
assign w8794 = pi20 & ~w8381;
assign w8795 = ~w8373 & w8794;
assign w8796 = w8373 & ~w8794;
assign v2665 = ~(w8795 | w8796);
assign w8797 = v2665;
assign w8798 = ~w8793 & w8797;
assign w8799 = w8375 & ~w8380;
assign v2666 = ~(w8381 | w8799);
assign w8800 = v2666;
assign w8801 = ~w3124 & w6236;
assign w8802 = ~w3162 & w5983;
assign v2667 = ~(w8801 | w8802);
assign w8803 = v2667;
assign w8804 = ~w3211 & w5764;
assign w8805 = w8803 & ~w8804;
assign w8806 = (w6641 & w29466) | (w6641 & w29467) | (w29466 & w29467);
assign w8807 = (~w6641 & w29468) | (~w6641 & w29469) | (w29468 & w29469);
assign v2668 = ~(w8806 | w8807);
assign w8808 = v2668;
assign w8809 = w8800 & ~w8808;
assign w8810 = w5765 & w6676;
assign w8811 = ~w3211 & w6236;
assign w8812 = ~w3332 & w5764;
assign w8813 = ~w3262 & w5983;
assign v2669 = ~(w8812 | w8813);
assign w8814 = v2669;
assign w8815 = ~w8811 & w8814;
assign w8816 = ~w8810 & w8815;
assign w8817 = (w5756 & ~w3331) | (w5756 & w29470) | (~w3331 & w29470);
assign w8818 = (~w3331 & w29650) | (~w3331 & w29651) | (w29650 & w29651);
assign w8819 = w5765 & ~w7309;
assign w8820 = (w6236 & ~w3261) | (w6236 & w29471) | (~w3261 & w29471);
assign w8821 = (w5983 & ~w3331) | (w5983 & w29472) | (~w3331 & w29472);
assign v2670 = ~(w8820 | w8821);
assign w8822 = v2670;
assign w8823 = ~w8819 & w8822;
assign w8824 = ~w8819 & w29246;
assign w8825 = w8816 & w29474;
assign w8826 = (~w8374 & ~w8816) | (~w8374 & w29475) | (~w8816 & w29475);
assign v2671 = ~(w8825 | w8826);
assign w8827 = v2671;
assign w8828 = ~w3162 & w6236;
assign w8829 = (w5764 & ~w3261) | (w5764 & w29843) | (~w3261 & w29843);
assign w8830 = (w5983 & ~w3210) | (w5983 & w29844) | (~w3210 & w29844);
assign v2672 = ~(w8829 | w8830);
assign w8831 = v2672;
assign w8832 = ~w8828 & w8831;
assign w8833 = (w6735 & w29652) | (w6735 & w29653) | (w29652 & w29653);
assign w8834 = (~w6735 & w29654) | (~w6735 & w29655) | (w29654 & w29655);
assign v2673 = ~(w8833 | w8834);
assign w8835 = v2673;
assign w8836 = w8827 & w8835;
assign w8837 = (~w8825 & ~w8827) | (~w8825 & w29656) | (~w8827 & w29656);
assign w8838 = ~w8800 & w8808;
assign v2674 = ~(w8809 | w8838);
assign w8839 = v2674;
assign w8840 = ~w8837 & w8839;
assign w8841 = (~w8809 & ~w8839) | (~w8809 & w29657) | (~w8839 & w29657);
assign w8842 = w8793 & ~w8797;
assign v2675 = ~(w8798 | w8842);
assign w8843 = v2675;
assign w8844 = ~w8841 & w8843;
assign v2676 = ~(w8798 | w8844);
assign w8845 = v2676;
assign w8846 = ~w8776 & w8784;
assign v2677 = ~(w8785 | w8846);
assign w8847 = v2677;
assign w8848 = ~w8845 & w8847;
assign w8849 = (~w8785 & w8845) | (~w8785 & w29845) | (w8845 & w29845);
assign w8850 = ~w8764 & w8773;
assign v2678 = ~(w8774 | w8850);
assign w8851 = v2678;
assign w8852 = ~w8849 & w8851;
assign v2679 = ~(w8774 | w8852);
assign w8853 = v2679;
assign w8854 = ~w8751 & w8761;
assign v2680 = ~(w8762 | w8854);
assign w8855 = v2680;
assign w8856 = ~w8853 & w8855;
assign w8857 = (~w8762 & w8853) | (~w8762 & w30018) | (w8853 & w30018);
assign w8858 = ~w8738 & w8748;
assign v2681 = ~(w8749 | w8858);
assign w8859 = v2681;
assign w8860 = ~w8857 & w8859;
assign v2682 = ~(w8749 | w8860);
assign w8861 = v2682;
assign w8862 = ~w8725 & w8735;
assign v2683 = ~(w8736 | w8862);
assign w8863 = v2683;
assign w8864 = ~w8861 & w8863;
assign w8865 = (~w8736 & w8861) | (~w8736 & w30156) | (w8861 & w30156);
assign w8866 = ~w8712 & w8722;
assign v2684 = ~(w8723 | w8866);
assign w8867 = v2684;
assign w8868 = ~w8865 & w8867;
assign v2685 = ~(w8723 | w8868);
assign w8869 = v2685;
assign v2686 = ~(w8699 | w8709);
assign w8870 = v2686;
assign v2687 = ~(w8710 | w8870);
assign w8871 = v2687;
assign w8872 = ~w8869 & w8871;
assign w8873 = (~w8710 & w8869) | (~w8710 & w30329) | (w8869 & w30329);
assign w8874 = w8697 & ~w8873;
assign v2688 = ~(w8695 | w8874);
assign w8875 = v2688;
assign v2689 = ~(w8671 | w8681);
assign w8876 = v2689;
assign v2690 = ~(w8682 | w8876);
assign w8877 = v2690;
assign w8878 = ~w8875 & w8877;
assign w8879 = (~w8682 & w8875) | (~w8682 & w30491) | (w8875 & w30491);
assign v2691 = ~(w8658 | w8668);
assign w8880 = v2691;
assign v2692 = ~(w8669 | w8880);
assign w8881 = v2692;
assign w8882 = ~w8879 & w8881;
assign v2693 = ~(w8669 | w8882);
assign w8883 = v2693;
assign w8884 = ~w8645 & w8655;
assign v2694 = ~(w8656 | w8884);
assign w8885 = v2694;
assign w8886 = ~w8883 & w8885;
assign w8887 = (~w8656 & w8883) | (~w8656 & w30608) | (w8883 & w30608);
assign v2695 = ~(w8632 | w8642);
assign w8888 = v2695;
assign v2696 = ~(w8643 | w8888);
assign w8889 = v2696;
assign w8890 = ~w8887 & w8889;
assign v2697 = ~(w8643 | w8890);
assign w8891 = v2697;
assign v2698 = ~(w8627 | w8629);
assign w8892 = v2698;
assign v2699 = ~(w8630 | w8892);
assign w8893 = v2699;
assign w8894 = ~w8891 & w8893;
assign w8895 = (~w8630 & w8891) | (~w8630 & w30804) | (w8891 & w30804);
assign v2700 = ~(w8606 | w8616);
assign w8896 = v2700;
assign v2701 = ~(w8617 | w8896);
assign w8897 = v2701;
assign w8898 = ~w8895 & w8897;
assign v2702 = ~(w8617 | w8898);
assign w8899 = v2702;
assign w8900 = ~w8898 & w31025;
assign v2703 = ~(w8603 | w8900);
assign w8901 = v2703;
assign w8902 = (~w8589 & ~w8901) | (~w8589 & w31174) | (~w8901 & w31174);
assign w8903 = ~w8576 & w8902;
assign v2704 = ~(w8575 | w8903);
assign w8904 = v2704;
assign w8905 = w8562 & w8904;
assign v2705 = ~(w8560 | w8905);
assign w8906 = v2705;
assign w8907 = w8545 & ~w8906;
assign w8908 = ~w8545 & w8906;
assign v2706 = ~(w8907 | w8908);
assign w8909 = v2706;
assign w8910 = w3758 & w7178;
assign w8911 = ~w3752 & w7765;
assign w8912 = ~w3587 & w7466;
assign v2707 = ~(w8911 | w8912);
assign w8913 = v2707;
assign w8914 = ~w3666 & w7177;
assign w8915 = w8913 & ~w8914;
assign w8916 = ~w8910 & w8915;
assign w8917 = pi11 & ~w8916;
assign w8918 = ~pi11 & w8916;
assign v2708 = ~(w8917 | w8918);
assign w8919 = v2708;
assign w8920 = w8909 & w8919;
assign v2709 = ~(w8907 | w8920);
assign w8921 = v2709;
assign w8922 = w8543 & ~w8921;
assign w8923 = ~w8543 & w8921;
assign v2710 = ~(w8922 | w8923);
assign w8924 = v2710;
assign w8925 = ~w4149 & w8141;
assign w8926 = w8132 & w8138;
assign w8927 = ~w4082 & w8926;
assign w8928 = ~w4134 & w8140;
assign w8929 = ~w4035 & w8526;
assign v2711 = ~(w8928 | w8929);
assign w8930 = v2711;
assign w8931 = ~w8927 & w8930;
assign w8932 = ~w8925 & w8931;
assign w8933 = pi08 & ~w8932;
assign w8934 = ~pi08 & w8932;
assign v2712 = ~(w8933 | w8934);
assign w8935 = v2712;
assign w8936 = w8924 & w8935;
assign v2713 = ~(w8922 | w8936);
assign w8937 = v2713;
assign w8938 = w4196 & w8141;
assign w8939 = ~w4082 & w8526;
assign w8940 = ~w4191 & w8926;
assign w8941 = ~w4035 & w8140;
assign v2714 = ~(w8940 | w8941);
assign w8942 = v2714;
assign w8943 = ~w8939 & w8942;
assign w8944 = ~w8938 & w8943;
assign w8945 = pi08 & ~w8944;
assign w8946 = ~pi08 & w8944;
assign v2715 = ~(w8945 | w8946);
assign w8947 = v2715;
assign w8948 = ~w8937 & w8947;
assign v2716 = ~(w8519 | w8521);
assign w8949 = v2716;
assign v2717 = ~(w8522 | w8949);
assign w8950 = v2717;
assign w8951 = w8937 & ~w8947;
assign v2718 = ~(w8948 | w8951);
assign w8952 = v2718;
assign w8953 = w8950 & w8952;
assign v2719 = ~(w8948 | w8953);
assign w8954 = v2719;
assign v2720 = ~(w8535 | w8537);
assign w8955 = v2720;
assign v2721 = ~(w8538 | w8955);
assign w8956 = v2721;
assign w8957 = ~w8954 & w8956;
assign w8958 = w8954 & ~w8956;
assign v2722 = ~(w8957 | w8958);
assign w8959 = v2722;
assign v2723 = ~(w8909 | w8919);
assign w8960 = v2723;
assign v2724 = ~(w8920 | w8960);
assign w8961 = v2724;
assign v2725 = ~(w8562 | w8904);
assign w8962 = v2725;
assign v2726 = ~(w8905 | w8962);
assign w8963 = v2726;
assign w8964 = w4291 & w7178;
assign w8965 = ~w3587 & w7765;
assign w8966 = ~w3666 & w7466;
assign w8967 = ~w1387 & w7177;
assign v2727 = ~(w8966 | w8967);
assign w8968 = v2727;
assign w8969 = ~w8965 & w8968;
assign w8970 = ~w8964 & w8969;
assign w8971 = pi11 & ~w8970;
assign w8972 = ~pi11 & w8970;
assign v2728 = ~(w8971 | w8972);
assign w8973 = v2728;
assign w8974 = w8963 & w8973;
assign v2729 = ~(w8963 | w8973);
assign w8975 = v2729;
assign v2730 = ~(w8974 | w8975);
assign w8976 = v2730;
assign w8977 = w4520 & w6389;
assign w8978 = ~w1795 & w6871;
assign w8979 = ~w1674 & w7004;
assign w8980 = ~w1860 & w6388;
assign v2731 = ~(w8979 | w8980);
assign w8981 = v2731;
assign w8982 = ~w8978 & w8981;
assign w8983 = ~w8977 & w8982;
assign w8984 = pi14 & ~w8983;
assign w8985 = ~pi14 & w8983;
assign v2732 = ~(w8984 | w8985);
assign w8986 = v2732;
assign v2733 = ~(w8589 | w8590);
assign w8987 = v2733;
assign v2734 = ~(w8901 | w8987);
assign w8988 = v2734;
assign w8989 = w8901 & w8987;
assign v2735 = ~(w8988 | w8989);
assign w8990 = v2735;
assign v2736 = ~(w8986 | w8990);
assign w8991 = v2736;
assign w8992 = w4538 & w6389;
assign w8993 = ~w1795 & w7004;
assign w8994 = ~w1942 & w6388;
assign w8995 = ~w1860 & w6871;
assign v2737 = ~(w8994 | w8995);
assign w8996 = v2737;
assign w8997 = ~w8993 & w8996;
assign w8998 = ~w8992 & w8997;
assign w8999 = pi14 & ~w8998;
assign w9000 = ~pi14 & w8998;
assign v2738 = ~(w8999 | w9000);
assign w9001 = v2738;
assign v2739 = ~(w8603 | w8604);
assign w9002 = v2739;
assign v2740 = ~(w8899 | w9002);
assign w9003 = v2740;
assign w9004 = w8899 & w9002;
assign v2741 = ~(w9003 | w9004);
assign w9005 = v2741;
assign w9006 = w9001 & ~w9005;
assign w9007 = ~w9001 & w9005;
assign v2742 = ~(w9006 | w9007);
assign w9008 = v2742;
assign w9009 = w4854 & w6389;
assign w9010 = ~w1860 & w7004;
assign w9011 = ~w1942 & w6871;
assign w9012 = ~w2038 & w6388;
assign v2743 = ~(w9011 | w9012);
assign w9013 = v2743;
assign w9014 = ~w9010 & w9013;
assign w9015 = ~w9009 & w9014;
assign w9016 = pi14 & ~w9015;
assign w9017 = ~pi14 & w9015;
assign v2744 = ~(w9016 | w9017);
assign w9018 = v2744;
assign w9019 = w8895 & ~w8897;
assign v2745 = ~(w8898 | w9019);
assign w9020 = v2745;
assign w9021 = w9018 & w9020;
assign v2746 = ~(w9018 | w9020);
assign w9022 = v2746;
assign w9023 = w8891 & ~w8893;
assign v2747 = ~(w8894 | w9023);
assign w9024 = v2747;
assign w9025 = w4702 & w6389;
assign w9026 = ~w1942 & w7004;
assign w9027 = ~w2038 & w6871;
assign w9028 = ~w2089 & w6388;
assign v2748 = ~(w9027 | w9028);
assign w9029 = v2748;
assign w9030 = ~w9026 & w9029;
assign w9031 = ~w9025 & w9030;
assign w9032 = pi14 & ~w9031;
assign w9033 = ~pi14 & w9031;
assign v2749 = ~(w9032 | w9033);
assign w9034 = v2749;
assign w9035 = w9024 & w9034;
assign w9036 = w8887 & ~w8889;
assign v2750 = ~(w8890 | w9036);
assign w9037 = v2750;
assign w9038 = w5049 & w6389;
assign w9039 = ~w2202 & w6388;
assign w9040 = ~w2089 & w6871;
assign w9041 = ~w2038 & w7004;
assign v2751 = ~(w9040 | w9041);
assign w9042 = v2751;
assign w9043 = ~w9039 & w9042;
assign w9044 = ~w9038 & w9043;
assign w9045 = pi14 & ~w9044;
assign w9046 = ~pi14 & w9044;
assign v2752 = ~(w9045 | w9046);
assign w9047 = v2752;
assign w9048 = w9037 & w9047;
assign v2753 = ~(w9037 | w9047);
assign w9049 = v2753;
assign v2754 = ~(w9048 | w9049);
assign w9050 = v2754;
assign w9051 = w8883 & ~w8885;
assign v2755 = ~(w8886 | w9051);
assign w9052 = v2755;
assign w9053 = w5033 & w6389;
assign w9054 = ~w2202 & w6871;
assign w9055 = ~w2089 & w7004;
assign v2756 = ~(w9054 | w9055);
assign w9056 = v2756;
assign w9057 = ~w2290 & w6388;
assign w9058 = w9056 & ~w9057;
assign w9059 = ~w9053 & w9058;
assign w9060 = ~pi14 & w9059;
assign w9061 = pi14 & ~w9059;
assign v2757 = ~(w9060 | w9061);
assign w9062 = v2757;
assign v2758 = ~(w9052 | w9062);
assign w9063 = v2758;
assign w9064 = w9052 & w9062;
assign w9065 = w5262 & w6389;
assign w9066 = ~w2202 & w7004;
assign w9067 = ~w2339 & w6388;
assign w9068 = ~w2290 & w6871;
assign v2759 = ~(w9067 | w9068);
assign w9069 = v2759;
assign w9070 = ~w9066 & w9069;
assign w9071 = ~w9065 & w9070;
assign w9072 = pi14 & ~w9071;
assign w9073 = ~pi14 & w9071;
assign v2760 = ~(w9072 | w9073);
assign w9074 = v2760;
assign w9075 = w8879 & ~w8881;
assign v2761 = ~(w8882 | w9075);
assign w9076 = v2761;
assign w9077 = w9074 & w9076;
assign v2762 = ~(w9074 | w9076);
assign w9078 = v2762;
assign v2763 = ~(w9077 | w9078);
assign w9079 = v2763;
assign w9080 = w8875 & ~w8877;
assign v2764 = ~(w8878 | w9080);
assign w9081 = v2764;
assign w9082 = w5280 & w6389;
assign w9083 = ~w2424 & w6388;
assign w9084 = ~w2339 & w6871;
assign v2765 = ~(w9083 | w9084);
assign w9085 = v2765;
assign w9086 = ~w2290 & w7004;
assign w9087 = w9085 & ~w9086;
assign w9088 = ~w9082 & w9087;
assign w9089 = pi14 & ~w9088;
assign w9090 = ~pi14 & w9088;
assign v2766 = ~(w9089 | w9090);
assign w9091 = v2766;
assign w9092 = w9081 & w9091;
assign w9093 = ~w8697 & w8873;
assign v2767 = ~(w8874 | w9093);
assign w9094 = v2767;
assign w9095 = ~w2492 & w6388;
assign w9096 = w5665 & w6389;
assign w9097 = ~w2424 & w6871;
assign w9098 = ~w2339 & w7004;
assign v2768 = ~(w9097 | w9098);
assign w9099 = v2768;
assign w9100 = ~w9096 & w9099;
assign w9101 = ~w9095 & w9100;
assign w9102 = pi14 & w9101;
assign v2769 = ~(pi14 | w9101);
assign w9103 = v2769;
assign v2770 = ~(w9102 | w9103);
assign w9104 = v2770;
assign w9105 = w9094 & ~w9104;
assign w9106 = w8869 & ~w8871;
assign v2771 = ~(w8872 | w9106);
assign w9107 = v2771;
assign w9108 = ~w2568 & w6388;
assign w9109 = w5449 & w6389;
assign w9110 = ~w2492 & w6871;
assign w9111 = ~w2424 & w7004;
assign v2772 = ~(w9110 | w9111);
assign w9112 = v2772;
assign w9113 = ~w9109 & w9112;
assign w9114 = ~w9108 & w9113;
assign w9115 = pi14 & w9114;
assign v2773 = ~(pi14 | w9114);
assign w9116 = v2773;
assign v2774 = ~(w9115 | w9116);
assign w9117 = v2774;
assign w9118 = w9107 & ~w9117;
assign w9119 = w8865 & ~w8867;
assign v2775 = ~(w8868 | w9119);
assign w9120 = v2775;
assign w9121 = w5898 & w6389;
assign w9122 = ~w2568 & w6871;
assign w9123 = ~w2596 & w6388;
assign w9124 = ~w2492 & w7004;
assign v2776 = ~(w9123 | w9124);
assign w9125 = v2776;
assign w9126 = ~w9122 & w9125;
assign w9127 = ~w9121 & w9126;
assign w9128 = pi14 & ~w9127;
assign w9129 = ~pi14 & w9127;
assign v2777 = ~(w9128 | w9129);
assign w9130 = v2777;
assign w9131 = w9120 & w9130;
assign w9132 = w8861 & ~w8863;
assign v2778 = ~(w8864 | w9132);
assign w9133 = v2778;
assign w9134 = w6031 & w6389;
assign w9135 = ~w2568 & w7004;
assign w9136 = ~w2596 & w6871;
assign v2779 = ~(w9135 | w9136);
assign w9137 = v2779;
assign w9138 = ~w2669 & w6388;
assign w9139 = w9137 & ~w9138;
assign w9140 = ~w9134 & w9139;
assign w9141 = pi14 & w9140;
assign v2780 = ~(pi14 | w9140);
assign w9142 = v2780;
assign v2781 = ~(w9141 | w9142);
assign w9143 = v2781;
assign w9144 = w9133 & ~w9143;
assign w9145 = w8857 & ~w8859;
assign v2782 = ~(w8860 | w9145);
assign w9146 = v2782;
assign w9147 = w5880 & w6389;
assign w9148 = ~w2669 & w6871;
assign w9149 = ~w2724 & w6388;
assign w9150 = ~w2596 & w7004;
assign v2783 = ~(w9149 | w9150);
assign w9151 = v2783;
assign w9152 = ~w9148 & w9151;
assign w9153 = ~w9147 & w9152;
assign w9154 = pi14 & ~w9153;
assign w9155 = ~pi14 & w9153;
assign v2784 = ~(w9154 | w9155);
assign w9156 = v2784;
assign w9157 = w9146 & w9156;
assign w9158 = w8853 & ~w8855;
assign v2785 = ~(w8856 | w9158);
assign w9159 = v2785;
assign w9160 = w6148 & w6389;
assign w9161 = ~w2669 & w7004;
assign w9162 = ~w2811 & w6388;
assign w9163 = ~w2724 & w6871;
assign v2786 = ~(w9162 | w9163);
assign w9164 = v2786;
assign w9165 = ~w9161 & w9164;
assign w9166 = ~w9160 & w9165;
assign w9167 = pi14 & ~w9166;
assign w9168 = ~pi14 & w9166;
assign v2787 = ~(w9167 | w9168);
assign w9169 = v2787;
assign w9170 = w9159 & w9169;
assign w9171 = w8849 & ~w8851;
assign v2788 = ~(w8852 | w9171);
assign w9172 = v2788;
assign w9173 = ~w2846 & w6388;
assign w9174 = w6389 & ~w6447;
assign w9175 = ~w2811 & w6871;
assign w9176 = ~w2724 & w7004;
assign v2789 = ~(w9175 | w9176);
assign w9177 = v2789;
assign w9178 = ~w9174 & w9177;
assign w9179 = ~w9173 & w9178;
assign w9180 = pi14 & w9179;
assign v2790 = ~(pi14 | w9179);
assign w9181 = v2790;
assign v2791 = ~(w9180 | w9181);
assign w9182 = v2791;
assign w9183 = w9172 & ~w9182;
assign w9184 = w8845 & ~w8847;
assign v2792 = ~(w8848 | w9184);
assign w9185 = v2792;
assign w9186 = w6389 & w6459;
assign w9187 = ~w2811 & w7004;
assign w9188 = ~w2846 & w6871;
assign w9189 = ~w2937 & w6388;
assign v2793 = ~(w9188 | w9189);
assign w9190 = v2793;
assign w9191 = ~w9187 & w9190;
assign w9192 = ~w9186 & w9191;
assign w9193 = pi14 & ~w9192;
assign w9194 = ~pi14 & w9192;
assign v2794 = ~(w9193 | w9194);
assign w9195 = v2794;
assign w9196 = w9185 & w9195;
assign w9197 = w8841 & ~w8843;
assign v2795 = ~(w8844 | w9197);
assign w9198 = v2795;
assign w9199 = w6130 & w6389;
assign w9200 = ~w2846 & w7004;
assign w9201 = ~w2937 & w6871;
assign v2796 = ~(w9200 | w9201);
assign w9202 = v2796;
assign w9203 = ~w3000 & w6388;
assign w9204 = w9202 & ~w9203;
assign w9205 = ~w9199 & w9204;
assign v2797 = ~(pi14 | w9205);
assign w9206 = v2797;
assign w9207 = pi14 & w9205;
assign v2798 = ~(w9206 | w9207);
assign w9208 = v2798;
assign w9209 = w9198 & ~w9208;
assign w9210 = w8837 & ~w8839;
assign v2799 = ~(w8840 | w9210);
assign w9211 = v2799;
assign w9212 = ~w3000 & w6871;
assign w9213 = ~w2937 & w7004;
assign v2800 = ~(w9212 | w9213);
assign w9214 = v2800;
assign w9215 = ~w3068 & w6388;
assign w9216 = w9214 & ~w9215;
assign w9217 = (w9216 & w6505) | (w9216 & w29658) | (w6505 & w29658);
assign w9218 = pi14 & w9217;
assign v2801 = ~(pi14 | w9217);
assign w9219 = v2801;
assign v2802 = ~(w9218 | w9219);
assign w9220 = v2802;
assign w9221 = w9211 & ~w9220;
assign v2803 = ~(w8827 | w8835);
assign w9222 = v2803;
assign v2804 = ~(w8836 | w9222);
assign w9223 = v2804;
assign w9224 = ~w3000 & w7004;
assign w9225 = ~w3068 & w6871;
assign v2805 = ~(w9224 | w9225);
assign w9226 = v2805;
assign w9227 = ~w3124 & w6388;
assign w9228 = w9226 & ~w9227;
assign w9229 = (w6551 & w29659) | (w6551 & w29660) | (w29659 & w29660);
assign w9230 = (~w6551 & w29661) | (~w6551 & w29662) | (w29661 & w29662);
assign v2806 = ~(w9229 | w9230);
assign w9231 = v2806;
assign w9232 = w9223 & ~w9231;
assign w9233 = ~w3124 & w6871;
assign w9234 = ~w3068 & w7004;
assign v2807 = ~(w9233 | w9234);
assign w9235 = v2807;
assign w9236 = ~w3162 & w6388;
assign w9237 = w9235 & ~w9236;
assign w9238 = (w6603 & w29247) | (w6603 & w29248) | (w29247 & w29248);
assign w9239 = (~w6603 & w29249) | (~w6603 & w29250) | (w29249 & w29250);
assign v2808 = ~(w9238 | w9239);
assign w9240 = v2808;
assign w9241 = pi17 & ~w8824;
assign w9242 = ~w8816 & w9241;
assign w9243 = w8816 & ~w9241;
assign v2809 = ~(w9242 | w9243);
assign w9244 = v2809;
assign w9245 = ~w9240 & w9244;
assign w9246 = w8818 & ~w8823;
assign v2810 = ~(w8824 | w9246);
assign w9247 = v2810;
assign w9248 = ~w3211 & w6388;
assign w9249 = ~w3124 & w7004;
assign w9250 = ~w3162 & w6871;
assign v2811 = ~(w9249 | w9250);
assign w9251 = v2811;
assign w9252 = ~w9248 & w9251;
assign w9253 = (~w6641 & w28959) | (~w6641 & w28960) | (w28959 & w28960);
assign w9254 = (w6641 & w28961) | (w6641 & w28962) | (w28961 & w28962);
assign v2812 = ~(w9253 | w9254);
assign w9255 = v2812;
assign w9256 = w9247 & w9255;
assign w9257 = ~w3262 & w6871;
assign w9258 = (w7004 & ~w3210) | (w7004 & w29251) | (~w3210 & w29251);
assign w9259 = (w6388 & ~w3331) | (w6388 & w29252) | (~w3331 & w29252);
assign v2813 = ~(w9258 | w9259);
assign w9260 = v2813;
assign w9261 = (~w6676 & w28963) | (~w6676 & w28964) | (w28963 & w28964);
assign w9262 = ~w3332 & w6383;
assign w9263 = (w28965 & ~w3331) | (w28965 & w29253) | (~w3331 & w29253);
assign w9264 = w6389 & ~w7309;
assign w9265 = (w6871 & ~w3331) | (w6871 & w28966) | (~w3331 & w28966);
assign w9266 = (w7004 & ~w3261) | (w7004 & w28967) | (~w3261 & w28967);
assign v2814 = ~(w9265 | w9266);
assign w9267 = v2814;
assign w9268 = ~w9264 & w9267;
assign w9269 = ~w9264 & w28694;
assign w9270 = ~w9264 & w28968;
assign w9271 = w9261 & w9270;
assign w9272 = w8817 & w9271;
assign v2815 = ~(w8817 | w9271);
assign w9273 = v2815;
assign v2816 = ~(w9272 | w9273);
assign w9274 = v2816;
assign w9275 = ~w3162 & w7004;
assign w9276 = (w6388 & ~w3261) | (w6388 & w29478) | (~w3261 & w29478);
assign v2817 = ~(w9275 | w9276);
assign w9277 = v2817;
assign w9278 = ~w3211 & w6871;
assign w9279 = (~w6735 & w29254) | (~w6735 & w29255) | (w29254 & w29255);
assign w9280 = (w6735 & w29256) | (w6735 & w29257) | (w29256 & w29257);
assign v2818 = ~(w9279 | w9280);
assign w9281 = v2818;
assign w9282 = w9274 & ~w9281;
assign w9283 = (~w9272 & ~w9274) | (~w9272 & w29258) | (~w9274 & w29258);
assign v2819 = ~(w9247 | w9255);
assign w9284 = v2819;
assign v2820 = ~(w9256 | w9284);
assign w9285 = v2820;
assign w9286 = ~w9283 & w9285;
assign w9287 = (~w9256 & ~w9285) | (~w9256 & w29259) | (~w9285 & w29259);
assign w9288 = w9240 & ~w9244;
assign v2821 = ~(w9245 | w9288);
assign w9289 = v2821;
assign w9290 = ~w9287 & w9289;
assign v2822 = ~(w9245 | w9290);
assign w9291 = v2822;
assign w9292 = ~w9223 & w9231;
assign v2823 = ~(w9232 | w9292);
assign w9293 = v2823;
assign w9294 = ~w9291 & w9293;
assign w9295 = (~w9232 & w9291) | (~w9232 & w29479) | (w9291 & w29479);
assign w9296 = ~w9211 & w9220;
assign v2824 = ~(w9221 | w9296);
assign w9297 = v2824;
assign w9298 = ~w9295 & w9297;
assign v2825 = ~(w9221 | w9298);
assign w9299 = v2825;
assign w9300 = ~w9198 & w9208;
assign v2826 = ~(w9209 | w9300);
assign w9301 = v2826;
assign w9302 = ~w9299 & w9301;
assign w9303 = (~w9209 & w9299) | (~w9209 & w29663) | (w9299 & w29663);
assign v2827 = ~(w9185 | w9195);
assign w9304 = v2827;
assign v2828 = ~(w9196 | w9304);
assign w9305 = v2828;
assign w9306 = ~w9303 & w9305;
assign v2829 = ~(w9196 | w9306);
assign w9307 = v2829;
assign w9308 = ~w9172 & w9182;
assign v2830 = ~(w9183 | w9308);
assign w9309 = v2830;
assign w9310 = ~w9307 & w9309;
assign w9311 = (~w9183 & w9307) | (~w9183 & w29846) | (w9307 & w29846);
assign v2831 = ~(w9159 | w9169);
assign w9312 = v2831;
assign v2832 = ~(w9170 | w9312);
assign w9313 = v2832;
assign w9314 = ~w9311 & w9313;
assign v2833 = ~(w9170 | w9314);
assign w9315 = v2833;
assign v2834 = ~(w9146 | w9156);
assign w9316 = v2834;
assign v2835 = ~(w9157 | w9316);
assign w9317 = v2835;
assign w9318 = ~w9315 & w9317;
assign w9319 = (~w9157 & w9315) | (~w9157 & w30019) | (w9315 & w30019);
assign w9320 = ~w9133 & w9143;
assign v2836 = ~(w9144 | w9320);
assign w9321 = v2836;
assign w9322 = ~w9319 & w9321;
assign v2837 = ~(w9144 | w9322);
assign w9323 = v2837;
assign v2838 = ~(w9120 | w9130);
assign w9324 = v2838;
assign v2839 = ~(w9131 | w9324);
assign w9325 = v2839;
assign w9326 = ~w9323 & w9325;
assign w9327 = (~w9131 & w9323) | (~w9131 & w30330) | (w9323 & w30330);
assign w9328 = ~w9107 & w9117;
assign v2840 = ~(w9118 | w9328);
assign w9329 = v2840;
assign w9330 = ~w9327 & w9329;
assign v2841 = ~(w9118 | w9330);
assign w9331 = v2841;
assign w9332 = ~w9094 & w9104;
assign v2842 = ~(w9105 | w9332);
assign w9333 = v2842;
assign w9334 = ~w9331 & w9333;
assign w9335 = (~w9105 & w9331) | (~w9105 & w30492) | (w9331 & w30492);
assign v2843 = ~(w9081 | w9091);
assign w9336 = v2843;
assign v2844 = ~(w9092 | w9336);
assign w9337 = v2844;
assign w9338 = ~w9335 & w9337;
assign v2845 = ~(w9092 | w9338);
assign w9339 = v2845;
assign w9340 = w9079 & ~w9339;
assign w9341 = (~w9077 & w9339) | (~w9077 & w30609) | (w9339 & w30609);
assign w9342 = (~w9063 & ~w9341) | (~w9063 & w30020) | (~w9341 & w30020);
assign w9343 = w9050 & w9342;
assign w9344 = (~w9048 & ~w9050) | (~w9048 & w30021) | (~w9050 & w30021);
assign v2846 = ~(w9024 | w9034);
assign w9345 = v2846;
assign w9346 = (~w9035 & w9344) | (~w9035 & w30805) | (w9344 & w30805);
assign w9347 = (~w9021 & w9346) | (~w9021 & w31026) | (w9346 & w31026);
assign w9348 = w9008 & ~w9347;
assign w9349 = (~w9006 & ~w9008) | (~w9006 & w30022) | (~w9008 & w30022);
assign w9350 = w8986 & w8990;
assign v2847 = ~(w8991 | w9350);
assign w9351 = v2847;
assign w9352 = w9349 & w9351;
assign v2848 = ~(w8991 | w9352);
assign w9353 = v2848;
assign w9354 = w3494 & w6389;
assign w9355 = ~w1609 & w7004;
assign w9356 = ~w1674 & w6871;
assign v2849 = ~(w9355 | w9356);
assign w9357 = v2849;
assign w9358 = ~w1795 & w6388;
assign w9359 = w9357 & ~w9358;
assign w9360 = ~w9354 & w9359;
assign w9361 = pi14 & ~w9360;
assign w9362 = ~pi14 & w9360;
assign v2850 = ~(w9361 | w9362);
assign w9363 = v2850;
assign v2851 = ~(w8575 | w8576);
assign w9364 = v2851;
assign w9365 = w8902 & ~w9364;
assign w9366 = ~w8902 & w9364;
assign v2852 = ~(w9365 | w9366);
assign w9367 = v2852;
assign w9368 = w9363 & ~w9367;
assign w9369 = ~w9363 & w9367;
assign v2853 = ~(w9368 | w9369);
assign w9370 = v2853;
assign v2854 = ~(w9353 | w9370);
assign w9371 = v2854;
assign v2855 = ~(w9363 | w9367);
assign w9372 = v2855;
assign v2856 = ~(w9371 | w9372);
assign w9373 = v2856;
assign w9374 = w8976 & w9373;
assign v2857 = ~(w8974 | w9374);
assign w9375 = v2857;
assign w9376 = w8961 & ~w9375;
assign w9377 = w4405 & w8141;
assign w9378 = ~w4035 & w8926;
assign w9379 = ~w3920 & w8140;
assign w9380 = ~w4134 & w8526;
assign v2858 = ~(w9379 | w9380);
assign w9381 = v2858;
assign w9382 = ~w9378 & w9381;
assign w9383 = ~w9377 & w9382;
assign w9384 = pi08 & ~w9383;
assign w9385 = ~pi08 & w9383;
assign v2859 = ~(w9384 | w9385);
assign w9386 = v2859;
assign w9387 = ~w8961 & w9375;
assign v2860 = ~(w9376 | w9387);
assign w9388 = v2860;
assign w9389 = w9386 & w9388;
assign v2861 = ~(w9376 | w9389);
assign w9390 = v2861;
assign w9391 = ~pi04 & pi05;
assign w9392 = pi04 & ~pi05;
assign v2862 = ~(w9391 | w9392);
assign w9393 = v2862;
assign v2863 = ~(pi02 | pi03);
assign w9394 = v2863;
assign w9395 = pi02 & pi03;
assign v2864 = ~(w9394 | w9395);
assign w9396 = v2864;
assign v2865 = ~(pi03 | pi04);
assign w9397 = v2865;
assign w9398 = pi03 & pi04;
assign v2866 = ~(w9397 | w9398);
assign w9399 = v2866;
assign v2867 = ~(w9396 | w9399);
assign w9400 = v2867;
assign w9401 = ~w9393 & w9400;
assign w9402 = ~w9393 & w9396;
assign w9403 = (w9402 & w4168) | (w9402 & w30023) | (w4168 & w30023);
assign v2868 = ~(w9401 | w9403);
assign w9404 = v2868;
assign v2869 = ~(w4191 | w9404);
assign w9405 = v2869;
assign w9406 = ~pi05 & w9405;
assign w9407 = pi05 & ~w9405;
assign v2870 = ~(w9406 | w9407);
assign w9408 = v2870;
assign v2871 = ~(w9390 | w9408);
assign w9409 = v2871;
assign v2872 = ~(w8924 | w8935);
assign w9410 = v2872;
assign v2873 = ~(w8936 | w9410);
assign w9411 = v2873;
assign w9412 = w9390 & w9408;
assign v2874 = ~(w9409 | w9412);
assign w9413 = v2874;
assign w9414 = w9411 & w9413;
assign v2875 = ~(w9409 | w9414);
assign w9415 = v2875;
assign v2876 = ~(w8950 | w8952);
assign w9416 = v2876;
assign v2877 = ~(w8953 | w9416);
assign w9417 = v2877;
assign w9418 = ~w9415 & w9417;
assign w9419 = w9415 & ~w9417;
assign v2878 = ~(w9418 | w9419);
assign w9420 = v2878;
assign v2879 = ~(w9411 | w9413);
assign w9421 = v2879;
assign v2880 = ~(w9414 | w9421);
assign w9422 = v2880;
assign v2881 = ~(w8976 | w9373);
assign w9423 = v2881;
assign v2882 = ~(w9374 | w9423);
assign w9424 = v2882;
assign w9425 = ~w3920 & w8526;
assign w9426 = ~w3752 & w8140;
assign w9427 = ~w4134 & w8926;
assign v2883 = ~(w9426 | w9427);
assign w9428 = v2883;
assign w9429 = ~w9425 & w9428;
assign w9430 = (w9429 & ~w4309) | (w9429 & w30024) | (~w4309 & w30024);
assign w9431 = pi08 & ~w9430;
assign w9432 = ~pi08 & w9430;
assign v2884 = ~(w9431 | w9432);
assign w9433 = v2884;
assign w9434 = w9424 & w9433;
assign v2885 = ~(w9424 | w9433);
assign w9435 = v2885;
assign v2886 = ~(w9434 | w9435);
assign w9436 = v2886;
assign w9437 = w3843 & w7178;
assign w9438 = ~w1496 & w7177;
assign w9439 = ~w3666 & w7765;
assign w9440 = ~w1387 & w7466;
assign v2887 = ~(w9439 | w9440);
assign w9441 = v2887;
assign w9442 = ~w9438 & w9441;
assign w9443 = ~w9437 & w9442;
assign w9444 = pi11 & ~w9443;
assign w9445 = ~pi11 & w9443;
assign v2888 = ~(w9444 | w9445);
assign w9446 = v2888;
assign w9447 = w9353 & ~w9370;
assign w9448 = ~w9353 & w9370;
assign v2889 = ~(w9447 | w9448);
assign w9449 = v2889;
assign w9450 = w9446 & w9449;
assign w9451 = w3397 & w7178;
assign w9452 = ~w1387 & w7765;
assign w9453 = ~w1609 & w7177;
assign w9454 = ~w1496 & w7466;
assign v2890 = ~(w9453 | w9454);
assign w9455 = v2890;
assign w9456 = ~w9452 & w9455;
assign w9457 = ~w9451 & w9456;
assign w9458 = pi11 & ~w9457;
assign w9459 = ~pi11 & w9457;
assign v2891 = ~(w9458 | w9459);
assign w9460 = v2891;
assign v2892 = ~(w9349 | w9351);
assign w9461 = v2892;
assign v2893 = ~(w9352 | w9461);
assign w9462 = v2893;
assign w9463 = ~w9460 & w9462;
assign w9464 = w7168 & w7172;
assign w9465 = ~w3510 & w9464;
assign w9466 = ~w1496 & w7765;
assign w9467 = ~w1674 & w7177;
assign w9468 = ~w1609 & w7466;
assign v2894 = ~(w9467 | w9468);
assign w9469 = v2894;
assign w9470 = ~w9466 & w9469;
assign w9471 = pi11 & ~w9470;
assign v2895 = ~(w9465 | w9471);
assign w9472 = v2895;
assign w9473 = ~w3510 & w7178;
assign w9474 = ~pi11 & w9470;
assign w9475 = ~w9473 & w9474;
assign w9476 = w9472 & ~w9475;
assign w9477 = ~w9008 & w9347;
assign v2896 = ~(w9348 | w9477);
assign w9478 = v2896;
assign w9479 = w9476 & w9478;
assign v2897 = ~(w9476 | w9478);
assign w9480 = v2897;
assign v2898 = ~(w9479 | w9480);
assign w9481 = v2898;
assign v2899 = ~(w9021 | w9022);
assign w9482 = v2899;
assign w9483 = w9346 & ~w9482;
assign w9484 = ~w9346 & w9482;
assign v2900 = ~(w9483 | w9484);
assign w9485 = v2900;
assign w9486 = w3494 & w7178;
assign w9487 = ~w1609 & w7765;
assign w9488 = ~w1674 & w7466;
assign v2901 = ~(w9487 | w9488);
assign w9489 = v2901;
assign w9490 = ~w1795 & w7177;
assign w9491 = w9489 & ~w9490;
assign w9492 = ~w9486 & w9491;
assign w9493 = ~pi11 & w9492;
assign w9494 = pi11 & ~w9492;
assign v2902 = ~(w9493 | w9494);
assign w9495 = v2902;
assign v2903 = ~(w9485 | w9495);
assign w9496 = v2903;
assign w9497 = w9485 & w9495;
assign w9498 = w4520 & w7178;
assign w9499 = ~w1795 & w7466;
assign w9500 = ~w1674 & w7765;
assign w9501 = ~w1860 & w7177;
assign v2904 = ~(w9500 | w9501);
assign w9502 = v2904;
assign w9503 = ~w9499 & w9502;
assign w9504 = ~w9498 & w9503;
assign w9505 = pi11 & ~w9504;
assign w9506 = ~pi11 & w9504;
assign v2905 = ~(w9505 | w9506);
assign w9507 = v2905;
assign v2906 = ~(w9035 | w9345);
assign w9508 = v2906;
assign w9509 = w9344 & ~w9508;
assign w9510 = ~w9344 & w9508;
assign v2907 = ~(w9509 | w9510);
assign w9511 = v2907;
assign w9512 = w9507 & ~w9511;
assign w9513 = ~w9507 & w9511;
assign v2908 = ~(w9512 | w9513);
assign w9514 = v2908;
assign w9515 = w4538 & w7178;
assign w9516 = ~w1795 & w7765;
assign w9517 = ~w1942 & w7177;
assign w9518 = ~w1860 & w7466;
assign v2909 = ~(w9517 | w9518);
assign w9519 = v2909;
assign w9520 = ~w9516 & w9519;
assign w9521 = ~w9515 & w9520;
assign w9522 = pi11 & ~w9521;
assign w9523 = ~pi11 & w9521;
assign v2910 = ~(w9522 | w9523);
assign w9524 = v2910;
assign v2911 = ~(w9050 | w9342);
assign w9525 = v2911;
assign v2912 = ~(w9343 | w9525);
assign w9526 = v2912;
assign v2913 = ~(w9524 | w9526);
assign w9527 = v2913;
assign w9528 = w9524 & w9526;
assign w9529 = w4854 & w7178;
assign w9530 = ~w1860 & w7765;
assign w9531 = ~w2038 & w7177;
assign w9532 = ~w1942 & w7466;
assign v2914 = ~(w9531 | w9532);
assign w9533 = v2914;
assign w9534 = ~w9530 & w9533;
assign w9535 = ~w9529 & w9534;
assign w9536 = pi11 & ~w9535;
assign w9537 = ~pi11 & w9535;
assign v2915 = ~(w9536 | w9537);
assign w9538 = v2915;
assign v2916 = ~(w9063 | w9064);
assign w9539 = v2916;
assign v2917 = ~(w9341 | w9539);
assign w9540 = v2917;
assign w9541 = w9341 & w9539;
assign v2918 = ~(w9540 | w9541);
assign w9542 = v2918;
assign w9543 = w9538 & ~w9542;
assign w9544 = ~w9538 & w9542;
assign v2919 = ~(w9543 | w9544);
assign w9545 = v2919;
assign w9546 = ~w9079 & w9339;
assign v2920 = ~(w9340 | w9546);
assign w9547 = v2920;
assign w9548 = w4702 & w7178;
assign w9549 = ~w2038 & w7466;
assign w9550 = ~w1942 & w7765;
assign w9551 = ~w2089 & w7177;
assign v2921 = ~(w9550 | w9551);
assign w9552 = v2921;
assign w9553 = ~w9549 & w9552;
assign w9554 = ~w9548 & w9553;
assign w9555 = pi11 & ~w9554;
assign w9556 = ~pi11 & w9554;
assign v2922 = ~(w9555 | w9556);
assign w9557 = v2922;
assign w9558 = w9547 & w9557;
assign v2923 = ~(w9547 | w9557);
assign w9559 = v2923;
assign w9560 = w9335 & ~w9337;
assign v2924 = ~(w9338 | w9560);
assign w9561 = v2924;
assign w9562 = w5049 & w7178;
assign w9563 = ~w2202 & w7177;
assign w9564 = ~w2089 & w7466;
assign w9565 = ~w2038 & w7765;
assign v2925 = ~(w9564 | w9565);
assign w9566 = v2925;
assign w9567 = ~w9563 & w9566;
assign w9568 = ~w9562 & w9567;
assign w9569 = pi11 & ~w9568;
assign w9570 = ~pi11 & w9568;
assign v2926 = ~(w9569 | w9570);
assign w9571 = v2926;
assign w9572 = w9561 & w9571;
assign v2927 = ~(w9561 | w9571);
assign w9573 = v2927;
assign v2928 = ~(w9572 | w9573);
assign w9574 = v2928;
assign w9575 = w9331 & ~w9333;
assign v2929 = ~(w9334 | w9575);
assign w9576 = v2929;
assign w9577 = w5033 & w7178;
assign w9578 = ~w2202 & w7466;
assign w9579 = ~w2089 & w7765;
assign v2930 = ~(w9578 | w9579);
assign w9580 = v2930;
assign w9581 = ~w2290 & w7177;
assign w9582 = w9580 & ~w9581;
assign w9583 = ~w9577 & w9582;
assign w9584 = ~pi11 & w9583;
assign w9585 = pi11 & ~w9583;
assign v2931 = ~(w9584 | w9585);
assign w9586 = v2931;
assign v2932 = ~(w9576 | w9586);
assign w9587 = v2932;
assign w9588 = w9576 & w9586;
assign w9589 = w5262 & w7178;
assign w9590 = ~w2202 & w7765;
assign w9591 = ~w2339 & w7177;
assign w9592 = ~w2290 & w7466;
assign v2933 = ~(w9591 | w9592);
assign w9593 = v2933;
assign w9594 = ~w9590 & w9593;
assign w9595 = ~w9589 & w9594;
assign w9596 = pi11 & ~w9595;
assign w9597 = ~pi11 & w9595;
assign v2934 = ~(w9596 | w9597);
assign w9598 = v2934;
assign w9599 = w9327 & ~w9329;
assign v2935 = ~(w9330 | w9599);
assign w9600 = v2935;
assign w9601 = w9598 & w9600;
assign w9602 = w9323 & ~w9325;
assign v2936 = ~(w9326 | w9602);
assign w9603 = v2936;
assign w9604 = w5280 & w7178;
assign w9605 = ~w2424 & w7177;
assign w9606 = ~w2339 & w7466;
assign v2937 = ~(w9605 | w9606);
assign w9607 = v2937;
assign w9608 = ~w2290 & w7765;
assign w9609 = w9607 & ~w9608;
assign w9610 = ~w9604 & w9609;
assign w9611 = pi11 & ~w9610;
assign w9612 = ~pi11 & w9610;
assign v2938 = ~(w9611 | w9612);
assign w9613 = v2938;
assign w9614 = w9603 & w9613;
assign w9615 = w9319 & ~w9321;
assign v2939 = ~(w9322 | w9615);
assign w9616 = v2939;
assign w9617 = w5665 & w7178;
assign w9618 = ~w2492 & w7177;
assign w9619 = ~w2424 & w7466;
assign w9620 = ~w2339 & w7765;
assign v2940 = ~(w9619 | w9620);
assign w9621 = v2940;
assign w9622 = ~w9618 & w9621;
assign w9623 = ~w9617 & w9622;
assign w9624 = pi11 & ~w9623;
assign w9625 = ~pi11 & w9623;
assign v2941 = ~(w9624 | w9625);
assign w9626 = v2941;
assign w9627 = w9616 & w9626;
assign w9628 = w9315 & ~w9317;
assign v2942 = ~(w9318 | w9628);
assign w9629 = v2942;
assign w9630 = w5449 & w7178;
assign w9631 = ~w2424 & w7765;
assign w9632 = ~w2492 & w7466;
assign w9633 = ~w2568 & w7177;
assign v2943 = ~(w9632 | w9633);
assign w9634 = v2943;
assign w9635 = ~w9631 & w9634;
assign w9636 = ~w9630 & w9635;
assign w9637 = pi11 & ~w9636;
assign w9638 = ~pi11 & w9636;
assign v2944 = ~(w9637 | w9638);
assign w9639 = v2944;
assign w9640 = w9629 & w9639;
assign w9641 = w9311 & ~w9313;
assign v2945 = ~(w9314 | w9641);
assign w9642 = v2945;
assign w9643 = w5898 & w7178;
assign w9644 = ~w2568 & w7466;
assign w9645 = ~w2596 & w7177;
assign w9646 = ~w2492 & w7765;
assign v2946 = ~(w9645 | w9646);
assign w9647 = v2946;
assign w9648 = ~w9644 & w9647;
assign w9649 = ~w9643 & w9648;
assign w9650 = pi11 & ~w9649;
assign w9651 = ~pi11 & w9649;
assign v2947 = ~(w9650 | w9651);
assign w9652 = v2947;
assign w9653 = w9642 & w9652;
assign w9654 = w9307 & ~w9309;
assign v2948 = ~(w9310 | w9654);
assign w9655 = v2948;
assign w9656 = w6031 & w7178;
assign w9657 = ~w2568 & w7765;
assign w9658 = ~w2669 & w7177;
assign w9659 = ~w2596 & w7466;
assign v2949 = ~(w9658 | w9659);
assign w9660 = v2949;
assign w9661 = ~w9657 & w9660;
assign w9662 = ~w9656 & w9661;
assign w9663 = pi11 & ~w9662;
assign w9664 = ~pi11 & w9662;
assign v2950 = ~(w9663 | w9664);
assign w9665 = v2950;
assign w9666 = w9655 & w9665;
assign w9667 = w9303 & ~w9305;
assign v2951 = ~(w9306 | w9667);
assign w9668 = v2951;
assign w9669 = w5880 & w7178;
assign w9670 = ~w2669 & w7466;
assign w9671 = ~w2724 & w7177;
assign w9672 = ~w2596 & w7765;
assign v2952 = ~(w9671 | w9672);
assign w9673 = v2952;
assign w9674 = ~w9670 & w9673;
assign w9675 = ~w9669 & w9674;
assign w9676 = pi11 & ~w9675;
assign w9677 = ~pi11 & w9675;
assign v2953 = ~(w9676 | w9677);
assign w9678 = v2953;
assign w9679 = w9668 & w9678;
assign w9680 = w9299 & ~w9301;
assign v2954 = ~(w9302 | w9680);
assign w9681 = v2954;
assign w9682 = w6148 & w7178;
assign w9683 = ~w2669 & w7765;
assign w9684 = ~w2811 & w7177;
assign w9685 = ~w2724 & w7466;
assign v2955 = ~(w9684 | w9685);
assign w9686 = v2955;
assign w9687 = ~w9683 & w9686;
assign w9688 = ~w9682 & w9687;
assign w9689 = pi11 & ~w9688;
assign w9690 = ~pi11 & w9688;
assign v2956 = ~(w9689 | w9690);
assign w9691 = v2956;
assign w9692 = w9681 & w9691;
assign w9693 = w9295 & ~w9297;
assign v2957 = ~(w9298 | w9693);
assign w9694 = v2957;
assign w9695 = ~w6447 & w7178;
assign w9696 = ~w2724 & w7765;
assign w9697 = ~w2811 & w7466;
assign v2958 = ~(w9696 | w9697);
assign w9698 = v2958;
assign w9699 = ~w2846 & w7177;
assign w9700 = w9698 & ~w9699;
assign w9701 = ~w9695 & w9700;
assign w9702 = ~pi11 & w9701;
assign w9703 = pi11 & ~w9701;
assign v2959 = ~(w9702 | w9703);
assign w9704 = v2959;
assign w9705 = w9694 & w9704;
assign w9706 = w9291 & ~w9293;
assign v2960 = ~(w9294 | w9706);
assign w9707 = v2960;
assign w9708 = w6459 & w7178;
assign w9709 = ~w2846 & w7466;
assign w9710 = ~w2811 & w7765;
assign w9711 = ~w2937 & w7177;
assign v2961 = ~(w9710 | w9711);
assign w9712 = v2961;
assign w9713 = ~w9709 & w9712;
assign w9714 = ~w9708 & w9713;
assign w9715 = pi11 & ~w9714;
assign w9716 = ~pi11 & w9714;
assign v2962 = ~(w9715 | w9716);
assign w9717 = v2962;
assign w9718 = w9707 & w9717;
assign w9719 = w9287 & ~w9289;
assign v2963 = ~(w9290 | w9719);
assign w9720 = v2963;
assign w9721 = w6130 & w7178;
assign w9722 = ~w2846 & w7765;
assign w9723 = ~w2937 & w7466;
assign v2964 = ~(w9722 | w9723);
assign w9724 = v2964;
assign w9725 = ~w3000 & w7177;
assign w9726 = w9724 & ~w9725;
assign w9727 = ~w9721 & w9726;
assign v2965 = ~(pi11 | w9727);
assign w9728 = v2965;
assign w9729 = pi11 & w9727;
assign v2966 = ~(w9728 | w9729);
assign w9730 = v2966;
assign w9731 = w9720 & ~w9730;
assign w9732 = w9283 & ~w9285;
assign v2967 = ~(w9286 | w9732);
assign w9733 = v2967;
assign w9734 = ~w3000 & w7466;
assign w9735 = ~w2937 & w7765;
assign v2968 = ~(w9734 | w9735);
assign w9736 = v2968;
assign w9737 = ~w3068 & w7177;
assign w9738 = w9736 & ~w9737;
assign w9739 = (w9738 & w6505) | (w9738 & w29480) | (w6505 & w29480);
assign v2969 = ~(pi11 | w9739);
assign w9740 = v2969;
assign w9741 = pi11 & w9739;
assign v2970 = ~(w9740 | w9741);
assign w9742 = v2970;
assign w9743 = w9733 & ~w9742;
assign w9744 = ~w9274 & w9281;
assign v2971 = ~(w9282 | w9744);
assign w9745 = v2971;
assign w9746 = ~w3124 & w7177;
assign w9747 = ~w3068 & w7466;
assign v2972 = ~(w9746 | w9747);
assign w9748 = v2972;
assign w9749 = ~w3000 & w7765;
assign w9750 = w9748 & ~w9749;
assign w9751 = (w6551 & w29481) | (w6551 & w29482) | (w29481 & w29482);
assign w9752 = (~w6551 & w29483) | (~w6551 & w29484) | (w29483 & w29484);
assign v2973 = ~(w9751 | w9752);
assign w9753 = v2973;
assign w9754 = w9745 & ~w9753;
assign w9755 = ~w3068 & w7765;
assign w9756 = ~w3162 & w7177;
assign w9757 = ~w3124 & w7466;
assign v2974 = ~(w9756 | w9757);
assign w9758 = v2974;
assign w9759 = ~w9755 & w9758;
assign w9760 = (w6603 & w28969) | (w6603 & w28970) | (w28969 & w28970);
assign w9761 = (~w6603 & w28971) | (~w6603 & w28972) | (w28971 & w28972);
assign v2975 = ~(w9760 | w9761);
assign w9762 = v2975;
assign w9763 = pi14 & ~w9269;
assign w9764 = ~w9261 & w9763;
assign w9765 = w9261 & ~w9763;
assign v2976 = ~(w9764 | w9765);
assign w9766 = v2976;
assign w9767 = w9762 & w9766;
assign w9768 = w9263 & ~w9268;
assign v2977 = ~(w9269 | w9768);
assign w9769 = v2977;
assign w9770 = ~w3162 & w7466;
assign w9771 = ~w3124 & w7765;
assign v2978 = ~(w9770 | w9771);
assign w9772 = v2978;
assign w9773 = ~w3211 & w7177;
assign w9774 = w9772 & ~w9773;
assign w9775 = (~w6641 & w28696) | (~w6641 & w28697) | (w28696 & w28697);
assign w9776 = (w6641 & w28698) | (w6641 & w28699) | (w28698 & w28699);
assign v2979 = ~(w9775 | w9776);
assign w9777 = v2979;
assign w9778 = w9769 & ~w9777;
assign w9779 = w6676 & w7178;
assign w9780 = ~w3211 & w7765;
assign w9781 = ~w3332 & w7177;
assign w9782 = ~w3262 & w7466;
assign v2980 = ~(w9781 | w9782);
assign w9783 = v2980;
assign w9784 = ~w9780 & w9783;
assign w9785 = ~w9779 & w9784;
assign w9786 = (w7172 & ~w3331) | (w7172 & w28700) | (~w3331 & w28700);
assign w9787 = (~w3331 & w28973) | (~w3331 & w28974) | (w28973 & w28974);
assign w9788 = w7178 & ~w7309;
assign w9789 = (w7466 & ~w3331) | (w7466 & w28701) | (~w3331 & w28701);
assign w9790 = (w7765 & ~w3261) | (w7765 & w28702) | (~w3261 & w28702);
assign v2981 = ~(w9789 | w9790);
assign w9791 = v2981;
assign w9792 = ~w9788 & w9791;
assign w9793 = ~w9788 & w28481;
assign w9794 = w9785 & w28704;
assign w9795 = (~w9262 & ~w9785) | (~w9262 & w28705) | (~w9785 & w28705);
assign v2982 = ~(w9794 | w9795);
assign w9796 = v2982;
assign w9797 = ~w3162 & w7765;
assign w9798 = (w7177 & ~w3261) | (w7177 & w29261) | (~w3261 & w29261);
assign v2983 = ~(w9797 | w9798);
assign w9799 = v2983;
assign w9800 = ~w3211 & w7466;
assign w9801 = (~w6735 & w28975) | (~w6735 & w28976) | (w28975 & w28976);
assign w9802 = (w6735 & w28977) | (w6735 & w28978) | (w28977 & w28978);
assign v2984 = ~(w9801 | w9802);
assign w9803 = v2984;
assign w9804 = w9796 & ~w9803;
assign w9805 = (~w9794 & ~w9796) | (~w9794 & w28979) | (~w9796 & w28979);
assign w9806 = ~w9769 & w9777;
assign v2985 = ~(w9778 | w9806);
assign w9807 = v2985;
assign w9808 = ~w9805 & w9807;
assign w9809 = (~w9778 & ~w9807) | (~w9778 & w28980) | (~w9807 & w28980);
assign v2986 = ~(w9762 | w9766);
assign w9810 = v2986;
assign v2987 = ~(w9767 | w9810);
assign w9811 = v2987;
assign w9812 = ~w9809 & w9811;
assign v2988 = ~(w9767 | w9812);
assign w9813 = v2988;
assign w9814 = ~w9745 & w9753;
assign v2989 = ~(w9754 | w9814);
assign w9815 = v2989;
assign w9816 = ~w9813 & w9815;
assign w9817 = (~w9754 & w9813) | (~w9754 & w29262) | (w9813 & w29262);
assign w9818 = ~w9733 & w9742;
assign v2990 = ~(w9743 | w9818);
assign w9819 = v2990;
assign w9820 = ~w9817 & w9819;
assign v2991 = ~(w9743 | w9820);
assign w9821 = v2991;
assign w9822 = ~w9720 & w9730;
assign v2992 = ~(w9731 | w9822);
assign w9823 = v2992;
assign w9824 = ~w9821 & w9823;
assign w9825 = (~w9731 & w9821) | (~w9731 & w29263) | (w9821 & w29263);
assign v2993 = ~(w9707 | w9717);
assign w9826 = v2993;
assign v2994 = ~(w9718 | w9826);
assign w9827 = v2994;
assign w9828 = ~w9825 & w9827;
assign v2995 = ~(w9718 | w9828);
assign w9829 = v2995;
assign v2996 = ~(w9694 | w9704);
assign w9830 = v2996;
assign v2997 = ~(w9705 | w9830);
assign w9831 = v2997;
assign w9832 = ~w9829 & w9831;
assign w9833 = (~w9705 & w9829) | (~w9705 & w29485) | (w9829 & w29485);
assign v2998 = ~(w9681 | w9691);
assign w9834 = v2998;
assign v2999 = ~(w9692 | w9834);
assign w9835 = v2999;
assign w9836 = ~w9833 & w9835;
assign v3000 = ~(w9692 | w9836);
assign w9837 = v3000;
assign v3001 = ~(w9668 | w9678);
assign w9838 = v3001;
assign v3002 = ~(w9679 | w9838);
assign w9839 = v3002;
assign w9840 = ~w9837 & w9839;
assign w9841 = (~w9679 & w9837) | (~w9679 & w29664) | (w9837 & w29664);
assign v3003 = ~(w9655 | w9665);
assign w9842 = v3003;
assign v3004 = ~(w9666 | w9842);
assign w9843 = v3004;
assign w9844 = ~w9841 & w9843;
assign v3005 = ~(w9666 | w9844);
assign w9845 = v3005;
assign v3006 = ~(w9642 | w9652);
assign w9846 = v3006;
assign v3007 = ~(w9653 | w9846);
assign w9847 = v3007;
assign w9848 = ~w9845 & w9847;
assign w9849 = (~w9653 & w9845) | (~w9653 & w29847) | (w9845 & w29847);
assign v3008 = ~(w9629 | w9639);
assign w9850 = v3008;
assign v3009 = ~(w9640 | w9850);
assign w9851 = v3009;
assign w9852 = ~w9849 & w9851;
assign v3010 = ~(w9640 | w9852);
assign w9853 = v3010;
assign v3011 = ~(w9616 | w9626);
assign w9854 = v3011;
assign v3012 = ~(w9627 | w9854);
assign w9855 = v3012;
assign w9856 = ~w9853 & w9855;
assign w9857 = (~w9627 & w9853) | (~w9627 & w30157) | (w9853 & w30157);
assign v3013 = ~(w9603 | w9613);
assign w9858 = v3013;
assign v3014 = ~(w9614 | w9858);
assign w9859 = v3014;
assign w9860 = ~w9857 & w9859;
assign v3015 = ~(w9614 | w9860);
assign w9861 = v3015;
assign v3016 = ~(w9598 | w9600);
assign w9862 = v3016;
assign v3017 = ~(w9601 | w9862);
assign w9863 = v3017;
assign w9864 = ~w9861 & w9863;
assign w9865 = (~w9601 & w9861) | (~w9601 & w30331) | (w9861 & w30331);
assign w9866 = (~w9587 & ~w9865) | (~w9587 & w29848) | (~w9865 & w29848);
assign w9867 = w9574 & w9866;
assign w9868 = (~w9572 & ~w9574) | (~w9572 & w29849) | (~w9574 & w29849);
assign w9869 = (~w9558 & w9868) | (~w9558 & w30610) | (w9868 & w30610);
assign w9870 = w9545 & ~w9869;
assign w9871 = (~w9543 & ~w9545) | (~w9543 & w29850) | (~w9545 & w29850);
assign w9872 = (w29850 & w30806) | (w29850 & w30807) | (w30806 & w30807);
assign v3018 = ~(w9527 | w9872);
assign w9873 = v3018;
assign w9874 = ~w9514 & w9873;
assign w9875 = ~w9510 & w29851;
assign w9876 = (~w9875 & w9514) | (~w9875 & w29264) | (w9514 & w29264);
assign w9877 = (~w9496 & ~w9876) | (~w9496 & w29852) | (~w9876 & w29852);
assign w9878 = w9481 & w9877;
assign w9879 = (~w9479 & ~w9481) | (~w9479 & w29853) | (~w9481 & w29853);
assign w9880 = w9460 & ~w9462;
assign v3019 = ~(w9463 | w9880);
assign w9881 = v3019;
assign w9882 = w9879 & w9881;
assign v3020 = ~(w9463 | w9882);
assign w9883 = v3020;
assign v3021 = ~(w9446 | w9449);
assign w9884 = v3021;
assign v3022 = ~(w9450 | w9884);
assign w9885 = v3022;
assign w9886 = w9883 & w9885;
assign v3023 = ~(w9450 | w9886);
assign w9887 = v3023;
assign w9888 = w9436 & ~w9887;
assign v3024 = ~(w9434 | w9888);
assign w9889 = v3024;
assign w9890 = ~w4082 & w9401;
assign w9891 = ~w9396 & w9399;
assign w9892 = ~w4191 & w9891;
assign v3025 = ~(w9890 | w9892);
assign w9893 = v3025;
assign w9894 = (~w4425 & w29854) | (~w4425 & w29855) | (w29854 & w29855);
assign w9895 = (w4425 & w29856) | (w4425 & w29857) | (w29856 & w29857);
assign v3026 = ~(w9894 | w9895);
assign w9896 = v3026;
assign w9897 = ~w9889 & w9896;
assign v3027 = ~(w9386 | w9388);
assign w9898 = v3027;
assign v3028 = ~(w9389 | w9898);
assign w9899 = v3028;
assign w9900 = w9889 & ~w9896;
assign v3029 = ~(w9897 | w9900);
assign w9901 = v3029;
assign w9902 = w9899 & w9901;
assign v3030 = ~(w9897 | w9902);
assign w9903 = v3030;
assign w9904 = w9422 & ~w9903;
assign w9905 = ~w9422 & w9903;
assign v3031 = ~(w9904 | w9905);
assign w9906 = v3031;
assign w9907 = ~w3928 & w8141;
assign w9908 = ~w3920 & w8926;
assign w9909 = ~w3752 & w8526;
assign w9910 = ~w3587 & w8140;
assign v3032 = ~(w9909 | w9910);
assign w9911 = v3032;
assign w9912 = ~w9908 & w9911;
assign w9913 = ~w9907 & w9912;
assign w9914 = pi08 & ~w9913;
assign w9915 = ~pi08 & w9913;
assign v3033 = ~(w9914 | w9915);
assign w9916 = v3033;
assign v3034 = ~(w9883 | w9885);
assign w9917 = v3034;
assign v3035 = ~(w9886 | w9917);
assign w9918 = v3035;
assign v3036 = ~(w9916 | w9918);
assign w9919 = v3036;
assign w9920 = w8130 & w8138;
assign w9921 = w3758 & w9920;
assign w9922 = ~w3752 & w8926;
assign w9923 = ~w3666 & w8140;
assign w9924 = ~w3587 & w8526;
assign v3037 = ~(w9923 | w9924);
assign w9925 = v3037;
assign w9926 = ~w9922 & w9925;
assign w9927 = pi08 & ~w9926;
assign v3038 = ~(w9921 | w9927);
assign w9928 = v3038;
assign w9929 = w3758 & w8141;
assign w9930 = ~pi08 & w9926;
assign w9931 = ~w9929 & w9930;
assign w9932 = w9928 & ~w9931;
assign v3039 = ~(w9879 | w9881);
assign w9933 = v3039;
assign v3040 = ~(w9882 | w9933);
assign w9934 = v3040;
assign w9935 = w9932 & ~w9934;
assign w9936 = ~w9932 & w9934;
assign v3041 = ~(w9935 | w9936);
assign w9937 = v3041;
assign w9938 = w4291 & w9920;
assign w9939 = ~w3666 & w8526;
assign w9940 = ~w1387 & w8140;
assign w9941 = ~w3587 & w8926;
assign v3042 = ~(w9940 | w9941);
assign w9942 = v3042;
assign w9943 = ~w9939 & w9942;
assign w9944 = pi08 & ~w9943;
assign v3043 = ~(w9938 | w9944);
assign w9945 = v3043;
assign w9946 = w4291 & w8141;
assign w9947 = ~pi08 & w9943;
assign w9948 = ~w9946 & w9947;
assign w9949 = w9945 & ~w9948;
assign v3044 = ~(w9481 | w9877);
assign w9950 = v3044;
assign v3045 = ~(w9878 | w9950);
assign w9951 = v3045;
assign v3046 = ~(w9949 | w9951);
assign w9952 = v3046;
assign w9953 = w9949 & w9951;
assign w9954 = ~w3666 & w8926;
assign w9955 = ~w1387 & w8526;
assign w9956 = ~w1496 & w8140;
assign v3047 = ~(w9955 | w9956);
assign w9957 = v3047;
assign w9958 = ~w9954 & w9957;
assign w9959 = pi08 & ~w9958;
assign w9960 = w3843 & w9920;
assign v3048 = ~(w9959 | w9960);
assign w9961 = v3048;
assign w9962 = w3843 & w8141;
assign w9963 = ~pi08 & w9958;
assign w9964 = ~w9962 & w9963;
assign w9965 = w9961 & ~w9964;
assign v3049 = ~(w9496 | w9497);
assign w9966 = v3049;
assign v3050 = ~(w9876 | w9966);
assign w9967 = v3050;
assign w9968 = w9876 & w9966;
assign v3051 = ~(w9967 | w9968);
assign w9969 = v3051;
assign w9970 = w9965 & ~w9969;
assign w9971 = ~w9965 & w9969;
assign v3052 = ~(w9970 | w9971);
assign w9972 = v3052;
assign w9973 = w3397 & w8141;
assign w9974 = ~w1609 & w8140;
assign w9975 = ~w1496 & w8526;
assign w9976 = ~w1387 & w8926;
assign v3053 = ~(w9975 | w9976);
assign w9977 = v3053;
assign w9978 = ~w9974 & w9977;
assign w9979 = ~w9973 & w9978;
assign w9980 = pi08 & ~w9979;
assign w9981 = ~pi08 & w9979;
assign v3054 = ~(w9980 | w9981);
assign w9982 = v3054;
assign w9983 = w9514 & ~w9873;
assign v3055 = ~(w9874 | w9983);
assign w9984 = v3055;
assign v3056 = ~(w9982 | w9984);
assign w9985 = v3056;
assign w9986 = ~w3510 & w9920;
assign w9987 = ~w1674 & w8140;
assign w9988 = ~w1609 & w8526;
assign w9989 = ~w1496 & w8926;
assign v3057 = ~(w9988 | w9989);
assign w9990 = v3057;
assign w9991 = ~w9987 & w9990;
assign w9992 = pi08 & ~w9991;
assign v3058 = ~(w9986 | w9992);
assign w9993 = v3058;
assign w9994 = ~w3510 & w8141;
assign w9995 = ~pi08 & w9991;
assign w9996 = ~w9994 & w9995;
assign w9997 = w9993 & ~w9996;
assign v3059 = ~(w9527 | w9528);
assign w9998 = v3059;
assign w9999 = w9871 & w9998;
assign v3060 = ~(w9871 | w9998);
assign w10000 = v3060;
assign v3061 = ~(w9999 | w10000);
assign w10001 = v3061;
assign w10002 = w9997 & ~w10001;
assign w10003 = ~w9997 & w10001;
assign v3062 = ~(w10002 | w10003);
assign w10004 = v3062;
assign w10005 = ~w9545 & w9869;
assign v3063 = ~(w9870 | w10005);
assign w10006 = v3063;
assign w10007 = w3494 & w8141;
assign w10008 = ~w1609 & w8926;
assign w10009 = ~w1674 & w8526;
assign v3064 = ~(w10008 | w10009);
assign w10010 = v3064;
assign w10011 = ~w1795 & w8140;
assign w10012 = w10010 & ~w10011;
assign w10013 = ~w10007 & w10012;
assign w10014 = pi08 & ~w10013;
assign w10015 = ~pi08 & w10013;
assign v3065 = ~(w10014 | w10015);
assign w10016 = v3065;
assign v3066 = ~(w10006 | w10016);
assign w10017 = v3066;
assign w10018 = w10006 & w10016;
assign w10019 = w4520 & w8141;
assign w10020 = ~w1795 & w8526;
assign w10021 = ~w1674 & w8926;
assign w10022 = ~w1860 & w8140;
assign v3067 = ~(w10021 | w10022);
assign w10023 = v3067;
assign w10024 = ~w10020 & w10023;
assign w10025 = ~w10019 & w10024;
assign w10026 = pi08 & ~w10025;
assign w10027 = ~pi08 & w10025;
assign v3068 = ~(w10026 | w10027);
assign w10028 = v3068;
assign v3069 = ~(w9558 | w9559);
assign w10029 = v3069;
assign w10030 = w9868 & ~w10029;
assign w10031 = ~w9868 & w10029;
assign v3070 = ~(w10030 | w10031);
assign w10032 = v3070;
assign w10033 = w10028 & ~w10032;
assign w10034 = ~w10028 & w10032;
assign v3071 = ~(w10033 | w10034);
assign w10035 = v3071;
assign w10036 = w4538 & w8141;
assign w10037 = ~w1795 & w8926;
assign w10038 = ~w1942 & w8140;
assign w10039 = ~w1860 & w8526;
assign v3072 = ~(w10038 | w10039);
assign w10040 = v3072;
assign w10041 = ~w10037 & w10040;
assign w10042 = ~w10036 & w10041;
assign w10043 = pi08 & ~w10042;
assign w10044 = ~pi08 & w10042;
assign v3073 = ~(w10043 | w10044);
assign w10045 = v3073;
assign v3074 = ~(w9574 | w9866);
assign w10046 = v3074;
assign v3075 = ~(w9867 | w10046);
assign w10047 = v3075;
assign v3076 = ~(w10045 | w10047);
assign w10048 = v3076;
assign w10049 = w10045 & w10047;
assign w10050 = w4854 & w8141;
assign w10051 = ~w1860 & w8926;
assign w10052 = ~w2038 & w8140;
assign w10053 = ~w1942 & w8526;
assign v3077 = ~(w10052 | w10053);
assign w10054 = v3077;
assign w10055 = ~w10051 & w10054;
assign w10056 = ~w10050 & w10055;
assign w10057 = pi08 & ~w10056;
assign w10058 = ~pi08 & w10056;
assign v3078 = ~(w10057 | w10058);
assign w10059 = v3078;
assign v3079 = ~(w9587 | w9588);
assign w10060 = v3079;
assign w10061 = w9865 & w10060;
assign v3080 = ~(w9865 | w10060);
assign w10062 = v3080;
assign v3081 = ~(w10061 | w10062);
assign w10063 = v3081;
assign w10064 = w10059 & ~w10063;
assign w10065 = ~w10059 & w10063;
assign v3082 = ~(w10064 | w10065);
assign w10066 = v3082;
assign w10067 = w9861 & ~w9863;
assign v3083 = ~(w9864 | w10067);
assign w10068 = v3083;
assign w10069 = w4702 & w8141;
assign w10070 = ~w2038 & w8526;
assign w10071 = ~w1942 & w8926;
assign w10072 = ~w2089 & w8140;
assign v3084 = ~(w10071 | w10072);
assign w10073 = v3084;
assign w10074 = ~w10070 & w10073;
assign w10075 = ~w10069 & w10074;
assign w10076 = pi08 & ~w10075;
assign w10077 = ~pi08 & w10075;
assign v3085 = ~(w10076 | w10077);
assign w10078 = v3085;
assign v3086 = ~(w10068 | w10078);
assign w10079 = v3086;
assign w10080 = w10068 & w10078;
assign w10081 = w9857 & ~w9859;
assign v3087 = ~(w9860 | w10081);
assign w10082 = v3087;
assign w10083 = ~w2202 & w8140;
assign w10084 = w5049 & w8141;
assign w10085 = ~w2089 & w8526;
assign w10086 = ~w2038 & w8926;
assign v3088 = ~(w10085 | w10086);
assign w10087 = v3088;
assign w10088 = ~w10084 & w10087;
assign w10089 = ~w10083 & w10088;
assign w10090 = pi08 & w10089;
assign v3089 = ~(pi08 | w10089);
assign w10091 = v3089;
assign v3090 = ~(w10090 | w10091);
assign w10092 = v3090;
assign w10093 = w10082 & ~w10092;
assign w10094 = ~w10082 & w10092;
assign v3091 = ~(w10093 | w10094);
assign w10095 = v3091;
assign w10096 = w9853 & ~w9855;
assign v3092 = ~(w9856 | w10096);
assign w10097 = v3092;
assign w10098 = w5033 & w8141;
assign w10099 = ~w2202 & w8526;
assign w10100 = ~w2089 & w8926;
assign w10101 = ~w2290 & w8140;
assign v3093 = ~(w10100 | w10101);
assign w10102 = v3093;
assign w10103 = ~w10099 & w10102;
assign w10104 = ~w10098 & w10103;
assign w10105 = pi08 & ~w10104;
assign w10106 = ~pi08 & w10104;
assign v3094 = ~(w10105 | w10106);
assign w10107 = v3094;
assign v3095 = ~(w10097 | w10107);
assign w10108 = v3095;
assign w10109 = w10097 & w10107;
assign w10110 = w9849 & ~w9851;
assign v3096 = ~(w9852 | w10110);
assign w10111 = v3096;
assign w10112 = w5262 & w8141;
assign w10113 = ~w2202 & w8926;
assign w10114 = ~w2339 & w8140;
assign w10115 = ~w2290 & w8526;
assign v3097 = ~(w10114 | w10115);
assign w10116 = v3097;
assign w10117 = ~w10113 & w10116;
assign w10118 = ~w10112 & w10117;
assign w10119 = pi08 & ~w10118;
assign w10120 = ~pi08 & w10118;
assign v3098 = ~(w10119 | w10120);
assign w10121 = v3098;
assign w10122 = w10111 & w10121;
assign w10123 = w9845 & ~w9847;
assign v3099 = ~(w9848 | w10123);
assign w10124 = v3099;
assign w10125 = w5280 & w8141;
assign w10126 = ~w2424 & w8140;
assign w10127 = ~w2339 & w8526;
assign v3100 = ~(w10126 | w10127);
assign w10128 = v3100;
assign w10129 = ~w2290 & w8926;
assign w10130 = w10128 & ~w10129;
assign w10131 = ~w10125 & w10130;
assign w10132 = ~pi08 & w10131;
assign w10133 = pi08 & ~w10131;
assign v3101 = ~(w10132 | w10133);
assign w10134 = v3101;
assign w10135 = w10124 & w10134;
assign w10136 = w9841 & ~w9843;
assign v3102 = ~(w9844 | w10136);
assign w10137 = v3102;
assign w10138 = ~w2492 & w8140;
assign w10139 = w5665 & w8141;
assign w10140 = ~w2424 & w8526;
assign w10141 = ~w2339 & w8926;
assign v3103 = ~(w10140 | w10141);
assign w10142 = v3103;
assign w10143 = ~w10139 & w10142;
assign w10144 = ~w10138 & w10143;
assign w10145 = pi08 & w10144;
assign v3104 = ~(pi08 | w10144);
assign w10146 = v3104;
assign v3105 = ~(w10145 | w10146);
assign w10147 = v3105;
assign w10148 = w10137 & ~w10147;
assign w10149 = w9837 & ~w9839;
assign v3106 = ~(w9840 | w10149);
assign w10150 = v3106;
assign w10151 = ~w2568 & w8140;
assign w10152 = w5449 & w8141;
assign w10153 = ~w2492 & w8526;
assign w10154 = ~w2424 & w8926;
assign v3107 = ~(w10153 | w10154);
assign w10155 = v3107;
assign w10156 = ~w10152 & w10155;
assign w10157 = ~w10151 & w10156;
assign w10158 = pi08 & w10157;
assign v3108 = ~(pi08 | w10157);
assign w10159 = v3108;
assign v3109 = ~(w10158 | w10159);
assign w10160 = v3109;
assign w10161 = w10150 & ~w10160;
assign w10162 = w9833 & ~w9835;
assign v3110 = ~(w9836 | w10162);
assign w10163 = v3110;
assign w10164 = w5898 & w8141;
assign w10165 = ~w2568 & w8526;
assign w10166 = ~w2596 & w8140;
assign w10167 = ~w2492 & w8926;
assign v3111 = ~(w10166 | w10167);
assign w10168 = v3111;
assign w10169 = ~w10165 & w10168;
assign w10170 = ~w10164 & w10169;
assign w10171 = pi08 & ~w10170;
assign w10172 = ~pi08 & w10170;
assign v3112 = ~(w10171 | w10172);
assign w10173 = v3112;
assign w10174 = w10163 & w10173;
assign w10175 = w9829 & ~w9831;
assign v3113 = ~(w9832 | w10175);
assign w10176 = v3113;
assign w10177 = w6031 & w8141;
assign w10178 = ~w2568 & w8926;
assign w10179 = ~w2669 & w8140;
assign w10180 = ~w2596 & w8526;
assign v3114 = ~(w10179 | w10180);
assign w10181 = v3114;
assign w10182 = ~w10178 & w10181;
assign w10183 = ~w10177 & w10182;
assign w10184 = pi08 & ~w10183;
assign w10185 = ~pi08 & w10183;
assign v3115 = ~(w10184 | w10185);
assign w10186 = v3115;
assign w10187 = w10176 & w10186;
assign w10188 = w9825 & ~w9827;
assign v3116 = ~(w9828 | w10188);
assign w10189 = v3116;
assign w10190 = w5880 & w8141;
assign w10191 = ~w2669 & w8526;
assign w10192 = ~w2724 & w8140;
assign w10193 = ~w2596 & w8926;
assign v3117 = ~(w10192 | w10193);
assign w10194 = v3117;
assign w10195 = ~w10191 & w10194;
assign w10196 = ~w10190 & w10195;
assign w10197 = pi08 & ~w10196;
assign w10198 = ~pi08 & w10196;
assign v3118 = ~(w10197 | w10198);
assign w10199 = v3118;
assign w10200 = w10189 & w10199;
assign w10201 = w9821 & ~w9823;
assign v3119 = ~(w9824 | w10201);
assign w10202 = v3119;
assign w10203 = ~w2811 & w8140;
assign w10204 = w6148 & w8141;
assign w10205 = ~w2669 & w8926;
assign w10206 = ~w2724 & w8526;
assign v3120 = ~(w10205 | w10206);
assign w10207 = v3120;
assign w10208 = ~w10204 & w10207;
assign w10209 = ~w10203 & w10208;
assign w10210 = pi08 & w10209;
assign v3121 = ~(pi08 | w10209);
assign w10211 = v3121;
assign v3122 = ~(w10210 | w10211);
assign w10212 = v3122;
assign w10213 = w10202 & ~w10212;
assign w10214 = w9817 & ~w9819;
assign v3123 = ~(w9820 | w10214);
assign w10215 = v3123;
assign w10216 = ~w2846 & w8140;
assign w10217 = ~w6447 & w8141;
assign w10218 = ~w2811 & w8526;
assign w10219 = ~w2724 & w8926;
assign v3124 = ~(w10218 | w10219);
assign w10220 = v3124;
assign w10221 = ~w10217 & w10220;
assign w10222 = ~w10216 & w10221;
assign w10223 = pi08 & w10222;
assign v3125 = ~(pi08 | w10222);
assign w10224 = v3125;
assign v3126 = ~(w10223 | w10224);
assign w10225 = v3126;
assign w10226 = w10215 & ~w10225;
assign w10227 = w9813 & ~w9815;
assign v3127 = ~(w9816 | w10227);
assign w10228 = v3127;
assign w10229 = ~w2937 & w8140;
assign w10230 = w6459 & w8141;
assign w10231 = ~w2846 & w8526;
assign w10232 = ~w2811 & w8926;
assign v3128 = ~(w10231 | w10232);
assign w10233 = v3128;
assign w10234 = ~w10230 & w10233;
assign w10235 = ~w10229 & w10234;
assign w10236 = ~pi08 & w10235;
assign w10237 = pi08 & ~w10235;
assign v3129 = ~(w10236 | w10237);
assign w10238 = v3129;
assign w10239 = w10228 & w10238;
assign w10240 = w9809 & ~w9811;
assign v3130 = ~(w9812 | w10240);
assign w10241 = v3130;
assign w10242 = w6130 & w8141;
assign w10243 = ~w2846 & w8926;
assign w10244 = ~w3000 & w8140;
assign w10245 = ~w2937 & w8526;
assign v3131 = ~(w10244 | w10245);
assign w10246 = v3131;
assign w10247 = ~w10243 & w10246;
assign w10248 = ~w10242 & w10247;
assign w10249 = pi08 & ~w10248;
assign w10250 = ~pi08 & w10248;
assign v3132 = ~(w10249 | w10250);
assign w10251 = v3132;
assign w10252 = w10241 & w10251;
assign w10253 = w9805 & ~w9807;
assign v3133 = ~(w9808 | w10253);
assign w10254 = v3133;
assign w10255 = ~w3068 & w8140;
assign w10256 = ~w2937 & w8926;
assign v3134 = ~(w10255 | w10256);
assign w10257 = v3134;
assign w10258 = ~w3000 & w8526;
assign w10259 = w10257 & ~w10258;
assign w10260 = (w10259 & w6505) | (w10259 & w28981) | (w6505 & w28981);
assign w10261 = pi08 & w10260;
assign v3135 = ~(pi08 | w10260);
assign w10262 = v3135;
assign v3136 = ~(w10261 | w10262);
assign w10263 = v3136;
assign w10264 = w10254 & ~w10263;
assign w10265 = ~w9796 & w9803;
assign v3137 = ~(w9804 | w10265);
assign w10266 = v3137;
assign w10267 = ~w3068 & w8526;
assign w10268 = ~w3124 & w8140;
assign w10269 = ~w3000 & w8926;
assign v3138 = ~(w10268 | w10269);
assign w10270 = v3138;
assign w10271 = ~w10267 & w10270;
assign w10272 = (w6551 & w28982) | (w6551 & w28983) | (w28982 & w28983);
assign w10273 = (~w6551 & w28984) | (~w6551 & w28985) | (w28984 & w28985);
assign v3139 = ~(w10272 | w10273);
assign w10274 = v3139;
assign w10275 = w10266 & w10274;
assign w10276 = ~w3068 & w8926;
assign w10277 = ~w3162 & w8140;
assign w10278 = ~w3124 & w8526;
assign v3140 = ~(w10277 | w10278);
assign w10279 = v3140;
assign w10280 = ~w10276 & w10279;
assign w10281 = (w6603 & w28707) | (w6603 & w28708) | (w28707 & w28708);
assign w10282 = (~w6603 & w28709) | (~w6603 & w28710) | (w28709 & w28710);
assign v3141 = ~(w10281 | w10282);
assign w10283 = v3141;
assign w10284 = pi11 & ~w9793;
assign w10285 = ~w9785 & w10284;
assign w10286 = w9785 & ~w10284;
assign v3142 = ~(w10285 | w10286);
assign w10287 = v3142;
assign w10288 = w10283 & w10287;
assign w10289 = w9787 & ~w9792;
assign v3143 = ~(w9793 | w10289);
assign w10290 = v3143;
assign w10291 = ~w3211 & w8140;
assign w10292 = ~w3124 & w8926;
assign w10293 = ~w3162 & w8526;
assign v3144 = ~(w10292 | w10293);
assign w10294 = v3144;
assign w10295 = ~w10291 & w10294;
assign w10296 = (~w6641 & w28483) | (~w6641 & w28484) | (w28483 & w28484);
assign w10297 = (w6641 & w28485) | (w6641 & w28486) | (w28485 & w28486);
assign v3145 = ~(w10296 | w10297);
assign w10298 = v3145;
assign w10299 = w10290 & w10298;
assign w10300 = ~w3332 & w8140;
assign w10301 = (w8526 & ~w3261) | (w8526 & w28487) | (~w3261 & w28487);
assign w10302 = (w8926 & ~w3210) | (w8926 & w28488) | (~w3210 & w28488);
assign v3146 = ~(w10301 | w10302);
assign w10303 = v3146;
assign w10304 = (~w6676 & w28279) | (~w6676 & w28280) | (w28279 & w28280);
assign w10305 = (w8926 & ~w3261) | (w8926 & w28159) | (~w3261 & w28159);
assign w10306 = (w8526 & ~w3331) | (w8526 & w28160) | (~w3331 & w28160);
assign v3147 = ~(w10305 | w10306);
assign w10307 = v3147;
assign w10308 = ~w7309 & w8141;
assign w10309 = (w10307 & w7309) | (w10307 & w28281) | (w7309 & w28281);
assign w10310 = (w8138 & ~w3331) | (w8138 & w28161) | (~w3331 & w28161);
assign w10311 = pi08 & ~w10310;
assign w10312 = w10309 & w10311;
assign w10313 = w10304 & w10312;
assign w10314 = w9786 & w10313;
assign v3148 = ~(w9786 | w10313);
assign w10315 = v3148;
assign v3149 = ~(w10314 | w10315);
assign w10316 = v3149;
assign w10317 = ~w3162 & w8926;
assign w10318 = (w8140 & ~w3261) | (w8140 & w28711) | (~w3261 & w28711);
assign v3150 = ~(w10317 | w10318);
assign w10319 = v3150;
assign w10320 = ~w3211 & w8526;
assign w10321 = (w6735 & w28489) | (w6735 & w28490) | (w28489 & w28490);
assign w10322 = (~w6735 & w28491) | (~w6735 & w28492) | (w28491 & w28492);
assign v3151 = ~(w10321 | w10322);
assign w10323 = v3151;
assign w10324 = w10316 & ~w10323;
assign w10325 = (~w10314 & ~w10316) | (~w10314 & w28493) | (~w10316 & w28493);
assign v3152 = ~(w10290 | w10298);
assign w10326 = v3152;
assign v3153 = ~(w10299 | w10326);
assign w10327 = v3153;
assign w10328 = ~w10325 & w10327;
assign w10329 = (~w10299 & ~w10327) | (~w10299 & w28282) | (~w10327 & w28282);
assign v3154 = ~(w10283 | w10287);
assign w10330 = v3154;
assign v3155 = ~(w10288 | w10330);
assign w10331 = v3155;
assign w10332 = ~w10329 & w10331;
assign w10333 = (~w10288 & ~w10331) | (~w10288 & w28283) | (~w10331 & w28283);
assign v3156 = ~(w10266 | w10274);
assign w10334 = v3156;
assign v3157 = ~(w10275 | w10334);
assign w10335 = v3157;
assign w10336 = ~w10333 & w10335;
assign w10337 = (~w10275 & w10333) | (~w10275 & w28712) | (w10333 & w28712);
assign w10338 = ~w10254 & w10263;
assign v3158 = ~(w10264 | w10338);
assign w10339 = v3158;
assign w10340 = ~w10337 & w10339;
assign v3159 = ~(w10264 | w10340);
assign w10341 = v3159;
assign v3160 = ~(w10241 | w10251);
assign w10342 = v3160;
assign v3161 = ~(w10252 | w10342);
assign w10343 = v3161;
assign w10344 = ~w10341 & w10343;
assign w10345 = (~w10252 & w10341) | (~w10252 & w28986) | (w10341 & w28986);
assign v3162 = ~(w10228 | w10238);
assign w10346 = v3162;
assign v3163 = ~(w10239 | w10346);
assign w10347 = v3163;
assign w10348 = ~w10345 & w10347;
assign v3164 = ~(w10239 | w10348);
assign w10349 = v3164;
assign w10350 = ~w10215 & w10225;
assign v3165 = ~(w10226 | w10350);
assign w10351 = v3165;
assign w10352 = ~w10349 & w10351;
assign w10353 = (~w10226 & w10349) | (~w10226 & w29486) | (w10349 & w29486);
assign w10354 = ~w10202 & w10212;
assign v3166 = ~(w10213 | w10354);
assign w10355 = v3166;
assign w10356 = ~w10353 & w10355;
assign v3167 = ~(w10213 | w10356);
assign w10357 = v3167;
assign v3168 = ~(w10189 | w10199);
assign w10358 = v3168;
assign v3169 = ~(w10200 | w10358);
assign w10359 = v3169;
assign w10360 = ~w10357 & w10359;
assign w10361 = (~w10200 & w10357) | (~w10200 & w29665) | (w10357 & w29665);
assign v3170 = ~(w10176 | w10186);
assign w10362 = v3170;
assign v3171 = ~(w10187 | w10362);
assign w10363 = v3171;
assign w10364 = ~w10361 & w10363;
assign v3172 = ~(w10187 | w10364);
assign w10365 = v3172;
assign v3173 = ~(w10163 | w10173);
assign w10366 = v3173;
assign v3174 = ~(w10174 | w10366);
assign w10367 = v3174;
assign w10368 = ~w10365 & w10367;
assign w10369 = (~w10174 & w10365) | (~w10174 & w29858) | (w10365 & w29858);
assign w10370 = ~w10150 & w10160;
assign v3175 = ~(w10161 | w10370);
assign w10371 = v3175;
assign w10372 = ~w10369 & w10371;
assign v3176 = ~(w10161 | w10372);
assign w10373 = v3176;
assign w10374 = ~w10137 & w10147;
assign v3177 = ~(w10148 | w10374);
assign w10375 = v3177;
assign w10376 = ~w10373 & w10375;
assign w10377 = (~w10148 & w10373) | (~w10148 & w30025) | (w10373 & w30025);
assign v3178 = ~(w10124 | w10134);
assign w10378 = v3178;
assign v3179 = ~(w10135 | w10378);
assign w10379 = v3179;
assign w10380 = ~w10377 & w10379;
assign v3180 = ~(w10135 | w10380);
assign w10381 = v3180;
assign v3181 = ~(w10111 | w10121);
assign w10382 = v3181;
assign v3182 = ~(w10122 | w10382);
assign w10383 = v3182;
assign w10384 = ~w10381 & w10383;
assign w10385 = (~w10122 & w10381) | (~w10122 & w30158) | (w10381 & w30158);
assign w10386 = (~w10108 & ~w10385) | (~w10108 & w28987) | (~w10385 & w28987);
assign w10387 = w10095 & w10386;
assign w10388 = (~w10093 & ~w10095) | (~w10093 & w28988) | (~w10095 & w28988);
assign w10389 = (~w10079 & ~w10388) | (~w10079 & w30332) | (~w10388 & w30332);
assign w10390 = w10066 & w10389;
assign w10391 = (~w10064 & ~w10066) | (~w10064 & w28989) | (~w10066 & w28989);
assign w10392 = (w28989 & w30493) | (w28989 & w30494) | (w30493 & w30494);
assign v3183 = ~(w10048 | w10392);
assign w10393 = v3183;
assign w10394 = ~w10035 & w10393;
assign w10395 = ~w10031 & w28990;
assign w10396 = (~w10395 & w10035) | (~w10395 & w28284) | (w10035 & w28284);
assign w10397 = (~w10017 & ~w10396) | (~w10017 & w28991) | (~w10396 & w28991);
assign w10398 = w10004 & w10397;
assign w10399 = (~w10002 & ~w10004) | (~w10002 & w28992) | (~w10004 & w28992);
assign w10400 = w9982 & w9984;
assign v3184 = ~(w9985 | w10400);
assign w10401 = v3184;
assign w10402 = w10399 & w10401;
assign w10403 = (~w9985 & ~w10401) | (~w9985 & w28993) | (~w10401 & w28993);
assign w10404 = w9972 & w10403;
assign w10405 = (~w9970 & ~w10403) | (~w9970 & w31027) | (~w10403 & w31027);
assign w10406 = (~w9952 & ~w10405) | (~w9952 & w29859) | (~w10405 & w29859);
assign w10407 = w9937 & w10406;
assign w10408 = (~w9935 & ~w9937) | (~w9935 & w28994) | (~w9937 & w28994);
assign w10409 = w9916 & w9918;
assign v3185 = ~(w9919 | w10409);
assign w10410 = v3185;
assign w10411 = w10408 & w10410;
assign w10412 = (~w9919 & ~w10410) | (~w9919 & w28995) | (~w10410 & w28995);
assign w10413 = ~w9436 & w9887;
assign v3186 = ~(w9888 | w10413);
assign w10414 = v3186;
assign w10415 = w10412 & w10414;
assign v3187 = ~(w10412 | w10414);
assign w10416 = v3187;
assign v3188 = ~(w10415 | w10416);
assign w10417 = v3188;
assign w10418 = ~w4082 & w9891;
assign w10419 = w9393 & w9396;
assign w10420 = ~w4191 & w10419;
assign w10421 = ~w4035 & w9401;
assign v3189 = ~(w10420 | w10421);
assign w10422 = v3189;
assign w10423 = ~w10418 & w10422;
assign w10424 = (w10423 & ~w4196) | (w10423 & w28996) | (~w4196 & w28996);
assign w10425 = pi05 & ~w10424;
assign w10426 = ~pi05 & w10424;
assign v3190 = ~(w10425 | w10426);
assign w10427 = v3190;
assign w10428 = w10417 & w10427;
assign v3191 = ~(w10415 | w10428);
assign w10429 = v3191;
assign v3192 = ~(w9899 | w9901);
assign w10430 = v3192;
assign v3193 = ~(w9902 | w10430);
assign w10431 = v3193;
assign w10432 = w10429 & ~w10431;
assign v3194 = ~(w9937 | w10406);
assign w10433 = v3194;
assign v3195 = ~(w10407 | w10433);
assign w10434 = v3195;
assign w10435 = ~w4035 & w10419;
assign w10436 = ~w3920 & w9401;
assign w10437 = ~w4134 & w9891;
assign v3196 = ~(w10436 | w10437);
assign w10438 = v3196;
assign w10439 = ~w10435 & w10438;
assign w10440 = (w10439 & ~w4405) | (w10439 & w28997) | (~w4405 & w28997);
assign w10441 = pi05 & ~w10440;
assign w10442 = ~pi05 & w10440;
assign v3197 = ~(w10441 | w10442);
assign w10443 = v3197;
assign w10444 = w10434 & w10443;
assign w10445 = w9391 & w9396;
assign w10446 = w4309 & w10445;
assign w10447 = w9392 & w9396;
assign w10448 = w4309 & w10447;
assign w10449 = ~w3920 & w9891;
assign w10450 = ~w4134 & w10419;
assign w10451 = ~w3752 & w9401;
assign v3198 = ~(w10450 | w10451);
assign w10452 = v3198;
assign w10453 = ~w10449 & w10452;
assign w10454 = pi05 & w10453;
assign v3199 = ~(pi05 | w10453);
assign w10455 = v3199;
assign v3200 = ~(w10454 | w10455);
assign w10456 = v3200;
assign w10457 = ~w10448 & w10456;
assign v3201 = ~(w10446 | w10457);
assign w10458 = v3201;
assign v3202 = ~(w9952 | w9953);
assign w10459 = v3202;
assign v3203 = ~(w10405 | w10459);
assign w10460 = v3203;
assign w10461 = w10405 & w10459;
assign v3204 = ~(w10460 | w10461);
assign w10462 = v3204;
assign w10463 = w10458 & ~w10462;
assign w10464 = ~w10458 & w10462;
assign v3205 = ~(w10463 | w10464);
assign w10465 = v3205;
assign v3206 = ~(w9972 | w10403);
assign w10466 = v3206;
assign v3207 = ~(w10404 | w10466);
assign w10467 = v3207;
assign w10468 = ~w3928 & w9402;
assign w10469 = ~w3920 & w10419;
assign w10470 = ~w3752 & w9891;
assign v3208 = ~(w10469 | w10470);
assign w10471 = v3208;
assign w10472 = ~w3587 & w9401;
assign w10473 = w10471 & ~w10472;
assign w10474 = ~w10468 & w10473;
assign w10475 = ~pi05 & w10474;
assign w10476 = pi05 & ~w10474;
assign v3209 = ~(w10475 | w10476);
assign w10477 = v3209;
assign v3210 = ~(w10467 | w10477);
assign w10478 = v3210;
assign w10479 = w10467 & w10477;
assign w10480 = w3758 & w10445;
assign w10481 = w3758 & w10447;
assign w10482 = ~w3666 & w9401;
assign w10483 = ~w3587 & w9891;
assign w10484 = ~w3752 & w10419;
assign v3211 = ~(w10483 | w10484);
assign w10485 = v3211;
assign w10486 = ~w10482 & w10485;
assign w10487 = pi05 & w10486;
assign v3212 = ~(pi05 | w10486);
assign w10488 = v3212;
assign v3213 = ~(w10487 | w10488);
assign w10489 = v3213;
assign w10490 = ~w10481 & w10489;
assign v3214 = ~(w10480 | w10490);
assign w10491 = v3214;
assign v3215 = ~(w10399 | w10401);
assign w10492 = v3215;
assign v3216 = ~(w10402 | w10492);
assign w10493 = v3216;
assign w10494 = w10491 & ~w10493;
assign w10495 = ~w10491 & w10493;
assign v3217 = ~(w10494 | w10495);
assign w10496 = v3217;
assign w10497 = w4291 & w10445;
assign w10498 = w4291 & w10447;
assign w10499 = ~w1387 & w9401;
assign w10500 = ~w3666 & w9891;
assign w10501 = ~w3587 & w10419;
assign v3218 = ~(w10500 | w10501);
assign w10502 = v3218;
assign w10503 = ~w10499 & w10502;
assign w10504 = pi05 & w10503;
assign v3219 = ~(pi05 | w10503);
assign w10505 = v3219;
assign v3220 = ~(w10504 | w10505);
assign w10506 = v3220;
assign w10507 = ~w10498 & w10506;
assign v3221 = ~(w10497 | w10507);
assign w10508 = v3221;
assign v3222 = ~(w10004 | w10397);
assign w10509 = v3222;
assign v3223 = ~(w10398 | w10509);
assign w10510 = v3223;
assign v3224 = ~(w10508 | w10510);
assign w10511 = v3224;
assign w10512 = w10508 & w10510;
assign w10513 = w3843 & w10445;
assign w10514 = w3843 & w10447;
assign w10515 = ~w3666 & w10419;
assign w10516 = ~w1387 & w9891;
assign w10517 = ~w1496 & w9401;
assign v3225 = ~(w10516 | w10517);
assign w10518 = v3225;
assign w10519 = ~w10515 & w10518;
assign w10520 = pi05 & w10519;
assign v3226 = ~(pi05 | w10519);
assign w10521 = v3226;
assign v3227 = ~(w10520 | w10521);
assign w10522 = v3227;
assign w10523 = ~w10514 & w10522;
assign v3228 = ~(w10513 | w10523);
assign w10524 = v3228;
assign v3229 = ~(w10017 | w10018);
assign w10525 = v3229;
assign v3230 = ~(w10396 | w10525);
assign w10526 = v3230;
assign w10527 = w10396 & w10525;
assign v3231 = ~(w10526 | w10527);
assign w10528 = v3231;
assign w10529 = w10524 & ~w10528;
assign w10530 = ~w10524 & w10528;
assign v3232 = ~(w10529 | w10530);
assign w10531 = v3232;
assign w10532 = w10035 & ~w10393;
assign v3233 = ~(w10394 | w10532);
assign w10533 = v3233;
assign w10534 = w3397 & w9402;
assign w10535 = ~w1609 & w9401;
assign w10536 = ~w1387 & w10419;
assign w10537 = ~w1496 & w9891;
assign v3234 = ~(w10536 | w10537);
assign w10538 = v3234;
assign w10539 = ~w10535 & w10538;
assign w10540 = ~w10534 & w10539;
assign w10541 = pi05 & ~w10540;
assign w10542 = ~pi05 & w10540;
assign v3235 = ~(w10541 | w10542);
assign w10543 = v3235;
assign v3236 = ~(w10533 | w10543);
assign w10544 = v3236;
assign w10545 = w10533 & w10543;
assign w10546 = ~w1674 & w9401;
assign w10547 = ~w3510 & w9402;
assign w10548 = ~w1609 & w9891;
assign w10549 = ~w1496 & w10419;
assign v3237 = ~(w10548 | w10549);
assign w10550 = v3237;
assign w10551 = ~w10547 & w10550;
assign w10552 = ~w10546 & w10551;
assign w10553 = pi05 & w10552;
assign v3238 = ~(pi05 | w10552);
assign w10554 = v3238;
assign v3239 = ~(w10553 | w10554);
assign w10555 = v3239;
assign v3240 = ~(w10048 | w10049);
assign w10556 = v3240;
assign w10557 = w10391 & w10556;
assign v3241 = ~(w10391 | w10556);
assign w10558 = v3241;
assign v3242 = ~(w10557 | w10558);
assign w10559 = v3242;
assign v3243 = ~(w10555 | w10559);
assign w10560 = v3243;
assign w10561 = w10555 & w10559;
assign v3244 = ~(w10560 | w10561);
assign w10562 = v3244;
assign v3245 = ~(w10066 | w10389);
assign w10563 = v3245;
assign v3246 = ~(w10390 | w10563);
assign w10564 = v3246;
assign w10565 = w3494 & w9402;
assign w10566 = ~w1609 & w10419;
assign w10567 = ~w1674 & w9891;
assign v3247 = ~(w10566 | w10567);
assign w10568 = v3247;
assign w10569 = ~w1795 & w9401;
assign w10570 = w10568 & ~w10569;
assign w10571 = ~w10565 & w10570;
assign w10572 = pi05 & ~w10571;
assign w10573 = ~pi05 & w10571;
assign v3248 = ~(w10572 | w10573);
assign w10574 = v3248;
assign v3249 = ~(w10564 | w10574);
assign w10575 = v3249;
assign w10576 = w10564 & w10574;
assign w10577 = w4520 & w9402;
assign w10578 = ~w1795 & w9891;
assign w10579 = ~w1674 & w10419;
assign w10580 = ~w1860 & w9401;
assign v3250 = ~(w10579 | w10580);
assign w10581 = v3250;
assign w10582 = ~w10578 & w10581;
assign w10583 = ~w10577 & w10582;
assign w10584 = pi05 & ~w10583;
assign w10585 = ~pi05 & w10583;
assign v3251 = ~(w10584 | w10585);
assign w10586 = v3251;
assign v3252 = ~(w10079 | w10080);
assign w10587 = v3252;
assign w10588 = w10388 & w10587;
assign v3253 = ~(w10388 | w10587);
assign w10589 = v3253;
assign v3254 = ~(w10588 | w10589);
assign w10590 = v3254;
assign w10591 = w10586 & ~w10590;
assign w10592 = ~w10586 & w10590;
assign v3255 = ~(w10591 | w10592);
assign w10593 = v3255;
assign v3256 = ~(w10095 | w10386);
assign w10594 = v3256;
assign v3257 = ~(w10387 | w10594);
assign w10595 = v3257;
assign w10596 = w4538 & w9402;
assign w10597 = ~w1795 & w10419;
assign w10598 = ~w1860 & w9891;
assign w10599 = ~w1942 & w9401;
assign v3258 = ~(w10598 | w10599);
assign w10600 = v3258;
assign w10601 = ~w10597 & w10600;
assign w10602 = ~w10596 & w10601;
assign w10603 = pi05 & ~w10602;
assign w10604 = ~pi05 & w10602;
assign v3259 = ~(w10603 | w10604);
assign w10605 = v3259;
assign v3260 = ~(w10595 | w10605);
assign w10606 = v3260;
assign w10607 = w10595 & w10605;
assign w10608 = w4854 & w9402;
assign w10609 = ~w1860 & w10419;
assign w10610 = ~w1942 & w9891;
assign w10611 = ~w2038 & w9401;
assign v3261 = ~(w10610 | w10611);
assign w10612 = v3261;
assign w10613 = ~w10609 & w10612;
assign w10614 = ~w10608 & w10613;
assign w10615 = pi05 & ~w10614;
assign w10616 = ~pi05 & w10614;
assign v3262 = ~(w10615 | w10616);
assign w10617 = v3262;
assign v3263 = ~(w10108 | w10109);
assign w10618 = v3263;
assign v3264 = ~(w10385 | w10618);
assign w10619 = v3264;
assign w10620 = w10385 & w10618;
assign v3265 = ~(w10619 | w10620);
assign w10621 = v3265;
assign w10622 = w10617 & ~w10621;
assign w10623 = w10381 & ~w10383;
assign v3266 = ~(w10384 | w10623);
assign w10624 = v3266;
assign w10625 = w4702 & w9402;
assign w10626 = ~w1942 & w10419;
assign w10627 = ~w2038 & w9891;
assign w10628 = ~w2089 & w9401;
assign v3267 = ~(w10627 | w10628);
assign w10629 = v3267;
assign w10630 = ~w10626 & w10629;
assign w10631 = ~w10625 & w10630;
assign w10632 = pi05 & ~w10631;
assign w10633 = ~pi05 & w10631;
assign v3268 = ~(w10632 | w10633);
assign w10634 = v3268;
assign w10635 = w10624 & w10634;
assign w10636 = w10377 & ~w10379;
assign v3269 = ~(w10380 | w10636);
assign w10637 = v3269;
assign w10638 = ~w2202 & w9401;
assign w10639 = w5049 & w9402;
assign w10640 = ~w2089 & w9891;
assign w10641 = ~w2038 & w10419;
assign v3270 = ~(w10640 | w10641);
assign w10642 = v3270;
assign w10643 = ~w10639 & w10642;
assign w10644 = ~w10638 & w10643;
assign w10645 = pi05 & w10644;
assign v3271 = ~(pi05 | w10644);
assign w10646 = v3271;
assign v3272 = ~(w10645 | w10646);
assign w10647 = v3272;
assign w10648 = w10637 & ~w10647;
assign w10649 = w10373 & ~w10375;
assign v3273 = ~(w10376 | w10649);
assign w10650 = v3273;
assign w10651 = w5033 & w9402;
assign w10652 = ~w2202 & w9891;
assign w10653 = ~w2089 & w10419;
assign v3274 = ~(w10652 | w10653);
assign w10654 = v3274;
assign w10655 = ~w2290 & w9401;
assign w10656 = w10654 & ~w10655;
assign w10657 = ~w10651 & w10656;
assign w10658 = pi05 & w10657;
assign v3275 = ~(pi05 | w10657);
assign w10659 = v3275;
assign v3276 = ~(w10658 | w10659);
assign w10660 = v3276;
assign w10661 = w10650 & ~w10660;
assign w10662 = w10369 & ~w10371;
assign v3277 = ~(w10372 | w10662);
assign w10663 = v3277;
assign w10664 = w5262 & w9402;
assign w10665 = ~w2202 & w10419;
assign w10666 = ~w2339 & w9401;
assign w10667 = ~w2290 & w9891;
assign v3278 = ~(w10666 | w10667);
assign w10668 = v3278;
assign w10669 = ~w10665 & w10668;
assign w10670 = ~w10664 & w10669;
assign w10671 = pi05 & ~w10670;
assign w10672 = ~pi05 & w10670;
assign v3279 = ~(w10671 | w10672);
assign w10673 = v3279;
assign w10674 = w10663 & w10673;
assign w10675 = w10365 & ~w10367;
assign v3280 = ~(w10368 | w10675);
assign w10676 = v3280;
assign w10677 = w5280 & w9402;
assign w10678 = ~w2290 & w10419;
assign w10679 = ~w2339 & w9891;
assign w10680 = ~w2424 & w9401;
assign v3281 = ~(w10679 | w10680);
assign w10681 = v3281;
assign w10682 = ~w10678 & w10681;
assign w10683 = ~w10677 & w10682;
assign w10684 = pi05 & ~w10683;
assign w10685 = ~pi05 & w10683;
assign v3282 = ~(w10684 | w10685);
assign w10686 = v3282;
assign w10687 = w10676 & w10686;
assign w10688 = w10361 & ~w10363;
assign v3283 = ~(w10364 | w10688);
assign w10689 = v3283;
assign w10690 = w5665 & w9402;
assign w10691 = ~w2492 & w9401;
assign w10692 = ~w2424 & w9891;
assign w10693 = ~w2339 & w10419;
assign v3284 = ~(w10692 | w10693);
assign w10694 = v3284;
assign w10695 = ~w10691 & w10694;
assign w10696 = ~w10690 & w10695;
assign w10697 = pi05 & ~w10696;
assign w10698 = ~pi05 & w10696;
assign v3285 = ~(w10697 | w10698);
assign w10699 = v3285;
assign w10700 = w10689 & w10699;
assign w10701 = w10357 & ~w10359;
assign v3286 = ~(w10360 | w10701);
assign w10702 = v3286;
assign w10703 = w5449 & w9402;
assign w10704 = ~w2424 & w10419;
assign w10705 = ~w2492 & w9891;
assign w10706 = ~w2568 & w9401;
assign v3287 = ~(w10705 | w10706);
assign w10707 = v3287;
assign w10708 = ~w10704 & w10707;
assign w10709 = ~w10703 & w10708;
assign w10710 = pi05 & ~w10709;
assign w10711 = ~pi05 & w10709;
assign v3288 = ~(w10710 | w10711);
assign w10712 = v3288;
assign w10713 = w10702 & w10712;
assign w10714 = w10353 & ~w10355;
assign v3289 = ~(w10356 | w10714);
assign w10715 = v3289;
assign w10716 = w5898 & w9402;
assign w10717 = ~w2568 & w9891;
assign w10718 = ~w2596 & w9401;
assign w10719 = ~w2492 & w10419;
assign v3290 = ~(w10718 | w10719);
assign w10720 = v3290;
assign w10721 = ~w10717 & w10720;
assign w10722 = ~w10716 & w10721;
assign w10723 = pi05 & ~w10722;
assign w10724 = ~pi05 & w10722;
assign v3291 = ~(w10723 | w10724);
assign w10725 = v3291;
assign w10726 = w10715 & w10725;
assign w10727 = w10349 & ~w10351;
assign v3292 = ~(w10352 | w10727);
assign w10728 = v3292;
assign w10729 = w6031 & w9402;
assign w10730 = ~w2568 & w10419;
assign w10731 = ~w2596 & w9891;
assign v3293 = ~(w10730 | w10731);
assign w10732 = v3293;
assign w10733 = ~w2669 & w9401;
assign w10734 = w10732 & ~w10733;
assign w10735 = ~w10729 & w10734;
assign w10736 = pi05 & ~w10735;
assign w10737 = ~pi05 & w10735;
assign v3294 = ~(w10736 | w10737);
assign w10738 = v3294;
assign w10739 = w10728 & w10738;
assign w10740 = w10345 & ~w10347;
assign v3295 = ~(w10348 | w10740);
assign w10741 = v3295;
assign w10742 = w5880 & w9402;
assign w10743 = ~w2669 & w9891;
assign w10744 = ~w2724 & w9401;
assign w10745 = ~w2596 & w10419;
assign v3296 = ~(w10744 | w10745);
assign w10746 = v3296;
assign w10747 = ~w10743 & w10746;
assign w10748 = ~w10742 & w10747;
assign w10749 = pi05 & ~w10748;
assign w10750 = ~pi05 & w10748;
assign v3297 = ~(w10749 | w10750);
assign w10751 = v3297;
assign w10752 = w10741 & w10751;
assign w10753 = w10341 & ~w10343;
assign v3298 = ~(w10344 | w10753);
assign w10754 = v3298;
assign w10755 = ~w2669 & w10419;
assign w10756 = w6148 & w9402;
assign w10757 = ~w2724 & w9891;
assign w10758 = ~w2811 & w9401;
assign v3299 = ~(w10757 | w10758);
assign w10759 = v3299;
assign w10760 = ~w10756 & w10759;
assign w10761 = ~w10755 & w10760;
assign w10762 = pi05 & w10761;
assign v3300 = ~(pi05 | w10761);
assign w10763 = v3300;
assign v3301 = ~(w10762 | w10763);
assign w10764 = v3301;
assign w10765 = w10754 & ~w10764;
assign w10766 = w10337 & ~w10339;
assign v3302 = ~(w10340 | w10766);
assign w10767 = v3302;
assign w10768 = ~w6447 & w9402;
assign w10769 = ~w2724 & w10419;
assign w10770 = ~w2811 & w9891;
assign v3303 = ~(w10769 | w10770);
assign w10771 = v3303;
assign w10772 = ~w2846 & w9401;
assign w10773 = w10771 & ~w10772;
assign w10774 = ~w10768 & w10773;
assign w10775 = ~pi05 & w10774;
assign w10776 = pi05 & ~w10774;
assign v3304 = ~(w10775 | w10776);
assign w10777 = v3304;
assign w10778 = w10767 & w10777;
assign w10779 = w10333 & ~w10335;
assign v3305 = ~(w10336 | w10779);
assign w10780 = v3305;
assign w10781 = w6459 & w9402;
assign w10782 = ~w2846 & w9891;
assign w10783 = ~w2811 & w10419;
assign w10784 = ~w2937 & w9401;
assign v3306 = ~(w10783 | w10784);
assign w10785 = v3306;
assign w10786 = ~w10782 & w10785;
assign w10787 = ~w10781 & w10786;
assign w10788 = pi05 & ~w10787;
assign w10789 = ~pi05 & w10787;
assign v3307 = ~(w10788 | w10789);
assign w10790 = v3307;
assign w10791 = w10780 & w10790;
assign w10792 = w10329 & ~w10331;
assign v3308 = ~(w10332 | w10792);
assign w10793 = v3308;
assign w10794 = ~w6129 & w29266;
assign w10795 = ~w2846 & w10419;
assign w10796 = ~w3000 & w9401;
assign w10797 = ~w2937 & w9891;
assign v3309 = ~(w10796 | w10797);
assign w10798 = v3309;
assign w10799 = ~w10795 & w10798;
assign w10800 = ~w10794 & w10799;
assign w10801 = pi05 & ~w10800;
assign w10802 = ~pi05 & w10800;
assign v3310 = ~(w10801 | w10802);
assign w10803 = v3310;
assign w10804 = w10793 & w10803;
assign w10805 = w10325 & ~w10327;
assign v3311 = ~(w10328 | w10805);
assign w10806 = v3311;
assign w10807 = ~w2937 & w10419;
assign w10808 = ~w3068 & w9401;
assign v3312 = ~(w10807 | w10808);
assign w10809 = v3312;
assign w10810 = ~w3000 & w9891;
assign w10811 = w10809 & ~w10810;
assign w10812 = (w10811 & w6505) | (w10811 & w28713) | (w6505 & w28713);
assign v3313 = ~(pi05 | w10812);
assign w10813 = v3313;
assign w10814 = pi05 & w10812;
assign v3314 = ~(w10813 | w10814);
assign w10815 = v3314;
assign w10816 = w10806 & ~w10815;
assign w10817 = ~w10316 & w10323;
assign v3315 = ~(w10324 | w10817);
assign w10818 = v3315;
assign w10819 = ~w3000 & w10419;
assign w10820 = ~w3068 & w9891;
assign v3316 = ~(w10819 | w10820);
assign w10821 = v3316;
assign w10822 = ~w3124 & w9401;
assign w10823 = w10821 & ~w10822;
assign w10824 = (~w6551 & w28714) | (~w6551 & w28715) | (w28714 & w28715);
assign w10825 = (w6551 & w28716) | (w6551 & w28717) | (w28716 & w28717);
assign v3317 = ~(w10824 | w10825);
assign w10826 = v3317;
assign w10827 = w10818 & ~w10826;
assign w10828 = w6603 & w10445;
assign w10829 = ~w3162 & w9401;
assign w10830 = (w9891 & ~w3112) | (w9891 & w28494) | (~w3112 & w28494);
assign w10831 = ~w3068 & w10419;
assign v3318 = ~(w10830 | w10831);
assign w10832 = v3318;
assign w10833 = w10832 & w28495;
assign w10834 = (pi05 & ~w10832) | (pi05 & w28496) | (~w10832 & w28496);
assign v3319 = ~(w10833 | w10834);
assign w10835 = v3319;
assign w10836 = (~w10835 & ~w6603) | (~w10835 & w28286) | (~w6603 & w28286);
assign v3320 = ~(w10828 | w10836);
assign w10837 = v3320;
assign w10838 = pi08 & ~w10312;
assign w10839 = ~w10304 & w10838;
assign w10840 = w10304 & ~w10838;
assign v3321 = ~(w10839 | w10840);
assign w10841 = v3321;
assign w10842 = w10837 & w10841;
assign w10843 = (w9401 & ~w3331) | (w9401 & w28287) | (~w3331 & w28287);
assign w10844 = (w10419 & ~w3210) | (w10419 & w28497) | (~w3210 & w28497);
assign w10845 = (w9891 & ~w3261) | (w9891 & w28288) | (~w3261 & w28288);
assign v3322 = ~(w10844 | w10845);
assign w10846 = v3322;
assign w10847 = (~w6676 & w28162) | (~w6676 & w28163) | (w28162 & w28163);
assign w10848 = ~w3332 & w9396;
assign w10849 = ~w7309 & w9402;
assign w10850 = (w10419 & ~w3261) | (w10419 & w28164) | (~w3261 & w28164);
assign w10851 = (w9891 & ~w3331) | (w9891 & w28165) | (~w3331 & w28165);
assign v3323 = ~(w10850 | w10851);
assign w10852 = v3323;
assign w10853 = (w10852 & w7309) | (w10852 & w28289) | (w7309 & w28289);
assign w10854 = ~w10849 & w28166;
assign w10855 = w10847 & w10854;
assign w10856 = w10310 & w10855;
assign v3324 = ~(w10310 | w10855);
assign w10857 = v3324;
assign v3325 = ~(w10856 | w10857);
assign w10858 = v3325;
assign w10859 = w6735 & w10445;
assign w10860 = w6735 & w10447;
assign w10861 = ~w3162 & w10419;
assign w10862 = ~w3211 & w9891;
assign w10863 = (w9401 & ~w3261) | (w9401 & w28290) | (~w3261 & w28290);
assign v3326 = ~(w10862 | w10863);
assign w10864 = v3326;
assign w10865 = w10864 & w28291;
assign w10866 = (~pi05 & ~w10864) | (~pi05 & w28292) | (~w10864 & w28292);
assign v3327 = ~(w10865 | w10866);
assign w10867 = v3327;
assign w10868 = ~w10860 & w10867;
assign v3328 = ~(w10859 | w10868);
assign w10869 = v3328;
assign w10870 = w10858 & w10869;
assign v3329 = ~(w10856 | w10870);
assign w10871 = v3329;
assign w10872 = ~w3162 & w9891;
assign w10873 = ~w3211 & w9401;
assign w10874 = ~w3124 & w10419;
assign v3330 = ~(w10873 | w10874);
assign w10875 = v3330;
assign w10876 = ~w10872 & w10875;
assign w10877 = (w10876 & w6641) | (w10876 & w28293) | (w6641 & w28293);
assign w10878 = w7308 & w9920;
assign w10879 = pi08 & w10310;
assign w10880 = ~w10307 & w10879;
assign w10881 = (~w10880 & w10308) | (~w10880 & w28167) | (w10308 & w28167);
assign w10882 = ~w10878 & w10881;
assign w10883 = (pi05 & ~w10881) | (pi05 & w28168) | (~w10881 & w28168);
assign w10884 = w10881 & w28169;
assign v3331 = ~(w10883 | w10884);
assign w10885 = v3331;
assign w10886 = w10877 & ~w10885;
assign w10887 = ~w10877 & w10885;
assign v3332 = ~(w10886 | w10887);
assign w10888 = v3332;
assign v3333 = ~(w10871 | w10888);
assign w10889 = v3333;
assign w10890 = w10882 & w10888;
assign v3334 = ~(w10889 | w10890);
assign w10891 = v3334;
assign v3335 = ~(w10837 | w10841);
assign w10892 = v3335;
assign v3336 = ~(w10842 | w10892);
assign w10893 = v3336;
assign w10894 = ~w10891 & w10893;
assign w10895 = (~w10842 & w10891) | (~w10842 & w28294) | (w10891 & w28294);
assign w10896 = ~w10818 & w10826;
assign v3337 = ~(w10827 | w10896);
assign w10897 = v3337;
assign w10898 = ~w10895 & w10897;
assign w10899 = (~w10827 & w10895) | (~w10827 & w28498) | (w10895 & w28498);
assign w10900 = ~w10806 & w10815;
assign v3338 = ~(w10816 | w10900);
assign w10901 = v3338;
assign w10902 = ~w10899 & w10901;
assign v3339 = ~(w10816 | w10902);
assign w10903 = v3339;
assign v3340 = ~(w10793 | w10803);
assign w10904 = v3340;
assign v3341 = ~(w10804 | w10904);
assign w10905 = v3341;
assign w10906 = ~w10903 & w10905;
assign w10907 = (~w10804 & w10903) | (~w10804 & w28718) | (w10903 & w28718);
assign v3342 = ~(w10780 | w10790);
assign w10908 = v3342;
assign v3343 = ~(w10791 | w10908);
assign w10909 = v3343;
assign w10910 = ~w10907 & w10909;
assign v3344 = ~(w10791 | w10910);
assign w10911 = v3344;
assign v3345 = ~(w10767 | w10777);
assign w10912 = v3345;
assign v3346 = ~(w10778 | w10912);
assign w10913 = v3346;
assign w10914 = ~w10911 & w10913;
assign w10915 = (~w10778 & w10911) | (~w10778 & w28719) | (w10911 & w28719);
assign w10916 = ~w10754 & w10764;
assign v3347 = ~(w10765 | w10916);
assign w10917 = v3347;
assign w10918 = ~w10915 & w10917;
assign w10919 = (~w10765 & ~w10917) | (~w10765 & w28720) | (~w10917 & w28720);
assign v3348 = ~(w10741 | w10751);
assign w10920 = v3348;
assign v3349 = ~(w10752 | w10920);
assign w10921 = v3349;
assign w10922 = ~w10919 & w10921;
assign w10923 = (~w10752 & w10919) | (~w10752 & w29267) | (w10919 & w29267);
assign v3350 = ~(w10728 | w10738);
assign w10924 = v3350;
assign v3351 = ~(w10739 | w10924);
assign w10925 = v3351;
assign w10926 = ~w10923 & w10925;
assign v3352 = ~(w10739 | w10926);
assign w10927 = v3352;
assign v3353 = ~(w10715 | w10725);
assign w10928 = v3353;
assign v3354 = ~(w10726 | w10928);
assign w10929 = v3354;
assign w10930 = ~w10927 & w10929;
assign w10931 = (~w10726 & w10927) | (~w10726 & w29487) | (w10927 & w29487);
assign v3355 = ~(w10702 | w10712);
assign w10932 = v3355;
assign v3356 = ~(w10713 | w10932);
assign w10933 = v3356;
assign w10934 = ~w10931 & w10933;
assign v3357 = ~(w10713 | w10934);
assign w10935 = v3357;
assign v3358 = ~(w10689 | w10699);
assign w10936 = v3358;
assign v3359 = ~(w10700 | w10936);
assign w10937 = v3359;
assign w10938 = ~w10935 & w10937;
assign w10939 = (~w10700 & w10935) | (~w10700 & w29666) | (w10935 & w29666);
assign v3360 = ~(w10676 | w10686);
assign w10940 = v3360;
assign v3361 = ~(w10687 | w10940);
assign w10941 = v3361;
assign w10942 = ~w10939 & w10941;
assign v3362 = ~(w10687 | w10942);
assign w10943 = v3362;
assign v3363 = ~(w10663 | w10673);
assign w10944 = v3363;
assign v3364 = ~(w10674 | w10944);
assign w10945 = v3364;
assign w10946 = ~w10943 & w10945;
assign w10947 = (~w10674 & w10943) | (~w10674 & w29860) | (w10943 & w29860);
assign w10948 = ~w10650 & w10660;
assign v3365 = ~(w10661 | w10948);
assign w10949 = v3365;
assign w10950 = ~w10947 & w10949;
assign v3366 = ~(w10661 | w10950);
assign w10951 = v3366;
assign w10952 = ~w10637 & w10647;
assign v3367 = ~(w10648 | w10952);
assign w10953 = v3367;
assign w10954 = ~w10951 & w10953;
assign w10955 = (~w10648 & w10951) | (~w10648 & w30026) | (w10951 & w30026);
assign v3368 = ~(w10624 | w10634);
assign w10956 = v3368;
assign v3369 = ~(w10635 | w10956);
assign w10957 = v3369;
assign w10958 = ~w10955 & w10957;
assign v3370 = ~(w10635 | w10958);
assign w10959 = v3370;
assign w10960 = ~w10617 & w10621;
assign v3371 = ~(w10622 | w10960);
assign w10961 = v3371;
assign w10962 = ~w10959 & w10961;
assign w10963 = (~w10622 & w10959) | (~w10622 & w30159) | (w10959 & w30159);
assign w10964 = (~w10606 & ~w10963) | (~w10606 & w28170) | (~w10963 & w28170);
assign w10965 = w10593 & w10964;
assign w10966 = (~w10591 & ~w10593) | (~w10591 & w28171) | (~w10593 & w28171);
assign w10967 = (w28171 & w30333) | (w28171 & w30334) | (w30333 & w30334);
assign v3372 = ~(w10575 | w10967);
assign w10968 = v3372;
assign w10969 = w10562 & w10968;
assign w10970 = (~w10560 & ~w10562) | (~w10560 & w28172) | (~w10562 & w28172);
assign w10971 = (w28172 & w30611) | (w28172 & w30612) | (w30611 & w30612);
assign w10972 = (~w10544 & ~w10970) | (~w10544 & w30335) | (~w10970 & w30335);
assign w10973 = w10531 & w10972;
assign w10974 = (~w10529 & ~w10531) | (~w10529 & w28173) | (~w10531 & w28173);
assign w10975 = (~w10511 & ~w10974) | (~w10511 & w28721) | (~w10974 & w28721);
assign w10976 = w10496 & w10975;
assign w10977 = (~w10494 & ~w10496) | (~w10494 & w28174) | (~w10496 & w28174);
assign w10978 = (~w10478 & ~w10977) | (~w10478 & w29861) | (~w10977 & w29861);
assign w10979 = w10465 & w10978;
assign w10980 = (~w10463 & ~w10465) | (~w10463 & w28175) | (~w10465 & w28175);
assign v3373 = ~(w10434 | w10443);
assign w10981 = v3373;
assign v3374 = ~(w10444 | w10981);
assign w10982 = v3374;
assign w10983 = ~w10980 & w10982;
assign w10984 = (~w10444 & w10980) | (~w10444 & w31028) | (w10980 & w31028);
assign w10985 = (w4147 & w29667) | (w4147 & w29668) | (w29667 & w29668);
assign v3375 = ~(pi00 | pi01);
assign w10986 = v3375;
assign w10987 = pi02 & w10986;
assign w10988 = ~pi02 & w4;
assign v3376 = ~(w1 | w10988);
assign w10989 = v3376;
assign w10990 = (w4145 & w29669) | (w4145 & w29670) | (w29669 & w29670);
assign v3377 = ~(w10987 | w10990);
assign w10991 = v3377;
assign v3378 = ~(w4191 | w10991);
assign w10992 = v3378;
assign v3379 = ~(w10985 | w10992);
assign w10993 = v3379;
assign w10994 = ~w4082 & w10419;
assign w10995 = ~w4134 & w9401;
assign w10996 = ~w4035 & w9891;
assign v3380 = ~(w10995 | w10996);
assign w10997 = v3380;
assign w10998 = ~w10994 & w10997;
assign w10999 = (~w4149 & w28726) | (~w4149 & w28727) | (w28726 & w28727);
assign w11000 = (w4149 & w28728) | (w4149 & w28729) | (w28728 & w28729);
assign v3381 = ~(w10999 | w11000);
assign w11001 = v3381;
assign w11002 = w10993 & w11001;
assign v3382 = ~(w10993 | w11001);
assign w11003 = v3382;
assign v3383 = ~(w11002 | w11003);
assign w11004 = v3383;
assign v3384 = ~(w10408 | w10410);
assign w11005 = v3384;
assign v3385 = ~(w10411 | w11005);
assign w11006 = v3385;
assign w11007 = w11004 & ~w11006;
assign w11008 = ~w11004 & w11006;
assign v3386 = ~(w11007 | w11008);
assign w11009 = v3386;
assign w11010 = ~w10984 & w11009;
assign v3387 = ~(w10417 | w10427);
assign w11011 = v3387;
assign v3388 = ~(w10428 | w11011);
assign w11012 = v3388;
assign v3389 = ~(w11002 | w11007);
assign w11013 = v3389;
assign v3390 = ~(w11012 | w11013);
assign w11014 = v3390;
assign w11015 = w11012 & w11013;
assign v3391 = ~(w11014 | w11015);
assign w11016 = v3391;
assign w11017 = w11010 & ~w11016;
assign w11018 = ~w11010 & w11016;
assign w11019 = w10984 & ~w11009;
assign v3392 = ~(w11010 | w11019);
assign w11020 = v3392;
assign w11021 = w10980 & ~w10982;
assign v3393 = ~(w10983 | w11021);
assign w11022 = v3393;
assign w11023 = ~pi00 & pi01;
assign w11024 = ~w4191 & w11023;
assign w11025 = (w4425 & w28730) | (w4425 & w28731) | (w28730 & w28731);
assign w11026 = ~w4082 & w10986;
assign w11027 = pi02 & ~w11026;
assign w11028 = (~w4425 & w28732) | (~w4425 & w28733) | (w28732 & w28733);
assign v3394 = ~(w11025 | w11028);
assign w11029 = v3394;
assign w11030 = ~w11022 & w11029;
assign v3395 = ~(w10465 | w10978);
assign w11031 = v3395;
assign v3396 = ~(w10979 | w11031);
assign w11032 = v3396;
assign w11033 = ~w4082 & w11023;
assign w11034 = pi00 & ~w2;
assign w11035 = ~w0 & w11034;
assign w11036 = ~w4191 & w11035;
assign v3397 = ~(w11033 | w11036);
assign w11037 = v3397;
assign w11038 = (w4196 & w28734) | (w4196 & w28735) | (w28734 & w28735);
assign w11039 = ~w4035 & w10986;
assign w11040 = pi02 & ~w11039;
assign w11041 = (~w4196 & w28736) | (~w4196 & w28737) | (w28736 & w28737);
assign v3398 = ~(w11038 | w11041);
assign w11042 = v3398;
assign w11043 = w11032 & ~w11042;
assign w11044 = ~w11032 & w11042;
assign v3399 = ~(w11043 | w11044);
assign w11045 = v3399;
assign v3400 = ~(w10478 | w10479);
assign w11046 = v3400;
assign v3401 = ~(w10977 | w11046);
assign w11047 = v3401;
assign w11048 = w10977 & w11046;
assign v3402 = ~(w11047 | w11048);
assign w11049 = v3402;
assign w11050 = ~w4035 & w11023;
assign w11051 = ~w4082 & w11035;
assign v3403 = ~(w11050 | w11051);
assign w11052 = v3403;
assign w11053 = (~w4149 & w29268) | (~w4149 & w29269) | (w29268 & w29269);
assign w11054 = ~w4134 & w10986;
assign w11055 = pi02 & ~w11054;
assign w11056 = (w4149 & w29270) | (w4149 & w29271) | (w29270 & w29271);
assign v3404 = ~(w11053 | w11056);
assign w11057 = v3404;
assign v3405 = ~(w11049 | w11057);
assign w11058 = v3405;
assign w11059 = w11049 & w11057;
assign v3406 = ~(w11058 | w11059);
assign w11060 = v3406;
assign v3407 = ~(w10496 | w10975);
assign w11061 = v3407;
assign v3408 = ~(w10976 | w11061);
assign w11062 = v3408;
assign w11063 = ~w4035 & w11035;
assign w11064 = ~w4134 & w11023;
assign v3409 = ~(w11063 | w11064);
assign w11065 = v3409;
assign w11066 = (w4405 & w29671) | (w4405 & w29672) | (w29671 & w29672);
assign w11067 = ~w3920 & w10986;
assign w11068 = pi02 & ~w11067;
assign w11069 = (~w4405 & w29673) | (~w4405 & w29674) | (w29673 & w29674);
assign v3410 = ~(w11066 | w11069);
assign w11070 = v3410;
assign w11071 = w11062 & ~w11070;
assign w11072 = ~w11062 & w11070;
assign w11073 = ~w4134 & w11035;
assign w11074 = ~w3920 & w11023;
assign v3411 = ~(w11073 | w11074);
assign w11075 = v3411;
assign w11076 = (w4309 & w29675) | (w4309 & w29676) | (w29675 & w29676);
assign w11077 = ~w3752 & w10986;
assign w11078 = pi02 & ~w11077;
assign w11079 = (~w4309 & w29677) | (~w4309 & w29678) | (w29677 & w29678);
assign v3412 = ~(w11076 | w11079);
assign w11080 = v3412;
assign v3413 = ~(w10511 | w10512);
assign w11081 = v3413;
assign v3414 = ~(w10974 | w11081);
assign w11082 = v3414;
assign w11083 = w10974 & w11081;
assign v3415 = ~(w11082 | w11083);
assign w11084 = v3415;
assign v3416 = ~(w11080 | w11084);
assign w11085 = v3416;
assign w11086 = w11080 & w11084;
assign v3417 = ~(w11085 | w11086);
assign w11087 = v3417;
assign w11088 = ~w3920 & w11035;
assign w11089 = ~w3752 & w11023;
assign v3418 = ~(w11088 | w11089);
assign w11090 = v3418;
assign w11091 = (~w3928 & w29679) | (~w3928 & w29680) | (w29679 & w29680);
assign w11092 = ~w3587 & w10986;
assign w11093 = pi02 & ~w11092;
assign w11094 = (w3928 & w29681) | (w3928 & w29682) | (w29681 & w29682);
assign v3419 = ~(w11091 | w11094);
assign w11095 = v3419;
assign v3420 = ~(w10531 | w10972);
assign w11096 = v3420;
assign v3421 = ~(w10973 | w11096);
assign w11097 = v3421;
assign w11098 = ~w11095 & w11097;
assign w11099 = w11095 & ~w11097;
assign v3422 = ~(w10544 | w10545);
assign w11100 = v3422;
assign v3423 = ~(w10970 | w11100);
assign w11101 = v3423;
assign w11102 = w10970 & w11100;
assign v3424 = ~(w11101 | w11102);
assign w11103 = v3424;
assign w11104 = ~w3587 & w11023;
assign w11105 = ~w3752 & w11035;
assign v3425 = ~(w11104 | w11105);
assign w11106 = v3425;
assign w11107 = (w3758 & w29683) | (w3758 & w29684) | (w29683 & w29684);
assign w11108 = ~w3666 & w10986;
assign w11109 = pi02 & ~w11108;
assign w11110 = (~w3758 & w29685) | (~w3758 & w29686) | (w29685 & w29686);
assign v3426 = ~(w11107 | w11110);
assign w11111 = v3426;
assign v3427 = ~(w11103 | w11111);
assign w11112 = v3427;
assign w11113 = w11103 & w11111;
assign v3428 = ~(w10562 | w10968);
assign w11114 = v3428;
assign v3429 = ~(w10969 | w11114);
assign w11115 = v3429;
assign w11116 = ~w3666 & w11023;
assign w11117 = ~w3587 & w11035;
assign v3430 = ~(w11116 | w11117);
assign w11118 = v3430;
assign w11119 = (w4291 & w29687) | (w4291 & w29688) | (w29687 & w29688);
assign w11120 = ~w1387 & w10986;
assign w11121 = pi02 & ~w11120;
assign w11122 = (~w4291 & w29689) | (~w4291 & w29690) | (w29689 & w29690);
assign v3431 = ~(w11119 | w11122);
assign w11123 = v3431;
assign w11124 = w11115 & ~w11123;
assign w11125 = ~w11115 & w11123;
assign w11126 = ~w3666 & w11035;
assign w11127 = ~w1387 & w11023;
assign v3432 = ~(w11126 | w11127);
assign w11128 = v3432;
assign w11129 = (w3843 & w29691) | (w3843 & w29692) | (w29691 & w29692);
assign w11130 = ~w1496 & w10986;
assign w11131 = pi02 & ~w11130;
assign w11132 = (~w3843 & w29693) | (~w3843 & w29694) | (w29693 & w29694);
assign v3433 = ~(w11129 | w11132);
assign w11133 = v3433;
assign v3434 = ~(w10575 | w10576);
assign w11134 = v3434;
assign w11135 = w10966 & w11134;
assign v3435 = ~(w10966 | w11134);
assign w11136 = v3435;
assign v3436 = ~(w11135 | w11136);
assign w11137 = v3436;
assign w11138 = w11133 & w11137;
assign w11139 = ~w1496 & w11023;
assign w11140 = ~w1387 & w11035;
assign v3437 = ~(w11139 | w11140);
assign w11141 = v3437;
assign w11142 = (w3397 & w29695) | (w3397 & w29696) | (w29695 & w29696);
assign w11143 = ~w1609 & w10986;
assign w11144 = pi02 & ~w11143;
assign w11145 = (~w3397 & w29697) | (~w3397 & w29698) | (w29697 & w29698);
assign v3438 = ~(w11142 | w11145);
assign w11146 = v3438;
assign v3439 = ~(w10593 | w10964);
assign w11147 = v3439;
assign v3440 = ~(w10965 | w11147);
assign w11148 = v3440;
assign w11149 = w11146 & ~w11148;
assign w11150 = ~w11146 & w11148;
assign w11151 = ~w1609 & w11023;
assign w11152 = ~w1496 & w11035;
assign v3441 = ~(w11151 | w11152);
assign w11153 = v3441;
assign w11154 = (~w3510 & w29699) | (~w3510 & w29700) | (w29699 & w29700);
assign w11155 = ~w1674 & w10986;
assign w11156 = pi02 & ~w11155;
assign w11157 = (w3510 & w29701) | (w3510 & w29702) | (w29701 & w29702);
assign v3442 = ~(w11154 | w11157);
assign w11158 = v3442;
assign v3443 = ~(w10606 | w10607);
assign w11159 = v3443;
assign v3444 = ~(w10963 | w11159);
assign w11160 = v3444;
assign w11161 = w10963 & w11159;
assign v3445 = ~(w11160 | w11161);
assign w11162 = v3445;
assign w11163 = w11158 & w11162;
assign w11164 = w10955 & ~w10957;
assign v3446 = ~(w10958 | w11164);
assign w11165 = v3446;
assign w11166 = ~w1795 & w11023;
assign w11167 = ~w1674 & w11035;
assign v3447 = ~(w11166 | w11167);
assign w11168 = v3447;
assign w11169 = (w11168 & ~w4520) | (w11168 & w29703) | (~w4520 & w29703);
assign v3448 = ~(pi02 | w11169);
assign w11170 = v3448;
assign w11171 = ~w1860 & w10986;
assign w11172 = pi02 & ~w11171;
assign w11173 = w11169 & w11172;
assign v3449 = ~(w11170 | w11173);
assign w11174 = v3449;
assign w11175 = w11165 & ~w11174;
assign w11176 = ~w11165 & w11174;
assign w11177 = w10951 & ~w10953;
assign v3450 = ~(w10954 | w11177);
assign w11178 = v3450;
assign w11179 = ~w1795 & w11035;
assign w11180 = ~w1860 & w11023;
assign v3451 = ~(w11179 | w11180);
assign w11181 = v3451;
assign w11182 = (w11181 & ~w4538) | (w11181 & w29704) | (~w4538 & w29704);
assign w11183 = pi02 & ~w11182;
assign w11184 = ~w1942 & w10986;
assign w11185 = pi02 & ~w11184;
assign w11186 = w11182 & ~w11185;
assign v3452 = ~(w11183 | w11186);
assign w11187 = v3452;
assign w11188 = w11178 & w11187;
assign w11189 = ~w1942 & w11023;
assign w11190 = ~w1860 & w11035;
assign v3453 = ~(w11189 | w11190);
assign w11191 = v3453;
assign w11192 = (w11191 & ~w4854) | (w11191 & w29705) | (~w4854 & w29705);
assign v3454 = ~(pi02 | w11192);
assign w11193 = v3454;
assign w11194 = ~w2038 & w10986;
assign w11195 = pi02 & ~w11194;
assign w11196 = w11192 & w11195;
assign v3455 = ~(w11193 | w11196);
assign w11197 = v3455;
assign w11198 = w10947 & ~w10949;
assign v3456 = ~(w10950 | w11198);
assign w11199 = v3456;
assign w11200 = ~w11197 & w11199;
assign w11201 = w11197 & ~w11199;
assign w11202 = ~w1942 & w11035;
assign w11203 = ~w2038 & w11023;
assign v3457 = ~(w11202 | w11203);
assign w11204 = v3457;
assign w11205 = (w11204 & ~w4702) | (w11204 & w29706) | (~w4702 & w29706);
assign v3458 = ~(pi02 | w11205);
assign w11206 = v3458;
assign w11207 = ~w2089 & w10986;
assign w11208 = pi02 & ~w11207;
assign w11209 = w11205 & w11208;
assign v3459 = ~(w11206 | w11209);
assign w11210 = v3459;
assign w11211 = w10943 & ~w10945;
assign v3460 = ~(w10946 | w11211);
assign w11212 = v3460;
assign w11213 = w11210 & ~w11212;
assign w11214 = ~w2202 & w10987;
assign w11215 = ~w2089 & w11023;
assign w11216 = ~w2038 & w11035;
assign v3461 = ~(w11215 | w11216);
assign w11217 = v3461;
assign w11218 = ~w11214 & w11217;
assign w11219 = (w11218 & ~w5049) | (w11218 & w29707) | (~w5049 & w29707);
assign w11220 = pi02 & ~w11219;
assign w11221 = ~pi02 & w11219;
assign v3462 = ~(w11220 | w11221);
assign w11222 = v3462;
assign w11223 = w10939 & ~w10941;
assign v3463 = ~(w10942 | w11223);
assign w11224 = v3463;
assign v3464 = ~(w11222 | w11224);
assign w11225 = v3464;
assign w11226 = w10931 & ~w10933;
assign v3465 = ~(w10934 | w11226);
assign w11227 = v3465;
assign w11228 = w10927 & ~w10929;
assign v3466 = ~(w10930 | w11228);
assign w11229 = v3466;
assign w11230 = ~w4 & w5280;
assign w11231 = ~w2339 & w11023;
assign w11232 = ~w2290 & w11035;
assign v3467 = ~(w11231 | w11232);
assign w11233 = v3467;
assign w11234 = ~w11230 & w11233;
assign w11235 = pi02 & ~w11234;
assign w11236 = ~w2424 & w10986;
assign w11237 = pi02 & ~w11236;
assign w11238 = w11234 & ~w11237;
assign v3468 = ~(w11235 | w11238);
assign w11239 = v3468;
assign v3469 = ~(w11229 | w11239);
assign w11240 = v3469;
assign w11241 = w10923 & ~w10925;
assign v3470 = ~(w10926 | w11241);
assign w11242 = v3470;
assign w11243 = ~w4 & w5665;
assign w11244 = ~w2492 & w10987;
assign w11245 = ~w2339 & w11035;
assign v3471 = ~(w11244 | w11245);
assign w11246 = v3471;
assign w11247 = ~w2424 & w11023;
assign w11248 = w11246 & ~w11247;
assign w11249 = ~w11243 & w11248;
assign w11250 = ~pi02 & w11249;
assign w11251 = pi02 & ~w11249;
assign v3472 = ~(w11250 | w11251);
assign w11252 = v3472;
assign w11253 = w11242 & w11252;
assign v3473 = ~(w11242 | w11252);
assign w11254 = v3473;
assign w11255 = ~w4 & w5449;
assign w11256 = ~w2568 & w10987;
assign w11257 = ~w2492 & w11023;
assign w11258 = ~w2424 & w11035;
assign v3474 = ~(w11257 | w11258);
assign w11259 = v3474;
assign w11260 = ~w11256 & w11259;
assign w11261 = ~w11255 & w11260;
assign w11262 = pi02 & ~w11261;
assign w11263 = ~pi02 & w11261;
assign v3475 = ~(w11262 | w11263);
assign w11264 = v3475;
assign w11265 = w10919 & ~w10921;
assign v3476 = ~(w10922 | w11265);
assign w11266 = v3476;
assign w11267 = w11264 & w11266;
assign v3477 = ~(w11264 | w11266);
assign w11268 = v3477;
assign w11269 = ~w2492 & w11035;
assign w11270 = ~w2568 & w11023;
assign v3478 = ~(w11269 | w11270);
assign w11271 = v3478;
assign v3479 = ~(pi02 | w11271);
assign w11272 = v3479;
assign v3480 = ~(pi02 | w5898);
assign w11273 = v3480;
assign w11274 = ~w2596 & w10987;
assign w11275 = ~w10988 & w11271;
assign w11276 = ~w11274 & w11275;
assign w11277 = ~w11273 & w11276;
assign v3481 = ~(w11272 | w11277);
assign w11278 = v3481;
assign w11279 = w1 & w5898;
assign v3482 = ~(w11278 | w11279);
assign w11280 = v3482;
assign w11281 = w10915 & ~w10917;
assign v3483 = ~(w10918 | w11281);
assign w11282 = v3483;
assign w11283 = w11280 & w11282;
assign v3484 = ~(w11280 | w11282);
assign w11284 = v3484;
assign w11285 = w10911 & ~w10913;
assign v3485 = ~(w10914 | w11285);
assign w11286 = v3485;
assign w11287 = ~w4 & w6031;
assign w11288 = ~w2568 & w11035;
assign w11289 = ~w2596 & w11023;
assign v3486 = ~(w11288 | w11289);
assign w11290 = v3486;
assign w11291 = ~w11287 & w11290;
assign v3487 = ~(pi02 | w11291);
assign w11292 = v3487;
assign w11293 = ~w2669 & w10986;
assign w11294 = pi02 & ~w11293;
assign w11295 = w11291 & w11294;
assign v3488 = ~(w11292 | w11295);
assign w11296 = v3488;
assign w11297 = w11286 & ~w11296;
assign w11298 = ~w11286 & w11296;
assign w11299 = w10907 & ~w10909;
assign v3489 = ~(w10910 | w11299);
assign w11300 = v3489;
assign w11301 = ~w4 & w5880;
assign w11302 = ~w2669 & w11023;
assign w11303 = ~w2596 & w11035;
assign v3490 = ~(w11302 | w11303);
assign w11304 = v3490;
assign w11305 = ~w11301 & w11304;
assign v3491 = ~(pi02 | w11305);
assign w11306 = v3491;
assign w11307 = ~w2724 & w10986;
assign w11308 = pi02 & ~w11307;
assign w11309 = w11305 & w11308;
assign v3492 = ~(w11306 | w11309);
assign w11310 = v3492;
assign w11311 = w11300 & ~w11310;
assign w11312 = ~w11300 & w11310;
assign w11313 = w10903 & ~w10905;
assign v3493 = ~(w10906 | w11313);
assign w11314 = v3493;
assign w11315 = ~w4 & w6459;
assign w11316 = ~w2937 & w10987;
assign w11317 = ~w2846 & w11023;
assign w11318 = ~w2811 & w11035;
assign v3494 = ~(w11317 | w11318);
assign w11319 = v3494;
assign w11320 = ~w11316 & w11319;
assign w11321 = ~w11315 & w11320;
assign w11322 = pi02 & ~w11321;
assign w11323 = ~pi02 & w11321;
assign v3495 = ~(w11322 | w11323);
assign w11324 = v3495;
assign w11325 = w10895 & ~w10897;
assign v3496 = ~(w10898 | w11325);
assign w11326 = v3496;
assign w11327 = w11324 & w11326;
assign v3497 = ~(w11324 | w11326);
assign w11328 = v3497;
assign w11329 = w3 & w6130;
assign w11330 = ~w2937 & w11023;
assign w11331 = ~w2846 & w11035;
assign v3498 = ~(w11330 | w11331);
assign w11332 = v3498;
assign w11333 = pi02 & ~w11332;
assign w11334 = ~w3000 & w10986;
assign w11335 = pi02 & ~w11334;
assign w11336 = w11332 & ~w11335;
assign v3499 = ~(w11333 | w11336);
assign w11337 = v3499;
assign v3500 = ~(w11329 | w11337);
assign w11338 = v3500;
assign w11339 = w1 & w6130;
assign v3501 = ~(w11338 | w11339);
assign w11340 = v3501;
assign w11341 = w10871 & w10888;
assign v3502 = ~(w10889 | w11341);
assign w11342 = v3502;
assign w11343 = ~w3000 & w11023;
assign w11344 = ~w2937 & w11035;
assign v3503 = ~(w11343 | w11344);
assign w11345 = v3503;
assign w11346 = (w11345 & w6505) | (w11345 & w28499) | (w6505 & w28499);
assign w11347 = pi02 & ~w11346;
assign w11348 = ~w3068 & w10986;
assign w11349 = pi02 & ~w11348;
assign w11350 = w11346 & ~w11349;
assign v3504 = ~(w11347 | w11350);
assign w11351 = v3504;
assign v3505 = ~(w11342 | w11351);
assign w11352 = v3505;
assign v3506 = ~(w10858 | w10869);
assign w11353 = v3506;
assign v3507 = ~(w10870 | w11353);
assign w11354 = v3507;
assign w11355 = ~w3068 & w11023;
assign w11356 = ~w3000 & w11035;
assign v3508 = ~(w11355 | w11356);
assign w11357 = v3508;
assign w11358 = (~w6551 & w28299) | (~w6551 & w28300) | (w28299 & w28300);
assign w11359 = ~w3124 & w10986;
assign w11360 = pi02 & ~w11359;
assign w11361 = (w6551 & w28301) | (w6551 & w28302) | (w28301 & w28302);
assign v3509 = ~(w11358 | w11361);
assign w11362 = v3509;
assign w11363 = w11354 & ~w11362;
assign w11364 = ~w11354 & w11362;
assign w11365 = pi05 & ~w10854;
assign w11366 = w10847 & w11365;
assign v3510 = ~(w10847 | w11365);
assign w11367 = v3510;
assign v3511 = ~(w11366 | w11367);
assign w11368 = v3511;
assign w11369 = ~w3124 & w11023;
assign w11370 = ~w3068 & w11035;
assign v3512 = ~(w11369 | w11370);
assign w11371 = v3512;
assign w11372 = (w6603 & w28303) | (w6603 & w28304) | (w28303 & w28304);
assign w11373 = ~w3162 & w10986;
assign w11374 = pi02 & ~w11373;
assign w11375 = (~w6603 & w28305) | (~w6603 & w28306) | (w28305 & w28306);
assign v3513 = ~(w11372 | w11375);
assign w11376 = v3513;
assign w11377 = ~w11368 & w11376;
assign w11378 = ~w3211 & w11023;
assign w11379 = ~w3162 & w11035;
assign v3514 = ~(w11378 | w11379);
assign w11380 = v3514;
assign w11381 = (~w6735 & w28307) | (~w6735 & w28308) | (w28307 & w28308);
assign w11382 = w1 & w6735;
assign v3515 = ~(w11381 | w11382);
assign w11383 = v3515;
assign w11384 = (w1 & ~w6674) | (w1 & w28001) | (~w6674 & w28001);
assign w11385 = (pi01 & ~w3261) | (pi01 & w28309) | (~w3261 & w28309);
assign w11386 = ~w3211 & w11035;
assign w11387 = (~w10848 & w11384) | (~w10848 & w28500) | (w11384 & w28500);
assign w11388 = ~w3262 & w10987;
assign w11389 = (~pi02 & ~w11380) | (~pi02 & w28310) | (~w11380 & w28310);
assign w11390 = w11380 & w28311;
assign v3516 = ~(w11389 | w11390);
assign w11391 = v3516;
assign v3517 = ~(w11387 | w11391);
assign w11392 = v3517;
assign w11393 = w11383 & w11392;
assign w11394 = pi05 & w9396;
assign w11395 = ~w3332 & w11394;
assign w11396 = w10853 & ~w11395;
assign w11397 = ~w10853 & w11395;
assign v3518 = ~(w11396 | w11397);
assign w11398 = v3518;
assign w11399 = w11393 & w11398;
assign w11400 = (~w11398 & ~w11383) | (~w11398 & w28003) | (~w11383 & w28003);
assign w11401 = ~w3162 & w11023;
assign w11402 = ~w3124 & w11035;
assign v3519 = ~(w11401 | w11402);
assign w11403 = v3519;
assign w11404 = (~w6641 & w28312) | (~w6641 & w28313) | (w28312 & w28313);
assign w11405 = ~w3211 & w10986;
assign w11406 = pi02 & ~w11405;
assign w11407 = (w6641 & w28314) | (w6641 & w28315) | (w28314 & w28315);
assign v3520 = ~(w11404 | w11407);
assign w11408 = v3520;
assign w11409 = ~w11400 & w11408;
assign v3521 = ~(w11399 | w11409);
assign w11410 = v3521;
assign w11411 = w11368 & ~w11376;
assign w11412 = (~w11377 & w11410) | (~w11377 & w28316) | (w11410 & w28316);
assign w11413 = (~w11363 & w11412) | (~w11363 & w28005) | (w11412 & w28005);
assign w11414 = w11342 & w11351;
assign w11415 = w11413 & ~w11414;
assign w11416 = ~w11415 & w28747;
assign w11417 = (~w11340 & w11415) | (~w11340 & w28501) | (w11415 & w28501);
assign w11418 = w10891 & ~w10893;
assign v3522 = ~(w10894 | w11418);
assign w11419 = v3522;
assign w11420 = ~w11417 & w11419;
assign v3523 = ~(w11416 | w11420);
assign w11421 = v3523;
assign w11422 = (~w11327 & w11421) | (~w11327 & w28502) | (w11421 & w28502);
assign w11423 = w10899 & ~w10901;
assign v3524 = ~(w10902 | w11423);
assign w11424 = v3524;
assign v3525 = ~(w4 | w6447);
assign w11425 = v3525;
assign w11426 = ~w2846 & w10987;
assign w11427 = ~w2724 & w11035;
assign v3526 = ~(w11426 | w11427);
assign w11428 = v3526;
assign w11429 = ~w2811 & w11023;
assign w11430 = w11428 & ~w11429;
assign w11431 = ~w11425 & w11430;
assign w11432 = pi02 & w11431;
assign v3527 = ~(pi02 | w11431);
assign w11433 = v3527;
assign v3528 = ~(w11432 | w11433);
assign w11434 = v3528;
assign w11435 = ~w11424 & w11434;
assign w11436 = w11424 & ~w11434;
assign w11437 = (~w11436 & w11422) | (~w11436 & w28748) | (w11422 & w28748);
assign w11438 = w11314 & ~w11437;
assign w11439 = ~w4 & w6148;
assign w11440 = ~w2724 & w11023;
assign w11441 = ~w2669 & w11035;
assign v3529 = ~(w11440 | w11441);
assign w11442 = v3529;
assign w11443 = ~w11439 & w11442;
assign w11444 = pi02 & ~w11443;
assign w11445 = ~w2811 & w10986;
assign w11446 = pi02 & ~w11445;
assign w11447 = w11443 & ~w11446;
assign v3530 = ~(w11444 | w11447);
assign w11448 = v3530;
assign w11449 = (w11448 & ~w11437) | (w11448 & w28998) | (~w11437 & w28998);
assign v3531 = ~(w11438 | w11449);
assign w11450 = v3531;
assign w11451 = (~w11311 & w11450) | (~w11311 & w29272) | (w11450 & w29272);
assign v3532 = ~(w11298 | w11451);
assign w11452 = v3532;
assign v3533 = ~(w11297 | w11452);
assign w11453 = v3533;
assign w11454 = (~w11283 & w11453) | (~w11283 & w29488) | (w11453 & w29488);
assign v3534 = ~(w11268 | w11454);
assign w11455 = v3534;
assign v3535 = ~(w11267 | w11455);
assign w11456 = v3535;
assign w11457 = (~w11253 & w11456) | (~w11253 & w29489) | (w11456 & w29489);
assign w11458 = w11229 & w11239;
assign w11459 = w11457 & ~w11458;
assign w11460 = ~w11459 & w29708;
assign w11461 = ~w4 & w5262;
assign w11462 = ~w2202 & w11035;
assign w11463 = ~w2290 & w11023;
assign v3536 = ~(w11462 | w11463);
assign w11464 = v3536;
assign w11465 = ~w11461 & w11464;
assign w11466 = pi02 & ~w11465;
assign w11467 = ~w2339 & w10986;
assign w11468 = pi02 & ~w11467;
assign w11469 = w11465 & ~w11468;
assign v3537 = ~(w11466 | w11469);
assign w11470 = v3537;
assign v3538 = ~(w11460 | w11470);
assign w11471 = v3538;
assign w11472 = w10935 & ~w10937;
assign v3539 = ~(w10938 | w11472);
assign w11473 = v3539;
assign w11474 = ~w2202 & w11023;
assign w11475 = ~w2089 & w11035;
assign v3540 = ~(w11474 | w11475);
assign w11476 = v3540;
assign w11477 = (w11476 & ~w5033) | (w11476 & w29490) | (~w5033 & w29490);
assign v3541 = ~(pi02 | w11477);
assign w11478 = v3541;
assign w11479 = ~w2290 & w10986;
assign w11480 = pi02 & ~w11479;
assign w11481 = w11477 & w11480;
assign v3542 = ~(w11478 | w11481);
assign w11482 = v3542;
assign w11483 = ~w11473 & w11482;
assign w11484 = (~w11227 & w11459) | (~w11227 & w29709) | (w11459 & w29709);
assign v3543 = ~(w11483 | w11484);
assign w11485 = v3543;
assign w11486 = ~w11471 & w11485;
assign w11487 = w11473 & ~w11482;
assign w11488 = (~w11487 & ~w11222) | (~w11487 & w28503) | (~w11222 & w28503);
assign w11489 = ~w11486 & w11488;
assign v3544 = ~(w11225 | w11489);
assign w11490 = v3544;
assign w11491 = ~w11210 & w11212;
assign w11492 = (~w11491 & ~w11490) | (~w11491 & w29710) | (~w11490 & w29710);
assign w11493 = (~w11200 & w11492) | (~w11200 & w30160) | (w11492 & w30160);
assign v3545 = ~(w11178 | w11187);
assign w11494 = v3545;
assign v3546 = ~(w11493 | w11494);
assign w11495 = v3546;
assign v3547 = ~(w11188 | w11495);
assign w11496 = v3547;
assign w11497 = (~w11175 & w11496) | (~w11175 & w30161) | (w11496 & w30161);
assign w11498 = w10959 & ~w10961;
assign v3548 = ~(w10962 | w11498);
assign w11499 = v3548;
assign w11500 = ~w1609 & w11035;
assign w11501 = ~w1674 & w11023;
assign v3549 = ~(w11500 | w11501);
assign w11502 = v3549;
assign w11503 = (w11502 & w3491) | (w11502 & w29491) | (w3491 & w29491);
assign w11504 = pi02 & ~w11503;
assign w11505 = ~w1795 & w10986;
assign w11506 = pi02 & ~w11505;
assign w11507 = w11503 & ~w11506;
assign v3550 = ~(w11504 | w11507);
assign w11508 = v3550;
assign v3551 = ~(w11499 | w11508);
assign w11509 = v3551;
assign v3552 = ~(w11497 | w11509);
assign w11510 = v3552;
assign w11511 = w11499 & w11508;
assign w11512 = (~w11511 & w11162) | (~w11511 & w29711) | (w11162 & w29711);
assign w11513 = (~w11163 & ~w11512) | (~w11163 & w28006) | (~w11512 & w28006);
assign w11514 = (~w11149 & w11513) | (~w11149 & w29712) | (w11513 & w29712);
assign w11515 = ~w11138 & w11514;
assign v3553 = ~(w11133 | w11137);
assign w11516 = v3553;
assign v3554 = ~(w11515 | w11516);
assign w11517 = v3554;
assign w11518 = (~w11124 & w11517) | (~w11124 & w30336) | (w11517 & w30336);
assign w11519 = (~w11112 & w11518) | (~w11112 & w29713) | (w11518 & w29713);
assign w11520 = (~w11098 & w11519) | (~w11098 & w30495) | (w11519 & w30495);
assign w11521 = w11087 & ~w11520;
assign w11522 = (~w11085 & ~w11087) | (~w11085 & w28007) | (~w11087 & w28007);
assign w11523 = (~w11071 & w11522) | (~w11071 & w30613) | (w11522 & w30613);
assign w11524 = w11060 & ~w11523;
assign w11525 = (~w11058 & ~w11060) | (~w11058 & w28008) | (~w11060 & w28008);
assign w11526 = w11045 & ~w11525;
assign w11527 = w11022 & ~w11029;
assign w11528 = (~w11043 & ~w11022) | (~w11043 & w28181) | (~w11022 & w28181);
assign w11529 = ~w11526 & w11528;
assign w11530 = (~w11030 & w11526) | (~w11030 & w31029) | (w11526 & w31029);
assign w11531 = ~w11529 & w11821;
assign w11532 = ~w11018 & w11531;
assign v3555 = ~(w11017 | w11532);
assign w11533 = v3555;
assign w11534 = ~w10429 & w10431;
assign w11535 = w11012 & ~w11013;
assign w11536 = (~w11535 & ~w10431) | (~w11535 & w28182) | (~w10431 & w28182);
assign w11537 = (~w11533 & w28184) | (~w11533 & w28185) | (w28184 & w28185);
assign w11538 = (~w11533 & w31265) | (~w11533 & w31266) | (w31265 & w31266);
assign w11539 = (~w11537 & w28505) | (~w11537 & w28506) | (w28505 & w28506);
assign w11540 = (w11537 & w28749) | (w11537 & w28750) | (w28749 & w28750);
assign w11541 = (~w28750 & w29273) | (~w28750 & w29274) | (w29273 & w29274);
assign w11542 = (w28750 & w29275) | (w28750 & w29276) | (w29275 & w29276);
assign w11543 = (w8157 & w11542) | (w8157 & w29492) | (w11542 & w29492);
assign w11544 = (w11542 & w29862) | (w11542 & w29863) | (w29862 & w29863);
assign w11545 = (w11542 & w30162) | (w11542 & w30163) | (w30162 & w30163);
assign v3556 = ~(w7480 | w11545);
assign w11546 = v3556;
assign w11547 = (w7196 & w11545) | (w7196 & w30337) | (w11545 & w30337);
assign w11548 = (~w11545 & w30496) | (~w11545 & w30497) | (w30496 & w30497);
assign w11549 = w7034 & ~w7036;
assign v3557 = ~(w7037 | w11549);
assign w11550 = v3557;
assign w11551 = (w11542 & w31175) | (w11542 & w31176) | (w31175 & w31176);
assign v3558 = ~(w7037 | w11551);
assign w11552 = v3558;
assign w11553 = w6409 & ~w6886;
assign w11554 = w11552 & ~w11553;
assign v3559 = ~(w6887 | w11554);
assign w11555 = v3559;
assign w11556 = w6407 & w11555;
assign v3560 = ~(w6405 | w11556);
assign w11557 = v3560;
assign w11558 = ~w5995 & w6264;
assign v3561 = ~(w6265 | w11558);
assign w11559 = v3561;
assign w11560 = ~w11557 & w11559;
assign v3562 = ~(w6265 | w11560);
assign w11561 = v3562;
assign w11562 = ~w5993 & w11561;
assign v3563 = ~(w5992 | w11562);
assign w11563 = v3563;
assign w11564 = w5783 & w11563;
assign v3564 = ~(w5781 | w11564);
assign w11565 = v3564;
assign w11566 = w5642 & ~w11565;
assign v3565 = ~(w5640 | w11566);
assign w11567 = v3565;
assign w11568 = ~w5541 & w11567;
assign v3566 = ~(w5540 | w11568);
assign w11569 = v3566;
assign w11570 = w5130 & w11569;
assign v3567 = ~(w5128 | w11570);
assign w11571 = v3567;
assign w11572 = w4943 & ~w4945;
assign v3568 = ~(w4946 | w11572);
assign w11573 = v3568;
assign w11574 = ~w11571 & w11573;
assign v3569 = ~(w4946 | w11574);
assign w11575 = v3569;
assign v3570 = ~(w4846 | w11575);
assign w11576 = v3570;
assign v3571 = ~(w4845 | w11576);
assign w11577 = v3571;
assign w11578 = w4782 & ~w11577;
assign v3572 = ~(w4780 | w11578);
assign w11579 = v3572;
assign w11580 = w4326 & ~w4436;
assign v3573 = ~(w4437 | w11580);
assign w11581 = v3573;
assign w11582 = ~w11579 & w11581;
assign v3574 = ~(w4437 | w11582);
assign w11583 = v3574;
assign v3575 = ~(w4419 | w4434);
assign w11584 = v3575;
assign v3576 = ~(w4401 | w4416);
assign w11585 = v3576;
assign v3577 = ~(w4387 | w4397);
assign w11586 = v3577;
assign w11587 = w619 & w1239;
assign w11588 = w2624 & w5862;
assign w11589 = w1056 & w2835;
assign w11590 = ~w978 & w3912;
assign w11591 = w11589 & w11590;
assign w11592 = w1514 & w11591;
assign w11593 = ~w107 & w6625;
assign w11594 = w1106 & w11593;
assign w11595 = w11592 & w11594;
assign w11596 = w11588 & w11595;
assign v3578 = ~(w135 | w370);
assign w11597 = v3578;
assign v3579 = ~(w202 | w235);
assign w11598 = v3579;
assign w11599 = ~w267 & w11598;
assign w11600 = w11597 & w11599;
assign w11601 = ~w195 & w565;
assign w11602 = ~w466 & w846;
assign w11603 = w11601 & w11602;
assign w11604 = w1999 & w4041;
assign w11605 = w1147 & w2904;
assign w11606 = w11604 & w11605;
assign w11607 = w11603 & w11606;
assign w11608 = w11600 & w11607;
assign w11609 = w11596 & w11608;
assign w11610 = w2318 & w6044;
assign v3580 = ~(w278 | w481);
assign w11611 = v3580;
assign w11612 = w181 & w11611;
assign w11613 = w3730 & w11612;
assign v3581 = ~(w143 | w260);
assign w11614 = v3581;
assign w11615 = w6089 & w11614;
assign w11616 = w11613 & w11615;
assign w11617 = ~w479 & w3300;
assign w11618 = w2920 & w11617;
assign w11619 = w3135 & w11618;
assign w11620 = w11616 & w11619;
assign w11621 = w11610 & w11620;
assign w11622 = w5003 & w11621;
assign w11623 = w11609 & w11622;
assign w11624 = w11587 & w11623;
assign w11625 = ~w4385 & w11624;
assign w11626 = w4385 & ~w11624;
assign v3582 = ~(w11625 | w11626);
assign w11627 = v3582;
assign w11628 = w928 & ~w3928;
assign w11629 = w3399 & ~w3587;
assign w11630 = w3402 & ~w3752;
assign v3583 = ~(w11629 | w11630);
assign w11631 = v3583;
assign w11632 = w3406 & ~w3920;
assign w11633 = w11631 & ~w11632;
assign w11634 = ~w11628 & w11633;
assign w11635 = w11627 & w11634;
assign v3584 = ~(w11627 | w11634);
assign w11636 = v3584;
assign v3585 = ~(w11635 | w11636);
assign w11637 = v3585;
assign v3586 = ~(w11586 | w11637);
assign w11638 = v3586;
assign w11639 = w11586 & w11637;
assign v3587 = ~(w11638 | w11639);
assign w11640 = v3587;
assign w11641 = ~w11585 & w11640;
assign w11642 = w11585 & ~w11640;
assign v3588 = ~(w11641 | w11642);
assign w11643 = v3588;
assign w11644 = w3529 & ~w4149;
assign w11645 = w3763 & ~w4035;
assign w11646 = w3767 & ~w4134;
assign v3589 = ~(w11645 | w11646);
assign w11647 = v3589;
assign w11648 = w3760 & ~w4082;
assign w11649 = w11647 & ~w11648;
assign w11650 = ~w11644 & w11649;
assign w11651 = ~pi29 & w11650;
assign w11652 = pi29 & ~w11650;
assign v3590 = ~(w11651 | w11652);
assign w11653 = v3590;
assign w11654 = w4153 & ~w4422;
assign w11655 = w2873 & ~w11654;
assign v3591 = ~(w4191 | w11655);
assign w11656 = v3591;
assign w11657 = ~pi26 & w11656;
assign w11658 = pi26 & ~w11656;
assign v3592 = ~(w11657 | w11658);
assign w11659 = v3592;
assign w11660 = w11653 & ~w11659;
assign w11661 = ~w11653 & w11659;
assign v3593 = ~(w11660 | w11661);
assign w11662 = v3593;
assign w11663 = w11643 & w11662;
assign v3594 = ~(w11643 | w11662);
assign w11664 = v3594;
assign v3595 = ~(w11663 | w11664);
assign w11665 = v3595;
assign w11666 = w11584 & ~w11665;
assign w11667 = ~w11584 & w11665;
assign v3596 = ~(w11666 | w11667);
assign w11668 = v3596;
assign w11669 = ~w11583 & w11668;
assign w11670 = w11583 & ~w11668;
assign v3597 = ~(w11669 | w11670);
assign w11671 = v3597;
assign w11672 = w11579 & ~w11581;
assign v3598 = ~(w11582 | w11672);
assign w11673 = v3598;
assign w11674 = w11671 & w11673;
assign v3599 = ~(w11671 | w11673);
assign w11675 = v3599;
assign v3600 = ~(w11674 | w11675);
assign w11676 = v3600;
assign w11677 = ~w4782 & w11577;
assign v3601 = ~(w11578 | w11677);
assign w11678 = v3601;
assign v3602 = ~(w11673 | w11678);
assign w11679 = v3602;
assign v3603 = ~(w4845 | w4846);
assign w11680 = v3603;
assign w11681 = w11575 & w11680;
assign v3604 = ~(w11575 | w11680);
assign w11682 = v3604;
assign v3605 = ~(w11681 | w11682);
assign w11683 = v3605;
assign w11684 = w11678 & ~w11683;
assign w11685 = w11571 & ~w11573;
assign v3606 = ~(w11574 | w11685);
assign w11686 = v3606;
assign w11687 = ~w11683 & w11686;
assign v3607 = ~(w5130 | w11569);
assign w11688 = v3607;
assign v3608 = ~(w11570 | w11688);
assign w11689 = v3608;
assign v3609 = ~(w11686 | w11689);
assign w11690 = v3609;
assign w11691 = w11686 & w11689;
assign v3610 = ~(w5540 | w5541);
assign w11692 = v3610;
assign v3611 = ~(w11567 | w11692);
assign w11693 = v3611;
assign w11694 = w11567 & w11692;
assign v3612 = ~(w11693 | w11694);
assign w11695 = v3612;
assign w11696 = w11689 & ~w11695;
assign w11697 = ~w11689 & w11695;
assign v3613 = ~(w11696 | w11697);
assign w11698 = v3613;
assign w11699 = ~w5642 & w11565;
assign v3614 = ~(w11566 | w11699);
assign w11700 = v3614;
assign w11701 = w11695 & ~w11700;
assign w11702 = ~w11695 & w11700;
assign v3615 = ~(w11701 | w11702);
assign w11703 = v3615;
assign v3616 = ~(w5992 | w5993);
assign w11704 = v3616;
assign w11705 = ~w11561 & w11704;
assign v3617 = ~(w5993 | w11705);
assign w11706 = v3617;
assign w11707 = ~w5783 & w11706;
assign v3618 = ~(w11564 | w11707);
assign w11708 = v3618;
assign w11709 = w11700 & w11708;
assign w11710 = w11561 & ~w11704;
assign v3619 = ~(w11705 | w11710);
assign w11711 = v3619;
assign w11712 = w11708 & w11711;
assign w11713 = w11557 & ~w11559;
assign v3620 = ~(w11560 | w11713);
assign w11714 = v3620;
assign w11715 = w11711 & w11714;
assign v3621 = ~(w6887 | w11553);
assign w11716 = v3621;
assign w11717 = ~w11552 & w11716;
assign v3622 = ~(w11553 | w11717);
assign w11718 = v3622;
assign w11719 = ~w6407 & w11718;
assign v3623 = ~(w11556 | w11719);
assign w11720 = v3623;
assign w11721 = w11714 & w11720;
assign w11722 = w11552 & ~w11716;
assign v3624 = ~(w11717 | w11722);
assign w11723 = v3624;
assign v3625 = ~(w11720 | w11723);
assign w11724 = v3625;
assign w11725 = w11548 & ~w11550;
assign v3626 = ~(w11551 | w11725);
assign w11726 = v3626;
assign v3627 = ~(w11723 | w11726);
assign w11727 = v3627;
assign w11728 = ~w7196 & w11546;
assign v3628 = ~(w11547 | w11728);
assign w11729 = v3628;
assign w11730 = w11726 & w11729;
assign v3629 = ~(w7480 | w7481);
assign w11731 = v3629;
assign w11732 = (w11542 & w30338) | (w11542 & w30339) | (w30338 & w30339);
assign w11733 = (~w11542 & w30340) | (~w11542 & w30341) | (w30340 & w30341);
assign v3630 = ~(w11732 | w11733);
assign w11734 = v3630;
assign w11735 = ~w11729 & w11734;
assign w11736 = (~w11542 & w30164) | (~w11542 & w30165) | (w30164 & w30165);
assign v3631 = ~(w11544 | w11736);
assign w11737 = v3631;
assign w11738 = ~w11734 & w11737;
assign w11739 = ~w11542 & w30029;
assign v3632 = ~(w11543 | w11739);
assign w11740 = v3632;
assign w11741 = w11737 & w11740;
assign v3633 = ~(w8540 | w8541);
assign w11742 = v3633;
assign v3634 = ~(w11541 | w11742);
assign w11743 = v3634;
assign w11744 = w11541 & w11742;
assign v3635 = ~(w11743 | w11744);
assign w11745 = v3635;
assign w11746 = ~w11740 & w11745;
assign w11747 = ~w8959 & w11539;
assign v3636 = ~(w11540 | w11747);
assign w11748 = v3636;
assign w11749 = ~w11745 & w11748;
assign w11750 = w11745 & ~w11748;
assign v3637 = ~(w11749 | w11750);
assign w11751 = v3637;
assign w11752 = (w11533 & w31267) | (w11533 & w31268) | (w31267 & w31268);
assign v3638 = ~(w8959 | w9418);
assign w11753 = v3638;
assign w11754 = w8959 & w9418;
assign v3639 = ~(w11753 | w11754);
assign w11755 = v3639;
assign w11756 = w11752 & ~w11755;
assign w11757 = ~w11752 & w11755;
assign v3640 = ~(w11756 | w11757);
assign w11758 = v3640;
assign v3641 = ~(w11538 | w11752);
assign w11759 = v3641;
assign w11760 = (w11533 & w29277) | (w11533 & w29278) | (w29277 & w29278);
assign v3642 = ~(w11537 | w11760);
assign w11761 = v3642;
assign w11762 = w11759 & w11761;
assign w11763 = w11759 & w28751;
assign v3643 = ~(w10432 | w11534);
assign w11764 = v3643;
assign w11765 = w11535 & ~w11764;
assign w11766 = (~w11765 & ~w28318) | (~w11765 & w31030) | (~w28318 & w31030);
assign w11767 = w11018 & ~w11531;
assign w11768 = w11533 & ~w11767;
assign w11769 = ~w11766 & w11768;
assign w11770 = (~w11764 & w11532) | (~w11764 & w30166) | (w11532 & w30166);
assign w11771 = w11766 & ~w11770;
assign w11772 = w11761 & ~w11771;
assign w11773 = ~w11761 & w11771;
assign v3644 = ~(w11017 | w11018);
assign w11774 = v3644;
assign v3645 = ~(w11020 | w11530);
assign w11775 = v3645;
assign v3646 = ~(w11531 | w11775);
assign w11776 = v3646;
assign w11777 = w11774 & w11776;
assign v3647 = ~(w11030 | w11527);
assign w11778 = v3647;
assign w11779 = w11043 & ~w11778;
assign w11780 = ~w11043 & w11778;
assign v3648 = ~(w11779 | w11780);
assign w11781 = v3648;
assign w11782 = ~w11526 & w11781;
assign w11783 = w11526 & w11778;
assign w11784 = (~w11783 & ~w11781) | (~w11783 & w28186) | (~w11781 & w28186);
assign w11785 = w11020 & ~w11527;
assign w11786 = ~w11020 & w11527;
assign v3649 = ~(w11785 | w11786);
assign w11787 = v3649;
assign w11788 = (~w11781 & w31031) | (~w11781 & w31032) | (w31031 & w31032);
assign w11789 = ~w11774 & w11775;
assign v3650 = ~(w11532 | w11789);
assign w11790 = v3650;
assign v3651 = ~(w11045 | w11058);
assign w11791 = v3651;
assign w11792 = ~w11045 & w29716;
assign v3652 = ~(w11526 | w11792);
assign w11793 = v3652;
assign w11794 = ~w11781 & w11793;
assign v3653 = ~(w11071 | w11072);
assign w11795 = v3653;
assign w11796 = w11522 & ~w11795;
assign w11797 = ~w11522 & w11795;
assign v3654 = ~(w11796 | w11797);
assign w11798 = v3654;
assign w11799 = ~w11087 & w11520;
assign v3655 = ~(w11521 | w11799);
assign w11800 = v3655;
assign w11801 = w11798 & ~w11800;
assign w11802 = ~w11060 & w11523;
assign v3656 = ~(w11524 | w11802);
assign w11803 = v3656;
assign w11804 = w11801 & ~w11803;
assign w11805 = (w11798 & w11803) | (w11798 & w28319) | (w11803 & w28319);
assign w11806 = w11045 & w11058;
assign v3657 = ~(w11791 | w11806);
assign w11807 = v3657;
assign w11808 = w11802 & ~w11807;
assign w11809 = ~w11802 & w11807;
assign v3658 = ~(w11808 | w11809);
assign w11810 = v3658;
assign w11811 = w11805 & w11810;
assign w11812 = w11803 & w11807;
assign w11813 = (~w11812 & ~w11810) | (~w11812 & w28010) | (~w11810 & w28010);
assign w11814 = ~w11794 & w11813;
assign w11815 = ~w11781 & w11792;
assign w11816 = w11781 & ~w11792;
assign v3659 = ~(w11815 | w11816);
assign w11817 = v3659;
assign w11818 = ~w11784 & w11817;
assign v3660 = ~(w11814 | w11818);
assign w11819 = v3660;
assign w11820 = ~w11020 & w11030;
assign w11821 = w11020 & ~w11030;
assign w11822 = (~w11781 & w31033) | (~w11781 & w31034) | (w31033 & w31034);
assign v3661 = ~(w11784 | w11822);
assign w11823 = v3661;
assign v3662 = ~(w11788 | w11823);
assign w11824 = v3662;
assign w11825 = w11819 & w11824;
assign w11826 = w11002 & w11010;
assign v3663 = ~(w11010 | w11012);
assign w11827 = v3663;
assign v3664 = ~(w11826 | w11827);
assign w11828 = v3664;
assign w11829 = ~w11531 & w11828;
assign w11830 = (~w11014 & ~w11530) | (~w11014 & w30808) | (~w11530 & w30808);
assign w11831 = (~w11764 & w11829) | (~w11764 & w31035) | (w11829 & w31035);
assign w11832 = ~w11829 & w31036;
assign v3665 = ~(w11831 | w11832);
assign w11833 = v3665;
assign w11834 = (w28011 & w29493) | (w28011 & w29494) | (w29493 & w29494);
assign w11835 = ~w11773 & w11834;
assign w11836 = ~w11835 & w28321;
assign v3666 = ~(w11759 | w11761);
assign w11837 = v3666;
assign v3667 = ~(w11762 | w11837);
assign w11838 = v3667;
assign w11839 = (w11838 & w11835) | (w11838 & w31269) | (w11835 & w31269);
assign v3668 = ~(w11758 | w11762);
assign w11840 = v3668;
assign w11841 = ~w11839 & w28322;
assign w11842 = (w11758 & w11839) | (w11758 & w29279) | (w11839 & w29279);
assign w11843 = ~w11538 & w11757;
assign w11844 = (~w11839 & w29280) | (~w11839 & w29281) | (w29280 & w29281);
assign w11845 = w11751 & ~w11844;
assign w11846 = (~w11749 & w11844) | (~w11749 & w29000) | (w11844 & w29000);
assign w11847 = w11740 & ~w11745;
assign w11848 = w11846 & ~w11847;
assign v3669 = ~(w11737 | w11740);
assign w11849 = v3669;
assign v3670 = ~(w11741 | w11849);
assign w11850 = v3670;
assign w11851 = ~w11848 & w29495;
assign w11852 = w11734 & ~w11737;
assign v3671 = ~(w11738 | w11852);
assign w11853 = v3671;
assign w11854 = (~w11848 & w30030) | (~w11848 & w30031) | (w30030 & w30031);
assign w11855 = (w11848 & w30167) | (w11848 & w30168) | (w30167 & w30168);
assign w11856 = w11729 & ~w11734;
assign v3672 = ~(w11735 | w11856);
assign w11857 = v3672;
assign w11858 = w11855 & w11857;
assign v3673 = ~(w11726 | w11729);
assign w11859 = v3673;
assign v3674 = ~(w11730 | w11859);
assign w11860 = v3674;
assign w11861 = (~w11855 & w30498) | (~w11855 & w30499) | (w30498 & w30499);
assign v3675 = ~(w11730 | w11861);
assign w11862 = v3675;
assign w11863 = w11723 & w11726;
assign v3676 = ~(w11727 | w11863);
assign w11864 = v3676;
assign w11865 = w11862 & w11864;
assign v3677 = ~(w11727 | w11865);
assign w11866 = v3677;
assign w11867 = w11720 & w11723;
assign v3678 = ~(w11724 | w11867);
assign w11868 = v3678;
assign w11869 = ~w11866 & w11868;
assign v3679 = ~(w11724 | w11869);
assign w11870 = v3679;
assign v3680 = ~(w11714 | w11720);
assign w11871 = v3680;
assign v3681 = ~(w11721 | w11871);
assign w11872 = v3681;
assign w11873 = w11870 & w11872;
assign v3682 = ~(w11721 | w11873);
assign w11874 = v3682;
assign v3683 = ~(w11711 | w11714);
assign w11875 = v3683;
assign v3684 = ~(w11715 | w11875);
assign w11876 = v3684;
assign w11877 = ~w11874 & w11876;
assign v3685 = ~(w11715 | w11877);
assign w11878 = v3685;
assign w11879 = ~w11712 & w11878;
assign v3686 = ~(w11708 | w11711);
assign w11880 = v3686;
assign v3687 = ~(w11700 | w11708);
assign w11881 = v3687;
assign v3688 = ~(w11709 | w11881);
assign w11882 = v3688;
assign w11883 = ~w11880 & w11882;
assign w11884 = ~w11879 & w11883;
assign w11885 = (~w11709 & ~w11883) | (~w11709 & w28323) | (~w11883 & w28323);
assign w11886 = w11703 & w11885;
assign v3689 = ~(w11701 | w11886);
assign w11887 = v3689;
assign w11888 = w11698 & w11887;
assign v3690 = ~(w11696 | w11888);
assign w11889 = v3690;
assign w11890 = ~w11691 & w11889;
assign v3691 = ~(w11690 | w11890);
assign w11891 = v3691;
assign w11892 = w11683 & ~w11686;
assign w11893 = ~w11678 & w11683;
assign v3692 = ~(w11684 | w11893);
assign w11894 = v3692;
assign w11895 = w11894 & w28324;
assign v3693 = ~(w11684 | w11895);
assign w11896 = v3693;
assign w11897 = w11673 & w11678;
assign w11898 = w11896 & ~w11897;
assign v3694 = ~(w11679 | w11898);
assign w11899 = v3694;
assign w11900 = w11676 & w11899;
assign v3695 = ~(w11660 | w11663);
assign w11901 = v3695;
assign w11902 = w3529 & w4196;
assign w11903 = w3763 & ~w4082;
assign w11904 = w3760 & ~w4191;
assign w11905 = w3767 & ~w4035;
assign v3696 = ~(w11904 | w11905);
assign w11906 = v3696;
assign w11907 = ~w11903 & w11906;
assign w11908 = ~w11902 & w11907;
assign w11909 = pi29 & ~w11908;
assign w11910 = ~pi29 & w11908;
assign v3697 = ~(w11909 | w11910);
assign w11911 = v3697;
assign v3698 = ~(w11638 | w11641);
assign w11912 = v3698;
assign v3699 = ~(w110 | w208);
assign w11913 = v3699;
assign w11914 = ~w27 & w11913;
assign w11915 = ~w234 & w11914;
assign w11916 = ~w410 & w11915;
assign w11917 = w6120 & w11916;
assign w11918 = w489 & w1476;
assign w11919 = w185 & w1641;
assign w11920 = w11918 & w11919;
assign w11921 = w6089 & w11920;
assign w11922 = w3982 & w5431;
assign w11923 = w2107 & w11922;
assign w11924 = ~w680 & w11923;
assign w11925 = w1354 & w11924;
assign w11926 = w11921 & w11925;
assign w11927 = w11917 & w11926;
assign w11928 = w4225 & w4995;
assign w11929 = w2507 & w11928;
assign w11930 = ~w494 & w1600;
assign w11931 = ~w474 & w11930;
assign w11932 = w4232 & w11931;
assign w11933 = w11929 & w11932;
assign w11934 = w91 & w6102;
assign w11935 = w2156 & w11934;
assign v3700 = ~(w73 | w179);
assign w11936 = v3700;
assign v3701 = ~(w125 | w666);
assign w11937 = v3701;
assign w11938 = w11936 & w11937;
assign w11939 = ~w111 & w11938;
assign w11940 = ~w1108 & w11939;
assign w11941 = w11935 & w11940;
assign w11942 = w279 & w1442;
assign w11943 = w1465 & ~w3816;
assign w11944 = w344 & w11943;
assign w11945 = w11942 & w11944;
assign w11946 = w2292 & w11945;
assign w11947 = w11941 & w11946;
assign w11948 = w11933 & w11947;
assign w11949 = w11927 & w11948;
assign w11950 = w3311 & w11949;
assign w11951 = w4385 & w11950;
assign v3702 = ~(w4385 | w11950);
assign w11952 = v3702;
assign v3703 = ~(w11951 | w11952);
assign w11953 = v3703;
assign w11954 = pi26 & w11953;
assign v3704 = ~(pi26 | w11953);
assign w11955 = v3704;
assign v3705 = ~(w11954 | w11955);
assign w11956 = v3705;
assign v3706 = ~(w11625 | w11635);
assign w11957 = v3706;
assign w11958 = ~w11956 & w11957;
assign w11959 = w11956 & ~w11957;
assign v3707 = ~(w11958 | w11959);
assign w11960 = v3707;
assign w11961 = w928 & w4309;
assign w11962 = w3402 & ~w3920;
assign w11963 = w3399 & ~w3752;
assign v3708 = ~(w11962 | w11963);
assign w11964 = v3708;
assign w11965 = w3406 & ~w4134;
assign w11966 = w11964 & ~w11965;
assign w11967 = ~w11961 & w11966;
assign w11968 = w11960 & ~w11967;
assign w11969 = ~w11960 & w11967;
assign v3709 = ~(w11968 | w11969);
assign w11970 = v3709;
assign w11971 = ~w11912 & w11970;
assign w11972 = w11912 & ~w11970;
assign v3710 = ~(w11971 | w11972);
assign w11973 = v3710;
assign w11974 = w11911 & w11973;
assign v3711 = ~(w11911 | w11973);
assign w11975 = v3711;
assign v3712 = ~(w11974 | w11975);
assign w11976 = v3712;
assign w11977 = ~w11901 & w11976;
assign w11978 = w11901 & ~w11976;
assign v3713 = ~(w11977 | w11978);
assign w11979 = v3713;
assign w11980 = (w28013 & w11579) | (w28013 & w28325) | (w11579 & w28325);
assign v3714 = ~(w11666 | w11980);
assign w11981 = v3714;
assign w11982 = w11979 & w11981;
assign w11983 = (w11583 & w28015) | (w11583 & w28016) | (w28015 & w28016);
assign v3715 = ~(w11982 | w11983);
assign w11984 = v3715;
assign w11985 = w11671 & w11984;
assign v3716 = ~(w11674 | w11985);
assign w11986 = v3716;
assign v3717 = ~(w11671 | w11984);
assign w11987 = v3717;
assign w11988 = w11986 & ~w11987;
assign w11989 = w11900 & w11988;
assign w11990 = w11673 & w11985;
assign v3718 = ~(w11900 | w11990);
assign w11991 = v3718;
assign w11992 = ~w11988 & w11991;
assign v3719 = ~(w11989 | w11992);
assign w11993 = v3719;
assign w11994 = w928 & w11993;
assign w11995 = w3406 & w11984;
assign w11996 = w3402 & w11671;
assign w11997 = w3399 & w11673;
assign v3720 = ~(w11996 | w11997);
assign w11998 = v3720;
assign w11999 = ~w11995 & w11998;
assign w12000 = ~w11994 & w11999;
assign w12001 = w926 & ~w12000;
assign v3721 = ~(w924 | w12001);
assign w12002 = v3721;
assign w12003 = w323 & ~w663;
assign v3722 = ~(w664 | w12003);
assign w12004 = v3722;
assign w12005 = w12002 & w12004;
assign v3723 = ~(w664 | w12005);
assign w12006 = v3723;
assign w12007 = w521 & w12006;
assign v3724 = ~(w521 | w12006);
assign w12008 = v3724;
assign v3725 = ~(w12007 | w12008);
assign w12009 = v3725;
assign v3726 = ~(w11951 | w11954);
assign w12010 = v3726;
assign w12011 = ~w63 & w4064;
assign w12012 = ~w162 & w426;
assign w12013 = w1967 & w12012;
assign w12014 = ~w70 & w1771;
assign w12015 = ~w103 & w136;
assign w12016 = w12014 & w12015;
assign v3727 = ~(w448 | w997);
assign w12017 = v3727;
assign w12018 = ~w194 & w12017;
assign w12019 = w5311 & w12018;
assign w12020 = w12016 & w12019;
assign w12021 = w1934 & w3451;
assign w12022 = w1262 & w12021;
assign w12023 = w12020 & w12022;
assign w12024 = w12013 & w12023;
assign w12025 = ~w302 & w1329;
assign w12026 = w12024 & w12025;
assign w12027 = w12011 & w12026;
assign w12028 = ~w145 & w6707;
assign w12029 = w1057 & w12028;
assign w12030 = ~w299 & w6520;
assign w12031 = w1689 & w2817;
assign w12032 = w12030 & w12031;
assign v3728 = ~(w172 | w307);
assign w12033 = v3728;
assign w12034 = w3644 & w12033;
assign w12035 = w1200 & w1947;
assign w12036 = w12034 & w12035;
assign w12037 = w12032 & w12036;
assign w12038 = ~w326 & w1049;
assign v3729 = ~(w337 | w685);
assign w12039 = v3729;
assign w12040 = w79 & w12039;
assign w12041 = w12038 & w12040;
assign w12042 = w12037 & w12041;
assign w12043 = w12029 & w12042;
assign w12044 = ~w418 & w990;
assign w12045 = ~w278 & w12044;
assign w12046 = w12043 & w12045;
assign w12047 = w4584 & w12046;
assign w12048 = w12027 & w12047;
assign w12049 = w12010 & w12048;
assign v3730 = ~(w12010 | w12048);
assign w12050 = v3730;
assign v3731 = ~(w12049 | w12050);
assign w12051 = v3731;
assign w12052 = w928 & w4405;
assign w12053 = w3406 & ~w4035;
assign w12054 = w3402 & ~w4134;
assign v3732 = ~(w12053 | w12054);
assign w12055 = v3732;
assign w12056 = w3399 & ~w3920;
assign w12057 = w12055 & ~w12056;
assign w12058 = ~w12052 & w12057;
assign w12059 = w12051 & ~w12058;
assign w12060 = ~w12051 & w12058;
assign v3733 = ~(w12059 | w12060);
assign w12061 = v3733;
assign v3734 = ~(w11958 | w11968);
assign w12062 = v3734;
assign w12063 = w12061 & ~w12062;
assign w12064 = ~w12061 & w12062;
assign v3735 = ~(w12063 | w12064);
assign w12065 = v3735;
assign w12066 = w3529 & w4425;
assign w12067 = w3767 & ~w4082;
assign w12068 = w3763 & ~w4191;
assign v3736 = ~(w12067 | w12068);
assign w12069 = v3736;
assign w12070 = ~w12066 & w12069;
assign w12071 = pi29 & ~w12070;
assign w12072 = ~pi29 & w12070;
assign v3737 = ~(w12071 | w12072);
assign w12073 = v3737;
assign w12074 = w12065 & w12073;
assign v3738 = ~(w12065 | w12073);
assign w12075 = v3738;
assign v3739 = ~(w12074 | w12075);
assign w12076 = v3739;
assign v3740 = ~(w11971 | w11974);
assign w12077 = v3740;
assign w12078 = w12076 & ~w12077;
assign w12079 = ~w12076 & w12077;
assign v3741 = ~(w12078 | w12079);
assign w12080 = v3741;
assign v3742 = ~(w11977 | w11982);
assign w12081 = v3742;
assign w12082 = w12080 & ~w12081;
assign w12083 = ~w12080 & w12081;
assign v3743 = ~(w12082 | w12083);
assign w12084 = v3743;
assign v3744 = ~(w12078 | w12082);
assign w12085 = v3744;
assign v3745 = ~(w12063 | w12074);
assign w12086 = v3745;
assign v3746 = ~(w12049 | w12059);
assign w12087 = v3746;
assign w12088 = ~w886 & w1547;
assign w12089 = ~w244 & w574;
assign w12090 = w12088 & w12089;
assign w12091 = w787 & w12090;
assign v3747 = ~(w220 | w499);
assign w12092 = v3747;
assign w12093 = w3544 & w12092;
assign w12094 = w401 & w12093;
assign w12095 = w3304 & w12094;
assign w12096 = w12091 & w12095;
assign w12097 = w1432 & w12096;
assign w12098 = ~w438 & w12097;
assign w12099 = w802 & w3133;
assign w12100 = w1014 & w12099;
assign w12101 = w489 & w1864;
assign w12102 = w1359 & w2634;
assign w12103 = w12101 & w12102;
assign w12104 = w12100 & w12103;
assign w12105 = w2442 & w12104;
assign w12106 = w5245 & w12105;
assign w12107 = w12098 & w12106;
assign w12108 = ~w195 & w1714;
assign w12109 = w2303 & w3086;
assign w12110 = ~w431 & w12109;
assign w12111 = w2026 & w12110;
assign w12112 = ~w159 & w12111;
assign w12113 = w12108 & w12112;
assign w12114 = w1325 & w4571;
assign w12115 = w2657 & w12114;
assign v3748 = ~(w127 | w298);
assign w12116 = v3748;
assign w12117 = ~w176 & w12116;
assign v3749 = ~(w143 | w179);
assign w12118 = v3749;
assign w12119 = ~w410 & w12118;
assign w12120 = w12117 & w12119;
assign w12121 = w4254 & w12120;
assign w12122 = w12115 & w12121;
assign w12123 = w12113 & w12122;
assign w12124 = w2087 & w12123;
assign w12125 = w12107 & w12124;
assign w12126 = ~w12048 & w12125;
assign w12127 = w12048 & ~w12125;
assign v3750 = ~(w12126 | w12127);
assign w12128 = v3750;
assign w12129 = w12087 & w12128;
assign v3751 = ~(w12087 | w12128);
assign w12130 = v3751;
assign v3752 = ~(w12129 | w12130);
assign w12131 = v3752;
assign w12132 = w3525 & w4422;
assign v3753 = ~(w3523 | w4191);
assign w12133 = v3753;
assign w12134 = ~w12132 & w12133;
assign w12135 = pi28 & w12134;
assign v3754 = ~(pi29 | w12135);
assign w12136 = v3754;
assign w12137 = w928 & ~w4149;
assign w12138 = w3402 & ~w4035;
assign w12139 = w3399 & ~w4134;
assign v3755 = ~(w12138 | w12139);
assign w12140 = v3755;
assign w12141 = w3406 & ~w4082;
assign w12142 = w12140 & ~w12141;
assign w12143 = ~w12137 & w12142;
assign v3756 = ~(w12136 | w12143);
assign w12144 = v3756;
assign w12145 = w12136 & w12143;
assign v3757 = ~(w12144 | w12145);
assign w12146 = v3757;
assign w12147 = ~w12131 & w12146;
assign w12148 = w12131 & ~w12146;
assign v3758 = ~(w12147 | w12148);
assign w12149 = v3758;
assign w12150 = w12086 & ~w12149;
assign w12151 = ~w12086 & w12149;
assign v3759 = ~(w12150 | w12151);
assign w12152 = v3759;
assign w12153 = ~w12085 & w12152;
assign w12154 = w12085 & ~w12152;
assign v3760 = ~(w12153 | w12154);
assign w12155 = v3760;
assign w12156 = w12084 & w12155;
assign v3761 = ~(w12084 | w12155);
assign w12157 = v3761;
assign v3762 = ~(w12156 | w12157);
assign w12158 = v3762;
assign w12159 = w11984 & w12084;
assign w12160 = w11986 & ~w11989;
assign v3763 = ~(w11984 | w12084);
assign w12161 = v3763;
assign v3764 = ~(w12159 | w12161);
assign w12162 = v3764;
assign w12163 = ~w12160 & w12162;
assign w12164 = (~w12159 & w12160) | (~w12159 & w28017) | (w12160 & w28017);
assign w12165 = w12158 & ~w12164;
assign w12166 = ~w12158 & w12164;
assign v3765 = ~(w12165 | w12166);
assign w12167 = v3765;
assign w12168 = w928 & w12167;
assign w12169 = w3406 & w12155;
assign w12170 = w3399 & w11984;
assign w12171 = w3402 & w12084;
assign v3766 = ~(w12170 | w12171);
assign w12172 = v3766;
assign w12173 = ~w12169 & w12172;
assign w12174 = ~w12168 & w12173;
assign w12175 = w12009 & ~w12174;
assign w12176 = ~w12009 & w12174;
assign v3767 = ~(w12175 | w12176);
assign w12177 = v3767;
assign v3768 = ~(w12002 | w12004);
assign w12178 = v3768;
assign v3769 = ~(w12005 | w12178);
assign w12179 = v3769;
assign w12180 = w12160 & ~w12162;
assign v3770 = ~(w12163 | w12180);
assign w12181 = v3770;
assign w12182 = w928 & w12181;
assign w12183 = w3406 & w12084;
assign w12184 = w3402 & w11984;
assign w12185 = w3399 & w11671;
assign v3771 = ~(w12184 | w12185);
assign w12186 = v3771;
assign w12187 = ~w12183 & w12186;
assign w12188 = ~w12182 & w12187;
assign v3772 = ~(w12179 | w12188);
assign w12189 = v3772;
assign w12190 = w12179 & w12188;
assign v3773 = ~(w12189 | w12190);
assign w12191 = v3773;
assign v3774 = ~(w12144 | w12147);
assign w12192 = v3774;
assign w12193 = w5216 & w6718;
assign w12194 = w4113 & w12193;
assign v3775 = ~(w381 | w685);
assign w12195 = v3775;
assign w12196 = w4075 & w12195;
assign w12197 = w4036 & w12196;
assign w12198 = w887 & w1888;
assign w12199 = w12197 & w12198;
assign w12200 = ~w187 & w2142;
assign w12201 = w4118 & w12200;
assign w12202 = w4014 & w12201;
assign w12203 = w681 & w3996;
assign w12204 = w12202 & w12203;
assign w12205 = w12199 & w12204;
assign w12206 = w2027 & w3970;
assign w12207 = w2443 & w12206;
assign w12208 = ~w584 & w12207;
assign w12209 = w12205 & w12208;
assign w12210 = w12194 & w12209;
assign w12211 = w12125 & w12210;
assign v3776 = ~(w12125 | w12210);
assign w12212 = v3776;
assign v3777 = ~(w12211 | w12212);
assign w12213 = v3777;
assign w12214 = pi29 & w12213;
assign v3778 = ~(pi29 | w12213);
assign w12215 = v3778;
assign v3779 = ~(w12214 | w12215);
assign w12216 = v3779;
assign v3780 = ~(w12127 | w12129);
assign w12217 = v3780;
assign w12218 = ~w12216 & w12217;
assign w12219 = w12216 & ~w12217;
assign v3781 = ~(w12218 | w12219);
assign w12220 = v3781;
assign w12221 = w928 & w4196;
assign w12222 = w3399 & ~w4035;
assign w12223 = w3402 & ~w4082;
assign v3782 = ~(w12222 | w12223);
assign w12224 = v3782;
assign w12225 = ~w12221 & w12224;
assign w12226 = w12220 & ~w12225;
assign w12227 = ~w12220 & w12225;
assign v3783 = ~(w12226 | w12227);
assign w12228 = v3783;
assign w12229 = ~w12192 & w12228;
assign w12230 = w12192 & ~w12228;
assign v3784 = ~(w12229 | w12230);
assign w12231 = v3784;
assign v3785 = ~(w12085 | w12150);
assign w12232 = v3785;
assign v3786 = ~(w12151 | w12232);
assign w12233 = v3786;
assign w12234 = w12231 & ~w12233;
assign v3787 = ~(w12151 | w12231);
assign w12235 = v3787;
assign w12236 = ~w12153 & w12235;
assign v3788 = ~(w12234 | w12236);
assign w12237 = v3788;
assign v3789 = ~(w12155 | w12237);
assign w12238 = v3789;
assign v3790 = ~(w12156 | w12165);
assign w12239 = v3790;
assign w12240 = w12155 & w12237;
assign v3791 = ~(w12238 | w12240);
assign w12241 = v3791;
assign w12242 = w12239 & w12241;
assign v3792 = ~(w12238 | w12242);
assign w12243 = v3792;
assign w12244 = w928 & w4425;
assign w12245 = w3402 & ~w4191;
assign v3793 = ~(w12244 | w12245);
assign w12246 = v3793;
assign v3794 = ~(w12211 | w12214);
assign w12247 = v3794;
assign w12248 = w4058 & w12202;
assign w12249 = w4174 & w12248;
assign w12250 = w2890 & w5378;
assign w12251 = ~w239 & w3998;
assign w12252 = w740 & w12251;
assign w12253 = w4102 & w12252;
assign w12254 = w3556 & w12253;
assign w12255 = w12250 & w12254;
assign w12256 = w3973 & w12255;
assign w12257 = w12249 & w12256;
assign w12258 = w12247 & w12257;
assign v3795 = ~(w12247 | w12257);
assign w12259 = v3795;
assign v3796 = ~(w12258 | w12259);
assign w12260 = v3796;
assign w12261 = ~w12246 & w12260;
assign w12262 = w12246 & ~w12260;
assign v3797 = ~(w12261 | w12262);
assign w12263 = v3797;
assign v3798 = ~(w12218 | w12226);
assign w12264 = v3798;
assign w12265 = w12263 & ~w12264;
assign w12266 = ~w12263 & w12264;
assign v3799 = ~(w12265 | w12266);
assign w12267 = v3799;
assign v3800 = ~(w12229 | w12234);
assign w12268 = v3800;
assign w12269 = w12267 & ~w12268;
assign w12270 = ~w12267 & w12268;
assign v3801 = ~(w12269 | w12270);
assign w12271 = v3801;
assign v3802 = ~(w12237 | w12271);
assign w12272 = v3802;
assign w12273 = w12237 & w12271;
assign v3803 = ~(w12272 | w12273);
assign w12274 = v3803;
assign w12275 = ~w12243 & w12274;
assign w12276 = w12243 & ~w12274;
assign v3804 = ~(w12275 | w12276);
assign w12277 = v3804;
assign w12278 = w3529 & ~w12277;
assign w12279 = w3763 & w12237;
assign w12280 = w3760 & w12271;
assign v3805 = ~(w12279 | w12280);
assign w12281 = v3805;
assign w12282 = w3767 & w12155;
assign w12283 = w12281 & ~w12282;
assign w12284 = ~w12278 & w12283;
assign w12285 = pi29 & w12284;
assign v3806 = ~(pi29 | w12284);
assign w12286 = v3806;
assign v3807 = ~(w12285 | w12286);
assign w12287 = v3807;
assign w12288 = w12191 & ~w12287;
assign v3808 = ~(w12189 | w12288);
assign w12289 = v3808;
assign w12290 = w12177 & ~w12289;
assign w12291 = ~w12177 & w12289;
assign v3809 = ~(w12290 | w12291);
assign w12292 = v3809;
assign v3810 = ~(w12258 | w12261);
assign w12293 = v3810;
assign w12294 = w2142 & w4119;
assign w12295 = w1647 & w12294;
assign w12296 = w12197 & w12295;
assign w12297 = ~w267 & w2465;
assign w12298 = ~w369 & w12297;
assign w12299 = w4177 & w12298;
assign w12300 = w12296 & w12299;
assign w12301 = w4061 & w12300;
assign w12302 = w12257 & ~w12301;
assign w12303 = ~w12257 & w12301;
assign v3811 = ~(w12302 | w12303);
assign w12304 = v3811;
assign w12305 = ~w12293 & w12304;
assign w12306 = w12293 & ~w12304;
assign v3812 = ~(w12305 | w12306);
assign w12307 = v3812;
assign v3813 = ~(w12265 | w12269);
assign w12308 = v3813;
assign w12309 = w12307 & ~w12308;
assign w12310 = ~w12307 & w12308;
assign v3814 = ~(w12309 | w12310);
assign w12311 = v3814;
assign w12312 = w12271 & w12311;
assign v3815 = ~(w12271 | w12311);
assign w12313 = v3815;
assign v3816 = ~(w12312 | w12313);
assign w12314 = v3816;
assign v3817 = ~(w12272 | w12275);
assign w12315 = v3817;
assign w12316 = w12314 & w12315;
assign v3818 = ~(w12314 | w12315);
assign w12317 = v3818;
assign v3819 = ~(w12316 | w12317);
assign w12318 = v3819;
assign w12319 = w3529 & w12318;
assign w12320 = w3760 & w12311;
assign w12321 = w3763 & w12271;
assign w12322 = w3767 & w12237;
assign v3820 = ~(w12321 | w12322);
assign w12323 = v3820;
assign w12324 = ~w12320 & w12323;
assign w12325 = ~w12319 & w12324;
assign w12326 = ~pi29 & w12325;
assign w12327 = pi29 & ~w12325;
assign v3821 = ~(w12326 | w12327);
assign w12328 = v3821;
assign w12329 = w12292 & w12328;
assign v3822 = ~(w12290 | w12329);
assign w12330 = v3822;
assign v3823 = ~(w12007 | w12175);
assign w12331 = v3823;
assign v3824 = ~(w516 | w519);
assign w12332 = v3824;
assign w12333 = w2349 & w3907;
assign w12334 = w1767 & w4017;
assign w12335 = ~w692 & w12334;
assign w12336 = ~w466 & w4092;
assign w12337 = w12335 & w12336;
assign w12338 = w6684 & w12337;
assign w12339 = w2141 & w2282;
assign w12340 = w12338 & w12339;
assign w12341 = w12333 & w12340;
assign w12342 = w2849 & w12202;
assign w12343 = ~w727 & w1786;
assign w12344 = w12342 & w12343;
assign w12345 = w12341 & w12344;
assign w12346 = w3721 & w12345;
assign w12347 = ~w12332 & w12346;
assign w12348 = w12332 & ~w12346;
assign v3825 = ~(w12347 | w12348);
assign w12349 = v3825;
assign v3826 = ~(w12239 | w12241);
assign w12350 = v3826;
assign v3827 = ~(w12242 | w12350);
assign w12351 = v3827;
assign w12352 = w928 & ~w12351;
assign w12353 = w3406 & w12237;
assign w12354 = w3399 & w12084;
assign w12355 = w3402 & w12155;
assign v3828 = ~(w12354 | w12355);
assign w12356 = v3828;
assign w12357 = ~w12353 & w12356;
assign w12358 = ~w12352 & w12357;
assign w12359 = w12349 & ~w12358;
assign w12360 = ~w12349 & w12358;
assign v3829 = ~(w12359 | w12360);
assign w12361 = v3829;
assign w12362 = ~w12331 & w12361;
assign w12363 = w12331 & ~w12361;
assign v3830 = ~(w12362 | w12363);
assign w12364 = v3830;
assign v3831 = ~(w12312 | w12316);
assign w12365 = v3831;
assign v3832 = ~(w12305 | w12309);
assign w12366 = v3832;
assign w12367 = w3973 & w4016;
assign w12368 = w3554 & w4102;
assign w12369 = w2139 & w4074;
assign w12370 = w12368 & w12369;
assign v3833 = ~(w456 | w697);
assign w12371 = v3833;
assign w12372 = ~w172 & w12371;
assign w12373 = w12370 & w12372;
assign w12374 = w12367 & w12373;
assign v3834 = ~(w12257 | w12374);
assign w12375 = v3834;
assign w12376 = w12257 & w12374;
assign w12377 = w12301 & w12376;
assign v3835 = ~(w12375 | w12377);
assign w12378 = v3835;
assign w12379 = w12366 & w12378;
assign v3836 = ~(w12366 | w12378);
assign w12380 = v3836;
assign v3837 = ~(w12379 | w12380);
assign w12381 = v3837;
assign v3838 = ~(w12311 | w12381);
assign w12382 = v3838;
assign w12383 = w12311 & w12381;
assign v3839 = ~(w12382 | w12383);
assign w12384 = v3839;
assign w12385 = w12365 & ~w12384;
assign w12386 = ~w12365 & w12384;
assign v3840 = ~(w12385 | w12386);
assign w12387 = v3840;
assign w12388 = w3529 & w12387;
assign w12389 = w3760 & w12381;
assign w12390 = w3767 & w12271;
assign w12391 = w3763 & w12311;
assign v3841 = ~(w12390 | w12391);
assign w12392 = v3841;
assign w12393 = ~w12389 & w12392;
assign w12394 = ~w12388 & w12393;
assign w12395 = ~pi29 & w12394;
assign w12396 = pi29 & ~w12394;
assign v3842 = ~(w12395 | w12396);
assign w12397 = v3842;
assign w12398 = w12364 & w12397;
assign v3843 = ~(w12364 | w12397);
assign w12399 = v3843;
assign v3844 = ~(w12398 | w12399);
assign w12400 = v3844;
assign w12401 = ~w12330 & w12400;
assign w12402 = w12330 & ~w12400;
assign v3845 = ~(w12401 | w12402);
assign w12403 = v3845;
assign w12404 = w4040 & ~w12376;
assign v3846 = ~(w12302 | w12380);
assign w12405 = v3846;
assign w12406 = ~w12404 & w12405;
assign v3847 = ~(w2873 | w12406);
assign w12407 = v3847;
assign v3848 = ~(w4027 | w12407);
assign w12408 = v3848;
assign w12409 = ~w4152 & w12408;
assign w12410 = pi26 & ~w12409;
assign w12411 = ~pi26 & w12409;
assign v3849 = ~(w12410 | w12411);
assign w12412 = v3849;
assign w12413 = w12403 & w12412;
assign v3850 = ~(w12403 | w12412);
assign w12414 = v3850;
assign v3851 = ~(w12413 | w12414);
assign w12415 = v3851;
assign w12416 = w919 & ~w921;
assign v3852 = ~(w922 | w12416);
assign w12417 = v3852;
assign w12418 = w1042 & w3615;
assign w12419 = w4611 & w12418;
assign w12420 = ~w169 & w12419;
assign w12421 = w2063 & w12420;
assign w12422 = w2640 & w12421;
assign w12423 = ~w107 & w1520;
assign w12424 = w2600 & w12423;
assign v3853 = ~(w593 | w630);
assign w12425 = v3853;
assign w12426 = w411 & w12425;
assign w12427 = w12424 & w12426;
assign w12428 = w1214 & w12427;
assign w12429 = w4342 & w12428;
assign w12430 = w12422 & w12429;
assign w12431 = w5335 & w12430;
assign w12432 = ~w309 & w1219;
assign w12433 = ~w132 & w694;
assign w12434 = w2341 & w12433;
assign v3854 = ~(w192 | w877);
assign w12435 = v3854;
assign w12436 = w2024 & w12435;
assign w12437 = ~w997 & w1960;
assign w12438 = w12436 & w12437;
assign w12439 = w12434 & w12438;
assign w12440 = w1780 & w3723;
assign w12441 = w12439 & w12440;
assign w12442 = w76 & w626;
assign w12443 = w2656 & w12442;
assign w12444 = w12441 & w12443;
assign w12445 = w12432 & w12444;
assign w12446 = w2319 & w12445;
assign w12447 = w12431 & w12446;
assign w12448 = ~w776 & w12447;
assign w12449 = w776 & ~w12447;
assign v3855 = ~(w12448 | w12449);
assign w12450 = v3855;
assign v3856 = ~(w11679 | w11897);
assign w12451 = v3856;
assign w12452 = ~w11896 & w12451;
assign w12453 = w11896 & ~w12451;
assign v3857 = ~(w12452 | w12453);
assign w12454 = v3857;
assign w12455 = w928 & w12454;
assign w12456 = w3406 & w11673;
assign w12457 = w3402 & w11678;
assign w12458 = w3399 & ~w11683;
assign v3858 = ~(w12457 | w12458);
assign w12459 = v3858;
assign w12460 = ~w12456 & w12459;
assign w12461 = ~w12455 & w12460;
assign w12462 = w12450 & w12461;
assign v3859 = ~(w12448 | w12462);
assign w12463 = v3859;
assign w12464 = w12417 & w12463;
assign v3860 = ~(w12417 | w12463);
assign w12465 = v3860;
assign v3861 = ~(w12464 | w12465);
assign w12466 = v3861;
assign v3862 = ~(w11897 | w12452);
assign w12467 = v3862;
assign w12468 = ~w11676 & w12467;
assign v3863 = ~(w11900 | w12468);
assign w12469 = v3863;
assign w12470 = w928 & w12469;
assign w12471 = w3406 & w11671;
assign w12472 = w3402 & w11673;
assign w12473 = w3399 & w11678;
assign v3864 = ~(w12472 | w12473);
assign w12474 = v3864;
assign w12475 = ~w12471 & w12474;
assign w12476 = ~w12470 & w12475;
assign w12477 = w12466 & ~w12476;
assign v3865 = ~(w12464 | w12477);
assign w12478 = v3865;
assign w12479 = ~w926 & w12000;
assign v3866 = ~(w12001 | w12479);
assign w12480 = v3866;
assign w12481 = ~w12478 & w12480;
assign w12482 = w12478 & ~w12480;
assign v3867 = ~(w12481 | w12482);
assign w12483 = v3867;
assign w12484 = w3529 & ~w12351;
assign w12485 = w3760 & w12237;
assign w12486 = w3763 & w12155;
assign w12487 = w3767 & w12084;
assign v3868 = ~(w12486 | w12487);
assign w12488 = v3868;
assign w12489 = ~w12485 & w12488;
assign w12490 = ~w12484 & w12489;
assign w12491 = ~pi29 & w12490;
assign w12492 = pi29 & ~w12490;
assign v3869 = ~(w12491 | w12492);
assign w12493 = v3869;
assign w12494 = w12483 & w12493;
assign v3870 = ~(w12481 | w12494);
assign w12495 = v3870;
assign w12496 = ~w12191 & w12287;
assign v3871 = ~(w12288 | w12496);
assign w12497 = v3871;
assign w12498 = ~w12495 & w12497;
assign w12499 = w12495 & ~w12497;
assign v3872 = ~(w12498 | w12499);
assign w12500 = v3872;
assign w12501 = w12381 & ~w12406;
assign w12502 = w12365 & ~w12383;
assign w12503 = w12501 & ~w12502;
assign w12504 = ~w12501 & w12502;
assign v3873 = ~(w12382 | w12504);
assign w12505 = v3873;
assign w12506 = ~w12503 & w12505;
assign w12507 = w4153 & ~w12506;
assign w12508 = w4155 & ~w12406;
assign w12509 = ~w2873 & w12311;
assign w12510 = w4158 & w12381;
assign v3874 = ~(w12509 | w12510);
assign w12511 = v3874;
assign w12512 = ~w12508 & w12511;
assign w12513 = ~w12507 & w12512;
assign w12514 = ~pi26 & w12513;
assign w12515 = pi26 & ~w12513;
assign v3875 = ~(w12514 | w12515);
assign w12516 = v3875;
assign w12517 = w12500 & w12516;
assign v3876 = ~(w12498 | w12517);
assign w12518 = v3876;
assign w12519 = ~w2873 & w12381;
assign w12520 = w4153 & w12505;
assign v3877 = ~(w4158 | w12520);
assign w12521 = v3877;
assign v3878 = ~(w12406 | w12521);
assign w12522 = v3878;
assign v3879 = ~(w4155 | w12522);
assign w12523 = v3879;
assign w12524 = ~w12519 & w12523;
assign w12525 = ~pi26 & w12524;
assign w12526 = pi26 & ~w12524;
assign v3880 = ~(w12525 | w12526);
assign w12527 = v3880;
assign w12528 = ~w12518 & w12527;
assign v3881 = ~(w12292 | w12328);
assign w12529 = v3881;
assign v3882 = ~(w12329 | w12529);
assign w12530 = v3882;
assign w12531 = w12518 & ~w12527;
assign v3883 = ~(w12528 | w12531);
assign w12532 = v3883;
assign w12533 = w12530 & w12532;
assign v3884 = ~(w12528 | w12533);
assign w12534 = v3884;
assign w12535 = w12415 & ~w12534;
assign w12536 = ~w12415 & w12534;
assign v3885 = ~(w12535 | w12536);
assign w12537 = v3885;
assign w12538 = ~w12466 & w12476;
assign v3886 = ~(w12477 | w12538);
assign w12539 = v3886;
assign w12540 = ~w326 & w3097;
assign w12541 = w5406 & w12540;
assign w12542 = ~w405 & w3620;
assign w12543 = w740 & w1359;
assign w12544 = w12542 & w12543;
assign w12545 = w12541 & w12544;
assign w12546 = w2986 & w12545;
assign v3887 = ~(w159 | w418);
assign w12547 = v3887;
assign w12548 = w3277 & w12547;
assign v3888 = ~(w299 | w308);
assign w12549 = v3888;
assign v3889 = ~(w281 | w888);
assign w12550 = v3889;
assign w12551 = w12549 & w12550;
assign w12552 = w12548 & w12551;
assign w12553 = ~w252 & w2517;
assign w12554 = ~w194 & w12553;
assign w12555 = w12552 & w12554;
assign v3890 = ~(w338 | w494);
assign w12556 = v3890;
assign w12557 = w1761 & w12556;
assign w12558 = w2223 & w6104;
assign w12559 = w12557 & w12558;
assign w12560 = w12555 & w12559;
assign w12561 = w1126 & w12560;
assign w12562 = w12546 & w12561;
assign w12563 = w368 & w6626;
assign v3891 = ~(w224 | w343);
assign w12564 = v3891;
assign w12565 = w2733 & w12564;
assign w12566 = w12563 & w12565;
assign w12567 = w2363 & w4575;
assign w12568 = w3291 & w12567;
assign w12569 = ~w245 & w12568;
assign w12570 = w714 & w3447;
assign w12571 = w12569 & w12570;
assign w12572 = w12566 & w12571;
assign w12573 = ~w277 & w1239;
assign w12574 = w3015 & w12573;
assign w12575 = w772 & w12574;
assign w12576 = w5011 & w12575;
assign w12577 = w12098 & w12576;
assign w12578 = w12572 & w12577;
assign v3892 = ~(w12562 | w12578);
assign w12579 = v3892;
assign w12580 = pi17 & ~w5760;
assign w12581 = ~pi14 & w5757;
assign v3893 = ~(w12580 | w12581);
assign w12582 = v3893;
assign w12583 = w12562 & w12578;
assign v3894 = ~(w12579 | w12583);
assign w12584 = v3894;
assign w12585 = ~w12582 & w12584;
assign v3895 = ~(w12579 | w12585);
assign w12586 = v3895;
assign w12587 = w776 & ~w12586;
assign w12588 = ~w776 & w12586;
assign v3896 = ~(w12587 | w12588);
assign w12589 = v3896;
assign v3897 = ~(w11687 | w11892);
assign w12590 = v3897;
assign w12591 = w11891 & w12590;
assign v3898 = ~(w11687 | w12591);
assign w12592 = v3898;
assign w12593 = ~w11894 & w12592;
assign v3899 = ~(w11895 | w12593);
assign w12594 = v3899;
assign w12595 = w928 & w12594;
assign w12596 = w3406 & w11678;
assign w12597 = w3399 & w11686;
assign w12598 = w3402 & ~w11683;
assign v3900 = ~(w12597 | w12598);
assign w12599 = v3900;
assign w12600 = ~w12596 & w12599;
assign w12601 = ~w12595 & w12600;
assign w12602 = w12589 & ~w12601;
assign v3901 = ~(w12587 | w12602);
assign w12603 = v3901;
assign v3902 = ~(w12450 | w12461);
assign w12604 = v3902;
assign v3903 = ~(w12462 | w12604);
assign w12605 = v3903;
assign v3904 = ~(w12603 | w12605);
assign w12606 = v3904;
assign w12607 = w12582 & ~w12584;
assign v3905 = ~(w12585 | w12607);
assign w12608 = v3905;
assign v3906 = ~(w11891 | w12590);
assign w12609 = v3906;
assign v3907 = ~(w12591 | w12609);
assign w12610 = v3907;
assign w12611 = w928 & w12610;
assign w12612 = w3406 & ~w11683;
assign w12613 = w3402 & w11686;
assign w12614 = w3399 & w11689;
assign v3908 = ~(w12613 | w12614);
assign w12615 = v3908;
assign w12616 = ~w12612 & w12615;
assign w12617 = ~w12611 & w12616;
assign w12618 = w12608 & ~w12617;
assign w12619 = ~w12608 & w12617;
assign v3909 = ~(w12618 | w12619);
assign w12620 = v3909;
assign w12621 = w75 & ~w739;
assign w12622 = w513 & w12621;
assign w12623 = w2174 & w4349;
assign w12624 = w790 & w2024;
assign w12625 = w1447 & w4554;
assign w12626 = w12624 & w12625;
assign w12627 = w2615 & w12626;
assign w12628 = w12623 & w12627;
assign w12629 = ~w263 & w1575;
assign w12630 = w641 & w3113;
assign w12631 = w12629 & w12630;
assign v3910 = ~(w252 | w405);
assign w12632 = v3910;
assign w12633 = w786 & w2134;
assign w12634 = w12632 & w12633;
assign w12635 = w12631 & w12634;
assign w12636 = w91 & w12635;
assign v3911 = ~(w167 | w525);
assign w12637 = v3911;
assign w12638 = w2363 & w3071;
assign w12639 = w12637 & w12638;
assign w12640 = ~w266 & w12639;
assign w12641 = w12636 & w12640;
assign w12642 = w3330 & w12641;
assign w12643 = w12628 & w12642;
assign w12644 = w12622 & w12643;
assign w12645 = ~w12562 & w12644;
assign w12646 = ~w274 & w5232;
assign w12647 = ~w221 & w3240;
assign w12648 = ~w457 & w3886;
assign w12649 = w5410 & w12648;
assign v3912 = ~(w179 | w505);
assign w12650 = v3912;
assign w12651 = w3679 & w12650;
assign w12652 = w12649 & w12651;
assign w12653 = w2012 & w12652;
assign v3913 = ~(w239 | w369);
assign w12654 = v3913;
assign w12655 = w2398 & w12425;
assign w12656 = w12654 & w12655;
assign w12657 = w12653 & w12656;
assign w12658 = w12647 & w12657;
assign w12659 = w12646 & w12658;
assign w12660 = w3612 & w12659;
assign w12661 = w121 & w3658;
assign v3914 = ~(w74 | w427);
assign w12662 = v3914;
assign v3915 = ~(w169 | w999);
assign w12663 = v3915;
assign w12664 = w12662 & w12663;
assign w12665 = w489 & w1603;
assign w12666 = w12664 & w12665;
assign w12667 = w4605 & w12666;
assign w12668 = w12661 & w12667;
assign w12669 = w6484 & w12668;
assign v3916 = ~(w111 | w753);
assign w12670 = v3916;
assign w12671 = ~w425 & w12670;
assign w12672 = w2504 & w12671;
assign v3917 = ~(w235 | w593);
assign w12673 = v3917;
assign w12674 = w540 & w12673;
assign w12675 = w1570 & w12674;
assign w12676 = w1045 & w12675;
assign w12677 = ~w456 & w12676;
assign w12678 = w12672 & w12677;
assign w12679 = w2539 & w4683;
assign w12680 = w12678 & w12679;
assign w12681 = w12669 & w12680;
assign v3918 = ~(w12660 | w12681);
assign w12682 = v3918;
assign w12683 = pi14 & ~w6387;
assign w12684 = ~pi11 & w6384;
assign v3919 = ~(w12683 | w12684);
assign w12685 = v3919;
assign w12686 = w12660 & w12681;
assign v3920 = ~(w12682 | w12686);
assign w12687 = v3920;
assign w12688 = ~w12685 & w12687;
assign v3921 = ~(w12682 | w12688);
assign w12689 = v3921;
assign w12690 = w12644 & ~w12689;
assign w12691 = ~w12644 & w12689;
assign v3922 = ~(w12690 | w12691);
assign w12692 = v3922;
assign v3923 = ~(w11698 | w11887);
assign w12693 = v3923;
assign v3924 = ~(w11888 | w12693);
assign w12694 = v3924;
assign w12695 = w928 & w12694;
assign w12696 = w3406 & w11689;
assign w12697 = w3399 & w11700;
assign w12698 = w3402 & ~w11695;
assign v3925 = ~(w12697 | w12698);
assign w12699 = v3925;
assign w12700 = ~w12696 & w12699;
assign w12701 = ~w12695 & w12700;
assign w12702 = w12692 & ~w12701;
assign v3926 = ~(w12690 | w12702);
assign w12703 = v3926;
assign w12704 = w12562 & ~w12644;
assign v3927 = ~(w12645 | w12704);
assign w12705 = v3927;
assign w12706 = w12703 & w12705;
assign v3928 = ~(w12645 | w12706);
assign w12707 = v3928;
assign w12708 = w12620 & w12707;
assign v3929 = ~(w12618 | w12708);
assign w12709 = v3929;
assign w12710 = ~w12589 & w12601;
assign v3930 = ~(w12602 | w12710);
assign w12711 = v3930;
assign w12712 = ~w12709 & w12711;
assign w12713 = w12709 & ~w12711;
assign v3931 = ~(w12712 | w12713);
assign w12714 = v3931;
assign w12715 = w3529 & w11993;
assign w12716 = w3763 & w11671;
assign w12717 = w3760 & w11984;
assign v3932 = ~(w12716 | w12717);
assign w12718 = v3932;
assign w12719 = w3767 & w11673;
assign w12720 = w12718 & ~w12719;
assign w12721 = ~w12715 & w12720;
assign w12722 = pi29 & w12721;
assign v3933 = ~(pi29 | w12721);
assign w12723 = v3933;
assign v3934 = ~(w12722 | w12723);
assign w12724 = v3934;
assign w12725 = w12714 & ~w12724;
assign v3935 = ~(w12712 | w12725);
assign w12726 = v3935;
assign w12727 = w12603 & w12605;
assign v3936 = ~(w12606 | w12727);
assign w12728 = v3936;
assign w12729 = ~w12726 & w12728;
assign v3937 = ~(w12606 | w12729);
assign w12730 = v3937;
assign w12731 = w12539 & ~w12730;
assign w12732 = ~w12539 & w12730;
assign v3938 = ~(w12731 | w12732);
assign w12733 = v3938;
assign w12734 = w3529 & w12167;
assign w12735 = w3767 & w11984;
assign w12736 = w3760 & w12155;
assign v3939 = ~(w12735 | w12736);
assign w12737 = v3939;
assign w12738 = w3763 & w12084;
assign w12739 = w12737 & ~w12738;
assign w12740 = ~w12734 & w12739;
assign w12741 = pi29 & w12740;
assign v3940 = ~(pi29 | w12740);
assign w12742 = v3940;
assign v3941 = ~(w12741 | w12742);
assign w12743 = v3941;
assign w12744 = w12733 & ~w12743;
assign v3942 = ~(w12731 | w12744);
assign w12745 = v3942;
assign v3943 = ~(w12483 | w12493);
assign w12746 = v3943;
assign v3944 = ~(w12494 | w12746);
assign w12747 = v3944;
assign w12748 = ~w12745 & w12747;
assign w12749 = w12745 & ~w12747;
assign v3945 = ~(w12748 | w12749);
assign w12750 = v3945;
assign w12751 = w4153 & w12387;
assign w12752 = w4155 & w12381;
assign w12753 = ~w2873 & w12271;
assign w12754 = w4158 & w12311;
assign v3946 = ~(w12753 | w12754);
assign w12755 = v3946;
assign w12756 = ~w12752 & w12755;
assign w12757 = ~w12751 & w12756;
assign w12758 = ~pi26 & w12757;
assign w12759 = pi26 & ~w12757;
assign v3947 = ~(w12758 | w12759);
assign w12760 = v3947;
assign w12761 = w12750 & w12760;
assign v3948 = ~(w12748 | w12761);
assign w12762 = v3948;
assign w12763 = w14 & ~w12762;
assign v3949 = ~(w12500 | w12516);
assign w12764 = v3949;
assign v3950 = ~(w12517 | w12764);
assign w12765 = v3950;
assign w12766 = ~w14 & w12762;
assign v3951 = ~(w12763 | w12766);
assign w12767 = v3951;
assign w12768 = w12765 & w12767;
assign v3952 = ~(w12763 | w12768);
assign w12769 = v3952;
assign v3953 = ~(w12530 | w12532);
assign w12770 = v3953;
assign v3954 = ~(w12533 | w12770);
assign w12771 = v3954;
assign w12772 = ~w12769 & w12771;
assign w12773 = w12769 & ~w12771;
assign v3955 = ~(w12772 | w12773);
assign w12774 = v3955;
assign v3956 = ~(w12765 | w12767);
assign w12775 = v3956;
assign v3957 = ~(w12768 | w12775);
assign w12776 = v3957;
assign v3958 = ~(w12750 | w12760);
assign w12777 = v3958;
assign v3959 = ~(w12761 | w12777);
assign w12778 = v3959;
assign w12779 = ~w12733 & w12743;
assign v3960 = ~(w12744 | w12779);
assign w12780 = v3960;
assign w12781 = w4153 & w12318;
assign w12782 = w4155 & w12311;
assign w12783 = ~w2873 & w12237;
assign w12784 = w4158 & w12271;
assign v3961 = ~(w12783 | w12784);
assign w12785 = v3961;
assign w12786 = ~w12782 & w12785;
assign w12787 = ~w12781 & w12786;
assign w12788 = ~pi26 & w12787;
assign w12789 = pi26 & ~w12787;
assign v3962 = ~(w12788 | w12789);
assign w12790 = v3962;
assign w12791 = w12780 & w12790;
assign w12792 = w12726 & ~w12728;
assign v3963 = ~(w12729 | w12792);
assign w12793 = v3963;
assign w12794 = w3529 & w12181;
assign w12795 = w3763 & w11984;
assign w12796 = w3760 & w12084;
assign v3964 = ~(w12795 | w12796);
assign w12797 = v3964;
assign w12798 = w3767 & w11671;
assign w12799 = w12797 & ~w12798;
assign w12800 = ~w12794 & w12799;
assign w12801 = pi29 & w12800;
assign v3965 = ~(pi29 | w12800);
assign w12802 = v3965;
assign v3966 = ~(w12801 | w12802);
assign w12803 = v3966;
assign w12804 = w12793 & ~w12803;
assign w12805 = ~w12793 & w12803;
assign v3967 = ~(w12804 | w12805);
assign w12806 = v3967;
assign w12807 = w4153 & ~w12277;
assign w12808 = w4155 & w12271;
assign w12809 = ~w2873 & w12155;
assign w12810 = w4158 & w12237;
assign v3968 = ~(w12809 | w12810);
assign w12811 = v3968;
assign w12812 = ~w12808 & w12811;
assign w12813 = ~w12807 & w12812;
assign w12814 = ~pi26 & w12813;
assign w12815 = pi26 & ~w12813;
assign v3969 = ~(w12814 | w12815);
assign w12816 = v3969;
assign w12817 = w12806 & w12816;
assign v3970 = ~(w12804 | w12817);
assign w12818 = v3970;
assign v3971 = ~(w12780 | w12790);
assign w12819 = v3971;
assign v3972 = ~(w12791 | w12819);
assign w12820 = v3972;
assign w12821 = ~w12818 & w12820;
assign v3973 = ~(w12791 | w12821);
assign w12822 = v3973;
assign w12823 = w12778 & ~w12822;
assign w12824 = ~w12778 & w12822;
assign v3974 = ~(w12823 | w12824);
assign w12825 = v3974;
assign w12826 = pi23 & w12406;
assign w12827 = pi22 & ~w12406;
assign v3975 = ~(w12826 | w12827);
assign w12828 = v3975;
assign w12829 = w11 & w12828;
assign v3976 = ~(w12 | w12829);
assign w12830 = v3976;
assign w12831 = w12825 & w12830;
assign v3977 = ~(w12823 | w12831);
assign w12832 = v3977;
assign w12833 = w12776 & ~w12832;
assign w12834 = ~w12776 & w12832;
assign v3978 = ~(w12825 | w12830);
assign w12835 = v3978;
assign v3979 = ~(w12831 | w12835);
assign w12836 = v3979;
assign v3980 = ~(w12703 | w12705);
assign w12837 = v3980;
assign v3981 = ~(w12706 | w12837);
assign w12838 = v3981;
assign v3982 = ~(w11690 | w11691);
assign w12839 = v3982;
assign w12840 = w11889 & w12839;
assign v3983 = ~(w11889 | w12839);
assign w12841 = v3983;
assign v3984 = ~(w12840 | w12841);
assign w12842 = v3984;
assign w12843 = w928 & ~w12842;
assign w12844 = w3406 & w11686;
assign w12845 = w3402 & w11689;
assign w12846 = w3399 & ~w11695;
assign v3985 = ~(w12845 | w12846);
assign w12847 = v3985;
assign w12848 = ~w12844 & w12847;
assign w12849 = ~w12843 & w12848;
assign v3986 = ~(w12838 | w12849);
assign w12850 = v3986;
assign w12851 = w12838 & w12849;
assign v3987 = ~(w12850 | w12851);
assign w12852 = v3987;
assign w12853 = w3529 & w12454;
assign w12854 = w3763 & w11678;
assign w12855 = w3760 & w11673;
assign v3988 = ~(w12854 | w12855);
assign w12856 = v3988;
assign w12857 = w3767 & ~w11683;
assign w12858 = w12856 & ~w12857;
assign w12859 = ~w12853 & w12858;
assign w12860 = pi29 & w12859;
assign v3989 = ~(pi29 | w12859);
assign w12861 = v3989;
assign v3990 = ~(w12860 | w12861);
assign w12862 = v3990;
assign w12863 = w12852 & ~w12862;
assign v3991 = ~(w12850 | w12863);
assign w12864 = v3991;
assign v3992 = ~(w12620 | w12707);
assign w12865 = v3992;
assign v3993 = ~(w12708 | w12865);
assign w12866 = v3993;
assign w12867 = ~w12864 & w12866;
assign w12868 = w12864 & ~w12866;
assign v3994 = ~(w12867 | w12868);
assign w12869 = v3994;
assign w12870 = w3529 & w12469;
assign w12871 = w3760 & w11671;
assign w12872 = w3763 & w11673;
assign w12873 = w3767 & w11678;
assign v3995 = ~(w12872 | w12873);
assign w12874 = v3995;
assign w12875 = ~w12871 & w12874;
assign w12876 = ~w12870 & w12875;
assign w12877 = pi29 & ~w12876;
assign w12878 = ~pi29 & w12876;
assign v3996 = ~(w12877 | w12878);
assign w12879 = v3996;
assign w12880 = w12869 & w12879;
assign v3997 = ~(w12867 | w12880);
assign w12881 = v3997;
assign w12882 = ~w12714 & w12724;
assign v3998 = ~(w12725 | w12882);
assign w12883 = v3998;
assign w12884 = ~w12881 & w12883;
assign w12885 = w12881 & ~w12883;
assign v3999 = ~(w12884 | w12885);
assign w12886 = v3999;
assign w12887 = w4153 & ~w12351;
assign w12888 = w4155 & w12237;
assign w12889 = ~w2873 & w12084;
assign w12890 = w4158 & w12155;
assign v4000 = ~(w12889 | w12890);
assign w12891 = v4000;
assign w12892 = ~w12888 & w12891;
assign w12893 = ~w12887 & w12892;
assign w12894 = ~pi26 & w12893;
assign w12895 = pi26 & ~w12893;
assign v4001 = ~(w12894 | w12895);
assign w12896 = v4001;
assign w12897 = w12886 & w12896;
assign v4002 = ~(w12884 | w12897);
assign w12898 = v4002;
assign v4003 = ~(w12806 | w12816);
assign w12899 = v4003;
assign v4004 = ~(w12817 | w12899);
assign w12900 = v4004;
assign w12901 = ~w12898 & w12900;
assign w12902 = w12898 & ~w12900;
assign v4005 = ~(w12901 | w12902);
assign w12903 = v4005;
assign w12904 = w4764 & ~w12506;
assign w12905 = w4913 & ~w12406;
assign w12906 = w4763 & w12311;
assign w12907 = w4836 & w12381;
assign v4006 = ~(w12906 | w12907);
assign w12908 = v4006;
assign w12909 = ~w12905 & w12908;
assign w12910 = ~w12904 & w12909;
assign w12911 = ~pi23 & w12910;
assign w12912 = pi23 & ~w12910;
assign v4007 = ~(w12911 | w12912);
assign w12913 = v4007;
assign w12914 = w12903 & w12913;
assign v4008 = ~(w12901 | w12914);
assign w12915 = v4008;
assign w12916 = w4763 & w12381;
assign w12917 = w4764 & w12505;
assign v4009 = ~(w4836 | w12917);
assign w12918 = v4009;
assign v4010 = ~(w12406 | w12918);
assign w12919 = v4010;
assign v4011 = ~(w4913 | w12919);
assign w12920 = v4011;
assign w12921 = ~w12916 & w12920;
assign w12922 = ~pi23 & w12921;
assign w12923 = pi23 & ~w12921;
assign v4012 = ~(w12922 | w12923);
assign w12924 = v4012;
assign w12925 = ~w12915 & w12924;
assign w12926 = w12818 & ~w12820;
assign v4013 = ~(w12821 | w12926);
assign w12927 = v4013;
assign w12928 = w12915 & ~w12924;
assign v4014 = ~(w12925 | w12928);
assign w12929 = v4014;
assign w12930 = w12927 & w12929;
assign v4015 = ~(w12925 | w12930);
assign w12931 = v4015;
assign w12932 = ~w12836 & w12931;
assign w12933 = w12836 & ~w12931;
assign v4016 = ~(w12886 | w12896);
assign w12934 = v4016;
assign v4017 = ~(w12897 | w12934);
assign w12935 = v4017;
assign v4018 = ~(w12869 | w12879);
assign w12936 = v4018;
assign v4019 = ~(w12880 | w12936);
assign w12937 = v4019;
assign w12938 = w4153 & w12167;
assign w12939 = ~w2873 & w11984;
assign w12940 = w4155 & w12155;
assign v4020 = ~(w12939 | w12940);
assign w12941 = v4020;
assign w12942 = w4158 & w12084;
assign w12943 = w12941 & ~w12942;
assign w12944 = ~w12938 & w12943;
assign w12945 = pi26 & w12944;
assign v4021 = ~(pi26 | w12944);
assign w12946 = v4021;
assign v4022 = ~(w12945 | w12946);
assign w12947 = v4022;
assign w12948 = w12937 & ~w12947;
assign w12949 = w12685 & ~w12687;
assign v4023 = ~(w12688 | w12949);
assign w12950 = v4023;
assign v4024 = ~(w143 | w447);
assign w12951 = v4024;
assign w12952 = w4336 & w12951;
assign w12953 = w585 & w1414;
assign w12954 = w12952 & w12953;
assign w12955 = w3655 & w12954;
assign w12956 = ~w997 & w1805;
assign v4025 = ~(w260 | w493);
assign w12957 = v4025;
assign w12958 = ~w37 & w12957;
assign w12959 = w12956 & w12958;
assign w12960 = w1767 & w12959;
assign w12961 = w1814 & w1956;
assign w12962 = ~w329 & w2681;
assign w12963 = w12961 & w12962;
assign w12964 = w12960 & w12963;
assign w12965 = w5394 & w12964;
assign w12966 = w12955 & w12965;
assign w12967 = ~w180 & w996;
assign v4026 = ~(w123 | w548);
assign w12968 = v4026;
assign w12969 = w1853 & w12968;
assign w12970 = ~w438 & w12969;
assign w12971 = ~w235 & w12970;
assign w12972 = w12967 & w12971;
assign w12973 = w2325 & w4456;
assign w12974 = w883 & w12973;
assign w12975 = w2684 & w12974;
assign w12976 = w3829 & w12975;
assign w12977 = w12972 & w12976;
assign w12978 = w12966 & w12977;
assign w12979 = ~w88 & w233;
assign w12980 = w4088 & w12979;
assign w12981 = w188 & ~w420;
assign w12982 = w3911 & w12981;
assign w12983 = w1156 & w12982;
assign w12984 = w12980 & w12983;
assign w12985 = w2590 & w12984;
assign w12986 = w2756 & w12985;
assign w12987 = w12978 & w12986;
assign w12988 = ~w12660 & w12987;
assign w12989 = w12660 & ~w12987;
assign v4027 = ~(w12988 | w12989);
assign w12990 = v4027;
assign w12991 = (~w11880 & w11877) | (~w11880 & w28018) | (w11877 & w28018);
assign v4028 = ~(w11712 | w12991);
assign w12992 = v4028;
assign w12993 = ~w11882 & w12992;
assign v4029 = ~(w11884 | w12993);
assign w12994 = v4029;
assign w12995 = w928 & w12994;
assign w12996 = w3406 & w11700;
assign w12997 = w3399 & w11711;
assign w12998 = w3402 & w11708;
assign v4030 = ~(w12997 | w12998);
assign w12999 = v4030;
assign w13000 = ~w12996 & w12999;
assign w13001 = ~w12995 & w13000;
assign w13002 = w12990 & w13001;
assign v4031 = ~(w12988 | w13002);
assign w13003 = v4031;
assign w13004 = w12950 & w13003;
assign v4032 = ~(w12950 | w13003);
assign w13005 = v4032;
assign v4033 = ~(w13004 | w13005);
assign w13006 = v4033;
assign v4034 = ~(w11703 | w11885);
assign w13007 = v4034;
assign v4035 = ~(w11886 | w13007);
assign w13008 = v4035;
assign w13009 = w928 & ~w13008;
assign w13010 = w3406 & ~w11695;
assign w13011 = w3402 & w11700;
assign w13012 = w3399 & w11708;
assign v4036 = ~(w13011 | w13012);
assign w13013 = v4036;
assign w13014 = ~w13010 & w13013;
assign w13015 = ~w13009 & w13014;
assign w13016 = w13006 & ~w13015;
assign v4037 = ~(w13004 | w13016);
assign w13017 = v4037;
assign w13018 = ~w12692 & w12701;
assign v4038 = ~(w12702 | w13018);
assign w13019 = v4038;
assign w13020 = ~w13017 & w13019;
assign w13021 = w13017 & ~w13019;
assign v4039 = ~(w13020 | w13021);
assign w13022 = v4039;
assign w13023 = w3529 & w12594;
assign w13024 = w3760 & w11678;
assign w13025 = w3763 & ~w11683;
assign w13026 = w3767 & w11686;
assign v4040 = ~(w13025 | w13026);
assign w13027 = v4040;
assign w13028 = ~w13024 & w13027;
assign w13029 = ~w13023 & w13028;
assign w13030 = pi29 & ~w13029;
assign w13031 = ~pi29 & w13029;
assign v4041 = ~(w13030 | w13031);
assign w13032 = v4041;
assign w13033 = w13022 & w13032;
assign v4042 = ~(w13020 | w13033);
assign w13034 = v4042;
assign w13035 = ~w12852 & w12862;
assign v4043 = ~(w12863 | w13035);
assign w13036 = v4043;
assign w13037 = ~w13034 & w13036;
assign w13038 = w13034 & ~w13036;
assign v4044 = ~(w13037 | w13038);
assign w13039 = v4044;
assign w13040 = w4153 & w12181;
assign w13041 = w4155 & w12084;
assign w13042 = ~w2873 & w11671;
assign w13043 = w4158 & w11984;
assign v4045 = ~(w13042 | w13043);
assign w13044 = v4045;
assign w13045 = ~w13041 & w13044;
assign w13046 = ~w13040 & w13045;
assign w13047 = pi26 & ~w13046;
assign w13048 = ~pi26 & w13046;
assign v4046 = ~(w13047 | w13048);
assign w13049 = v4046;
assign w13050 = w13039 & w13049;
assign v4047 = ~(w13037 | w13050);
assign w13051 = v4047;
assign w13052 = ~w12937 & w12947;
assign v4048 = ~(w12948 | w13052);
assign w13053 = v4048;
assign w13054 = ~w13051 & w13053;
assign v4049 = ~(w12948 | w13054);
assign w13055 = v4049;
assign w13056 = w12935 & ~w13055;
assign w13057 = ~w12935 & w13055;
assign v4050 = ~(w13056 | w13057);
assign w13058 = v4050;
assign w13059 = w4764 & w12387;
assign w13060 = w4913 & w12381;
assign w13061 = w4763 & w12271;
assign w13062 = w4836 & w12311;
assign v4051 = ~(w13061 | w13062);
assign w13063 = v4051;
assign w13064 = ~w13060 & w13063;
assign w13065 = ~w13059 & w13064;
assign w13066 = ~pi23 & w13065;
assign w13067 = pi23 & ~w13065;
assign v4052 = ~(w13066 | w13067);
assign w13068 = v4052;
assign w13069 = w13058 & w13068;
assign v4053 = ~(w13056 | w13069);
assign w13070 = v4053;
assign w13071 = w919 & ~w13070;
assign v4054 = ~(w12903 | w12913);
assign w13072 = v4054;
assign v4055 = ~(w12914 | w13072);
assign w13073 = v4055;
assign w13074 = ~w919 & w13070;
assign v4056 = ~(w13071 | w13074);
assign w13075 = v4056;
assign w13076 = w13073 & w13075;
assign v4057 = ~(w13071 | w13076);
assign w13077 = v4057;
assign v4058 = ~(w12927 | w12929);
assign w13078 = v4058;
assign v4059 = ~(w12930 | w13078);
assign w13079 = v4059;
assign w13080 = ~w13077 & w13079;
assign w13081 = w13077 & ~w13079;
assign v4060 = ~(w13080 | w13081);
assign w13082 = v4060;
assign v4061 = ~(w13073 | w13075);
assign w13083 = v4061;
assign v4062 = ~(w13076 | w13083);
assign w13084 = v4062;
assign v4063 = ~(w13058 | w13068);
assign w13085 = v4063;
assign v4064 = ~(w13069 | w13085);
assign w13086 = v4064;
assign w13087 = w13051 & ~w13053;
assign v4065 = ~(w13054 | w13087);
assign w13088 = v4065;
assign w13089 = w4764 & w12318;
assign w13090 = w4836 & w12271;
assign w13091 = w4913 & w12311;
assign v4066 = ~(w13090 | w13091);
assign w13092 = v4066;
assign w13093 = w4763 & w12237;
assign w13094 = w13092 & ~w13093;
assign w13095 = ~w13089 & w13094;
assign w13096 = pi23 & w13095;
assign v4067 = ~(pi23 | w13095);
assign w13097 = v4067;
assign v4068 = ~(w13096 | w13097);
assign w13098 = v4068;
assign w13099 = w13088 & ~w13098;
assign v4069 = ~(w13039 | w13049);
assign w13100 = v4069;
assign v4070 = ~(w13050 | w13100);
assign w13101 = v4070;
assign w13102 = ~w13006 & w13015;
assign v4071 = ~(w13016 | w13102);
assign w13103 = v4071;
assign w13104 = w3529 & w12610;
assign w13105 = w3763 & w11686;
assign w13106 = w3760 & ~w11683;
assign v4072 = ~(w13105 | w13106);
assign w13107 = v4072;
assign w13108 = w3767 & w11689;
assign w13109 = w13107 & ~w13108;
assign w13110 = ~w13104 & w13109;
assign v4073 = ~(pi29 | w13110);
assign w13111 = v4073;
assign w13112 = pi29 & w13110;
assign v4074 = ~(w13111 | w13112);
assign w13113 = v4074;
assign w13114 = w13103 & ~w13113;
assign w13115 = w576 & w2905;
assign w13116 = ~w666 & w5216;
assign w13117 = w13115 & w13116;
assign w13118 = w1330 & w2681;
assign w13119 = w12117 & w13118;
assign w13120 = w13117 & w13119;
assign w13121 = ~w215 & w449;
assign v4075 = ~(w56 | w235);
assign w13122 = v4075;
assign w13123 = w13121 & w13122;
assign w13124 = w2125 & w13123;
assign v4076 = ~(w324 | w566);
assign w13125 = v4076;
assign w13126 = w5007 & w13125;
assign w13127 = w2803 & w13126;
assign w13128 = ~w238 & w13127;
assign w13129 = w13124 & w13128;
assign w13130 = w13120 & w13129;
assign w13131 = w2693 & w13130;
assign v4077 = ~(w431 | w484);
assign w13132 = v4077;
assign w13133 = w2282 & w13132;
assign w13134 = ~w107 & w6661;
assign w13135 = w13133 & w13134;
assign w13136 = w4497 & w13135;
assign w13137 = w740 & w3737;
assign w13138 = ~w711 & w13137;
assign w13139 = ~w303 & w13138;
assign w13140 = w13136 & w13139;
assign w13141 = w13131 & w13140;
assign w13142 = w3311 & w6099;
assign w13143 = w13141 & w13142;
assign v4078 = ~(w192 | w244);
assign w13144 = v4078;
assign w13145 = w2929 & w13144;
assign w13146 = w1981 & w13145;
assign w13147 = ~w179 & w13146;
assign w13148 = w1827 & w13147;
assign v4079 = ~(w239 | w739);
assign w13149 = v4079;
assign w13150 = w2951 & w13149;
assign w13151 = ~w343 & w13150;
assign w13152 = w13148 & w13151;
assign w13153 = w5836 & w13152;
assign w13154 = w1963 & w3696;
assign v4080 = ~(w581 | w978);
assign w13155 = v4080;
assign w13156 = w1799 & w13155;
assign w13157 = w1989 & w13156;
assign w13158 = w665 & w13157;
assign w13159 = w3133 & w13158;
assign w13160 = w3609 & w13159;
assign w13161 = w1403 & w13160;
assign w13162 = w13154 & w13161;
assign w13163 = w13153 & w13162;
assign v4081 = ~(w13143 | w13163);
assign w13164 = v4081;
assign w13165 = pi11 & ~w7176;
assign w13166 = ~pi08 & w7173;
assign v4082 = ~(w13165 | w13166);
assign w13167 = v4082;
assign w13168 = w13143 & w13163;
assign v4083 = ~(w13164 | w13168);
assign w13169 = v4083;
assign w13170 = ~w13167 & w13169;
assign v4084 = ~(w13164 | w13170);
assign w13171 = v4084;
assign w13172 = w12660 & ~w13171;
assign w13173 = ~w12660 & w13171;
assign v4085 = ~(w13172 | w13173);
assign w13174 = v4085;
assign v4086 = ~(w11712 | w11880);
assign w13175 = v4086;
assign w13176 = w11878 & ~w13175;
assign w13177 = ~w11878 & w13175;
assign v4087 = ~(w13176 | w13177);
assign w13178 = v4087;
assign w13179 = w928 & w13178;
assign w13180 = w3406 & w11708;
assign w13181 = w3399 & w11714;
assign w13182 = w3402 & w11711;
assign v4088 = ~(w13181 | w13182);
assign w13183 = v4088;
assign w13184 = ~w13180 & w13183;
assign w13185 = ~w13179 & w13184;
assign w13186 = w13174 & ~w13185;
assign v4089 = ~(w13172 | w13186);
assign w13187 = v4089;
assign v4090 = ~(w12990 | w13001);
assign w13188 = v4090;
assign v4091 = ~(w13002 | w13188);
assign w13189 = v4091;
assign v4092 = ~(w13187 | w13189);
assign w13190 = v4092;
assign w13191 = w13167 & ~w13169;
assign v4093 = ~(w13170 | w13191);
assign w13192 = v4093;
assign w13193 = ~w11873 & w28019;
assign v4094 = ~(w11877 | w13193);
assign w13194 = v4094;
assign w13195 = w928 & w13194;
assign w13196 = w3406 & w11711;
assign w13197 = w3402 & w11714;
assign w13198 = w3399 & w11720;
assign v4095 = ~(w13197 | w13198);
assign w13199 = v4095;
assign w13200 = ~w13196 & w13199;
assign w13201 = ~w13195 & w13200;
assign w13202 = w13192 & ~w13201;
assign w13203 = ~w13192 & w13201;
assign v4096 = ~(w13202 | w13203);
assign w13204 = v4096;
assign w13205 = ~w49 & w442;
assign w13206 = w2107 & w4661;
assign w13207 = w13205 & w13206;
assign w13208 = ~w418 & w6478;
assign w13209 = w1542 & w13208;
assign w13210 = w3204 & w13209;
assign w13211 = w13207 & w13210;
assign w13212 = ~w245 & w1081;
assign w13213 = ~w533 & w13212;
assign v4097 = ~(w82 | w179);
assign w13214 = v4097;
assign w13215 = ~w624 & w13214;
assign w13216 = w13213 & w13215;
assign w13217 = w887 & w3015;
assign w13218 = w222 & w13217;
assign w13219 = w1455 & w13218;
assign w13220 = w13216 & w13219;
assign w13221 = w2610 & w13220;
assign w13222 = w13211 & w13221;
assign v4098 = ~(w128 | w522);
assign w13223 = v4098;
assign w13224 = w3965 & w13223;
assign w13225 = w2342 & w13224;
assign w13226 = w2824 & w5174;
assign w13227 = w1647 & w5222;
assign w13228 = w13226 & w13227;
assign w13229 = ~w215 & w684;
assign w13230 = w2052 & w13229;
assign w13231 = w13228 & w13230;
assign w13232 = w13225 & w13231;
assign w13233 = ~w642 & w1768;
assign w13234 = w1449 & w13233;
assign v4099 = ~(w103 | w280);
assign w13235 = v4099;
assign w13236 = w12953 & w13235;
assign w13237 = w13234 & w13236;
assign w13238 = w1252 & w5012;
assign w13239 = w13237 & w13238;
assign w13240 = w13232 & w13239;
assign w13241 = w4560 & w13240;
assign w13242 = w13222 & w13241;
assign w13243 = w13143 & ~w13242;
assign w13244 = ~w640 & w2433;
assign w13245 = w2159 & w4480;
assign w13246 = w13244 & w13245;
assign w13247 = ~w201 & w2757;
assign w13248 = w883 & w1120;
assign w13249 = w13247 & w13248;
assign w13250 = w3861 & w13249;
assign w13251 = w13246 & w13250;
assign w13252 = w395 & w13251;
assign v4100 = ~(w742 | w1108);
assign w13253 = v4100;
assign w13254 = w1340 & w13253;
assign w13255 = w101 & w4491;
assign w13256 = w13254 & w13255;
assign w13257 = w532 & w2382;
assign w13258 = w13256 & w13257;
assign w13259 = w1042 & w13258;
assign w13260 = w708 & w6583;
assign w13261 = w13259 & w13260;
assign w13262 = w13252 & w13261;
assign v4101 = ~(w179 | w312);
assign w13263 = v4101;
assign w13264 = w1076 & w13263;
assign v4102 = ~(w216 | w749);
assign w13265 = v4102;
assign w13266 = w13264 & w13265;
assign w13267 = w1380 & w13266;
assign w13268 = w290 & w2671;
assign w13269 = w3637 & w13268;
assign w13270 = w13267 & w13269;
assign w13271 = w13262 & w13270;
assign w13272 = w1006 & w13271;
assign w13273 = w852 & w1121;
assign w13274 = w11927 & w13273;
assign w13275 = w1177 & w1759;
assign w13276 = w836 & w13275;
assign v4103 = ~(w162 | w484);
assign w13277 = v4103;
assign w13278 = w449 & w13277;
assign w13279 = w2718 & w13278;
assign w13280 = w13276 & w13279;
assign w13281 = w1413 & w13280;
assign w13282 = ~w652 & w2571;
assign w13283 = w5203 & w13282;
assign w13284 = ~w441 & w1202;
assign v4104 = ~(w82 | w307);
assign w13285 = v4104;
assign w13286 = w3115 & w13285;
assign w13287 = w1626 & w13286;
assign w13288 = w13284 & w13287;
assign w13289 = w3952 & w4651;
assign v4105 = ~(w317 | w388);
assign w13290 = v4105;
assign w13291 = ~w1134 & w13290;
assign w13292 = w13289 & w13291;
assign w13293 = w13288 & w13292;
assign w13294 = w13283 & w13293;
assign w13295 = w13281 & w13294;
assign w13296 = w2021 & w13295;
assign w13297 = w13274 & w13296;
assign v4106 = ~(w13272 | w13297);
assign w13298 = v4106;
assign w13299 = pi08 & ~w8139;
assign w13300 = ~pi07 & w8136;
assign v4107 = ~(w13299 | w13300);
assign w13301 = v4107;
assign w13302 = w13272 & w13297;
assign v4108 = ~(w13298 | w13302);
assign w13303 = v4108;
assign w13304 = ~w13301 & w13303;
assign v4109 = ~(w13298 | w13304);
assign w13305 = v4109;
assign w13306 = w13143 & ~w13305;
assign w13307 = ~w13143 & w13305;
assign v4110 = ~(w13306 | w13307);
assign w13308 = v4110;
assign w13309 = ~w11865 & w28020;
assign v4111 = ~(w11869 | w13309);
assign w13310 = v4111;
assign w13311 = w928 & ~w13310;
assign w13312 = w3406 & w11720;
assign w13313 = w3402 & w11723;
assign w13314 = w3399 & w11726;
assign v4112 = ~(w13313 | w13314);
assign w13315 = v4112;
assign w13316 = ~w13312 & w13315;
assign w13317 = ~w13311 & w13316;
assign w13318 = w13308 & ~w13317;
assign v4113 = ~(w13306 | w13318);
assign w13319 = v4113;
assign w13320 = ~w13143 & w13242;
assign v4114 = ~(w13243 | w13320);
assign w13321 = v4114;
assign w13322 = ~w13319 & w13321;
assign v4115 = ~(w13243 | w13322);
assign w13323 = v4115;
assign w13324 = w13204 & ~w13323;
assign v4116 = ~(w13202 | w13324);
assign w13325 = v4116;
assign w13326 = ~w13174 & w13185;
assign v4117 = ~(w13186 | w13326);
assign w13327 = v4117;
assign w13328 = ~w13325 & w13327;
assign w13329 = w13325 & ~w13327;
assign v4118 = ~(w13328 | w13329);
assign w13330 = v4118;
assign w13331 = w3529 & w12694;
assign w13332 = w3760 & w11689;
assign w13333 = w3767 & w11700;
assign w13334 = w3763 & ~w11695;
assign v4119 = ~(w13333 | w13334);
assign w13335 = v4119;
assign w13336 = ~w13332 & w13335;
assign w13337 = ~w13331 & w13336;
assign w13338 = pi29 & w13337;
assign v4120 = ~(pi29 | w13337);
assign w13339 = v4120;
assign v4121 = ~(w13338 | w13339);
assign w13340 = v4121;
assign w13341 = w13330 & ~w13340;
assign v4122 = ~(w13328 | w13341);
assign w13342 = v4122;
assign w13343 = w13187 & w13189;
assign v4123 = ~(w13190 | w13343);
assign w13344 = v4123;
assign w13345 = ~w13342 & w13344;
assign v4124 = ~(w13190 | w13345);
assign w13346 = v4124;
assign w13347 = ~w13103 & w13113;
assign v4125 = ~(w13114 | w13347);
assign w13348 = v4125;
assign w13349 = ~w13346 & w13348;
assign v4126 = ~(w13114 | w13349);
assign w13350 = v4126;
assign v4127 = ~(w13022 | w13032);
assign w13351 = v4127;
assign v4128 = ~(w13033 | w13351);
assign w13352 = v4128;
assign w13353 = ~w13350 & w13352;
assign w13354 = w13350 & ~w13352;
assign v4129 = ~(w13353 | w13354);
assign w13355 = v4129;
assign w13356 = w4153 & w11993;
assign w13357 = w4155 & w11984;
assign w13358 = w4158 & w11671;
assign w13359 = ~w2873 & w11673;
assign v4130 = ~(w13358 | w13359);
assign w13360 = v4130;
assign w13361 = ~w13357 & w13360;
assign w13362 = ~w13356 & w13361;
assign w13363 = ~pi26 & w13362;
assign w13364 = pi26 & ~w13362;
assign v4131 = ~(w13363 | w13364);
assign w13365 = v4131;
assign w13366 = w13355 & w13365;
assign v4132 = ~(w13353 | w13366);
assign w13367 = v4132;
assign w13368 = w13101 & ~w13367;
assign w13369 = ~w13101 & w13367;
assign v4133 = ~(w13368 | w13369);
assign w13370 = v4133;
assign w13371 = w4764 & ~w12277;
assign w13372 = w4836 & w12237;
assign w13373 = w4913 & w12271;
assign v4134 = ~(w13372 | w13373);
assign w13374 = v4134;
assign w13375 = w4763 & w12155;
assign w13376 = w13374 & ~w13375;
assign w13377 = ~w13371 & w13376;
assign w13378 = pi23 & w13377;
assign v4135 = ~(pi23 | w13377);
assign w13379 = v4135;
assign v4136 = ~(w13378 | w13379);
assign w13380 = v4136;
assign w13381 = w13370 & ~w13380;
assign v4137 = ~(w13368 | w13381);
assign w13382 = v4137;
assign w13383 = ~w13088 & w13098;
assign v4138 = ~(w13099 | w13383);
assign w13384 = v4138;
assign w13385 = ~w13382 & w13384;
assign v4139 = ~(w13099 | w13385);
assign w13386 = v4139;
assign w13387 = w13086 & ~w13386;
assign w13388 = ~w13086 & w13386;
assign v4140 = ~(w13387 | w13388);
assign w13389 = v4140;
assign w13390 = pi20 & w12406;
assign w13391 = pi19 & ~w12406;
assign v4141 = ~(w13390 | w13391);
assign w13392 = v4141;
assign w13393 = w916 & w13392;
assign v4142 = ~(w917 | w13393);
assign w13394 = v4142;
assign w13395 = w13389 & w13394;
assign v4143 = ~(w13387 | w13395);
assign w13396 = v4143;
assign w13397 = ~w13084 & w13396;
assign w13398 = w13084 & ~w13396;
assign v4144 = ~(w13389 | w13394);
assign w13399 = v4144;
assign v4145 = ~(w13395 | w13399);
assign w13400 = v4145;
assign w13401 = ~w13370 & w13380;
assign v4146 = ~(w13381 | w13401);
assign w13402 = v4146;
assign v4147 = ~(w13355 | w13365);
assign w13403 = v4147;
assign v4148 = ~(w13366 | w13403);
assign w13404 = v4148;
assign w13405 = w13346 & ~w13348;
assign v4149 = ~(w13349 | w13405);
assign w13406 = v4149;
assign w13407 = w4153 & w12469;
assign w13408 = ~w2873 & w11678;
assign w13409 = w4155 & w11671;
assign v4150 = ~(w13408 | w13409);
assign w13410 = v4150;
assign w13411 = w4158 & w11673;
assign w13412 = w13410 & ~w13411;
assign w13413 = ~w13407 & w13412;
assign v4151 = ~(pi26 | w13413);
assign w13414 = v4151;
assign w13415 = pi26 & w13413;
assign v4152 = ~(w13414 | w13415);
assign w13416 = v4152;
assign w13417 = w13406 & ~w13416;
assign w13418 = ~w13406 & w13416;
assign v4153 = ~(w13417 | w13418);
assign w13419 = v4153;
assign w13420 = w13342 & ~w13344;
assign v4154 = ~(w13345 | w13420);
assign w13421 = v4154;
assign w13422 = w3529 & ~w12842;
assign w13423 = w3760 & w11686;
assign w13424 = w3763 & w11689;
assign w13425 = w3767 & ~w11695;
assign v4155 = ~(w13424 | w13425);
assign w13426 = v4155;
assign w13427 = ~w13423 & w13426;
assign w13428 = ~w13422 & w13427;
assign w13429 = pi29 & w13428;
assign v4156 = ~(pi29 | w13428);
assign w13430 = v4156;
assign v4157 = ~(w13429 | w13430);
assign w13431 = v4157;
assign w13432 = w13421 & ~w13431;
assign w13433 = ~w13421 & w13431;
assign v4158 = ~(w13432 | w13433);
assign w13434 = v4158;
assign w13435 = w4153 & w12454;
assign w13436 = w4155 & w11673;
assign v4159 = ~(w2873 | w11683);
assign w13437 = v4159;
assign w13438 = w4158 & w11678;
assign v4160 = ~(w13437 | w13438);
assign w13439 = v4160;
assign w13440 = ~w13436 & w13439;
assign w13441 = ~w13435 & w13440;
assign w13442 = ~pi26 & w13441;
assign w13443 = pi26 & ~w13441;
assign v4161 = ~(w13442 | w13443);
assign w13444 = v4161;
assign w13445 = w13434 & w13444;
assign v4162 = ~(w13432 | w13445);
assign w13446 = v4162;
assign w13447 = w13419 & ~w13446;
assign v4163 = ~(w13417 | w13447);
assign w13448 = v4163;
assign w13449 = w13404 & ~w13448;
assign w13450 = ~w13404 & w13448;
assign v4164 = ~(w13449 | w13450);
assign w13451 = v4164;
assign w13452 = w4764 & ~w12351;
assign w13453 = w4836 & w12155;
assign w13454 = w4913 & w12237;
assign v4165 = ~(w13453 | w13454);
assign w13455 = v4165;
assign w13456 = w4763 & w12084;
assign w13457 = w13455 & ~w13456;
assign w13458 = ~w13452 & w13457;
assign w13459 = pi23 & w13458;
assign v4166 = ~(pi23 | w13458);
assign w13460 = v4166;
assign v4167 = ~(w13459 | w13460);
assign w13461 = v4167;
assign w13462 = w13451 & ~w13461;
assign v4168 = ~(w13449 | w13462);
assign w13463 = v4168;
assign w13464 = w13402 & ~w13463;
assign w13465 = ~w13402 & w13463;
assign v4169 = ~(w13464 | w13465);
assign w13466 = v4169;
assign w13467 = w5114 & ~w12506;
assign w13468 = w5610 & ~w12406;
assign w13469 = w5113 & w12311;
assign w13470 = w5531 & w12381;
assign v4170 = ~(w13469 | w13470);
assign w13471 = v4170;
assign w13472 = ~w13468 & w13471;
assign w13473 = ~w13467 & w13472;
assign w13474 = ~pi20 & w13473;
assign w13475 = pi20 & ~w13473;
assign v4171 = ~(w13474 | w13475);
assign w13476 = v4171;
assign w13477 = w13466 & w13476;
assign v4172 = ~(w13464 | w13477);
assign w13478 = v4172;
assign w13479 = w5113 & w12381;
assign w13480 = w5114 & w12505;
assign v4173 = ~(w5531 | w13480);
assign w13481 = v4173;
assign v4174 = ~(w12406 | w13481);
assign w13482 = v4174;
assign v4175 = ~(w5610 | w13482);
assign w13483 = v4175;
assign w13484 = ~w13479 & w13483;
assign w13485 = ~pi20 & w13484;
assign w13486 = pi20 & ~w13484;
assign v4176 = ~(w13485 | w13486);
assign w13487 = v4176;
assign w13488 = ~w13478 & w13487;
assign w13489 = w13382 & ~w13384;
assign v4177 = ~(w13385 | w13489);
assign w13490 = v4177;
assign w13491 = w13478 & ~w13487;
assign v4178 = ~(w13488 | w13491);
assign w13492 = v4178;
assign w13493 = w13490 & w13492;
assign v4179 = ~(w13488 | w13493);
assign w13494 = v4179;
assign w13495 = w13400 & ~w13494;
assign w13496 = ~w13451 & w13461;
assign v4180 = ~(w13462 | w13496);
assign w13497 = v4180;
assign w13498 = ~w13419 & w13446;
assign v4181 = ~(w13447 | w13498);
assign w13499 = v4181;
assign w13500 = w4764 & w12167;
assign w13501 = w4913 & w12155;
assign w13502 = w4763 & w11984;
assign w13503 = w4836 & w12084;
assign v4182 = ~(w13502 | w13503);
assign w13504 = v4182;
assign w13505 = ~w13501 & w13504;
assign w13506 = ~w13500 & w13505;
assign w13507 = ~pi23 & w13506;
assign w13508 = pi23 & ~w13506;
assign v4183 = ~(w13507 | w13508);
assign w13509 = v4183;
assign w13510 = w13499 & w13509;
assign w13511 = w13319 & ~w13321;
assign v4184 = ~(w13322 | w13511);
assign w13512 = v4184;
assign w13513 = (~w11872 & w11869) | (~w11872 & w28021) | (w11869 & w28021);
assign v4185 = ~(w11873 | w13513);
assign w13514 = v4185;
assign w13515 = w928 & w13514;
assign w13516 = w3406 & w11714;
assign w13517 = w3402 & w11720;
assign w13518 = w3399 & w11723;
assign v4186 = ~(w13517 | w13518);
assign w13519 = v4186;
assign w13520 = ~w13516 & w13519;
assign w13521 = ~w13515 & w13520;
assign w13522 = w13512 & ~w13521;
assign w13523 = ~w13512 & w13521;
assign v4187 = ~(w13522 | w13523);
assign w13524 = v4187;
assign w13525 = w3529 & w12994;
assign w13526 = w3760 & w11700;
assign w13527 = w3767 & w11711;
assign w13528 = w3763 & w11708;
assign v4188 = ~(w13527 | w13528);
assign w13529 = v4188;
assign w13530 = ~w13526 & w13529;
assign w13531 = ~w13525 & w13530;
assign w13532 = pi29 & ~w13531;
assign w13533 = ~pi29 & w13531;
assign v4189 = ~(w13532 | w13533);
assign w13534 = v4189;
assign w13535 = w13524 & w13534;
assign v4190 = ~(w13522 | w13535);
assign w13536 = v4190;
assign w13537 = ~w13204 & w13323;
assign v4191 = ~(w13324 | w13537);
assign w13538 = v4191;
assign w13539 = ~w13536 & w13538;
assign w13540 = w13536 & ~w13538;
assign v4192 = ~(w13539 | w13540);
assign w13541 = v4192;
assign w13542 = w3529 & ~w13008;
assign w13543 = w3760 & ~w11695;
assign w13544 = w3763 & w11700;
assign w13545 = w3767 & w11708;
assign v4193 = ~(w13544 | w13545);
assign w13546 = v4193;
assign w13547 = ~w13543 & w13546;
assign w13548 = ~w13542 & w13547;
assign w13549 = pi29 & w13548;
assign v4194 = ~(pi29 | w13548);
assign w13550 = v4194;
assign v4195 = ~(w13549 | w13550);
assign w13551 = v4195;
assign w13552 = w13541 & ~w13551;
assign v4196 = ~(w13539 | w13552);
assign w13553 = v4196;
assign w13554 = ~w13330 & w13340;
assign v4197 = ~(w13341 | w13554);
assign w13555 = v4197;
assign w13556 = ~w13553 & w13555;
assign w13557 = w13553 & ~w13555;
assign v4198 = ~(w13556 | w13557);
assign w13558 = v4198;
assign w13559 = w4153 & w12594;
assign w13560 = w4155 & w11678;
assign w13561 = ~w2873 & w11686;
assign w13562 = w4158 & ~w11683;
assign v4199 = ~(w13561 | w13562);
assign w13563 = v4199;
assign w13564 = ~w13560 & w13563;
assign w13565 = ~w13559 & w13564;
assign w13566 = ~pi26 & w13565;
assign w13567 = pi26 & ~w13565;
assign v4200 = ~(w13566 | w13567);
assign w13568 = v4200;
assign w13569 = w13558 & w13568;
assign v4201 = ~(w13556 | w13569);
assign w13570 = v4201;
assign v4202 = ~(w13434 | w13444);
assign w13571 = v4202;
assign v4203 = ~(w13445 | w13571);
assign w13572 = v4203;
assign w13573 = ~w13570 & w13572;
assign w13574 = w13570 & ~w13572;
assign v4204 = ~(w13573 | w13574);
assign w13575 = v4204;
assign w13576 = w4764 & w12181;
assign w13577 = w4836 & w11984;
assign w13578 = w4913 & w12084;
assign v4205 = ~(w13577 | w13578);
assign w13579 = v4205;
assign w13580 = w4763 & w11671;
assign w13581 = w13579 & ~w13580;
assign w13582 = ~w13576 & w13581;
assign v4206 = ~(pi23 | w13582);
assign w13583 = v4206;
assign w13584 = pi23 & w13582;
assign v4207 = ~(w13583 | w13584);
assign w13585 = v4207;
assign w13586 = w13575 & ~w13585;
assign v4208 = ~(w13573 | w13586);
assign w13587 = v4208;
assign v4209 = ~(w13499 | w13509);
assign w13588 = v4209;
assign v4210 = ~(w13510 | w13588);
assign w13589 = v4210;
assign w13590 = ~w13587 & w13589;
assign v4211 = ~(w13510 | w13590);
assign w13591 = v4211;
assign w13592 = w13497 & ~w13591;
assign w13593 = ~w13497 & w13591;
assign v4212 = ~(w13592 | w13593);
assign w13594 = v4212;
assign w13595 = w5114 & w12387;
assign w13596 = w5610 & w12381;
assign w13597 = w5113 & w12271;
assign w13598 = w5531 & w12311;
assign v4213 = ~(w13597 | w13598);
assign w13599 = v4213;
assign w13600 = ~w13596 & w13599;
assign w13601 = ~w13595 & w13600;
assign w13602 = ~pi20 & w13601;
assign w13603 = pi20 & ~w13601;
assign v4214 = ~(w13602 | w13603);
assign w13604 = v4214;
assign w13605 = w13594 & w13604;
assign v4215 = ~(w13592 | w13605);
assign w13606 = v4215;
assign w13607 = w12582 & ~w13606;
assign v4216 = ~(w13466 | w13476);
assign w13608 = v4216;
assign v4217 = ~(w13477 | w13608);
assign w13609 = v4217;
assign w13610 = ~w12582 & w13606;
assign v4218 = ~(w13607 | w13610);
assign w13611 = v4218;
assign w13612 = w13609 & w13611;
assign v4219 = ~(w13607 | w13612);
assign w13613 = v4219;
assign v4220 = ~(w13490 | w13492);
assign w13614 = v4220;
assign v4221 = ~(w13493 | w13614);
assign w13615 = v4221;
assign w13616 = ~w13613 & w13615;
assign w13617 = w13613 & ~w13615;
assign v4222 = ~(w13616 | w13617);
assign w13618 = v4222;
assign v4223 = ~(w13609 | w13611);
assign w13619 = v4223;
assign v4224 = ~(w13612 | w13619);
assign w13620 = v4224;
assign v4225 = ~(w13594 | w13604);
assign w13621 = v4225;
assign v4226 = ~(w13605 | w13621);
assign w13622 = v4226;
assign w13623 = w13587 & ~w13589;
assign v4227 = ~(w13590 | w13623);
assign w13624 = v4227;
assign w13625 = w5114 & w12318;
assign w13626 = w5531 & w12271;
assign w13627 = w5610 & w12311;
assign v4228 = ~(w13626 | w13627);
assign w13628 = v4228;
assign w13629 = w5113 & w12237;
assign w13630 = w13628 & ~w13629;
assign w13631 = ~w13625 & w13630;
assign w13632 = pi20 & w13631;
assign v4229 = ~(pi20 | w13631);
assign w13633 = v4229;
assign v4230 = ~(w13632 | w13633);
assign w13634 = v4230;
assign w13635 = w13624 & ~w13634;
assign w13636 = ~w13575 & w13585;
assign v4231 = ~(w13586 | w13636);
assign w13637 = v4231;
assign v4232 = ~(w13558 | w13568);
assign w13638 = v4232;
assign v4233 = ~(w13569 | w13638);
assign w13639 = v4233;
assign w13640 = ~w13541 & w13551;
assign v4234 = ~(w13552 | w13640);
assign w13641 = v4234;
assign w13642 = w4153 & w12610;
assign w13643 = w4155 & ~w11683;
assign w13644 = ~w2873 & w11689;
assign w13645 = w4158 & w11686;
assign v4235 = ~(w13644 | w13645);
assign w13646 = v4235;
assign w13647 = ~w13643 & w13646;
assign w13648 = ~w13642 & w13647;
assign w13649 = pi26 & ~w13648;
assign w13650 = ~pi26 & w13648;
assign v4236 = ~(w13649 | w13650);
assign w13651 = v4236;
assign w13652 = w13641 & w13651;
assign w13653 = ~w13308 & w13317;
assign v4237 = ~(w13318 | w13653);
assign w13654 = v4237;
assign w13655 = w13301 & ~w13303;
assign v4238 = ~(w13304 | w13655);
assign w13656 = v4238;
assign v4239 = ~(pi02 | w10986);
assign w13657 = v4239;
assign w13658 = w1405 & w12661;
assign w13659 = w2878 & w13658;
assign w13660 = w724 & w13659;
assign w13661 = ~w338 & w1220;
assign w13662 = w1026 & w13661;
assign w13663 = w11613 & w13662;
assign w13664 = ~w299 & w13663;
assign w13665 = w13660 & w13664;
assign w13666 = w1436 & ~w3816;
assign w13667 = w386 & w3107;
assign w13668 = w13666 & w13667;
assign w13669 = w1127 & w2444;
assign w13670 = w313 & w13669;
assign w13671 = w13668 & w13670;
assign v4240 = ~(w99 | w135);
assign w13672 = v4240;
assign w13673 = ~w224 & w13672;
assign w13674 = w3533 & w13673;
assign w13675 = w13671 & w13674;
assign w13676 = ~w292 & w658;
assign w13677 = ~w522 & w13676;
assign w13678 = w13213 & w13677;
assign w13679 = w779 & w13678;
assign w13680 = w13675 & w13679;
assign w13681 = w13665 & w13680;
assign w13682 = w895 & w3475;
assign w13683 = ~w211 & w1398;
assign w13684 = w743 & w13683;
assign w13685 = w6111 & w13684;
assign w13686 = w13682 & w13685;
assign w13687 = ~w280 & w1425;
assign w13688 = w2319 & w13687;
assign w13689 = w6634 & w13688;
assign w13690 = w4259 & w13689;
assign w13691 = w13686 & w13690;
assign w13692 = w13129 & w13691;
assign w13693 = w13681 & w13692;
assign v4241 = ~(w13657 | w13693);
assign w13694 = v4241;
assign w13695 = pi05 & ~w9400;
assign w13696 = ~pi02 & w9397;
assign v4242 = ~(w13695 | w13696);
assign w13697 = v4242;
assign w13698 = w13657 & w13693;
assign v4243 = ~(w13694 | w13698);
assign w13699 = v4243;
assign w13700 = ~w13697 & w13699;
assign v4244 = ~(w13694 | w13700);
assign w13701 = v4244;
assign w13702 = (~w11857 & w11854) | (~w11857 & w28022) | (w11854 & w28022);
assign v4245 = ~(w11858 | w13702);
assign w13703 = v4245;
assign w13704 = w928 & ~w13703;
assign w13705 = w3406 & w11729;
assign w13706 = w3399 & w11737;
assign w13707 = w3402 & ~w11734;
assign v4246 = ~(w13706 | w13707);
assign w13708 = v4246;
assign w13709 = ~w13705 & w13708;
assign w13710 = ~w13704 & w13709;
assign v4247 = ~(w13701 | w13710);
assign w13711 = v4247;
assign v4248 = ~(w13272 | w13711);
assign w13712 = v4248;
assign w13713 = w13701 & w13710;
assign w13714 = w13272 & ~w13713;
assign w13715 = w3575 & w4335;
assign w13716 = w1165 & w3268;
assign w13717 = w2835 & w13716;
assign w13718 = w4065 & w13717;
assign w13719 = w2805 & w13718;
assign w13720 = w13715 & w13719;
assign w13721 = ~w353 & w4641;
assign w13722 = w3285 & w13721;
assign w13723 = w5356 & w13722;
assign v4249 = ~(w159 | w640);
assign w13724 = v4249;
assign w13725 = w1390 & w13724;
assign w13726 = w13723 & w13725;
assign w13727 = w13720 & w13726;
assign w13728 = w2521 & w13727;
assign w13729 = w1440 & w2629;
assign w13730 = w13728 & w13729;
assign w13731 = ~w13714 & w13730;
assign v4250 = ~(w13712 | w13731);
assign w13732 = v4250;
assign w13733 = w13656 & w13732;
assign v4251 = ~(w13656 | w13732);
assign w13734 = v4251;
assign v4252 = ~(w13733 | w13734);
assign w13735 = v4252;
assign w13736 = (~w11864 & w11861) | (~w11864 & w28023) | (w11861 & w28023);
assign v4253 = ~(w11865 | w13736);
assign w13737 = v4253;
assign w13738 = w928 & ~w13737;
assign w13739 = w3406 & w11723;
assign w13740 = w3399 & w11729;
assign w13741 = w3402 & w11726;
assign v4254 = ~(w13740 | w13741);
assign w13742 = v4254;
assign w13743 = ~w13739 & w13742;
assign w13744 = ~w13738 & w13743;
assign w13745 = w13735 & ~w13744;
assign v4255 = ~(w13733 | w13745);
assign w13746 = v4255;
assign w13747 = w13654 & ~w13746;
assign w13748 = ~w13654 & w13746;
assign v4256 = ~(w13747 | w13748);
assign w13749 = v4256;
assign w13750 = w3529 & w13178;
assign w13751 = w3760 & w11708;
assign w13752 = w3767 & w11714;
assign w13753 = w3763 & w11711;
assign v4257 = ~(w13752 | w13753);
assign w13754 = v4257;
assign w13755 = ~w13751 & w13754;
assign w13756 = ~w13750 & w13755;
assign w13757 = ~pi29 & w13756;
assign w13758 = pi29 & ~w13756;
assign v4258 = ~(w13757 | w13758);
assign w13759 = v4258;
assign w13760 = w13749 & w13759;
assign v4259 = ~(w13747 | w13760);
assign w13761 = v4259;
assign v4260 = ~(w13524 | w13534);
assign w13762 = v4260;
assign v4261 = ~(w13535 | w13762);
assign w13763 = v4261;
assign w13764 = ~w13761 & w13763;
assign w13765 = w13761 & ~w13763;
assign v4262 = ~(w13764 | w13765);
assign w13766 = v4262;
assign w13767 = w4153 & ~w12842;
assign w13768 = w4155 & w11686;
assign v4263 = ~(w2873 | w11695);
assign w13769 = v4263;
assign w13770 = w4158 & w11689;
assign v4264 = ~(w13769 | w13770);
assign w13771 = v4264;
assign w13772 = ~w13768 & w13771;
assign w13773 = ~w13767 & w13772;
assign w13774 = ~pi26 & w13773;
assign w13775 = pi26 & ~w13773;
assign v4265 = ~(w13774 | w13775);
assign w13776 = v4265;
assign w13777 = w13766 & w13776;
assign v4266 = ~(w13764 | w13777);
assign w13778 = v4266;
assign v4267 = ~(w13641 | w13651);
assign w13779 = v4267;
assign v4268 = ~(w13652 | w13779);
assign w13780 = v4268;
assign w13781 = ~w13778 & w13780;
assign v4269 = ~(w13652 | w13781);
assign w13782 = v4269;
assign w13783 = w13639 & ~w13782;
assign w13784 = ~w13639 & w13782;
assign v4270 = ~(w13783 | w13784);
assign w13785 = v4270;
assign w13786 = w4764 & w11993;
assign w13787 = w4913 & w11984;
assign w13788 = w4836 & w11671;
assign w13789 = w4763 & w11673;
assign v4271 = ~(w13788 | w13789);
assign w13790 = v4271;
assign w13791 = ~w13787 & w13790;
assign w13792 = ~w13786 & w13791;
assign w13793 = ~pi23 & w13792;
assign w13794 = pi23 & ~w13792;
assign v4272 = ~(w13793 | w13794);
assign w13795 = v4272;
assign w13796 = w13785 & w13795;
assign v4273 = ~(w13783 | w13796);
assign w13797 = v4273;
assign w13798 = w13637 & ~w13797;
assign w13799 = ~w13637 & w13797;
assign v4274 = ~(w13798 | w13799);
assign w13800 = v4274;
assign w13801 = w5114 & ~w12277;
assign w13802 = w5531 & w12237;
assign w13803 = w5610 & w12271;
assign v4275 = ~(w13802 | w13803);
assign w13804 = v4275;
assign w13805 = w5113 & w12155;
assign w13806 = w13804 & ~w13805;
assign w13807 = ~w13801 & w13806;
assign w13808 = pi20 & w13807;
assign v4276 = ~(pi20 | w13807);
assign w13809 = v4276;
assign v4277 = ~(w13808 | w13809);
assign w13810 = v4277;
assign w13811 = w13800 & ~w13810;
assign v4278 = ~(w13798 | w13811);
assign w13812 = v4278;
assign w13813 = ~w13624 & w13634;
assign v4279 = ~(w13635 | w13813);
assign w13814 = v4279;
assign w13815 = ~w13812 & w13814;
assign v4280 = ~(w13635 | w13815);
assign w13816 = v4280;
assign w13817 = w13622 & ~w13816;
assign w13818 = ~w13622 & w13816;
assign v4281 = ~(w13817 | w13818);
assign w13819 = v4281;
assign w13820 = pi17 & w12406;
assign w13821 = pi16 & ~w12406;
assign v4282 = ~(w13820 | w13821);
assign w13822 = v4282;
assign w13823 = w5760 & w13822;
assign v4283 = ~(w12580 | w13823);
assign w13824 = v4283;
assign w13825 = w13819 & w13824;
assign v4284 = ~(w13817 | w13825);
assign w13826 = v4284;
assign w13827 = ~w13620 & w13826;
assign v4285 = ~(w13819 | w13824);
assign w13828 = v4285;
assign v4286 = ~(w13825 | w13828);
assign w13829 = v4286;
assign w13830 = ~w13800 & w13810;
assign v4287 = ~(w13811 | w13830);
assign w13831 = v4287;
assign v4288 = ~(w13785 | w13795);
assign w13832 = v4288;
assign v4289 = ~(w13796 | w13832);
assign w13833 = v4289;
assign w13834 = w13778 & ~w13780;
assign v4290 = ~(w13781 | w13834);
assign w13835 = v4290;
assign w13836 = w4764 & w12469;
assign w13837 = w4913 & w11671;
assign w13838 = w4836 & w11673;
assign w13839 = w4763 & w11678;
assign v4291 = ~(w13838 | w13839);
assign w13840 = v4291;
assign w13841 = ~w13837 & w13840;
assign w13842 = ~w13836 & w13841;
assign w13843 = pi23 & ~w13842;
assign w13844 = ~pi23 & w13842;
assign v4292 = ~(w13843 | w13844);
assign w13845 = v4292;
assign w13846 = w13835 & w13845;
assign v4293 = ~(w13766 | w13776);
assign w13847 = v4293;
assign v4294 = ~(w13777 | w13847);
assign w13848 = v4294;
assign w13849 = ~w13735 & w13744;
assign v4295 = ~(w13745 | w13849);
assign w13850 = v4295;
assign w13851 = w3529 & w13194;
assign w13852 = w3763 & w11714;
assign w13853 = w3760 & w11711;
assign v4296 = ~(w13852 | w13853);
assign w13854 = v4296;
assign w13855 = w3767 & w11720;
assign w13856 = w13854 & ~w13855;
assign w13857 = ~w13851 & w13856;
assign v4297 = ~(pi29 | w13857);
assign w13858 = v4297;
assign w13859 = pi29 & w13857;
assign v4298 = ~(w13858 | w13859);
assign w13860 = v4298;
assign w13861 = ~w13850 & w13860;
assign w13862 = (~w11735 & ~w11855) | (~w11735 & w28024) | (~w11855 & w28024);
assign v4299 = ~(w11860 | w13862);
assign w13863 = v4299;
assign v4300 = ~(w11861 | w13863);
assign w13864 = v4300;
assign w13865 = w928 & w13864;
assign w13866 = w3406 & w11726;
assign w13867 = w3402 & w11729;
assign w13868 = w3399 & ~w11734;
assign v4301 = ~(w13867 | w13868);
assign w13869 = v4301;
assign w13870 = ~w13866 & w13869;
assign w13871 = ~w13865 & w13870;
assign v4302 = ~(w13712 | w13714);
assign w13872 = v4302;
assign v4303 = ~(w13730 | w13872);
assign w13873 = v4303;
assign w13874 = w13730 & w13872;
assign v4304 = ~(w13873 | w13874);
assign w13875 = v4304;
assign v4305 = ~(w13871 | w13875);
assign w13876 = v4305;
assign w13877 = w13871 & w13875;
assign v4306 = ~(w13876 | w13877);
assign w13878 = v4306;
assign w13879 = w13697 & ~w13699;
assign v4307 = ~(w13700 | w13879);
assign w13880 = v4307;
assign w13881 = ~w11851 & w28025;
assign v4308 = ~(w11854 | w13881);
assign w13882 = v4308;
assign w13883 = w928 & w13882;
assign w13884 = w3406 & ~w11734;
assign w13885 = w3402 & w11737;
assign w13886 = w3399 & w11740;
assign v4309 = ~(w13885 | w13886);
assign w13887 = v4309;
assign w13888 = ~w13884 & w13887;
assign w13889 = ~w13883 & w13888;
assign w13890 = ~w13880 & w13889;
assign w13891 = w777 & w2072;
assign v4310 = ~(w244 | w566);
assign w13892 = v4310;
assign w13893 = w2350 & w13892;
assign w13894 = w13891 & w13893;
assign w13895 = ~w454 & w2803;
assign w13896 = ~w674 & w708;
assign w13897 = w13895 & w13896;
assign w13898 = w1164 & w4019;
assign w13899 = w13897 & w13898;
assign w13900 = w3322 & w13899;
assign w13901 = w13894 & w13900;
assign w13902 = w4345 & w13901;
assign w13903 = w3824 & w3860;
assign w13904 = w13902 & w13903;
assign w13905 = w13657 & ~w13904;
assign w13906 = ~w13657 & w13904;
assign v4311 = ~(w13905 | w13906);
assign w13907 = v4311;
assign v4312 = ~(w303 | w479);
assign w13908 = v4312;
assign w13909 = ~w173 & w13908;
assign w13910 = w2927 & w4503;
assign w13911 = w13909 & w13910;
assign w13912 = w2292 & w13911;
assign w13913 = ~w369 & w13912;
assign w13914 = ~w999 & w4276;
assign w13915 = w2488 & w13914;
assign w13916 = w13913 & w13915;
assign w13917 = w667 & w2374;
assign w13918 = w3075 & w13917;
assign w13919 = w1406 & w2185;
assign w13920 = w13918 & w13919;
assign w13921 = w5245 & w13920;
assign w13922 = w13916 & w13921;
assign w13923 = w524 & w13922;
assign v4313 = ~(w95 | w211);
assign w13924 = v4313;
assign w13925 = w13149 & w13924;
assign w13926 = w5320 & w13925;
assign w13927 = w13923 & w13926;
assign v4314 = ~(w697 | w870);
assign w13928 = v4314;
assign w13929 = w2453 & w13928;
assign w13930 = ~w125 & w2233;
assign w13931 = w6573 & w13930;
assign w13932 = w13929 & w13931;
assign w13933 = w594 & w2475;
assign w13934 = w13932 & w13933;
assign v4315 = ~(w131 | w162);
assign w13935 = v4315;
assign w13936 = w752 & w3277;
assign w13937 = w13935 & w13936;
assign w13938 = w13934 & w13937;
assign w13939 = w2330 & w2767;
assign w13940 = w13213 & w13939;
assign v4316 = ~(w241 | w541);
assign w13941 = v4316;
assign w13942 = w13940 & w13941;
assign w13943 = w1730 & w13942;
assign w13944 = w13938 & w13943;
assign w13945 = w12444 & w13944;
assign w13946 = w13927 & w13945;
assign w13947 = ~w11842 & w28026;
assign v4317 = ~(w11845 | w13947);
assign w13948 = v4317;
assign w13949 = w928 & w13948;
assign w13950 = w3406 & ~w11745;
assign w13951 = w3402 & w11748;
assign w13952 = w3399 & w11759;
assign v4318 = ~(w13951 | w13952);
assign w13953 = v4318;
assign w13954 = ~w13950 & w13953;
assign w13955 = ~w13949 & w13954;
assign w13956 = w13946 & w13955;
assign w13957 = w13657 & ~w13956;
assign v4319 = ~(w13946 | w13955);
assign w13958 = v4319;
assign v4320 = ~(w13657 | w13958);
assign w13959 = v4320;
assign v4321 = ~(w13957 | w13959);
assign w13960 = v4321;
assign w13961 = w478 & w6585;
assign w13962 = w1476 & w13961;
assign w13963 = w4456 & w12195;
assign w13964 = w2545 & w13963;
assign w13965 = w646 & w13964;
assign w13966 = w13962 & w13965;
assign w13967 = ~w272 & w2452;
assign w13968 = w2635 & w13967;
assign w13969 = w1239 & w2661;
assign w13970 = ~w680 & w2186;
assign w13971 = ~w141 & w13970;
assign w13972 = w13969 & w13971;
assign w13973 = w13968 & w13972;
assign w13974 = w1524 & w1714;
assign w13975 = w13973 & w13974;
assign w13976 = w13966 & w13975;
assign w13977 = w13681 & w13976;
assign w13978 = w13960 & ~w13977;
assign v4322 = ~(w13957 | w13978);
assign w13979 = v4322;
assign w13980 = w13907 & ~w13979;
assign v4323 = ~(w13905 | w13980);
assign w13981 = v4323;
assign w13982 = w13880 & ~w13889;
assign v4324 = ~(w13890 | w13982);
assign w13983 = v4324;
assign w13984 = w13981 & w13983;
assign v4325 = ~(w13890 | w13984);
assign w13985 = v4325;
assign v4326 = ~(w13711 | w13713);
assign w13986 = v4326;
assign v4327 = ~(w13272 | w13986);
assign w13987 = v4327;
assign w13988 = ~w13711 & w13714;
assign v4328 = ~(w13987 | w13988);
assign w13989 = v4328;
assign v4329 = ~(w13985 | w13989);
assign w13990 = v4329;
assign w13991 = w13985 & w13989;
assign v4330 = ~(w13990 | w13991);
assign w13992 = v4330;
assign w13993 = w3529 & ~w13310;
assign w13994 = w3760 & w11720;
assign w13995 = w3763 & w11723;
assign w13996 = w3767 & w11726;
assign v4331 = ~(w13995 | w13996);
assign w13997 = v4331;
assign w13998 = ~w13994 & w13997;
assign w13999 = ~w13993 & w13998;
assign w14000 = ~pi29 & w13999;
assign w14001 = pi29 & ~w13999;
assign v4332 = ~(w14000 | w14001);
assign w14002 = v4332;
assign w14003 = w13992 & ~w14002;
assign v4333 = ~(w13990 | w14003);
assign w14004 = v4333;
assign w14005 = w13878 & w14004;
assign v4334 = ~(w13876 | w14005);
assign w14006 = v4334;
assign w14007 = w13850 & ~w13860;
assign v4335 = ~(w13861 | w14007);
assign w14008 = v4335;
assign w14009 = w14006 & w14008;
assign v4336 = ~(w13861 | w14009);
assign w14010 = v4336;
assign v4337 = ~(w13749 | w13759);
assign w14011 = v4337;
assign v4338 = ~(w13760 | w14011);
assign w14012 = v4338;
assign w14013 = w14010 & w14012;
assign v4339 = ~(w14010 | w14012);
assign w14014 = v4339;
assign v4340 = ~(w14013 | w14014);
assign w14015 = v4340;
assign w14016 = w4153 & w12694;
assign w14017 = w4155 & w11689;
assign w14018 = ~w2873 & w11700;
assign w14019 = w4158 & ~w11695;
assign v4341 = ~(w14018 | w14019);
assign w14020 = v4341;
assign w14021 = ~w14017 & w14020;
assign w14022 = ~w14016 & w14021;
assign w14023 = ~pi26 & w14022;
assign w14024 = pi26 & ~w14022;
assign v4342 = ~(w14023 | w14024);
assign w14025 = v4342;
assign w14026 = w14015 & w14025;
assign v4343 = ~(w14013 | w14026);
assign w14027 = v4343;
assign w14028 = w13848 & ~w14027;
assign w14029 = ~w13848 & w14027;
assign v4344 = ~(w14028 | w14029);
assign w14030 = v4344;
assign w14031 = w4764 & w12454;
assign w14032 = w4836 & w11678;
assign w14033 = w4913 & w11673;
assign v4345 = ~(w14032 | w14033);
assign w14034 = v4345;
assign w14035 = w4763 & ~w11683;
assign w14036 = w14034 & ~w14035;
assign w14037 = ~w14031 & w14036;
assign w14038 = pi23 & w14037;
assign v4346 = ~(pi23 | w14037);
assign w14039 = v4346;
assign v4347 = ~(w14038 | w14039);
assign w14040 = v4347;
assign w14041 = w14030 & ~w14040;
assign v4348 = ~(w14028 | w14041);
assign w14042 = v4348;
assign v4349 = ~(w13835 | w13845);
assign w14043 = v4349;
assign v4350 = ~(w13846 | w14043);
assign w14044 = v4350;
assign w14045 = ~w14042 & w14044;
assign v4351 = ~(w13846 | w14045);
assign w14046 = v4351;
assign w14047 = w13833 & ~w14046;
assign w14048 = ~w13833 & w14046;
assign v4352 = ~(w14047 | w14048);
assign w14049 = v4352;
assign w14050 = w5114 & ~w12351;
assign w14051 = w5610 & w12237;
assign w14052 = w5531 & w12155;
assign w14053 = w5113 & w12084;
assign v4353 = ~(w14052 | w14053);
assign w14054 = v4353;
assign w14055 = ~w14051 & w14054;
assign w14056 = ~w14050 & w14055;
assign w14057 = ~pi20 & w14056;
assign w14058 = pi20 & ~w14056;
assign v4354 = ~(w14057 | w14058);
assign w14059 = v4354;
assign w14060 = w14049 & w14059;
assign v4355 = ~(w14047 | w14060);
assign w14061 = v4355;
assign w14062 = w13831 & ~w14061;
assign w14063 = ~w13831 & w14061;
assign v4356 = ~(w14062 | w14063);
assign w14064 = v4356;
assign w14065 = w5765 & ~w12506;
assign w14066 = w6236 & ~w12406;
assign w14067 = w5764 & w12311;
assign w14068 = w5983 & w12381;
assign v4357 = ~(w14067 | w14068);
assign w14069 = v4357;
assign w14070 = ~w14066 & w14069;
assign w14071 = ~w14065 & w14070;
assign w14072 = ~pi17 & w14071;
assign w14073 = pi17 & ~w14071;
assign v4358 = ~(w14072 | w14073);
assign w14074 = v4358;
assign w14075 = w14064 & w14074;
assign v4359 = ~(w14062 | w14075);
assign w14076 = v4359;
assign w14077 = w5764 & w12381;
assign w14078 = w5765 & w12505;
assign v4360 = ~(w5983 | w14078);
assign w14079 = v4360;
assign v4361 = ~(w12406 | w14079);
assign w14080 = v4361;
assign v4362 = ~(w6236 | w14080);
assign w14081 = v4362;
assign w14082 = ~w14077 & w14081;
assign w14083 = ~pi17 & w14082;
assign w14084 = pi17 & ~w14082;
assign v4363 = ~(w14083 | w14084);
assign w14085 = v4363;
assign w14086 = ~w14076 & w14085;
assign w14087 = w13812 & ~w13814;
assign v4364 = ~(w13815 | w14087);
assign w14088 = v4364;
assign w14089 = w14076 & ~w14085;
assign v4365 = ~(w14086 | w14089);
assign w14090 = v4365;
assign w14091 = w14088 & w14090;
assign v4366 = ~(w14086 | w14091);
assign w14092 = v4366;
assign w14093 = w13829 & ~w14092;
assign w14094 = ~w13829 & w14092;
assign v4367 = ~(w14093 | w14094);
assign w14095 = v4367;
assign v4368 = ~(w14049 | w14059);
assign w14096 = v4368;
assign v4369 = ~(w14060 | w14096);
assign w14097 = v4369;
assign w14098 = w14042 & ~w14044;
assign v4370 = ~(w14045 | w14098);
assign w14099 = v4370;
assign w14100 = w5114 & w12167;
assign w14101 = w5610 & w12155;
assign w14102 = w5113 & w11984;
assign w14103 = w5531 & w12084;
assign v4371 = ~(w14102 | w14103);
assign w14104 = v4371;
assign w14105 = ~w14101 & w14104;
assign w14106 = ~w14100 & w14105;
assign w14107 = ~pi20 & w14106;
assign w14108 = pi20 & ~w14106;
assign v4372 = ~(w14107 | w14108);
assign w14109 = v4372;
assign w14110 = w14099 & w14109;
assign w14111 = ~w14030 & w14040;
assign v4373 = ~(w14041 | w14111);
assign w14112 = v4373;
assign v4374 = ~(w14015 | w14025);
assign w14113 = v4374;
assign v4375 = ~(w14026 | w14113);
assign w14114 = v4375;
assign v4376 = ~(w14006 | w14008);
assign w14115 = v4376;
assign v4377 = ~(w14009 | w14115);
assign w14116 = v4377;
assign w14117 = w4153 & ~w13008;
assign w14118 = w4155 & ~w11695;
assign w14119 = ~w2873 & w11708;
assign w14120 = w4158 & w11700;
assign v4378 = ~(w14119 | w14120);
assign w14121 = v4378;
assign w14122 = ~w14118 & w14121;
assign w14123 = ~w14117 & w14122;
assign w14124 = ~pi26 & w14123;
assign w14125 = pi26 & ~w14123;
assign v4379 = ~(w14124 | w14125);
assign w14126 = v4379;
assign w14127 = ~w14116 & w14126;
assign w14128 = w3529 & w13514;
assign w14129 = w3763 & w11720;
assign w14130 = w3760 & w11714;
assign v4380 = ~(w14129 | w14130);
assign w14131 = v4380;
assign w14132 = w3767 & w11723;
assign w14133 = w14131 & ~w14132;
assign w14134 = ~w14128 & w14133;
assign w14135 = pi29 & w14134;
assign v4381 = ~(pi29 | w14134);
assign w14136 = v4381;
assign v4382 = ~(w14135 | w14136);
assign w14137 = v4382;
assign w14138 = w4153 & w12994;
assign w14139 = w4155 & w11700;
assign w14140 = ~w2873 & w11711;
assign w14141 = w4158 & w11708;
assign v4383 = ~(w14140 | w14141);
assign w14142 = v4383;
assign w14143 = ~w14139 & w14142;
assign w14144 = ~w14138 & w14143;
assign w14145 = ~pi26 & w14144;
assign w14146 = pi26 & ~w14144;
assign v4384 = ~(w14145 | w14146);
assign w14147 = v4384;
assign w14148 = ~w14137 & w14147;
assign v4385 = ~(w13878 | w14004);
assign w14149 = v4385;
assign v4386 = ~(w14005 | w14149);
assign w14150 = v4386;
assign w14151 = w14137 & ~w14147;
assign v4387 = ~(w14148 | w14151);
assign w14152 = v4387;
assign w14153 = w14150 & w14152;
assign v4388 = ~(w14148 | w14153);
assign w14154 = v4388;
assign w14155 = w14116 & ~w14126;
assign v4389 = ~(w14127 | w14155);
assign w14156 = v4389;
assign w14157 = ~w14154 & w14156;
assign v4390 = ~(w14127 | w14157);
assign w14158 = v4390;
assign w14159 = w14114 & ~w14158;
assign w14160 = ~w14114 & w14158;
assign v4391 = ~(w14159 | w14160);
assign w14161 = v4391;
assign w14162 = w4764 & w12594;
assign w14163 = w4836 & ~w11683;
assign w14164 = w4913 & w11678;
assign v4392 = ~(w14163 | w14164);
assign w14165 = v4392;
assign w14166 = w4763 & w11686;
assign w14167 = w14165 & ~w14166;
assign w14168 = ~w14162 & w14167;
assign w14169 = pi23 & w14168;
assign v4393 = ~(pi23 | w14168);
assign w14170 = v4393;
assign v4394 = ~(w14169 | w14170);
assign w14171 = v4394;
assign w14172 = w14161 & ~w14171;
assign v4395 = ~(w14159 | w14172);
assign w14173 = v4395;
assign w14174 = w14112 & ~w14173;
assign w14175 = ~w14112 & w14173;
assign v4396 = ~(w14174 | w14175);
assign w14176 = v4396;
assign w14177 = w5114 & w12181;
assign w14178 = w5531 & w11984;
assign w14179 = w5610 & w12084;
assign v4397 = ~(w14178 | w14179);
assign w14180 = v4397;
assign w14181 = w5113 & w11671;
assign w14182 = w14180 & ~w14181;
assign w14183 = ~w14177 & w14182;
assign w14184 = pi20 & w14183;
assign v4398 = ~(pi20 | w14183);
assign w14185 = v4398;
assign v4399 = ~(w14184 | w14185);
assign w14186 = v4399;
assign w14187 = w14176 & ~w14186;
assign v4400 = ~(w14174 | w14187);
assign w14188 = v4400;
assign v4401 = ~(w14099 | w14109);
assign w14189 = v4401;
assign v4402 = ~(w14110 | w14189);
assign w14190 = v4402;
assign w14191 = ~w14188 & w14190;
assign v4403 = ~(w14110 | w14191);
assign w14192 = v4403;
assign w14193 = w14097 & ~w14192;
assign w14194 = ~w14097 & w14192;
assign v4404 = ~(w14193 | w14194);
assign w14195 = v4404;
assign w14196 = w5765 & w12387;
assign w14197 = w6236 & w12381;
assign w14198 = w5764 & w12271;
assign w14199 = w5983 & w12311;
assign v4405 = ~(w14198 | w14199);
assign w14200 = v4405;
assign w14201 = ~w14197 & w14200;
assign w14202 = ~w14196 & w14201;
assign w14203 = ~pi17 & w14202;
assign w14204 = pi17 & ~w14202;
assign v4406 = ~(w14203 | w14204);
assign w14205 = v4406;
assign w14206 = w14195 & w14205;
assign v4407 = ~(w14193 | w14206);
assign w14207 = v4407;
assign w14208 = w12685 & ~w14207;
assign v4408 = ~(w14064 | w14074);
assign w14209 = v4408;
assign v4409 = ~(w14075 | w14209);
assign w14210 = v4409;
assign w14211 = ~w12685 & w14207;
assign v4410 = ~(w14208 | w14211);
assign w14212 = v4410;
assign w14213 = w14210 & w14212;
assign v4411 = ~(w14208 | w14213);
assign w14214 = v4411;
assign v4412 = ~(w14088 | w14090);
assign w14215 = v4412;
assign v4413 = ~(w14091 | w14215);
assign w14216 = v4413;
assign w14217 = ~w14214 & w14216;
assign w14218 = w14214 & ~w14216;
assign v4414 = ~(w14217 | w14218);
assign w14219 = v4414;
assign v4415 = ~(w14210 | w14212);
assign w14220 = v4415;
assign v4416 = ~(w14213 | w14220);
assign w14221 = v4416;
assign v4417 = ~(w14195 | w14205);
assign w14222 = v4417;
assign v4418 = ~(w14206 | w14222);
assign w14223 = v4418;
assign w14224 = w14188 & ~w14190;
assign v4419 = ~(w14191 | w14224);
assign w14225 = v4419;
assign w14226 = w5765 & w12318;
assign w14227 = w5983 & w12271;
assign w14228 = w6236 & w12311;
assign v4420 = ~(w14227 | w14228);
assign w14229 = v4420;
assign w14230 = w5764 & w12237;
assign w14231 = w14229 & ~w14230;
assign w14232 = ~w14226 & w14231;
assign w14233 = pi17 & w14232;
assign v4421 = ~(pi17 | w14232);
assign w14234 = v4421;
assign v4422 = ~(w14233 | w14234);
assign w14235 = v4422;
assign w14236 = w14225 & ~w14235;
assign w14237 = ~w14176 & w14186;
assign v4423 = ~(w14187 | w14237);
assign w14238 = v4423;
assign w14239 = ~w14161 & w14171;
assign v4424 = ~(w14172 | w14239);
assign w14240 = v4424;
assign w14241 = w14154 & ~w14156;
assign v4425 = ~(w14157 | w14241);
assign w14242 = v4425;
assign w14243 = w4764 & w12610;
assign w14244 = w4913 & ~w11683;
assign w14245 = w4836 & w11686;
assign w14246 = w4763 & w11689;
assign v4426 = ~(w14245 | w14246);
assign w14247 = v4426;
assign w14248 = ~w14244 & w14247;
assign w14249 = ~w14243 & w14248;
assign w14250 = ~pi23 & w14249;
assign w14251 = pi23 & ~w14249;
assign v4427 = ~(w14250 | w14251);
assign w14252 = v4427;
assign w14253 = w14242 & w14252;
assign v4428 = ~(w14242 | w14252);
assign w14254 = v4428;
assign v4429 = ~(w14253 | w14254);
assign w14255 = v4429;
assign w14256 = ~w13992 & w14002;
assign v4430 = ~(w14003 | w14256);
assign w14257 = v4430;
assign w14258 = w4153 & w13178;
assign w14259 = w4155 & w11708;
assign w14260 = ~w2873 & w11714;
assign w14261 = w4158 & w11711;
assign v4431 = ~(w14260 | w14261);
assign w14262 = v4431;
assign w14263 = ~w14259 & w14262;
assign w14264 = ~w14258 & w14263;
assign w14265 = ~pi26 & w14264;
assign w14266 = pi26 & ~w14264;
assign v4432 = ~(w14265 | w14266);
assign w14267 = v4432;
assign w14268 = w14257 & ~w14267;
assign v4433 = ~(w13981 | w13983);
assign w14269 = v4433;
assign v4434 = ~(w13984 | w14269);
assign w14270 = v4434;
assign w14271 = w3529 & ~w13737;
assign w14272 = w3760 & w11723;
assign w14273 = w3767 & w11729;
assign w14274 = w3763 & w11726;
assign v4435 = ~(w14273 | w14274);
assign w14275 = v4435;
assign w14276 = ~w14272 & w14275;
assign w14277 = ~w14271 & w14276;
assign w14278 = pi29 & ~w14277;
assign w14279 = ~pi29 & w14277;
assign v4436 = ~(w14278 | w14279);
assign w14280 = v4436;
assign w14281 = w14270 & ~w14280;
assign w14282 = ~w13907 & w13979;
assign v4437 = ~(w13980 | w14282);
assign w14283 = v4437;
assign v4438 = ~(w11746 | w11847);
assign w14284 = v4438;
assign w14285 = (w14284 & w11845) | (w14284 & w28027) | (w11845 & w28027);
assign w14286 = (~w11845 & w30169) | (~w11845 & w30170) | (w30169 & w30170);
assign w14287 = ~w11847 & w14286;
assign v4439 = ~(w11851 | w14287);
assign w14288 = v4439;
assign w14289 = w928 & w14288;
assign w14290 = w3406 & w11737;
assign w14291 = w3399 & ~w11745;
assign w14292 = w3402 & w11740;
assign v4440 = ~(w14291 | w14292);
assign w14293 = v4440;
assign w14294 = ~w14290 & w14293;
assign w14295 = ~w14289 & w14294;
assign w14296 = w14283 & ~w14295;
assign w14297 = ~w13960 & w13977;
assign v4441 = ~(w13978 | w14297);
assign w14298 = v4441;
assign w14299 = ~w11845 & w28028;
assign v4442 = ~(w14285 | w14299);
assign w14300 = v4442;
assign w14301 = w928 & w14300;
assign w14302 = w3406 & w11740;
assign w14303 = w3402 & ~w11745;
assign w14304 = w3399 & w11748;
assign v4443 = ~(w14303 | w14304);
assign w14305 = v4443;
assign w14306 = ~w14302 & w14305;
assign w14307 = ~w14301 & w14306;
assign w14308 = w14298 & ~w14307;
assign w14309 = ~w14298 & w14307;
assign v4444 = ~(w14308 | w14309);
assign w14310 = v4444;
assign w14311 = ~w640 & w1293;
assign w14312 = ~w245 & w11617;
assign v4445 = ~(w253 | w499);
assign w14313 = v4445;
assign w14314 = w878 & w14313;
assign w14315 = w14312 & w14314;
assign w14316 = w14311 & w14315;
assign v4446 = ~(w259 | w711);
assign w14317 = v4446;
assign w14318 = w13117 & w14317;
assign v4447 = ~(w162 | w463);
assign w14319 = v4447;
assign w14320 = w14318 & w14319;
assign w14321 = w14316 & w14320;
assign w14322 = w5011 & w14321;
assign w14323 = w971 & w2922;
assign w14324 = w1163 & w3325;
assign w14325 = w4368 & w14324;
assign w14326 = w3267 & w14325;
assign w14327 = w14323 & w14326;
assign w14328 = w1672 & w14327;
assign w14329 = w14322 & w14328;
assign w14330 = ~w11836 & w29282;
assign v4448 = ~(w11841 | w14330);
assign w14331 = v4448;
assign w14332 = w928 & ~w14331;
assign w14333 = w3406 & w11748;
assign w14334 = w3402 & w11759;
assign w14335 = w3399 & w11761;
assign v4449 = ~(w14334 | w14335);
assign w14336 = v4449;
assign w14337 = ~w14333 & w14336;
assign w14338 = ~w14332 & w14337;
assign v4450 = ~(w14329 | w14338);
assign w14339 = v4450;
assign w14340 = w1170 & w6052;
assign w14341 = ~w656 & w14340;
assign w14342 = w406 & w767;
assign w14343 = ~w288 & w4485;
assign w14344 = w712 & w14343;
assign w14345 = w14342 & w14344;
assign w14346 = ~w252 & w14345;
assign w14347 = w14341 & w14346;
assign w14348 = w1927 & w14347;
assign w14349 = w4046 & w6657;
assign w14350 = w3047 & w14349;
assign w14351 = w4037 & w14350;
assign w14352 = w12037 & w14351;
assign w14353 = w1568 & w14352;
assign w14354 = w14348 & w14353;
assign w14355 = w11836 & ~w11838;
assign v4451 = ~(w11839 | w14355);
assign w14356 = v4451;
assign w14357 = w928 & w14356;
assign w14358 = w3399 & ~w11771;
assign v4452 = ~(w14357 | w14358);
assign w14359 = v4452;
assign w14360 = w3406 & w11759;
assign w14361 = w3402 & w11761;
assign v4453 = ~(w14360 | w14361);
assign w14362 = v4453;
assign w14363 = w14359 & w14362;
assign v4454 = ~(w14354 | w14363);
assign w14364 = v4454;
assign w14365 = w2451 & w3946;
assign v4455 = ~(w145 | w886);
assign w14366 = v4455;
assign w14367 = w808 & w14366;
assign w14368 = ~w88 & w14367;
assign w14369 = w3139 & w14368;
assign v4456 = ~(w107 | w548);
assign w14370 = v4456;
assign w14371 = w2401 & w14370;
assign w14372 = w1934 & w14371;
assign w14373 = w665 & w738;
assign w14374 = w1814 & w14373;
assign w14375 = w14372 & w14374;
assign w14376 = w14369 & w14375;
assign w14377 = w14365 & w14376;
assign w14378 = w13927 & w14377;
assign v4457 = ~(w11772 | w11773);
assign w14379 = v4457;
assign w14380 = (~w29494 & w30032) | (~w29494 & w30033) | (w30032 & w30033);
assign w14381 = w14379 & w14380;
assign v4458 = ~(w14379 | w14380);
assign w14382 = v4458;
assign v4459 = ~(w14381 | w14382);
assign w14383 = v4459;
assign w14384 = w928 & ~w14383;
assign w14385 = w3402 & ~w11771;
assign w14386 = w3406 & w11761;
assign w14387 = w3399 & w11768;
assign v4460 = ~(w14386 | w14387);
assign w14388 = v4460;
assign w14389 = ~w14385 & w14388;
assign w14390 = ~w14384 & w14389;
assign v4461 = ~(w14378 | w14390);
assign w14391 = v4461;
assign v4462 = ~(w379 | w727);
assign w14392 = v4462;
assign v4463 = ~(w488 | w652);
assign w14393 = v4463;
assign w14394 = w14392 & w14393;
assign w14395 = w339 & w1239;
assign w14396 = w14394 & w14395;
assign w14397 = w2657 & w14396;
assign w14398 = w808 & w2719;
assign w14399 = w6539 & w14398;
assign w14400 = w14397 & w14399;
assign w14401 = w1199 & w14400;
assign w14402 = w4619 & w6707;
assign w14403 = w2117 & w14402;
assign w14404 = w3032 & w14403;
assign w14405 = w14401 & w14404;
assign w14406 = w3704 & w14405;
assign w14407 = w4252 & w14406;
assign w14408 = (~w28011 & w29496) | (~w28011 & w29497) | (w29496 & w29497);
assign v4464 = ~(w11834 | w14408);
assign w14409 = v4464;
assign w14410 = w928 & w14409;
assign w14411 = w3402 & w11768;
assign v4465 = ~(w14410 | w14411);
assign w14412 = v4465;
assign w14413 = w3406 & ~w11771;
assign w14414 = w3399 & w11776;
assign v4466 = ~(w14413 | w14414);
assign w14415 = v4466;
assign w14416 = w14412 & w14415;
assign v4467 = ~(w14407 | w14416);
assign w14417 = v4467;
assign v4468 = ~(w31 | w309);
assign w14418 = v4468;
assign w14419 = w740 & w14418;
assign w14420 = w12663 & w14419;
assign w14421 = w938 & w14420;
assign w14422 = w12984 & w14421;
assign w14423 = ~w127 & w1173;
assign v4469 = ~(w292 | w692);
assign w14424 = v4469;
assign w14425 = ~w558 & w14424;
assign w14426 = ~w259 & w14425;
assign w14427 = w14423 & w14426;
assign w14428 = w6566 & w14427;
assign w14429 = w1848 & w3724;
assign w14430 = w6115 & w14429;
assign w14431 = w1870 & w2246;
assign w14432 = w12973 & w14431;
assign w14433 = w14430 & w14432;
assign w14434 = w14428 & w14433;
assign w14435 = ~w899 & w2128;
assign w14436 = w3251 & w14435;
assign w14437 = w4366 & w6534;
assign w14438 = w13969 & w14437;
assign w14439 = w675 & w3298;
assign w14440 = w14438 & w14439;
assign w14441 = w6486 & w14440;
assign w14442 = w14436 & w14441;
assign w14443 = w419 & ~w731;
assign w14444 = w2927 & w14443;
assign w14445 = ~w202 & w3659;
assign w14446 = w14444 & w14445;
assign w14447 = w6707 & w13254;
assign w14448 = w5366 & w12654;
assign w14449 = w14447 & w14448;
assign w14450 = w14446 & w14449;
assign w14451 = w3941 & w3963;
assign w14452 = w3950 & w14451;
assign w14453 = w14450 & w14452;
assign w14454 = w14442 & w14453;
assign w14455 = w14434 & w14454;
assign w14456 = w14422 & w14455;
assign w14457 = ~w11777 & w11790;
assign w14458 = (~w11788 & ~w11824) | (~w11788 & w28029) | (~w11824 & w28029);
assign w14459 = ~w14457 & w14458;
assign w14460 = w14457 & ~w14458;
assign v4470 = ~(w14459 | w14460);
assign w14461 = v4470;
assign w14462 = w928 & w14461;
assign w14463 = w3406 & w11768;
assign w14464 = w3399 & w11784;
assign w14465 = w3402 & w11776;
assign v4471 = ~(w14464 | w14465);
assign w14466 = v4471;
assign w14467 = ~w14463 & w14466;
assign w14468 = ~w14462 & w14467;
assign v4472 = ~(w14456 | w14468);
assign w14469 = v4472;
assign w14470 = ~w331 & w1398;
assign w14471 = w11914 & w14470;
assign w14472 = w12297 & w14471;
assign w14473 = w1157 & w11614;
assign w14474 = w2621 & w14473;
assign w14475 = w14472 & w14474;
assign w14476 = w13280 & w14475;
assign w14477 = w1026 & w2076;
assign w14478 = ~w749 & w14477;
assign w14479 = w1263 & w14478;
assign w14480 = w585 & w14479;
assign w14481 = w2146 & w14480;
assign w14482 = w14476 & w14481;
assign v4473 = ~(w624 | w1108);
assign w14483 = v4473;
assign w14484 = w1179 & w14483;
assign w14485 = w4474 & w14484;
assign w14486 = w1292 & w2525;
assign w14487 = w14485 & w14486;
assign w14488 = ~w680 & w2147;
assign w14489 = ~w639 & w2681;
assign w14490 = w14488 & w14489;
assign w14491 = w1905 & w2188;
assign w14492 = w1087 & w1864;
assign w14493 = w14491 & w14492;
assign w14494 = w14490 & w14493;
assign w14495 = w289 & w3952;
assign w14496 = w217 & w14495;
assign v4474 = ~(w264 | w505);
assign w14497 = v4474;
assign w14498 = w14496 & w14497;
assign w14499 = w14494 & w14498;
assign w14500 = w14487 & w14499;
assign w14501 = w11596 & w14500;
assign w14502 = w14482 & w14501;
assign v4475 = ~(w11819 | w11824);
assign w14503 = v4475;
assign v4476 = ~(w11825 | w14503);
assign w14504 = v4476;
assign w14505 = w3399 & w11793;
assign w14506 = (~w14505 & ~w14504) | (~w14505 & w31270) | (~w14504 & w31270);
assign w14507 = w3406 & w11776;
assign w14508 = w3402 & w11784;
assign v4477 = ~(w14507 | w14508);
assign w14509 = v4477;
assign w14510 = w14506 & w14509;
assign v4478 = ~(w14502 | w14510);
assign w14511 = v4478;
assign w14512 = w801 & w1584;
assign w14513 = ~w299 & w2901;
assign w14514 = w2239 & w14513;
assign w14515 = w2950 & w14514;
assign v4479 = ~(w563 | w605);
assign w14516 = v4479;
assign w14517 = ~w88 & w649;
assign w14518 = w14516 & w14517;
assign w14519 = ~w465 & w2134;
assign w14520 = w1001 & w14519;
assign w14521 = w14518 & w14520;
assign w14522 = w434 & w14521;
assign w14523 = w14515 & w14522;
assign w14524 = w14512 & w14523;
assign w14525 = w476 & w3684;
assign v4480 = ~(w326 | w739);
assign w14526 = v4480;
assign w14527 = ~w420 & w14526;
assign w14528 = w14525 & w14527;
assign v4481 = ~(w300 | w564);
assign w14529 = v4481;
assign w14530 = w965 & w14529;
assign w14531 = ~w53 & w14530;
assign w14532 = w14528 & w14531;
assign w14533 = w1337 & w3438;
assign w14534 = ~w758 & w14533;
assign w14535 = w12673 & w14534;
assign w14536 = ~w200 & w14535;
assign w14537 = w14532 & w14536;
assign w14538 = w1690 & w12556;
assign w14539 = ~w550 & w14538;
assign w14540 = w290 & w13231;
assign w14541 = w14539 & w14540;
assign w14542 = w14537 & w14541;
assign w14543 = w2337 & w14542;
assign w14544 = w14524 & w14543;
assign w14545 = w11813 & w11817;
assign v4482 = ~(w11813 | w11817);
assign w14546 = v4482;
assign v4483 = ~(w14545 | w14546);
assign w14547 = v4483;
assign w14548 = w3402 & w11793;
assign w14549 = (~w14548 & ~w14547) | (~w14548 & w31271) | (~w14547 & w31271);
assign w14550 = w3406 & w11784;
assign w14551 = w3399 & w11803;
assign v4484 = ~(w14550 | w14551);
assign w14552 = v4484;
assign w14553 = w14549 & w14552;
assign v4485 = ~(w14544 | w14553);
assign w14554 = v4485;
assign w14555 = w3986 & w6523;
assign w14556 = w3202 & w14555;
assign w14557 = w12024 & w14556;
assign w14558 = w1260 & w1364;
assign w14559 = w5426 & w14558;
assign w14560 = w12096 & w14559;
assign w14561 = ~w131 & w2749;
assign w14562 = w3422 & w14561;
assign w14563 = w725 & w14562;
assign w14564 = ~w317 & w14563;
assign w14565 = w14560 & w14564;
assign w14566 = w1248 & w14565;
assign w14567 = w14557 & w14566;
assign v4486 = ~(w11805 | w11810);
assign w14568 = v4486;
assign v4487 = ~(w11811 | w14568);
assign w14569 = v4487;
assign w14570 = w3399 & w11798;
assign w14571 = (~w14570 & ~w14569) | (~w14570 & w31272) | (~w14569 & w31272);
assign w14572 = w3406 & w11793;
assign w14573 = w3402 & w11803;
assign v4488 = ~(w14572 | w14573);
assign w14574 = v4488;
assign w14575 = w14571 & w14574;
assign v4489 = ~(w14567 | w14575);
assign w14576 = v4489;
assign w14577 = w14567 & w14575;
assign v4490 = ~(w14576 | w14577);
assign w14578 = v4490;
assign w14579 = w2781 & w2837;
assign w14580 = w3880 & w14579;
assign w14581 = w6618 & w14580;
assign w14582 = w2746 & w14581;
assign w14583 = w332 & w1066;
assign w14584 = w1869 & w2348;
assign w14585 = ~w550 & w14584;
assign w14586 = w14583 & w14585;
assign w14587 = w2967 & w14586;
assign w14588 = w14582 & w14587;
assign w14589 = w4100 & w14396;
assign w14590 = w109 & w2704;
assign w14591 = w14589 & w14590;
assign v4491 = ~(w27 | w447);
assign w14592 = v4491;
assign w14593 = w265 & w14592;
assign v4492 = ~(w134 | w466);
assign w14594 = v4492;
assign w14595 = w1073 & w14594;
assign w14596 = w2028 & w14595;
assign w14597 = w14593 & w14596;
assign w14598 = w726 & w14597;
assign w14599 = w14591 & w14598;
assign v4493 = ~(w112 | w457);
assign w14600 = v4493;
assign w14601 = ~w541 & w14600;
assign w14602 = w966 & w14601;
assign w14603 = w11938 & w14602;
assign w14604 = w6059 & w14603;
assign w14605 = w14599 & w14604;
assign w14606 = w3066 & w14605;
assign w14607 = w14588 & w14606;
assign w14608 = ~w11798 & w11800;
assign v4494 = ~(w11801 | w14608);
assign w14609 = v4494;
assign w14610 = w928 & ~w14609;
assign w14611 = w3406 & w11798;
assign w14612 = w3402 & w11800;
assign v4495 = ~(w14611 | w14612);
assign w14613 = v4495;
assign w14614 = ~w14610 & w14613;
assign v4496 = ~(w14607 | w14614);
assign w14615 = v4496;
assign v4497 = ~(w172 | w186);
assign w14616 = v4497;
assign v4498 = ~(w247 | w317);
assign w14617 = v4498;
assign w14618 = w11930 & w14617;
assign w14619 = w14616 & w14618;
assign w14620 = ~w253 & w375;
assign w14621 = w606 & w14620;
assign w14622 = w14619 & w14621;
assign w14623 = ~w168 & w1106;
assign v4499 = ~(w74 | w673);
assign w14624 = v4499;
assign w14625 = w14623 & w14624;
assign w14626 = w1654 & w2681;
assign w14627 = w1315 & w14626;
assign w14628 = w14625 & w14627;
assign w14629 = ~w566 & w5245;
assign w14630 = w14628 & w14629;
assign w14631 = w14622 & w14630;
assign w14632 = w351 & w13932;
assign w14633 = w14631 & w14632;
assign w14634 = w13222 & w14633;
assign w14635 = w14615 & ~w14634;
assign w14636 = ~w14615 & w14634;
assign v4500 = ~(w14635 | w14636);
assign w14637 = v4500;
assign w14638 = ~w11801 & w11803;
assign v4501 = ~(w11804 | w14638);
assign w14639 = v4501;
assign w14640 = w928 & ~w14639;
assign w14641 = w3399 & w11800;
assign v4502 = ~(w14640 | w14641);
assign w14642 = v4502;
assign w14643 = w3406 & w11803;
assign w14644 = w3402 & w11798;
assign v4503 = ~(w14643 | w14644);
assign w14645 = v4503;
assign w14646 = w14642 & w14645;
assign w14647 = w14637 & ~w14646;
assign v4504 = ~(w14635 | w14647);
assign w14648 = v4504;
assign w14649 = w14578 & ~w14648;
assign v4505 = ~(w14576 | w14649);
assign w14650 = v4505;
assign w14651 = w14544 & w14553;
assign v4506 = ~(w14554 | w14651);
assign w14652 = v4506;
assign w14653 = ~w14650 & w14652;
assign v4507 = ~(w14554 | w14653);
assign w14654 = v4507;
assign w14655 = w14502 & w14510;
assign v4508 = ~(w14511 | w14655);
assign w14656 = v4508;
assign w14657 = ~w14654 & w14656;
assign v4509 = ~(w14511 | w14657);
assign w14658 = v4509;
assign w14659 = w14456 & w14468;
assign v4510 = ~(w14469 | w14659);
assign w14660 = v4510;
assign w14661 = ~w14658 & w14660;
assign v4511 = ~(w14469 | w14661);
assign w14662 = v4511;
assign w14663 = w14407 & w14416;
assign v4512 = ~(w14417 | w14663);
assign w14664 = v4512;
assign w14665 = ~w14662 & w14664;
assign v4513 = ~(w14417 | w14665);
assign w14666 = v4513;
assign w14667 = w14378 & w14390;
assign v4514 = ~(w14391 | w14667);
assign w14668 = v4514;
assign w14669 = ~w14666 & w14668;
assign v4515 = ~(w14391 | w14669);
assign w14670 = v4515;
assign w14671 = w14354 & w14363;
assign v4516 = ~(w14364 | w14671);
assign w14672 = v4516;
assign w14673 = ~w14670 & w14672;
assign v4517 = ~(w14364 | w14673);
assign w14674 = v4517;
assign w14675 = w14329 & w14338;
assign v4518 = ~(w14339 | w14675);
assign w14676 = v4518;
assign w14677 = ~w14674 & w14676;
assign v4519 = ~(w14339 | w14677);
assign w14678 = v4519;
assign w14679 = w3529 & w13882;
assign w14680 = w3760 & ~w11734;
assign w14681 = w3763 & w11737;
assign w14682 = w3767 & w11740;
assign v4520 = ~(w14681 | w14682);
assign w14683 = v4520;
assign w14684 = ~w14680 & w14683;
assign w14685 = ~w14679 & w14684;
assign w14686 = ~pi29 & w14685;
assign w14687 = pi29 & ~w14685;
assign v4521 = ~(w14686 | w14687);
assign w14688 = v4521;
assign w14689 = w14678 & ~w14688;
assign w14690 = ~w14678 & w14688;
assign v4522 = ~(w14689 | w14690);
assign w14691 = v4522;
assign v4523 = ~(w13956 | w13958);
assign w14692 = v4523;
assign w14693 = w13657 & ~w14692;
assign w14694 = ~w13657 & w14692;
assign v4524 = ~(w14693 | w14694);
assign w14695 = v4524;
assign w14696 = w14691 & w14695;
assign v4525 = ~(w14689 | w14696);
assign w14697 = v4525;
assign w14698 = w14310 & w14697;
assign v4526 = ~(w14308 | w14698);
assign w14699 = v4526;
assign w14700 = ~w14283 & w14295;
assign v4527 = ~(w14296 | w14700);
assign w14701 = v4527;
assign w14702 = ~w14699 & w14701;
assign v4528 = ~(w14296 | w14702);
assign w14703 = v4528;
assign w14704 = ~w14270 & w14280;
assign v4529 = ~(w14281 | w14704);
assign w14705 = v4529;
assign w14706 = w14703 & w14705;
assign v4530 = ~(w14281 | w14706);
assign w14707 = v4530;
assign w14708 = ~w14257 & w14267;
assign v4531 = ~(w14268 | w14708);
assign w14709 = v4531;
assign w14710 = ~w14707 & w14709;
assign v4532 = ~(w14268 | w14710);
assign w14711 = v4532;
assign v4533 = ~(w14150 | w14152);
assign w14712 = v4533;
assign v4534 = ~(w14153 | w14712);
assign w14713 = v4534;
assign v4535 = ~(w14711 | w14713);
assign w14714 = v4535;
assign w14715 = w14711 & w14713;
assign v4536 = ~(w14714 | w14715);
assign w14716 = v4536;
assign w14717 = w4764 & ~w12842;
assign w14718 = w4913 & w11686;
assign w14719 = w4836 & w11689;
assign w14720 = w4763 & ~w11695;
assign v4537 = ~(w14719 | w14720);
assign w14721 = v4537;
assign w14722 = ~w14718 & w14721;
assign w14723 = ~w14717 & w14722;
assign w14724 = pi23 & w14723;
assign v4538 = ~(pi23 | w14723);
assign w14725 = v4538;
assign v4539 = ~(w14724 | w14725);
assign w14726 = v4539;
assign w14727 = w14716 & w14726;
assign v4540 = ~(w14714 | w14727);
assign w14728 = v4540;
assign w14729 = w14255 & w14728;
assign v4541 = ~(w14253 | w14729);
assign w14730 = v4541;
assign w14731 = w14240 & ~w14730;
assign w14732 = ~w14240 & w14730;
assign v4542 = ~(w14731 | w14732);
assign w14733 = v4542;
assign w14734 = w5114 & w11993;
assign w14735 = w5610 & w11984;
assign w14736 = w5531 & w11671;
assign w14737 = w5113 & w11673;
assign v4543 = ~(w14736 | w14737);
assign w14738 = v4543;
assign w14739 = ~w14735 & w14738;
assign w14740 = ~w14734 & w14739;
assign w14741 = pi20 & ~w14740;
assign w14742 = ~pi20 & w14740;
assign v4544 = ~(w14741 | w14742);
assign w14743 = v4544;
assign w14744 = w14733 & w14743;
assign v4545 = ~(w14731 | w14744);
assign w14745 = v4545;
assign w14746 = w14238 & ~w14745;
assign w14747 = ~w14238 & w14745;
assign v4546 = ~(w14746 | w14747);
assign w14748 = v4546;
assign w14749 = w5765 & ~w12277;
assign w14750 = w5983 & w12237;
assign w14751 = w6236 & w12271;
assign v4547 = ~(w14750 | w14751);
assign w14752 = v4547;
assign w14753 = w5764 & w12155;
assign w14754 = w14752 & ~w14753;
assign w14755 = ~w14749 & w14754;
assign w14756 = pi17 & w14755;
assign v4548 = ~(pi17 | w14755);
assign w14757 = v4548;
assign v4549 = ~(w14756 | w14757);
assign w14758 = v4549;
assign w14759 = w14748 & ~w14758;
assign v4550 = ~(w14746 | w14759);
assign w14760 = v4550;
assign w14761 = ~w14225 & w14235;
assign v4551 = ~(w14236 | w14761);
assign w14762 = v4551;
assign w14763 = ~w14760 & w14762;
assign v4552 = ~(w14236 | w14763);
assign w14764 = v4552;
assign w14765 = w14223 & ~w14764;
assign w14766 = ~w14223 & w14764;
assign v4553 = ~(w14765 | w14766);
assign w14767 = v4553;
assign w14768 = pi14 & w12406;
assign w14769 = pi13 & ~w12406;
assign v4554 = ~(w14768 | w14769);
assign w14770 = v4554;
assign w14771 = w6387 & w14770;
assign v4555 = ~(w12683 | w14771);
assign w14772 = v4555;
assign w14773 = w14767 & w14772;
assign v4556 = ~(w14765 | w14773);
assign w14774 = v4556;
assign w14775 = w14221 & ~w14774;
assign w14776 = ~w14221 & w14774;
assign v4557 = ~(w14767 | w14772);
assign w14777 = v4557;
assign v4558 = ~(w14773 | w14777);
assign w14778 = v4558;
assign w14779 = ~w14748 & w14758;
assign v4559 = ~(w14759 | w14779);
assign w14780 = v4559;
assign v4560 = ~(w14733 | w14743);
assign w14781 = v4560;
assign v4561 = ~(w14744 | w14781);
assign w14782 = v4561;
assign v4562 = ~(w14255 | w14728);
assign w14783 = v4562;
assign v4563 = ~(w14729 | w14783);
assign w14784 = v4563;
assign w14785 = w5114 & w12469;
assign w14786 = w5610 & w11671;
assign w14787 = w5531 & w11673;
assign w14788 = w5113 & w11678;
assign v4564 = ~(w14787 | w14788);
assign w14789 = v4564;
assign w14790 = ~w14786 & w14789;
assign w14791 = ~w14785 & w14790;
assign w14792 = pi20 & ~w14791;
assign w14793 = ~pi20 & w14791;
assign v4565 = ~(w14792 | w14793);
assign w14794 = v4565;
assign w14795 = w14784 & w14794;
assign w14796 = w14707 & ~w14709;
assign v4566 = ~(w14710 | w14796);
assign w14797 = v4566;
assign v4567 = ~(w14703 | w14705);
assign w14798 = v4567;
assign v4568 = ~(w14706 | w14798);
assign w14799 = v4568;
assign w14800 = w4153 & w13194;
assign w14801 = w4155 & w11711;
assign w14802 = ~w2873 & w11720;
assign w14803 = w4158 & w11714;
assign v4569 = ~(w14802 | w14803);
assign w14804 = v4569;
assign w14805 = ~w14801 & w14804;
assign w14806 = ~w14800 & w14805;
assign w14807 = pi26 & w14806;
assign v4570 = ~(pi26 | w14806);
assign w14808 = v4570;
assign v4571 = ~(w14807 | w14808);
assign w14809 = v4571;
assign w14810 = w14799 & w14809;
assign v4572 = ~(w14799 | w14809);
assign w14811 = v4572;
assign v4573 = ~(w14810 | w14811);
assign w14812 = v4573;
assign w14813 = w3529 & w13864;
assign w14814 = w3763 & w11729;
assign w14815 = w3760 & w11726;
assign v4574 = ~(w14814 | w14815);
assign w14816 = v4574;
assign w14817 = w3767 & ~w11734;
assign w14818 = w14816 & ~w14817;
assign w14819 = ~w14813 & w14818;
assign v4575 = ~(pi29 | w14819);
assign w14820 = v4575;
assign w14821 = pi29 & w14819;
assign v4576 = ~(w14820 | w14821);
assign w14822 = v4576;
assign w14823 = w4153 & w13514;
assign w14824 = w4155 & w11714;
assign w14825 = ~w2873 & w11723;
assign w14826 = w4158 & w11720;
assign v4577 = ~(w14825 | w14826);
assign w14827 = v4577;
assign w14828 = ~w14824 & w14827;
assign w14829 = ~w14823 & w14828;
assign w14830 = ~pi26 & w14829;
assign w14831 = pi26 & ~w14829;
assign v4578 = ~(w14830 | w14831);
assign w14832 = v4578;
assign w14833 = w14822 & ~w14832;
assign w14834 = w14699 & ~w14701;
assign v4579 = ~(w14702 | w14834);
assign w14835 = v4579;
assign w14836 = ~w14822 & w14832;
assign v4580 = ~(w14833 | w14836);
assign w14837 = v4580;
assign w14838 = ~w14835 & w14837;
assign v4581 = ~(w14833 | w14838);
assign w14839 = v4581;
assign w14840 = w14812 & ~w14839;
assign v4582 = ~(w14810 | w14840);
assign w14841 = v4582;
assign w14842 = ~w14797 & w14841;
assign w14843 = w14797 & ~w14841;
assign v4583 = ~(w14842 | w14843);
assign w14844 = v4583;
assign w14845 = w4764 & w12694;
assign w14846 = w4913 & w11689;
assign w14847 = w4763 & w11700;
assign w14848 = w4836 & ~w11695;
assign v4584 = ~(w14847 | w14848);
assign w14849 = v4584;
assign w14850 = ~w14846 & w14849;
assign w14851 = ~w14845 & w14850;
assign w14852 = pi23 & w14851;
assign v4585 = ~(pi23 | w14851);
assign w14853 = v4585;
assign v4586 = ~(w14852 | w14853);
assign w14854 = v4586;
assign w14855 = w14844 & ~w14854;
assign v4587 = ~(w14842 | w14855);
assign w14856 = v4587;
assign v4588 = ~(w14716 | w14726);
assign w14857 = v4588;
assign v4589 = ~(w14727 | w14857);
assign w14858 = v4589;
assign v4590 = ~(w14856 | w14858);
assign w14859 = v4590;
assign w14860 = w14856 & w14858;
assign v4591 = ~(w14859 | w14860);
assign w14861 = v4591;
assign w14862 = w5114 & w12454;
assign w14863 = w5531 & w11678;
assign w14864 = w5610 & w11673;
assign v4592 = ~(w14863 | w14864);
assign w14865 = v4592;
assign w14866 = w5113 & ~w11683;
assign w14867 = w14865 & ~w14866;
assign w14868 = ~w14862 & w14867;
assign w14869 = pi20 & w14868;
assign v4593 = ~(pi20 | w14868);
assign w14870 = v4593;
assign v4594 = ~(w14869 | w14870);
assign w14871 = v4594;
assign w14872 = w14861 & ~w14871;
assign v4595 = ~(w14859 | w14872);
assign w14873 = v4595;
assign v4596 = ~(w14784 | w14794);
assign w14874 = v4596;
assign v4597 = ~(w14795 | w14874);
assign w14875 = v4597;
assign w14876 = ~w14873 & w14875;
assign v4598 = ~(w14795 | w14876);
assign w14877 = v4598;
assign w14878 = w14782 & ~w14877;
assign w14879 = ~w14782 & w14877;
assign v4599 = ~(w14878 | w14879);
assign w14880 = v4599;
assign w14881 = w5765 & ~w12351;
assign w14882 = w5983 & w12155;
assign w14883 = w6236 & w12237;
assign v4600 = ~(w14882 | w14883);
assign w14884 = v4600;
assign w14885 = w5764 & w12084;
assign w14886 = w14884 & ~w14885;
assign w14887 = ~w14881 & w14886;
assign w14888 = pi17 & w14887;
assign v4601 = ~(pi17 | w14887);
assign w14889 = v4601;
assign v4602 = ~(w14888 | w14889);
assign w14890 = v4602;
assign w14891 = w14880 & ~w14890;
assign v4603 = ~(w14878 | w14891);
assign w14892 = v4603;
assign w14893 = w14780 & ~w14892;
assign w14894 = ~w14780 & w14892;
assign v4604 = ~(w14893 | w14894);
assign w14895 = v4604;
assign w14896 = w6389 & ~w12506;
assign w14897 = w7004 & ~w12406;
assign w14898 = w6388 & w12311;
assign w14899 = w6871 & w12381;
assign v4605 = ~(w14898 | w14899);
assign w14900 = v4605;
assign w14901 = ~w14897 & w14900;
assign w14902 = ~w14896 & w14901;
assign w14903 = pi14 & ~w14902;
assign w14904 = ~pi14 & w14902;
assign v4606 = ~(w14903 | w14904);
assign w14905 = v4606;
assign w14906 = w14895 & w14905;
assign v4607 = ~(w14893 | w14906);
assign w14907 = v4607;
assign w14908 = w6388 & w12381;
assign w14909 = w6389 & w12505;
assign v4608 = ~(w6871 | w14909);
assign w14910 = v4608;
assign v4609 = ~(w12406 | w14910);
assign w14911 = v4609;
assign v4610 = ~(w7004 | w14911);
assign w14912 = v4610;
assign w14913 = ~w14908 & w14912;
assign w14914 = ~pi14 & w14913;
assign w14915 = pi14 & ~w14913;
assign v4611 = ~(w14914 | w14915);
assign w14916 = v4611;
assign w14917 = ~w14907 & w14916;
assign w14918 = w14760 & ~w14762;
assign v4612 = ~(w14763 | w14918);
assign w14919 = v4612;
assign w14920 = w14907 & ~w14916;
assign v4613 = ~(w14917 | w14920);
assign w14921 = v4613;
assign w14922 = w14919 & w14921;
assign v4614 = ~(w14917 | w14922);
assign w14923 = v4614;
assign w14924 = w14778 & ~w14923;
assign w14925 = ~w14880 & w14890;
assign v4615 = ~(w14891 | w14925);
assign w14926 = v4615;
assign w14927 = w14873 & ~w14875;
assign v4616 = ~(w14876 | w14927);
assign w14928 = v4616;
assign w14929 = w5765 & w12167;
assign w14930 = w6236 & w12155;
assign w14931 = w5764 & w11984;
assign w14932 = w5983 & w12084;
assign v4617 = ~(w14931 | w14932);
assign w14933 = v4617;
assign w14934 = ~w14930 & w14933;
assign w14935 = ~w14929 & w14934;
assign w14936 = ~pi17 & w14935;
assign w14937 = pi17 & ~w14935;
assign v4618 = ~(w14936 | w14937);
assign w14938 = v4618;
assign w14939 = w14928 & w14938;
assign w14940 = ~w14812 & w14839;
assign v4619 = ~(w14840 | w14940);
assign w14941 = v4619;
assign w14942 = w4764 & ~w13008;
assign w14943 = w4836 & w11700;
assign w14944 = w4913 & ~w11695;
assign v4620 = ~(w14943 | w14944);
assign w14945 = v4620;
assign w14946 = w4763 & w11708;
assign w14947 = w14945 & ~w14946;
assign w14948 = ~w14942 & w14947;
assign w14949 = pi23 & w14948;
assign v4621 = ~(pi23 | w14948);
assign w14950 = v4621;
assign v4622 = ~(w14949 | w14950);
assign w14951 = v4622;
assign v4623 = ~(w14941 | w14951);
assign w14952 = v4623;
assign v4624 = ~(w14310 | w14697);
assign w14953 = v4624;
assign v4625 = ~(w14698 | w14953);
assign w14954 = v4625;
assign w14955 = w3529 & ~w13703;
assign w14956 = w3763 & ~w11734;
assign w14957 = w3760 & w11729;
assign v4626 = ~(w14956 | w14957);
assign w14958 = v4626;
assign w14959 = w3767 & w11737;
assign w14960 = w14958 & ~w14959;
assign w14961 = ~w14955 & w14960;
assign w14962 = pi29 & w14961;
assign v4627 = ~(pi29 | w14961);
assign w14963 = v4627;
assign v4628 = ~(w14962 | w14963);
assign w14964 = v4628;
assign w14965 = ~w14954 & w14964;
assign w14966 = w14954 & ~w14964;
assign v4629 = ~(w14965 | w14966);
assign w14967 = v4629;
assign w14968 = w4153 & ~w13310;
assign w14969 = w4155 & w11720;
assign w14970 = w4158 & w11723;
assign w14971 = ~w2873 & w11726;
assign v4630 = ~(w14970 | w14971);
assign w14972 = v4630;
assign w14973 = ~w14969 & w14972;
assign w14974 = ~w14968 & w14973;
assign w14975 = ~pi26 & w14974;
assign w14976 = pi26 & ~w14974;
assign v4631 = ~(w14975 | w14976);
assign w14977 = v4631;
assign w14978 = w14967 & ~w14977;
assign v4632 = ~(w14965 | w14978);
assign w14979 = v4632;
assign w14980 = w4764 & w12994;
assign w14981 = w4913 & w11700;
assign w14982 = w4763 & w11711;
assign w14983 = w4836 & w11708;
assign v4633 = ~(w14982 | w14983);
assign w14984 = v4633;
assign w14985 = ~w14981 & w14984;
assign w14986 = ~w14980 & w14985;
assign w14987 = ~pi23 & w14986;
assign w14988 = pi23 & ~w14986;
assign v4634 = ~(w14987 | w14988);
assign w14989 = v4634;
assign v4635 = ~(w14979 | w14989);
assign w14990 = v4635;
assign w14991 = w14835 & ~w14837;
assign v4636 = ~(w14838 | w14991);
assign w14992 = v4636;
assign w14993 = w14979 & w14989;
assign v4637 = ~(w14990 | w14993);
assign w14994 = v4637;
assign w14995 = w14992 & w14994;
assign v4638 = ~(w14990 | w14995);
assign w14996 = v4638;
assign w14997 = w14941 & w14951;
assign v4639 = ~(w14952 | w14997);
assign w14998 = v4639;
assign w14999 = w14996 & w14998;
assign v4640 = ~(w14952 | w14999);
assign w15000 = v4640;
assign w15001 = w5114 & w12594;
assign w15002 = w5610 & w11678;
assign w15003 = w5531 & ~w11683;
assign w15004 = w5113 & w11686;
assign v4641 = ~(w15003 | w15004);
assign w15005 = v4641;
assign w15006 = ~w15002 & w15005;
assign w15007 = ~w15001 & w15006;
assign w15008 = pi20 & ~w15007;
assign w15009 = ~pi20 & w15007;
assign v4642 = ~(w15008 | w15009);
assign w15010 = v4642;
assign w15011 = ~w15000 & w15010;
assign w15012 = ~w14844 & w14854;
assign v4643 = ~(w14855 | w15012);
assign w15013 = v4643;
assign w15014 = w15000 & ~w15010;
assign v4644 = ~(w15011 | w15014);
assign w15015 = v4644;
assign w15016 = w15013 & w15015;
assign v4645 = ~(w15011 | w15016);
assign w15017 = v4645;
assign w15018 = w5765 & w12181;
assign w15019 = w5983 & w11984;
assign w15020 = w6236 & w12084;
assign v4646 = ~(w15019 | w15020);
assign w15021 = v4646;
assign w15022 = w5764 & w11671;
assign w15023 = w15021 & ~w15022;
assign w15024 = ~w15018 & w15023;
assign v4647 = ~(pi17 | w15024);
assign w15025 = v4647;
assign w15026 = pi17 & w15024;
assign v4648 = ~(w15025 | w15026);
assign w15027 = v4648;
assign v4649 = ~(w15017 | w15027);
assign w15028 = v4649;
assign w15029 = ~w14861 & w14871;
assign v4650 = ~(w14872 | w15029);
assign w15030 = v4650;
assign w15031 = w15017 & w15027;
assign v4651 = ~(w15028 | w15031);
assign w15032 = v4651;
assign w15033 = w15030 & w15032;
assign v4652 = ~(w15028 | w15033);
assign w15034 = v4652;
assign v4653 = ~(w14928 | w14938);
assign w15035 = v4653;
assign v4654 = ~(w14939 | w15035);
assign w15036 = v4654;
assign w15037 = ~w15034 & w15036;
assign v4655 = ~(w14939 | w15037);
assign w15038 = v4655;
assign w15039 = w14926 & ~w15038;
assign w15040 = ~w14926 & w15038;
assign v4656 = ~(w15039 | w15040);
assign w15041 = v4656;
assign w15042 = w6389 & w12387;
assign w15043 = w6388 & w12271;
assign w15044 = w7004 & w12381;
assign v4657 = ~(w15043 | w15044);
assign w15045 = v4657;
assign w15046 = w6871 & w12311;
assign w15047 = w15045 & ~w15046;
assign w15048 = ~w15042 & w15047;
assign v4658 = ~(pi14 | w15048);
assign w15049 = v4658;
assign w15050 = pi14 & w15048;
assign v4659 = ~(w15049 | w15050);
assign w15051 = v4659;
assign w15052 = w15041 & ~w15051;
assign v4660 = ~(w15039 | w15052);
assign w15053 = v4660;
assign w15054 = w13167 & ~w15053;
assign v4661 = ~(w14895 | w14905);
assign w15055 = v4661;
assign v4662 = ~(w14906 | w15055);
assign w15056 = v4662;
assign w15057 = ~w13167 & w15053;
assign v4663 = ~(w15054 | w15057);
assign w15058 = v4663;
assign w15059 = w15056 & w15058;
assign v4664 = ~(w15054 | w15059);
assign w15060 = v4664;
assign v4665 = ~(w14919 | w14921);
assign w15061 = v4665;
assign v4666 = ~(w14922 | w15061);
assign w15062 = v4666;
assign w15063 = ~w15060 & w15062;
assign w15064 = w15060 & ~w15062;
assign v4667 = ~(w15063 | w15064);
assign w15065 = v4667;
assign v4668 = ~(w15056 | w15058);
assign w15066 = v4668;
assign v4669 = ~(w15059 | w15066);
assign w15067 = v4669;
assign w15068 = ~w15041 & w15051;
assign v4670 = ~(w15052 | w15068);
assign w15069 = v4670;
assign w15070 = w15034 & ~w15036;
assign v4671 = ~(w15037 | w15070);
assign w15071 = v4671;
assign w15072 = w6389 & w12318;
assign w15073 = w6871 & w12271;
assign w15074 = w7004 & w12311;
assign v4672 = ~(w15073 | w15074);
assign w15075 = v4672;
assign w15076 = w6388 & w12237;
assign w15077 = w15075 & ~w15076;
assign w15078 = ~w15072 & w15077;
assign w15079 = pi14 & w15078;
assign v4673 = ~(pi14 | w15078);
assign w15080 = v4673;
assign v4674 = ~(w15079 | w15080);
assign w15081 = v4674;
assign w15082 = w15071 & ~w15081;
assign v4675 = ~(w15030 | w15032);
assign w15083 = v4675;
assign v4676 = ~(w15033 | w15083);
assign w15084 = v4676;
assign v4677 = ~(w14996 | w14998);
assign w15085 = v4677;
assign v4678 = ~(w14999 | w15085);
assign w15086 = v4678;
assign w15087 = w5114 & w12610;
assign w15088 = w5610 & ~w11683;
assign w15089 = w5531 & w11686;
assign w15090 = w5113 & w11689;
assign v4679 = ~(w15089 | w15090);
assign w15091 = v4679;
assign w15092 = ~w15088 & w15091;
assign w15093 = ~w15087 & w15092;
assign w15094 = ~pi20 & w15093;
assign w15095 = pi20 & ~w15093;
assign v4680 = ~(w15094 | w15095);
assign w15096 = v4680;
assign w15097 = w15086 & w15096;
assign w15098 = w14674 & ~w14676;
assign v4681 = ~(w14677 | w15098);
assign w15099 = v4681;
assign w15100 = w3529 & w14288;
assign w15101 = w3760 & w11737;
assign w15102 = w3767 & ~w11745;
assign w15103 = w3763 & w11740;
assign v4682 = ~(w15102 | w15103);
assign w15104 = v4682;
assign w15105 = ~w15101 & w15104;
assign w15106 = ~w15100 & w15105;
assign w15107 = ~pi29 & w15106;
assign w15108 = pi29 & ~w15106;
assign v4683 = ~(w15107 | w15108);
assign w15109 = v4683;
assign w15110 = w15099 & w15109;
assign w15111 = w14670 & ~w14672;
assign v4684 = ~(w14673 | w15111);
assign w15112 = v4684;
assign w15113 = w3529 & w14300;
assign w15114 = w3763 & ~w11745;
assign w15115 = w3760 & w11740;
assign v4685 = ~(w15114 | w15115);
assign w15116 = v4685;
assign w15117 = w3767 & w11748;
assign w15118 = w15116 & ~w15117;
assign w15119 = ~w15113 & w15118;
assign w15120 = pi29 & w15119;
assign v4686 = ~(pi29 | w15119);
assign w15121 = v4686;
assign v4687 = ~(w15120 | w15121);
assign w15122 = v4687;
assign w15123 = w15112 & ~w15122;
assign w15124 = w14666 & ~w14668;
assign v4688 = ~(w14669 | w15124);
assign w15125 = v4688;
assign w15126 = w3529 & w13948;
assign w15127 = w3763 & w11748;
assign w15128 = w3760 & ~w11745;
assign v4689 = ~(w15127 | w15128);
assign w15129 = v4689;
assign w15130 = w3767 & w11759;
assign w15131 = w15129 & ~w15130;
assign w15132 = ~w15126 & w15131;
assign w15133 = pi29 & w15132;
assign v4690 = ~(pi29 | w15132);
assign w15134 = v4690;
assign v4691 = ~(w15133 | w15134);
assign w15135 = v4691;
assign w15136 = w15125 & ~w15135;
assign w15137 = w14662 & ~w14664;
assign v4692 = ~(w14665 | w15137);
assign w15138 = v4692;
assign w15139 = w3529 & ~w14331;
assign w15140 = w3760 & w11748;
assign w15141 = w3763 & w11759;
assign w15142 = w3767 & w11761;
assign v4693 = ~(w15141 | w15142);
assign w15143 = v4693;
assign w15144 = ~w15140 & w15143;
assign w15145 = ~w15139 & w15144;
assign w15146 = ~pi29 & w15145;
assign w15147 = pi29 & ~w15145;
assign v4694 = ~(w15146 | w15147);
assign w15148 = v4694;
assign w15149 = w15138 & w15148;
assign w15150 = w14658 & ~w14660;
assign v4695 = ~(w14661 | w15150);
assign w15151 = v4695;
assign w15152 = w3529 & w14356;
assign w15153 = w3767 & ~w11771;
assign w15154 = w3760 & w11759;
assign w15155 = w3763 & w11761;
assign v4696 = ~(w15154 | w15155);
assign w15156 = v4696;
assign w15157 = ~w15153 & w15156;
assign w15158 = ~w15152 & w15157;
assign w15159 = pi29 & ~w15158;
assign w15160 = ~pi29 & w15158;
assign v4697 = ~(w15159 | w15160);
assign w15161 = v4697;
assign w15162 = w15151 & w15161;
assign w15163 = w14654 & ~w14656;
assign v4698 = ~(w14657 | w15163);
assign w15164 = v4698;
assign w15165 = w3763 & ~w11771;
assign w15166 = w3760 & w11761;
assign w15167 = w3767 & w11768;
assign v4699 = ~(w15166 | w15167);
assign w15168 = v4699;
assign w15169 = ~w15165 & w15168;
assign w15170 = (w15169 & w14383) | (w15169 & w31273) | (w14383 & w31273);
assign w15171 = ~pi29 & w15170;
assign w15172 = pi29 & ~w15170;
assign v4700 = ~(w15171 | w15172);
assign w15173 = v4700;
assign w15174 = w15164 & w15173;
assign w15175 = w14650 & ~w14652;
assign v4701 = ~(w14653 | w15175);
assign w15176 = v4701;
assign w15177 = w3529 & w14409;
assign w15178 = w3763 & w11768;
assign w15179 = w3760 & ~w11771;
assign v4702 = ~(w15178 | w15179);
assign w15180 = v4702;
assign w15181 = w3767 & w11776;
assign w15182 = w15180 & ~w15181;
assign w15183 = ~w15177 & w31274;
assign w15184 = (~pi29 & w15177) | (~pi29 & w31275) | (w15177 & w31275);
assign v4703 = ~(w15183 | w15184);
assign w15185 = v4703;
assign w15186 = w15176 & ~w15185;
assign w15187 = ~w14578 & w14648;
assign v4704 = ~(w14649 | w15187);
assign w15188 = v4704;
assign w15189 = w3767 & w11784;
assign w15190 = w3760 & w11768;
assign v4705 = ~(w15189 | w15190);
assign w15191 = v4705;
assign w15192 = w3763 & w11776;
assign w15193 = (~w14461 & w31177) | (~w14461 & w31178) | (w31177 & w31178);
assign w15194 = (w14461 & w31179) | (w14461 & w31180) | (w31179 & w31180);
assign v4706 = ~(w15193 | w15194);
assign w15195 = v4706;
assign w15196 = w15188 & ~w15195;
assign w15197 = ~w14637 & w14646;
assign v4707 = ~(w14647 | w15197);
assign w15198 = v4707;
assign w15199 = w3763 & w11784;
assign w15200 = w3760 & w11776;
assign v4708 = ~(w15199 | w15200);
assign w15201 = v4708;
assign w15202 = w3767 & w11793;
assign w15203 = w15201 & ~w15202;
assign w15204 = (w14504 & w31037) | (w14504 & w31038) | (w31037 & w31038);
assign w15205 = (~w14504 & w31039) | (~w14504 & w31040) | (w31039 & w31040);
assign v4709 = ~(w15204 | w15205);
assign w15206 = v4709;
assign w15207 = w15198 & ~w15206;
assign w15208 = w14607 & w14614;
assign v4710 = ~(w14615 | w15208);
assign w15209 = v4710;
assign w15210 = w3529 & w14547;
assign w15211 = w3763 & w11793;
assign w15212 = w3760 & w11784;
assign w15213 = w3767 & w11803;
assign v4711 = ~(w15212 | w15213);
assign w15214 = v4711;
assign w15215 = (pi29 & w15210) | (pi29 & w30617) | (w15210 & w30617);
assign w15216 = ~w15210 & w30618;
assign v4712 = ~(w15215 | w15216);
assign w15217 = v4712;
assign w15218 = w15209 & w15217;
assign w15219 = ~w3405 & w11800;
assign w15220 = w3525 & w11800;
assign w15221 = pi29 & w15220;
assign w15222 = w3529 & ~w14609;
assign w15223 = w3760 & w11798;
assign w15224 = w3763 & w11800;
assign v4713 = ~(w15223 | w15224);
assign w15225 = v4713;
assign w15226 = ~w15222 & w15225;
assign w15227 = ~w15222 & w31181;
assign w15228 = pi29 & ~w15227;
assign w15229 = w3767 & w11800;
assign w15230 = (~w15229 & w14639) | (~w15229 & w31182) | (w14639 & w31182);
assign w15231 = w3760 & w11803;
assign w15232 = w3763 & w11798;
assign v4714 = ~(w15231 | w15232);
assign w15233 = v4714;
assign w15234 = w15230 & w15233;
assign w15235 = ~w15228 & w15234;
assign w15236 = pi29 & w15235;
assign w15237 = w15219 & w15236;
assign v4715 = ~(w15219 | w15236);
assign w15238 = v4715;
assign v4716 = ~(w15237 | w15238);
assign w15239 = v4716;
assign w15240 = w3529 & w14569;
assign w15241 = w3767 & w11798;
assign w15242 = w3760 & w11793;
assign w15243 = w3763 & w11803;
assign v4717 = ~(w15242 | w15243);
assign w15244 = v4717;
assign w15245 = ~w15241 & w15244;
assign w15246 = (pi29 & w15240) | (pi29 & w31183) | (w15240 & w31183);
assign w15247 = ~w15240 & w31184;
assign v4718 = ~(w15246 | w15247);
assign w15248 = v4718;
assign w15249 = w15239 & w15248;
assign v4719 = ~(w15237 | w15249);
assign w15250 = v4719;
assign v4720 = ~(w15209 | w15217);
assign w15251 = v4720;
assign v4721 = ~(w15218 | w15251);
assign w15252 = v4721;
assign w15253 = ~w15250 & w15252;
assign w15254 = (~w15218 & ~w15252) | (~w15218 & w31041) | (~w15252 & w31041);
assign w15255 = ~w15198 & w15206;
assign v4722 = ~(w15207 | w15255);
assign w15256 = v4722;
assign w15257 = ~w15254 & w15256;
assign v4723 = ~(w15207 | w15257);
assign w15258 = v4723;
assign w15259 = ~w15188 & w15195;
assign v4724 = ~(w15196 | w15259);
assign w15260 = v4724;
assign w15261 = ~w15258 & w15260;
assign w15262 = (~w15196 & w15258) | (~w15196 & w31185) | (w15258 & w31185);
assign w15263 = ~w15176 & w15185;
assign v4725 = ~(w15186 | w15263);
assign w15264 = v4725;
assign w15265 = ~w15262 & w15264;
assign w15266 = (~w15186 & w15262) | (~w15186 & w31276) | (w15262 & w31276);
assign v4726 = ~(w15164 | w15173);
assign w15267 = v4726;
assign v4727 = ~(w15174 | w15267);
assign w15268 = v4727;
assign w15269 = ~w15266 & w15268;
assign v4728 = ~(w15174 | w15269);
assign w15270 = v4728;
assign v4729 = ~(w15151 | w15161);
assign w15271 = v4729;
assign v4730 = ~(w15162 | w15271);
assign w15272 = v4730;
assign w15273 = ~w15270 & w15272;
assign v4731 = ~(w15162 | w15273);
assign w15274 = v4731;
assign v4732 = ~(w15138 | w15148);
assign w15275 = v4732;
assign v4733 = ~(w15149 | w15275);
assign w15276 = v4733;
assign w15277 = ~w15274 & w15276;
assign v4734 = ~(w15149 | w15277);
assign w15278 = v4734;
assign w15279 = ~w15125 & w15135;
assign v4735 = ~(w15136 | w15279);
assign w15280 = v4735;
assign w15281 = ~w15278 & w15280;
assign v4736 = ~(w15136 | w15281);
assign w15282 = v4736;
assign w15283 = ~w15112 & w15122;
assign v4737 = ~(w15123 | w15283);
assign w15284 = v4737;
assign w15285 = ~w15282 & w15284;
assign v4738 = ~(w15123 | w15285);
assign w15286 = v4738;
assign v4739 = ~(w15099 | w15109);
assign w15287 = v4739;
assign v4740 = ~(w15110 | w15287);
assign w15288 = v4740;
assign w15289 = ~w15286 & w15288;
assign v4741 = ~(w15110 | w15289);
assign w15290 = v4741;
assign w15291 = w4153 & ~w13737;
assign w15292 = ~w2873 & w11729;
assign w15293 = w4155 & w11723;
assign v4742 = ~(w15292 | w15293);
assign w15294 = v4742;
assign w15295 = w4158 & w11726;
assign w15296 = w15294 & ~w15295;
assign w15297 = ~w15291 & w15296;
assign w15298 = pi26 & w15297;
assign v4743 = ~(pi26 | w15297);
assign w15299 = v4743;
assign v4744 = ~(w15298 | w15299);
assign w15300 = v4744;
assign v4745 = ~(w15290 | w15300);
assign w15301 = v4745;
assign w15302 = w15290 & w15300;
assign v4746 = ~(w15301 | w15302);
assign w15303 = v4746;
assign v4747 = ~(w14691 | w14695);
assign w15304 = v4747;
assign v4748 = ~(w14696 | w15304);
assign w15305 = v4748;
assign w15306 = w15303 & ~w15305;
assign v4749 = ~(w15301 | w15306);
assign w15307 = v4749;
assign w15308 = w4764 & w13178;
assign w15309 = w4913 & w11708;
assign w15310 = w4763 & w11714;
assign w15311 = w4836 & w11711;
assign v4750 = ~(w15310 | w15311);
assign w15312 = v4750;
assign w15313 = ~w15309 & w15312;
assign w15314 = ~w15308 & w15313;
assign w15315 = ~pi23 & w15314;
assign w15316 = pi23 & ~w15314;
assign v4751 = ~(w15315 | w15316);
assign w15317 = v4751;
assign w15318 = ~w15307 & w15317;
assign w15319 = w15307 & ~w15317;
assign v4752 = ~(w15318 | w15319);
assign w15320 = v4752;
assign w15321 = ~w14967 & w14977;
assign v4753 = ~(w14978 | w15321);
assign w15322 = v4753;
assign w15323 = w15320 & ~w15322;
assign v4754 = ~(w15318 | w15323);
assign w15324 = v4754;
assign w15325 = w5114 & ~w12842;
assign w15326 = w5610 & w11686;
assign w15327 = w5531 & w11689;
assign w15328 = w5113 & ~w11695;
assign v4755 = ~(w15327 | w15328);
assign w15329 = v4755;
assign w15330 = ~w15326 & w15329;
assign w15331 = ~w15325 & w15330;
assign w15332 = ~pi20 & w15331;
assign w15333 = pi20 & ~w15331;
assign v4756 = ~(w15332 | w15333);
assign w15334 = v4756;
assign w15335 = w15324 & ~w15334;
assign w15336 = ~w15324 & w15334;
assign v4757 = ~(w15335 | w15336);
assign w15337 = v4757;
assign v4758 = ~(w14992 | w14994);
assign w15338 = v4758;
assign v4759 = ~(w14995 | w15338);
assign w15339 = v4759;
assign w15340 = w15337 & w15339;
assign v4760 = ~(w15335 | w15340);
assign w15341 = v4760;
assign v4761 = ~(w15086 | w15096);
assign w15342 = v4761;
assign v4762 = ~(w15097 | w15342);
assign w15343 = v4762;
assign w15344 = w15341 & w15343;
assign v4763 = ~(w15097 | w15344);
assign w15345 = v4763;
assign w15346 = w5765 & w11993;
assign w15347 = w5983 & w11671;
assign w15348 = w6236 & w11984;
assign v4764 = ~(w15347 | w15348);
assign w15349 = v4764;
assign w15350 = w5764 & w11673;
assign w15351 = w15349 & ~w15350;
assign w15352 = ~w15346 & w15351;
assign w15353 = pi17 & w15352;
assign v4765 = ~(pi17 | w15352);
assign w15354 = v4765;
assign v4766 = ~(w15353 | w15354);
assign w15355 = v4766;
assign v4767 = ~(w15345 | w15355);
assign w15356 = v4767;
assign v4768 = ~(w15013 | w15015);
assign w15357 = v4768;
assign v4769 = ~(w15016 | w15357);
assign w15358 = v4769;
assign w15359 = w15345 & w15355;
assign v4770 = ~(w15356 | w15359);
assign w15360 = v4770;
assign w15361 = w15358 & w15360;
assign v4771 = ~(w15356 | w15361);
assign w15362 = v4771;
assign w15363 = w15084 & ~w15362;
assign w15364 = ~w15084 & w15362;
assign v4772 = ~(w15363 | w15364);
assign w15365 = v4772;
assign w15366 = w6389 & ~w12277;
assign w15367 = w7004 & w12271;
assign w15368 = w6388 & w12155;
assign w15369 = w6871 & w12237;
assign v4773 = ~(w15368 | w15369);
assign w15370 = v4773;
assign w15371 = ~w15367 & w15370;
assign w15372 = ~w15366 & w15371;
assign w15373 = pi14 & w15372;
assign v4774 = ~(pi14 | w15372);
assign w15374 = v4774;
assign v4775 = ~(w15373 | w15374);
assign w15375 = v4775;
assign w15376 = w15365 & ~w15375;
assign v4776 = ~(w15363 | w15376);
assign w15377 = v4776;
assign w15378 = ~w15071 & w15081;
assign v4777 = ~(w15082 | w15378);
assign w15379 = v4777;
assign w15380 = ~w15377 & w15379;
assign v4778 = ~(w15082 | w15380);
assign w15381 = v4778;
assign w15382 = w15069 & ~w15381;
assign w15383 = ~w15069 & w15381;
assign v4779 = ~(w15382 | w15383);
assign w15384 = v4779;
assign w15385 = pi11 & w12406;
assign w15386 = pi10 & ~w12406;
assign v4780 = ~(w15385 | w15386);
assign w15387 = v4780;
assign w15388 = w7176 & w15387;
assign v4781 = ~(w13165 | w15388);
assign w15389 = v4781;
assign w15390 = w15384 & w15389;
assign v4782 = ~(w15382 | w15390);
assign w15391 = v4782;
assign w15392 = ~w15067 & w15391;
assign v4783 = ~(w15384 | w15389);
assign w15393 = v4783;
assign v4784 = ~(w15390 | w15393);
assign w15394 = v4784;
assign w15395 = w15377 & ~w15379;
assign v4785 = ~(w15380 | w15395);
assign w15396 = v4785;
assign w15397 = w7177 & w12381;
assign w15398 = w7178 & w12505;
assign v4786 = ~(w7466 | w15398);
assign w15399 = v4786;
assign v4787 = ~(w12406 | w15399);
assign w15400 = v4787;
assign v4788 = ~(w7765 | w15400);
assign w15401 = v4788;
assign w15402 = ~w15397 & w15401;
assign w15403 = ~pi11 & w15402;
assign w15404 = pi11 & ~w15402;
assign v4789 = ~(w15403 | w15404);
assign w15405 = v4789;
assign w15406 = w15396 & w15405;
assign w15407 = ~w15365 & w15375;
assign v4790 = ~(w15376 | w15407);
assign w15408 = v4790;
assign v4791 = ~(w15341 | w15343);
assign w15409 = v4791;
assign v4792 = ~(w15344 | w15409);
assign w15410 = v4792;
assign w15411 = w5765 & w12469;
assign w15412 = w5983 & w11673;
assign w15413 = w6236 & w11671;
assign v4793 = ~(w15412 | w15413);
assign w15414 = v4793;
assign w15415 = w5764 & w11678;
assign w15416 = w15414 & ~w15415;
assign w15417 = ~w15411 & w15416;
assign v4794 = ~(pi17 | w15417);
assign w15418 = v4794;
assign w15419 = pi17 & w15417;
assign v4795 = ~(w15418 | w15419);
assign w15420 = v4795;
assign w15421 = w15410 & ~w15420;
assign w15422 = w15286 & ~w15288;
assign v4796 = ~(w15289 | w15422);
assign w15423 = v4796;
assign w15424 = w4153 & w13864;
assign w15425 = w4155 & w11726;
assign v4797 = ~(w2873 | w11734);
assign w15426 = v4797;
assign w15427 = w4158 & w11729;
assign v4798 = ~(w15426 | w15427);
assign w15428 = v4798;
assign w15429 = ~w15425 & w15428;
assign w15430 = ~w15424 & w15429;
assign w15431 = ~pi26 & w15430;
assign w15432 = pi26 & ~w15430;
assign v4799 = ~(w15431 | w15432);
assign w15433 = v4799;
assign w15434 = w15423 & w15433;
assign w15435 = w15282 & ~w15284;
assign v4800 = ~(w15285 | w15435);
assign w15436 = v4800;
assign w15437 = w4153 & ~w13703;
assign w15438 = w4155 & w11729;
assign w15439 = w4158 & ~w11734;
assign w15440 = ~w2873 & w11737;
assign v4801 = ~(w15439 | w15440);
assign w15441 = v4801;
assign w15442 = ~w15438 & w15441;
assign w15443 = ~w15437 & w15442;
assign w15444 = ~pi26 & w15443;
assign w15445 = pi26 & ~w15443;
assign v4802 = ~(w15444 | w15445);
assign w15446 = v4802;
assign w15447 = w15436 & w15446;
assign w15448 = w15278 & ~w15280;
assign v4803 = ~(w15281 | w15448);
assign w15449 = v4803;
assign w15450 = w4153 & w13882;
assign w15451 = ~w2873 & w11740;
assign w15452 = w4155 & ~w11734;
assign v4804 = ~(w15451 | w15452);
assign w15453 = v4804;
assign w15454 = w4158 & w11737;
assign w15455 = w15453 & ~w15454;
assign w15456 = ~w15450 & w15455;
assign w15457 = pi26 & w15456;
assign v4805 = ~(pi26 | w15456);
assign w15458 = v4805;
assign v4806 = ~(w15457 | w15458);
assign w15459 = v4806;
assign w15460 = w15449 & ~w15459;
assign w15461 = w15274 & ~w15276;
assign v4807 = ~(w15277 | w15461);
assign w15462 = v4807;
assign w15463 = w4153 & w14288;
assign w15464 = w4155 & w11737;
assign v4808 = ~(w2873 | w11745);
assign w15465 = v4808;
assign w15466 = w4158 & w11740;
assign v4809 = ~(w15465 | w15466);
assign w15467 = v4809;
assign w15468 = ~w15464 & w15467;
assign w15469 = ~w15463 & w15468;
assign w15470 = pi26 & ~w15469;
assign w15471 = ~pi26 & w15469;
assign v4810 = ~(w15470 | w15471);
assign w15472 = v4810;
assign w15473 = w15462 & w15472;
assign w15474 = w15270 & ~w15272;
assign v4811 = ~(w15273 | w15474);
assign w15475 = v4811;
assign w15476 = w4153 & w14300;
assign w15477 = w4155 & w11740;
assign w15478 = ~w2873 & w11748;
assign w15479 = w4158 & ~w11745;
assign v4812 = ~(w15478 | w15479);
assign w15480 = v4812;
assign w15481 = ~w15477 & w15480;
assign w15482 = ~w15476 & w15481;
assign w15483 = ~pi26 & w15482;
assign w15484 = pi26 & ~w15482;
assign v4813 = ~(w15483 | w15484);
assign w15485 = v4813;
assign w15486 = w15475 & w15485;
assign w15487 = w15266 & ~w15268;
assign v4814 = ~(w15269 | w15487);
assign w15488 = v4814;
assign w15489 = w4153 & w13948;
assign w15490 = w4155 & ~w11745;
assign w15491 = ~w2873 & w11759;
assign w15492 = w4158 & w11748;
assign v4815 = ~(w15491 | w15492);
assign w15493 = v4815;
assign w15494 = ~w15490 & w15493;
assign w15495 = ~w15489 & w15494;
assign w15496 = ~pi26 & w15495;
assign w15497 = pi26 & ~w15495;
assign v4816 = ~(w15496 | w15497);
assign w15498 = v4816;
assign w15499 = w15488 & w15498;
assign w15500 = w15262 & ~w15264;
assign v4817 = ~(w15265 | w15500);
assign w15501 = v4817;
assign w15502 = w4153 & ~w14331;
assign w15503 = w4155 & w11748;
assign w15504 = ~w2873 & w11761;
assign w15505 = w4158 & w11759;
assign v4818 = ~(w15504 | w15505);
assign w15506 = v4818;
assign w15507 = ~w15503 & w15506;
assign w15508 = ~w15502 & w15507;
assign w15509 = ~pi26 & w15508;
assign w15510 = pi26 & ~w15508;
assign v4819 = ~(w15509 | w15510);
assign w15511 = v4819;
assign w15512 = w15501 & w15511;
assign w15513 = w15258 & ~w15260;
assign v4820 = ~(w15261 | w15513);
assign w15514 = v4820;
assign v4821 = ~(w2873 | w11771);
assign w15515 = v4821;
assign w15516 = w4155 & w11759;
assign w15517 = w4158 & w11761;
assign v4822 = ~(w15516 | w15517);
assign w15518 = v4822;
assign w15519 = ~w15515 & w15518;
assign w15520 = (w15519 & ~w14356) | (w15519 & w31186) | (~w14356 & w31186);
assign w15521 = pi26 & ~w15520;
assign w15522 = ~pi26 & w15520;
assign v4823 = ~(w15521 | w15522);
assign w15523 = v4823;
assign w15524 = w15514 & w15523;
assign w15525 = w15254 & ~w15256;
assign v4824 = ~(w15257 | w15525);
assign w15526 = v4824;
assign w15527 = w4158 & ~w11771;
assign w15528 = w4155 & w11761;
assign w15529 = ~w2873 & w11768;
assign v4825 = ~(w15528 | w15529);
assign w15530 = v4825;
assign w15531 = ~w15527 & w15530;
assign w15532 = (w14383 & w31187) | (w14383 & w31188) | (w31187 & w31188);
assign w15533 = (~w14383 & w31189) | (~w14383 & w31190) | (w31189 & w31190);
assign v4826 = ~(w15532 | w15533);
assign w15534 = v4826;
assign w15535 = w15526 & w15534;
assign w15536 = w15250 & ~w15252;
assign v4827 = ~(w15253 | w15536);
assign w15537 = v4827;
assign w15538 = w4153 & w14409;
assign w15539 = ~w2873 & w11776;
assign w15540 = w4155 & ~w11771;
assign w15541 = w4158 & w11768;
assign v4828 = ~(w15540 | w15541);
assign w15542 = v4828;
assign w15543 = (pi26 & w15538) | (pi26 & w30619) | (w15538 & w30619);
assign w15544 = ~w15538 & w30620;
assign v4829 = ~(w15543 | w15544);
assign w15545 = v4829;
assign w15546 = w15537 & w15545;
assign v4830 = ~(w15239 | w15248);
assign w15547 = v4830;
assign v4831 = ~(w15249 | w15547);
assign w15548 = v4831;
assign w15549 = w4155 & w11768;
assign w15550 = ~w2873 & w11784;
assign w15551 = w4158 & w11776;
assign v4832 = ~(w15550 | w15551);
assign w15552 = v4832;
assign w15553 = ~w15549 & w15552;
assign w15554 = (~w14461 & w30621) | (~w14461 & w30622) | (w30621 & w30622);
assign w15555 = (w14461 & w30623) | (w14461 & w30624) | (w30623 & w30624);
assign v4833 = ~(w15554 | w15555);
assign w15556 = v4833;
assign w15557 = w15548 & w15556;
assign w15558 = w15228 & ~w15234;
assign v4834 = ~(w15235 | w15558);
assign w15559 = v4834;
assign w15560 = w4158 & w11784;
assign w15561 = w4155 & w11776;
assign v4835 = ~(w15560 | w15561);
assign w15562 = v4835;
assign w15563 = ~w2873 & w11793;
assign w15564 = (w14504 & w30500) | (w14504 & w30501) | (w30500 & w30501);
assign w15565 = (~w14504 & w30502) | (~w14504 & w30503) | (w30502 & w30503);
assign v4836 = ~(w15564 | w15565);
assign w15566 = v4836;
assign w15567 = w15559 & ~w15566;
assign w15568 = w15221 & ~w15226;
assign v4837 = ~(w15227 | w15568);
assign w15569 = v4837;
assign w15570 = w4153 & w14547;
assign w15571 = w4158 & w11793;
assign w15572 = w4155 & w11784;
assign w15573 = ~w2873 & w11803;
assign v4838 = ~(w15572 | w15573);
assign w15574 = v4838;
assign w15575 = (pi26 & w15570) | (pi26 & w30344) | (w15570 & w30344);
assign w15576 = ~w15570 & w30345;
assign v4839 = ~(w15575 | w15576);
assign w15577 = v4839;
assign w15578 = w15569 & w15577;
assign w15579 = w4152 & w11800;
assign w15580 = pi26 & w15579;
assign w15581 = w4153 & ~w14609;
assign w15582 = w4155 & w11798;
assign w15583 = w4158 & w11800;
assign v4840 = ~(w15582 | w15583);
assign w15584 = v4840;
assign w15585 = ~w15581 & w15584;
assign w15586 = ~w15580 & w15585;
assign w15587 = ~w2873 & w11800;
assign w15588 = (~w15587 & w14639) | (~w15587 & w31043) | (w14639 & w31043);
assign w15589 = w4155 & w11803;
assign w15590 = w4158 & w11798;
assign v4841 = ~(w15589 | w15590);
assign w15591 = v4841;
assign w15592 = w15588 & w15591;
assign w15593 = pi26 & w15592;
assign w15594 = w15586 & w15593;
assign w15595 = w15220 & w15594;
assign v4842 = ~(w15220 | w15594);
assign w15596 = v4842;
assign v4843 = ~(w15595 | w15596);
assign w15597 = v4843;
assign w15598 = w4158 & w11803;
assign w15599 = w4155 & w11793;
assign w15600 = ~w2873 & w11798;
assign v4844 = ~(w15599 | w15600);
assign w15601 = v4844;
assign w15602 = ~w15598 & w15601;
assign w15603 = (w15602 & ~w14569) | (w15602 & w30625) | (~w14569 & w30625);
assign w15604 = pi26 & ~w15603;
assign w15605 = ~pi26 & w15603;
assign v4845 = ~(w15604 | w15605);
assign w15606 = v4845;
assign w15607 = w15597 & w15606;
assign v4846 = ~(w15595 | w15607);
assign w15608 = v4846;
assign v4847 = ~(w15569 | w15577);
assign w15609 = v4847;
assign v4848 = ~(w15578 | w15609);
assign w15610 = v4848;
assign w15611 = ~w15608 & w15610;
assign w15612 = (~w15578 & ~w15610) | (~w15578 & w30504) | (~w15610 & w30504);
assign w15613 = ~w15559 & w15566;
assign v4849 = ~(w15567 | w15613);
assign w15614 = v4849;
assign w15615 = ~w15612 & w15614;
assign v4850 = ~(w15567 | w15615);
assign w15616 = v4850;
assign v4851 = ~(w15548 | w15556);
assign w15617 = v4851;
assign v4852 = ~(w15557 | w15617);
assign w15618 = v4852;
assign w15619 = ~w15616 & w15618;
assign w15620 = (~w15557 & w15616) | (~w15557 & w30626) | (w15616 & w30626);
assign v4853 = ~(w15537 | w15545);
assign w15621 = v4853;
assign v4854 = ~(w15546 | w15621);
assign w15622 = v4854;
assign w15623 = ~w15620 & w15622;
assign w15624 = (~w15546 & w15620) | (~w15546 & w30810) | (w15620 & w30810);
assign v4855 = ~(w15526 | w15534);
assign w15625 = v4855;
assign v4856 = ~(w15535 | w15625);
assign w15626 = v4856;
assign w15627 = ~w15624 & w15626;
assign w15628 = (~w15535 & w15624) | (~w15535 & w31044) | (w15624 & w31044);
assign v4857 = ~(w15514 | w15523);
assign w15629 = v4857;
assign v4858 = ~(w15524 | w15629);
assign w15630 = v4858;
assign w15631 = ~w15628 & w15630;
assign v4859 = ~(w15524 | w15631);
assign w15632 = v4859;
assign v4860 = ~(w15501 | w15511);
assign w15633 = v4860;
assign v4861 = ~(w15512 | w15633);
assign w15634 = v4861;
assign w15635 = ~w15632 & w15634;
assign w15636 = (~w15512 & w15632) | (~w15512 & w31191) | (w15632 & w31191);
assign v4862 = ~(w15488 | w15498);
assign w15637 = v4862;
assign v4863 = ~(w15499 | w15637);
assign w15638 = v4863;
assign w15639 = ~w15636 & w15638;
assign w15640 = (~w15499 & w15636) | (~w15499 & w31277) | (w15636 & w31277);
assign v4864 = ~(w15475 | w15485);
assign w15641 = v4864;
assign v4865 = ~(w15486 | w15641);
assign w15642 = v4865;
assign w15643 = ~w15640 & w15642;
assign v4866 = ~(w15486 | w15643);
assign w15644 = v4866;
assign v4867 = ~(w15462 | w15472);
assign w15645 = v4867;
assign v4868 = ~(w15473 | w15645);
assign w15646 = v4868;
assign w15647 = ~w15644 & w15646;
assign v4869 = ~(w15473 | w15647);
assign w15648 = v4869;
assign w15649 = ~w15449 & w15459;
assign v4870 = ~(w15460 | w15649);
assign w15650 = v4870;
assign w15651 = ~w15648 & w15650;
assign v4871 = ~(w15460 | w15651);
assign w15652 = v4871;
assign v4872 = ~(w15436 | w15446);
assign w15653 = v4872;
assign v4873 = ~(w15447 | w15653);
assign w15654 = v4873;
assign w15655 = ~w15652 & w15654;
assign v4874 = ~(w15447 | w15655);
assign w15656 = v4874;
assign v4875 = ~(w15423 | w15433);
assign w15657 = v4875;
assign v4876 = ~(w15434 | w15657);
assign w15658 = v4876;
assign w15659 = ~w15656 & w15658;
assign v4877 = ~(w15434 | w15659);
assign w15660 = v4877;
assign w15661 = w4764 & w13194;
assign w15662 = w4836 & w11714;
assign w15663 = w4913 & w11711;
assign v4878 = ~(w15662 | w15663);
assign w15664 = v4878;
assign w15665 = w4763 & w11720;
assign w15666 = w15664 & ~w15665;
assign w15667 = ~w15661 & w15666;
assign w15668 = pi23 & w15667;
assign v4879 = ~(pi23 | w15667);
assign w15669 = v4879;
assign v4880 = ~(w15668 | w15669);
assign w15670 = v4880;
assign w15671 = w15660 & w15670;
assign w15672 = ~w15303 & w15305;
assign v4881 = ~(w15306 | w15672);
assign w15673 = v4881;
assign v4882 = ~(w15660 | w15670);
assign w15674 = v4882;
assign v4883 = ~(w15671 | w15674);
assign w15675 = v4883;
assign w15676 = ~w15673 & w15675;
assign v4884 = ~(w15671 | w15676);
assign w15677 = v4884;
assign w15678 = w5114 & w12694;
assign w15679 = w5610 & w11689;
assign w15680 = w5113 & w11700;
assign w15681 = w5531 & ~w11695;
assign v4885 = ~(w15680 | w15681);
assign w15682 = v4885;
assign w15683 = ~w15679 & w15682;
assign w15684 = ~w15678 & w15683;
assign w15685 = ~pi20 & w15684;
assign w15686 = pi20 & ~w15684;
assign v4886 = ~(w15685 | w15686);
assign w15687 = v4886;
assign v4887 = ~(w15677 | w15687);
assign w15688 = v4887;
assign w15689 = ~w15320 & w15322;
assign v4888 = ~(w15323 | w15689);
assign w15690 = v4888;
assign w15691 = w15677 & w15687;
assign v4889 = ~(w15688 | w15691);
assign w15692 = v4889;
assign w15693 = ~w15690 & w15692;
assign v4890 = ~(w15688 | w15693);
assign w15694 = v4890;
assign w15695 = w5765 & w12454;
assign w15696 = w5983 & w11678;
assign w15697 = w6236 & w11673;
assign v4891 = ~(w15696 | w15697);
assign w15698 = v4891;
assign w15699 = w5764 & ~w11683;
assign w15700 = w15698 & ~w15699;
assign w15701 = ~w15695 & w15700;
assign w15702 = pi17 & w15701;
assign v4892 = ~(pi17 | w15701);
assign w15703 = v4892;
assign v4893 = ~(w15702 | w15703);
assign w15704 = v4893;
assign w15705 = w15694 & ~w15704;
assign v4894 = ~(w15337 | w15339);
assign w15706 = v4894;
assign v4895 = ~(w15340 | w15706);
assign w15707 = v4895;
assign w15708 = ~w15694 & w15704;
assign v4896 = ~(w15705 | w15708);
assign w15709 = v4896;
assign w15710 = ~w15707 & w15709;
assign v4897 = ~(w15705 | w15710);
assign w15711 = v4897;
assign w15712 = ~w15410 & w15420;
assign v4898 = ~(w15421 | w15712);
assign w15713 = v4898;
assign w15714 = ~w15711 & w15713;
assign v4899 = ~(w15421 | w15714);
assign w15715 = v4899;
assign w15716 = w6389 & ~w12351;
assign w15717 = w6871 & w12155;
assign w15718 = w7004 & w12237;
assign v4900 = ~(w15717 | w15718);
assign w15719 = v4900;
assign w15720 = w6388 & w12084;
assign w15721 = w15719 & ~w15720;
assign w15722 = ~w15716 & w15721;
assign w15723 = pi14 & w15722;
assign v4901 = ~(pi14 | w15722);
assign w15724 = v4901;
assign v4902 = ~(w15723 | w15724);
assign w15725 = v4902;
assign v4903 = ~(w15715 | w15725);
assign w15726 = v4903;
assign v4904 = ~(w15358 | w15360);
assign w15727 = v4904;
assign v4905 = ~(w15361 | w15727);
assign w15728 = v4905;
assign w15729 = w15715 & w15725;
assign v4906 = ~(w15726 | w15729);
assign w15730 = v4906;
assign w15731 = w15728 & w15730;
assign v4907 = ~(w15726 | w15731);
assign w15732 = v4907;
assign w15733 = ~w15408 & w15732;
assign w15734 = w15408 & ~w15732;
assign v4908 = ~(w15733 | w15734);
assign w15735 = v4908;
assign w15736 = w7178 & ~w12506;
assign w15737 = w7765 & ~w12406;
assign w15738 = w7466 & w12381;
assign v4909 = ~(w15737 | w15738);
assign w15739 = v4909;
assign w15740 = w7177 & w12311;
assign w15741 = w15739 & ~w15740;
assign w15742 = ~w15736 & w15741;
assign w15743 = pi11 & w15742;
assign v4910 = ~(pi11 | w15742);
assign w15744 = v4910;
assign v4911 = ~(w15743 | w15744);
assign w15745 = v4911;
assign w15746 = w15735 & w15745;
assign v4912 = ~(w15733 | w15746);
assign w15747 = v4912;
assign v4913 = ~(w15396 | w15405);
assign w15748 = v4913;
assign v4914 = ~(w15406 | w15748);
assign w15749 = v4914;
assign w15750 = w15747 & w15749;
assign v4915 = ~(w15406 | w15750);
assign w15751 = v4915;
assign w15752 = w15394 & ~w15751;
assign w15753 = w15711 & ~w15713;
assign v4916 = ~(w15714 | w15753);
assign w15754 = v4916;
assign w15755 = w6389 & w12167;
assign w15756 = w6388 & w11984;
assign w15757 = w7004 & w12155;
assign v4917 = ~(w15756 | w15757);
assign w15758 = v4917;
assign w15759 = w6871 & w12084;
assign w15760 = w15758 & ~w15759;
assign w15761 = ~w15755 & w15760;
assign w15762 = pi14 & w15761;
assign v4918 = ~(pi14 | w15761);
assign w15763 = v4918;
assign v4919 = ~(w15762 | w15763);
assign w15764 = v4919;
assign w15765 = w15754 & ~w15764;
assign w15766 = w15656 & ~w15658;
assign v4920 = ~(w15659 | w15766);
assign w15767 = v4920;
assign w15768 = w4764 & w13514;
assign w15769 = w4836 & w11720;
assign w15770 = w4913 & w11714;
assign v4921 = ~(w15769 | w15770);
assign w15771 = v4921;
assign w15772 = w4763 & w11723;
assign w15773 = w15771 & ~w15772;
assign w15774 = ~w15768 & w15773;
assign w15775 = pi23 & w15774;
assign v4922 = ~(pi23 | w15774);
assign w15776 = v4922;
assign v4923 = ~(w15775 | w15776);
assign w15777 = v4923;
assign w15778 = w15767 & ~w15777;
assign w15779 = w15652 & ~w15654;
assign v4924 = ~(w15655 | w15779);
assign w15780 = v4924;
assign w15781 = w4764 & ~w13310;
assign w15782 = w4913 & w11720;
assign w15783 = w4836 & w11723;
assign w15784 = w4763 & w11726;
assign v4925 = ~(w15783 | w15784);
assign w15785 = v4925;
assign w15786 = ~w15782 & w15785;
assign w15787 = ~w15781 & w15786;
assign w15788 = ~pi23 & w15787;
assign w15789 = pi23 & ~w15787;
assign v4926 = ~(w15788 | w15789);
assign w15790 = v4926;
assign w15791 = w15780 & w15790;
assign v4927 = ~(w15780 | w15790);
assign w15792 = v4927;
assign v4928 = ~(w15791 | w15792);
assign w15793 = v4928;
assign w15794 = w15648 & ~w15650;
assign v4929 = ~(w15651 | w15794);
assign w15795 = v4929;
assign w15796 = w4764 & ~w13737;
assign w15797 = w4913 & w11723;
assign w15798 = w4763 & w11729;
assign w15799 = w4836 & w11726;
assign v4930 = ~(w15798 | w15799);
assign w15800 = v4930;
assign w15801 = ~w15797 & w15800;
assign w15802 = ~w15796 & w15801;
assign w15803 = pi23 & ~w15802;
assign w15804 = ~pi23 & w15802;
assign v4931 = ~(w15803 | w15804);
assign w15805 = v4931;
assign w15806 = w15795 & w15805;
assign v4932 = ~(w15795 | w15805);
assign w15807 = v4932;
assign w15808 = w15644 & ~w15646;
assign v4933 = ~(w15647 | w15808);
assign w15809 = v4933;
assign w15810 = w4764 & w13864;
assign w15811 = w4836 & w11729;
assign w15812 = w4913 & w11726;
assign v4934 = ~(w15811 | w15812);
assign w15813 = v4934;
assign w15814 = w4763 & ~w11734;
assign w15815 = w15813 & ~w15814;
assign w15816 = ~w15810 & w15815;
assign w15817 = pi23 & w15816;
assign v4935 = ~(pi23 | w15816);
assign w15818 = v4935;
assign v4936 = ~(w15817 | w15818);
assign w15819 = v4936;
assign w15820 = w15809 & ~w15819;
assign w15821 = ~w15809 & w15819;
assign w15822 = w15640 & ~w15642;
assign v4937 = ~(w15643 | w15822);
assign w15823 = v4937;
assign w15824 = w4764 & ~w13703;
assign w15825 = w4913 & w11729;
assign w15826 = w4836 & ~w11734;
assign w15827 = w4763 & w11737;
assign v4938 = ~(w15826 | w15827);
assign w15828 = v4938;
assign w15829 = ~w15825 & w15828;
assign w15830 = ~w15824 & w15829;
assign w15831 = ~pi23 & w15830;
assign w15832 = pi23 & ~w15830;
assign v4939 = ~(w15831 | w15832);
assign w15833 = v4939;
assign v4940 = ~(w15823 | w15833);
assign w15834 = v4940;
assign w15835 = w15823 & w15833;
assign w15836 = w15636 & ~w15638;
assign v4941 = ~(w15639 | w15836);
assign w15837 = v4941;
assign w15838 = w4764 & w13882;
assign w15839 = w4836 & w11737;
assign w15840 = w4913 & ~w11734;
assign v4942 = ~(w15839 | w15840);
assign w15841 = v4942;
assign w15842 = w4763 & w11740;
assign w15843 = w15841 & ~w15842;
assign w15844 = ~w15838 & w15843;
assign w15845 = pi23 & w15844;
assign v4943 = ~(pi23 | w15844);
assign w15846 = v4943;
assign v4944 = ~(w15845 | w15846);
assign w15847 = v4944;
assign w15848 = w15837 & ~w15847;
assign w15849 = ~w15837 & w15847;
assign v4945 = ~(w15848 | w15849);
assign w15850 = v4945;
assign w15851 = w15632 & ~w15634;
assign v4946 = ~(w15635 | w15851);
assign w15852 = v4946;
assign w15853 = w4764 & w14288;
assign w15854 = w4913 & w11737;
assign w15855 = w4763 & ~w11745;
assign w15856 = w4836 & w11740;
assign v4947 = ~(w15855 | w15856);
assign w15857 = v4947;
assign w15858 = ~w15854 & w15857;
assign w15859 = ~w15853 & w15858;
assign w15860 = ~pi23 & w15859;
assign w15861 = pi23 & ~w15859;
assign v4948 = ~(w15860 | w15861);
assign w15862 = v4948;
assign v4949 = ~(w15852 | w15862);
assign w15863 = v4949;
assign w15864 = w15852 & w15862;
assign w15865 = w15628 & ~w15630;
assign v4950 = ~(w15631 | w15865);
assign w15866 = v4950;
assign w15867 = w4764 & w14300;
assign w15868 = w4836 & ~w11745;
assign w15869 = w4913 & w11740;
assign v4951 = ~(w15868 | w15869);
assign w15870 = v4951;
assign w15871 = w4763 & w11748;
assign w15872 = w15870 & ~w15871;
assign w15873 = ~w15867 & w15872;
assign w15874 = pi23 & w15873;
assign v4952 = ~(pi23 | w15873);
assign w15875 = v4952;
assign v4953 = ~(w15874 | w15875);
assign w15876 = v4953;
assign w15877 = w15866 & ~w15876;
assign w15878 = w15624 & ~w15626;
assign v4954 = ~(w15627 | w15878);
assign w15879 = v4954;
assign w15880 = w4764 & w13948;
assign w15881 = w4836 & w11748;
assign w15882 = w4913 & ~w11745;
assign v4955 = ~(w15881 | w15882);
assign w15883 = v4955;
assign w15884 = w4763 & w11759;
assign w15885 = w15883 & ~w15884;
assign w15886 = ~w15880 & w15885;
assign w15887 = pi23 & w15886;
assign v4956 = ~(pi23 | w15886);
assign w15888 = v4956;
assign v4957 = ~(w15887 | w15888);
assign w15889 = v4957;
assign w15890 = w15879 & ~w15889;
assign w15891 = w15620 & ~w15622;
assign v4958 = ~(w15623 | w15891);
assign w15892 = v4958;
assign w15893 = (w4764 & w11841) | (w4764 & w30627) | (w11841 & w30627);
assign w15894 = w4913 & w11748;
assign w15895 = w4836 & w11759;
assign w15896 = w4763 & w11761;
assign v4959 = ~(w15895 | w15896);
assign w15897 = v4959;
assign w15898 = ~w15894 & w15897;
assign w15899 = ~w15893 & w15898;
assign w15900 = pi23 & w15899;
assign v4960 = ~(pi23 | w15899);
assign w15901 = v4960;
assign v4961 = ~(w15900 | w15901);
assign w15902 = v4961;
assign w15903 = w15892 & ~w15902;
assign w15904 = w15616 & ~w15618;
assign v4962 = ~(w15619 | w15904);
assign w15905 = v4962;
assign w15906 = w4763 & ~w11771;
assign w15907 = w4913 & w11759;
assign v4963 = ~(w15906 | w15907);
assign w15908 = v4963;
assign w15909 = w4836 & w11761;
assign w15910 = w15908 & ~w15909;
assign w15911 = (~w14356 & w30628) | (~w14356 & w30629) | (w30628 & w30629);
assign w15912 = (w14356 & w30630) | (w14356 & w30631) | (w30630 & w30631);
assign v4964 = ~(w15911 | w15912);
assign w15913 = v4964;
assign w15914 = w15905 & ~w15913;
assign w15915 = w15612 & ~w15614;
assign v4965 = ~(w15615 | w15915);
assign w15916 = v4965;
assign w15917 = w4836 & ~w11771;
assign w15918 = w4913 & w11761;
assign w15919 = w4763 & w11768;
assign v4966 = ~(w15918 | w15919);
assign w15920 = v4966;
assign w15921 = ~w15917 & w15920;
assign w15922 = (w14383 & w30632) | (w14383 & w30633) | (w30632 & w30633);
assign w15923 = (~w14383 & w30634) | (~w14383 & w30635) | (w30634 & w30635);
assign v4967 = ~(w15922 | w15923);
assign w15924 = v4967;
assign w15925 = w15916 & w15924;
assign w15926 = w15608 & ~w15610;
assign v4968 = ~(w15611 | w15926);
assign w15927 = v4968;
assign w15928 = w4764 & w14409;
assign w15929 = w4836 & w11768;
assign w15930 = (w4913 & ~w11766) | (w4913 & w30507) | (~w11766 & w30507);
assign v4969 = ~(w15929 | w15930);
assign w15931 = v4969;
assign w15932 = w4763 & w11776;
assign w15933 = w15931 & ~w15932;
assign w15934 = ~w15928 & w30346;
assign w15935 = (w14409 & w30508) | (w14409 & w30509) | (w30508 & w30509);
assign v4970 = ~(w15934 | w15935);
assign w15936 = v4970;
assign w15937 = w15927 & ~w15936;
assign v4971 = ~(w15597 | w15606);
assign w15938 = v4971;
assign v4972 = ~(w15607 | w15938);
assign w15939 = v4972;
assign w15940 = w11533 & w30510;
assign w15941 = w4763 & w11784;
assign w15942 = w4836 & w11776;
assign v4973 = ~(w15941 | w15942);
assign w15943 = v4973;
assign w15944 = ~w15940 & w15943;
assign w15945 = (~w14461 & w30348) | (~w14461 & w30349) | (w30348 & w30349);
assign w15946 = (w14461 & w30350) | (w14461 & w30351) | (w30350 & w30351);
assign v4974 = ~(w15945 | w15946);
assign w15947 = v4974;
assign w15948 = w15939 & w15947;
assign w15949 = pi26 & ~w15586;
assign v4975 = ~(w15592 | w15949);
assign w15950 = v4975;
assign w15951 = w15592 & w15949;
assign v4976 = ~(w15950 | w15951);
assign w15952 = v4976;
assign w15953 = w4836 & w11784;
assign w15954 = w4913 & w11776;
assign v4977 = ~(w15953 | w15954);
assign w15955 = v4977;
assign w15956 = w4763 & w11793;
assign w15957 = (w14504 & w30171) | (w14504 & w30172) | (w30171 & w30172);
assign w15958 = (~w14504 & w30173) | (~w14504 & w30174) | (w30173 & w30174);
assign v4978 = ~(w15957 | w15958);
assign w15959 = v4978;
assign v4979 = ~(w15952 | w15959);
assign w15960 = v4979;
assign w15961 = w15580 & ~w15585;
assign v4980 = ~(w15586 | w15961);
assign w15962 = v4980;
assign w15963 = w4764 & w14547;
assign w15964 = w4763 & w11803;
assign w15965 = w4913 & w11784;
assign w15966 = w4836 & w11793;
assign v4981 = ~(w15965 | w15966);
assign w15967 = v4981;
assign w15968 = (pi23 & w15963) | (pi23 & w30035) | (w15963 & w30035);
assign w15969 = ~w15963 & w30036;
assign v4982 = ~(w15968 | w15969);
assign w15970 = v4982;
assign w15971 = w15962 & w15970;
assign w15972 = w10 & w11800;
assign w15973 = pi23 & w15972;
assign w15974 = w4764 & ~w14609;
assign w15975 = w4913 & w11798;
assign w15976 = w4836 & w11800;
assign v4983 = ~(w15975 | w15976);
assign w15977 = v4983;
assign w15978 = ~w15974 & w15977;
assign w15979 = ~w15973 & w15978;
assign w15980 = w4763 & w11800;
assign w15981 = (~w15980 & w14639) | (~w15980 & w30511) | (w14639 & w30511);
assign w15982 = w4913 & w11803;
assign w15983 = w4836 & w11798;
assign v4984 = ~(w15982 | w15983);
assign w15984 = v4984;
assign w15985 = w15981 & w15984;
assign w15986 = pi23 & w15985;
assign w15987 = w15979 & w15986;
assign w15988 = w15579 & w15987;
assign v4985 = ~(w15579 | w15987);
assign w15989 = v4985;
assign v4986 = ~(w15988 | w15989);
assign w15990 = v4986;
assign w15991 = w4763 & w11798;
assign w15992 = ~w11792 & w30512;
assign w15993 = w4836 & w11803;
assign v4987 = ~(w15992 | w15993);
assign w15994 = v4987;
assign w15995 = ~w15991 & w15994;
assign w15996 = (w15995 & ~w14569) | (w15995 & w30352) | (~w14569 & w30352);
assign w15997 = pi23 & ~w15996;
assign w15998 = ~pi23 & w15996;
assign v4988 = ~(w15997 | w15998);
assign w15999 = v4988;
assign w16000 = w15990 & w15999;
assign v4989 = ~(w15988 | w16000);
assign w16001 = v4989;
assign v4990 = ~(w15962 | w15970);
assign w16002 = v4990;
assign v4991 = ~(w15971 | w16002);
assign w16003 = v4991;
assign w16004 = ~w16001 & w16003;
assign w16005 = (~w15971 & ~w16003) | (~w15971 & w30175) | (~w16003 & w30175);
assign w16006 = w15952 & w15959;
assign v4992 = ~(w15960 | w16006);
assign w16007 = v4992;
assign w16008 = ~w16005 & w16007;
assign v4993 = ~(w15960 | w16008);
assign w16009 = v4993;
assign v4994 = ~(w15939 | w15947);
assign w16010 = v4994;
assign v4995 = ~(w15948 | w16010);
assign w16011 = v4995;
assign w16012 = ~w16009 & w16011;
assign w16013 = (~w15948 & w16009) | (~w15948 & w30353) | (w16009 & w30353);
assign w16014 = ~w15927 & w15936;
assign v4996 = ~(w15937 | w16014);
assign w16015 = v4996;
assign w16016 = ~w16013 & w16015;
assign w16017 = (~w15937 & w16013) | (~w15937 & w30811) | (w16013 & w30811);
assign v4997 = ~(w15916 | w15924);
assign w16018 = v4997;
assign v4998 = ~(w15925 | w16018);
assign w16019 = v4998;
assign w16020 = ~w16017 & w16019;
assign w16021 = (~w15925 & w16017) | (~w15925 & w30513) | (w16017 & w30513);
assign w16022 = ~w15905 & w15913;
assign v4999 = ~(w15914 | w16022);
assign w16023 = v4999;
assign w16024 = ~w16021 & w16023;
assign v5000 = ~(w15914 | w16024);
assign w16025 = v5000;
assign w16026 = ~w15892 & w15902;
assign v5001 = ~(w15903 | w16026);
assign w16027 = v5001;
assign w16028 = ~w16025 & w16027;
assign w16029 = (~w15903 & w16025) | (~w15903 & w30636) | (w16025 & w30636);
assign w16030 = ~w15879 & w15889;
assign v5002 = ~(w15890 | w16030);
assign w16031 = v5002;
assign w16032 = ~w16029 & w16031;
assign w16033 = (~w15890 & w16029) | (~w15890 & w30812) | (w16029 & w30812);
assign w16034 = ~w15866 & w15876;
assign v5003 = ~(w15877 | w16034);
assign w16035 = v5003;
assign w16036 = ~w16033 & w16035;
assign w16037 = (~w15877 & w16033) | (~w15877 & w31045) | (w16033 & w31045);
assign w16038 = (~w15863 & ~w16037) | (~w15863 & w31192) | (~w16037 & w31192);
assign w16039 = w15850 & w16038;
assign v5004 = ~(w15848 | w16039);
assign w16040 = v5004;
assign w16041 = ~w16039 & w31278;
assign v5005 = ~(w15834 | w16041);
assign w16042 = v5005;
assign w16043 = ~w15821 & w16042;
assign v5006 = ~(w15820 | w16043);
assign w16044 = v5006;
assign v5007 = ~(w15807 | w16044);
assign w16045 = v5007;
assign v5008 = ~(w15806 | w16045);
assign w16046 = v5008;
assign w16047 = w15793 & ~w16046;
assign v5009 = ~(w15791 | w16047);
assign w16048 = v5009;
assign w16049 = ~w15767 & w15777;
assign v5010 = ~(w15778 | w16049);
assign w16050 = v5010;
assign w16051 = ~w16048 & w16050;
assign v5011 = ~(w15778 | w16051);
assign w16052 = v5011;
assign w16053 = w15673 & ~w15675;
assign v5012 = ~(w15676 | w16053);
assign w16054 = v5012;
assign w16055 = w16052 & w16054;
assign v5013 = ~(w16052 | w16054);
assign w16056 = v5013;
assign v5014 = ~(w16055 | w16056);
assign w16057 = v5014;
assign w16058 = w5114 & ~w13008;
assign w16059 = w5610 & ~w11695;
assign w16060 = w5531 & w11700;
assign w16061 = w5113 & w11708;
assign v5015 = ~(w16060 | w16061);
assign w16062 = v5015;
assign w16063 = ~w16059 & w16062;
assign w16064 = ~w16058 & w16063;
assign w16065 = ~pi20 & w16064;
assign w16066 = pi20 & ~w16064;
assign v5016 = ~(w16065 | w16066);
assign w16067 = v5016;
assign w16068 = w16057 & ~w16067;
assign v5017 = ~(w16055 | w16068);
assign w16069 = v5017;
assign w16070 = w5765 & w12594;
assign w16071 = w6236 & w11678;
assign w16072 = w5983 & ~w11683;
assign w16073 = w5764 & w11686;
assign v5018 = ~(w16072 | w16073);
assign w16074 = v5018;
assign w16075 = ~w16071 & w16074;
assign w16076 = ~w16070 & w16075;
assign w16077 = pi17 & w16076;
assign v5019 = ~(pi17 | w16076);
assign w16078 = v5019;
assign v5020 = ~(w16077 | w16078);
assign w16079 = v5020;
assign w16080 = w16069 & ~w16079;
assign w16081 = w15690 & ~w15692;
assign v5021 = ~(w15693 | w16081);
assign w16082 = v5021;
assign w16083 = ~w16069 & w16079;
assign v5022 = ~(w16080 | w16083);
assign w16084 = v5022;
assign w16085 = ~w16082 & w16084;
assign v5023 = ~(w16080 | w16085);
assign w16086 = v5023;
assign w16087 = w6389 & w12181;
assign w16088 = w6871 & w11984;
assign w16089 = w7004 & w12084;
assign v5024 = ~(w16088 | w16089);
assign w16090 = v5024;
assign w16091 = w6388 & w11671;
assign w16092 = w16090 & ~w16091;
assign w16093 = ~w16087 & w16092;
assign w16094 = pi14 & w16093;
assign v5025 = ~(pi14 | w16093);
assign w16095 = v5025;
assign v5026 = ~(w16094 | w16095);
assign w16096 = v5026;
assign w16097 = w16086 & w16096;
assign w16098 = w15707 & ~w15709;
assign v5027 = ~(w15710 | w16098);
assign w16099 = v5027;
assign v5028 = ~(w16086 | w16096);
assign w16100 = v5028;
assign v5029 = ~(w16097 | w16100);
assign w16101 = v5029;
assign w16102 = ~w16099 & w16101;
assign v5030 = ~(w16097 | w16102);
assign w16103 = v5030;
assign w16104 = ~w15754 & w15764;
assign v5031 = ~(w15765 | w16104);
assign w16105 = v5031;
assign w16106 = w16103 & w16105;
assign v5032 = ~(w15765 | w16106);
assign w16107 = v5032;
assign w16108 = w7178 & w12387;
assign w16109 = w7765 & w12381;
assign w16110 = w7177 & w12271;
assign w16111 = w7466 & w12311;
assign v5033 = ~(w16110 | w16111);
assign w16112 = v5033;
assign w16113 = ~w16109 & w16112;
assign w16114 = ~w16108 & w16113;
assign w16115 = ~pi11 & w16114;
assign w16116 = pi11 & ~w16114;
assign v5034 = ~(w16115 | w16116);
assign w16117 = v5034;
assign w16118 = ~w16107 & w16117;
assign v5035 = ~(w15728 | w15730);
assign w16119 = v5035;
assign v5036 = ~(w15731 | w16119);
assign w16120 = v5036;
assign w16121 = w16107 & ~w16117;
assign v5037 = ~(w16118 | w16121);
assign w16122 = v5037;
assign w16123 = w16120 & w16122;
assign v5038 = ~(w16118 | w16123);
assign w16124 = v5038;
assign w16125 = w13301 & ~w16124;
assign w16126 = ~w13301 & w16124;
assign v5039 = ~(w16125 | w16126);
assign w16127 = v5039;
assign v5040 = ~(w15735 | w15745);
assign w16128 = v5040;
assign v5041 = ~(w15746 | w16128);
assign w16129 = v5041;
assign w16130 = w16127 & ~w16129;
assign v5042 = ~(w16125 | w16130);
assign w16131 = v5042;
assign v5043 = ~(w15747 | w15749);
assign w16132 = v5043;
assign v5044 = ~(w15750 | w16132);
assign w16133 = v5044;
assign w16134 = ~w16131 & w16133;
assign w16135 = w16131 & ~w16133;
assign v5045 = ~(w16134 | w16135);
assign w16136 = v5045;
assign w16137 = ~w16127 & w16129;
assign v5046 = ~(w16130 | w16137);
assign w16138 = v5046;
assign v5047 = ~(w16103 | w16105);
assign w16139 = v5047;
assign v5048 = ~(w16106 | w16139);
assign w16140 = v5048;
assign w16141 = w7178 & w12318;
assign w16142 = w7466 & w12271;
assign w16143 = w7765 & w12311;
assign v5049 = ~(w16142 | w16143);
assign w16144 = v5049;
assign w16145 = w7177 & w12237;
assign w16146 = w16144 & ~w16145;
assign w16147 = ~w16141 & w16146;
assign w16148 = pi11 & w16147;
assign v5050 = ~(pi11 | w16147);
assign w16149 = v5050;
assign v5051 = ~(w16148 | w16149);
assign w16150 = v5051;
assign w16151 = w16140 & ~w16150;
assign w16152 = w16048 & ~w16050;
assign v5052 = ~(w16051 | w16152);
assign w16153 = v5052;
assign w16154 = w5114 & w12994;
assign w16155 = w5610 & w11700;
assign w16156 = w5113 & w11711;
assign w16157 = w5531 & w11708;
assign v5053 = ~(w16156 | w16157);
assign w16158 = v5053;
assign w16159 = ~w16155 & w16158;
assign w16160 = ~w16154 & w16159;
assign w16161 = pi20 & ~w16160;
assign w16162 = ~pi20 & w16160;
assign v5054 = ~(w16161 | w16162);
assign w16163 = v5054;
assign w16164 = w16153 & w16163;
assign w16165 = ~w15793 & w16046;
assign v5055 = ~(w16047 | w16165);
assign w16166 = v5055;
assign w16167 = w5114 & w13178;
assign w16168 = w5610 & w11708;
assign w16169 = w5113 & w11714;
assign w16170 = w5531 & w11711;
assign v5056 = ~(w16169 | w16170);
assign w16171 = v5056;
assign w16172 = ~w16168 & w16171;
assign w16173 = ~w16167 & w16172;
assign w16174 = ~pi20 & w16173;
assign w16175 = pi20 & ~w16173;
assign v5057 = ~(w16174 | w16175);
assign w16176 = v5057;
assign w16177 = w16166 & w16176;
assign v5058 = ~(w16166 | w16176);
assign w16178 = v5058;
assign v5059 = ~(w16177 | w16178);
assign w16179 = v5059;
assign w16180 = w5114 & w13194;
assign w16181 = w5610 & w11711;
assign w16182 = w5531 & w11714;
assign w16183 = w5113 & w11720;
assign v5060 = ~(w16182 | w16183);
assign w16184 = v5060;
assign w16185 = ~w16181 & w16184;
assign w16186 = ~w16180 & w16185;
assign w16187 = ~pi20 & w16186;
assign w16188 = pi20 & ~w16186;
assign v5061 = ~(w16187 | w16188);
assign w16189 = v5061;
assign v5062 = ~(w15806 | w15807);
assign w16190 = v5062;
assign w16191 = w16044 & ~w16190;
assign w16192 = ~w16044 & w16190;
assign v5063 = ~(w16191 | w16192);
assign w16193 = v5063;
assign v5064 = ~(w16189 | w16193);
assign w16194 = v5064;
assign w16195 = w16189 & w16193;
assign v5065 = ~(w15820 | w15821);
assign w16196 = v5065;
assign v5066 = ~(w16042 | w16196);
assign w16197 = v5066;
assign w16198 = w16042 & w16196;
assign v5067 = ~(w16197 | w16198);
assign w16199 = v5067;
assign w16200 = w5114 & w13514;
assign w16201 = w5531 & w11720;
assign w16202 = w5610 & w11714;
assign v5068 = ~(w16201 | w16202);
assign w16203 = v5068;
assign w16204 = w5113 & w11723;
assign w16205 = w16203 & ~w16204;
assign w16206 = ~w16200 & w16205;
assign w16207 = pi20 & w16206;
assign v5069 = ~(pi20 | w16206);
assign w16208 = v5069;
assign v5070 = ~(w16207 | w16208);
assign w16209 = v5070;
assign w16210 = ~w16199 & w16209;
assign w16211 = w5114 & ~w13310;
assign w16212 = w5610 & w11720;
assign w16213 = w5531 & w11723;
assign w16214 = w5113 & w11726;
assign v5071 = ~(w16213 | w16214);
assign w16215 = v5071;
assign w16216 = ~w16212 & w16215;
assign w16217 = ~w16211 & w16216;
assign w16218 = ~pi20 & w16217;
assign w16219 = pi20 & ~w16217;
assign v5072 = ~(w16218 | w16219);
assign w16220 = v5072;
assign v5073 = ~(w15834 | w15835);
assign w16221 = v5073;
assign w16222 = w16040 & w16221;
assign v5074 = ~(w16040 | w16221);
assign w16223 = v5074;
assign v5075 = ~(w16222 | w16223);
assign w16224 = v5075;
assign w16225 = w16220 & ~w16224;
assign w16226 = ~w16220 & w16224;
assign v5076 = ~(w16225 | w16226);
assign w16227 = v5076;
assign v5077 = ~(w15850 | w16038);
assign w16228 = v5077;
assign v5078 = ~(w16039 | w16228);
assign w16229 = v5078;
assign w16230 = w5114 & ~w13737;
assign w16231 = w5610 & w11723;
assign w16232 = w5113 & w11729;
assign w16233 = w5531 & w11726;
assign v5079 = ~(w16232 | w16233);
assign w16234 = v5079;
assign w16235 = ~w16231 & w16234;
assign w16236 = ~w16230 & w16235;
assign w16237 = pi20 & ~w16236;
assign w16238 = ~pi20 & w16236;
assign v5080 = ~(w16237 | w16238);
assign w16239 = v5080;
assign v5081 = ~(w16229 | w16239);
assign w16240 = v5081;
assign w16241 = w16229 & w16239;
assign w16242 = w5114 & w13864;
assign w16243 = w5531 & w11729;
assign w16244 = w5610 & w11726;
assign v5082 = ~(w16243 | w16244);
assign w16245 = v5082;
assign w16246 = w5113 & ~w11734;
assign w16247 = w16245 & ~w16246;
assign w16248 = ~w16242 & w16247;
assign w16249 = pi20 & w16248;
assign v5083 = ~(pi20 | w16248);
assign w16250 = v5083;
assign v5084 = ~(w16249 | w16250);
assign w16251 = v5084;
assign v5085 = ~(w15863 | w15864);
assign w16252 = v5085;
assign w16253 = w16037 & w16252;
assign v5086 = ~(w16037 | w16252);
assign w16254 = v5086;
assign v5087 = ~(w16253 | w16254);
assign w16255 = v5087;
assign v5088 = ~(w16251 | w16255);
assign w16256 = v5088;
assign w16257 = w16251 & w16255;
assign v5089 = ~(w16256 | w16257);
assign w16258 = v5089;
assign w16259 = w16033 & ~w16035;
assign v5090 = ~(w16036 | w16259);
assign w16260 = v5090;
assign w16261 = w5114 & ~w13703;
assign w16262 = w5610 & w11729;
assign w16263 = w5531 & ~w11734;
assign w16264 = w5113 & w11737;
assign v5091 = ~(w16263 | w16264);
assign w16265 = v5091;
assign w16266 = ~w16262 & w16265;
assign w16267 = ~w16261 & w16266;
assign w16268 = pi20 & w16267;
assign v5092 = ~(pi20 | w16267);
assign w16269 = v5092;
assign v5093 = ~(w16268 | w16269);
assign w16270 = v5093;
assign w16271 = ~w16260 & w16270;
assign w16272 = w16260 & ~w16270;
assign w16273 = w16029 & ~w16031;
assign v5094 = ~(w16032 | w16273);
assign w16274 = v5094;
assign w16275 = w5114 & w13882;
assign w16276 = w5610 & ~w11734;
assign w16277 = w5531 & w11737;
assign w16278 = w5113 & w11740;
assign v5095 = ~(w16277 | w16278);
assign w16279 = v5095;
assign w16280 = ~w16276 & w16279;
assign w16281 = ~w16275 & w16280;
assign w16282 = ~pi20 & w16281;
assign w16283 = pi20 & ~w16281;
assign v5096 = ~(w16282 | w16283);
assign w16284 = v5096;
assign w16285 = w16274 & w16284;
assign v5097 = ~(w16274 | w16284);
assign w16286 = v5097;
assign v5098 = ~(w16285 | w16286);
assign w16287 = v5098;
assign w16288 = w16025 & ~w16027;
assign v5099 = ~(w16028 | w16288);
assign w16289 = v5099;
assign w16290 = w5114 & w14288;
assign w16291 = w5610 & w11737;
assign w16292 = w5113 & ~w11745;
assign w16293 = w5531 & w11740;
assign v5100 = ~(w16292 | w16293);
assign w16294 = v5100;
assign w16295 = ~w16291 & w16294;
assign w16296 = ~w16290 & w16295;
assign w16297 = pi20 & ~w16296;
assign w16298 = ~pi20 & w16296;
assign v5101 = ~(w16297 | w16298);
assign w16299 = v5101;
assign v5102 = ~(w16289 | w16299);
assign w16300 = v5102;
assign w16301 = w16289 & w16299;
assign w16302 = w16021 & ~w16023;
assign v5103 = ~(w16024 | w16302);
assign w16303 = v5103;
assign w16304 = w5610 & w11740;
assign w16305 = w5531 & ~w11745;
assign w16306 = w5113 & w11748;
assign v5104 = ~(w16305 | w16306);
assign w16307 = v5104;
assign w16308 = ~w16304 & w16307;
assign w16309 = (w16308 & ~w14300) | (w16308 & w30637) | (~w14300 & w30637);
assign w16310 = ~pi20 & w16309;
assign w16311 = pi20 & ~w16309;
assign v5105 = ~(w16310 | w16311);
assign w16312 = v5105;
assign w16313 = w16303 & w16312;
assign w16314 = w16017 & ~w16019;
assign v5106 = ~(w16020 | w16314);
assign w16315 = v5106;
assign w16316 = w5610 & ~w11745;
assign w16317 = w5531 & w11748;
assign w16318 = w5113 & w11759;
assign v5107 = ~(w16317 | w16318);
assign w16319 = v5107;
assign w16320 = ~w16316 & w16319;
assign w16321 = (w16320 & ~w13948) | (w16320 & w30514) | (~w13948 & w30514);
assign w16322 = pi20 & w16321;
assign v5108 = ~(pi20 | w16321);
assign w16323 = v5108;
assign v5109 = ~(w16322 | w16323);
assign w16324 = v5109;
assign w16325 = w16315 & ~w16324;
assign w16326 = w16013 & ~w16015;
assign v5110 = ~(w16016 | w16326);
assign w16327 = v5110;
assign w16328 = (w5114 & w11841) | (w5114 & w30354) | (w11841 & w30354);
assign w16329 = w5610 & w11748;
assign w16330 = w5531 & w11759;
assign w16331 = w5113 & w11761;
assign v5111 = ~(w16330 | w16331);
assign w16332 = v5111;
assign w16333 = ~w16329 & w16332;
assign w16334 = ~w16328 & w30515;
assign w16335 = (pi20 & w16328) | (pi20 & w30516) | (w16328 & w30516);
assign v5112 = ~(w16334 | w16335);
assign w16336 = v5112;
assign w16337 = w16327 & w16336;
assign w16338 = w16009 & ~w16011;
assign v5113 = ~(w16012 | w16338);
assign w16339 = v5113;
assign w16340 = w5113 & ~w11771;
assign w16341 = w5610 & w11759;
assign w16342 = w5531 & w11761;
assign v5114 = ~(w16341 | w16342);
assign w16343 = v5114;
assign w16344 = ~w16340 & w16343;
assign w16345 = (w14356 & w30355) | (w14356 & w30356) | (w30355 & w30356);
assign w16346 = (~w14356 & w30357) | (~w14356 & w30358) | (w30357 & w30358);
assign v5115 = ~(w16345 | w16346);
assign w16347 = v5115;
assign w16348 = w16339 & w16347;
assign w16349 = w16005 & ~w16007;
assign v5116 = ~(w16008 | w16349);
assign w16350 = v5116;
assign w16351 = w5531 & ~w11771;
assign w16352 = w5610 & w11761;
assign w16353 = w5113 & w11768;
assign v5117 = ~(w16352 | w16353);
assign w16354 = v5117;
assign w16355 = ~w16351 & w16354;
assign w16356 = (w14383 & w30359) | (w14383 & w30360) | (w30359 & w30360);
assign w16357 = (~w14383 & w30361) | (~w14383 & w30362) | (w30361 & w30362);
assign v5118 = ~(w16356 | w16357);
assign w16358 = v5118;
assign w16359 = w16350 & w16358;
assign w16360 = w16001 & ~w16003;
assign v5119 = ~(w16004 | w16360);
assign w16361 = v5119;
assign w16362 = w5114 & w14409;
assign w16363 = w5531 & w11768;
assign w16364 = (w5610 & ~w11766) | (w5610 & w30178) | (~w11766 & w30178);
assign v5120 = ~(w16363 | w16364);
assign w16365 = v5120;
assign w16366 = w5113 & w11776;
assign w16367 = w16365 & ~w16366;
assign w16368 = ~w16362 & w30037;
assign w16369 = (w14409 & w30179) | (w14409 & w30180) | (w30179 & w30180);
assign v5121 = ~(w16368 | w16369);
assign w16370 = v5121;
assign w16371 = w16361 & ~w16370;
assign v5122 = ~(w15990 | w15999);
assign w16372 = v5122;
assign v5123 = ~(w16000 | w16372);
assign w16373 = v5123;
assign w16374 = w11533 & w30181;
assign w16375 = w5113 & w11784;
assign w16376 = w5531 & w11776;
assign v5124 = ~(w16375 | w16376);
assign w16377 = v5124;
assign w16378 = ~w16374 & w16377;
assign w16379 = (~w14461 & w30039) | (~w14461 & w30040) | (w30039 & w30040);
assign w16380 = (w14461 & w30041) | (w14461 & w30042) | (w30041 & w30042);
assign v5125 = ~(w16379 | w16380);
assign w16381 = v5125;
assign w16382 = w16373 & w16381;
assign w16383 = pi23 & ~w15979;
assign v5126 = ~(w15985 | w16383);
assign w16384 = v5126;
assign w16385 = w15985 & w16383;
assign v5127 = ~(w16384 | w16385);
assign w16386 = v5127;
assign w16387 = w5531 & w11784;
assign w16388 = w5610 & w11776;
assign v5128 = ~(w16387 | w16388);
assign w16389 = v5128;
assign w16390 = w5113 & w11793;
assign w16391 = (w14504 & w29864) | (w14504 & w29865) | (w29864 & w29865);
assign w16392 = (~w14504 & w29866) | (~w14504 & w29867) | (w29866 & w29867);
assign v5129 = ~(w16391 | w16392);
assign w16393 = v5129;
assign v5130 = ~(w16386 | w16393);
assign w16394 = v5130;
assign w16395 = w15973 & ~w15978;
assign v5131 = ~(w15979 | w16395);
assign w16396 = v5131;
assign w16397 = w5114 & w14547;
assign w16398 = w5113 & w11803;
assign w16399 = (~w11781 & w29868) | (~w11781 & w29869) | (w29868 & w29869);
assign w16400 = w5531 & w11793;
assign v5132 = ~(w16399 | w16400);
assign w16401 = v5132;
assign w16402 = ~w16398 & w16401;
assign w16403 = (pi20 & w16397) | (pi20 & w29719) | (w16397 & w29719);
assign w16404 = ~w16397 & w29720;
assign v5133 = ~(w16403 | w16404);
assign w16405 = v5133;
assign w16406 = w16396 & w16405;
assign w16407 = w912 & w11800;
assign w16408 = pi20 & w16407;
assign w16409 = w5114 & ~w14609;
assign w16410 = w5610 & w11798;
assign w16411 = w5531 & w11800;
assign v5134 = ~(w16410 | w16411);
assign w16412 = v5134;
assign w16413 = ~w16409 & w16412;
assign w16414 = ~w16408 & w16413;
assign w16415 = w5113 & w11800;
assign w16416 = (~w16415 & w14639) | (~w16415 & w30517) | (w14639 & w30517);
assign w16417 = w5610 & w11803;
assign w16418 = w5531 & w11798;
assign v5135 = ~(w16417 | w16418);
assign w16419 = v5135;
assign w16420 = w16416 & w16419;
assign w16421 = pi20 & w16420;
assign w16422 = w16414 & w16421;
assign w16423 = w15972 & w16422;
assign v5136 = ~(w15972 | w16422);
assign w16424 = v5136;
assign v5137 = ~(w16423 | w16424);
assign w16425 = v5137;
assign w16426 = w5113 & w11798;
assign w16427 = ~w11792 & w30518;
assign w16428 = w5531 & w11803;
assign v5138 = ~(w16427 | w16428);
assign w16429 = v5138;
assign w16430 = ~w16426 & w16429;
assign w16431 = (w16430 & ~w14569) | (w16430 & w30043) | (~w14569 & w30043);
assign w16432 = pi20 & ~w16431;
assign w16433 = ~pi20 & w16431;
assign v5139 = ~(w16432 | w16433);
assign w16434 = v5139;
assign w16435 = w16425 & w16434;
assign v5140 = ~(w16423 | w16435);
assign w16436 = v5140;
assign v5141 = ~(w16396 | w16405);
assign w16437 = v5141;
assign v5142 = ~(w16406 | w16437);
assign w16438 = v5142;
assign w16439 = ~w16436 & w16438;
assign w16440 = (~w16406 & ~w16438) | (~w16406 & w29870) | (~w16438 & w29870);
assign w16441 = w16386 & w16393;
assign v5143 = ~(w16394 | w16441);
assign w16442 = v5143;
assign w16443 = ~w16440 & w16442;
assign v5144 = ~(w16394 | w16443);
assign w16444 = v5144;
assign v5145 = ~(w16373 | w16381);
assign w16445 = v5145;
assign v5146 = ~(w16382 | w16445);
assign w16446 = v5146;
assign w16447 = ~w16444 & w16446;
assign w16448 = (~w16382 & w16444) | (~w16382 & w30044) | (w16444 & w30044);
assign w16449 = ~w16361 & w16370;
assign v5147 = ~(w16371 | w16449);
assign w16450 = v5147;
assign w16451 = ~w16448 & w16450;
assign w16452 = (~w16371 & w16448) | (~w16371 & w30813) | (w16448 & w30813);
assign v5148 = ~(w16350 | w16358);
assign w16453 = v5148;
assign v5149 = ~(w16359 | w16453);
assign w16454 = v5149;
assign w16455 = ~w16452 & w16454;
assign w16456 = (~w16359 & w16452) | (~w16359 & w30182) | (w16452 & w30182);
assign v5150 = ~(w16339 | w16347);
assign w16457 = v5150;
assign v5151 = ~(w16348 | w16457);
assign w16458 = v5151;
assign w16459 = ~w16456 & w16458;
assign v5152 = ~(w16348 | w16459);
assign w16460 = v5152;
assign v5153 = ~(w16327 | w16336);
assign w16461 = v5153;
assign v5154 = ~(w16337 | w16461);
assign w16462 = v5154;
assign w16463 = ~w16460 & w16462;
assign w16464 = (~w16337 & w16460) | (~w16337 & w30363) | (w16460 & w30363);
assign w16465 = ~w16315 & w16324;
assign v5155 = ~(w16325 | w16465);
assign w16466 = v5155;
assign w16467 = ~w16464 & w16466;
assign w16468 = (~w16325 & w16464) | (~w16325 & w30814) | (w16464 & w30814);
assign v5156 = ~(w16303 | w16312);
assign w16469 = v5156;
assign v5157 = ~(w16313 | w16469);
assign w16470 = v5157;
assign w16471 = ~w16468 & w16470;
assign w16472 = (~w16313 & w16468) | (~w16313 & w30519) | (w16468 & w30519);
assign w16473 = (~w16300 & ~w16472) | (~w16300 & w30638) | (~w16472 & w30638);
assign w16474 = w16287 & w16473;
assign w16475 = (~w16285 & ~w16287) | (~w16285 & w30815) | (~w16287 & w30815);
assign w16476 = (~w16271 & ~w16475) | (~w16271 & w31046) | (~w16475 & w31046);
assign w16477 = w16258 & w16476;
assign v5158 = ~(w16256 | w16477);
assign w16478 = v5158;
assign w16479 = ~w16477 & w31193;
assign v5159 = ~(w16240 | w16479);
assign w16480 = v5159;
assign w16481 = w16227 & w16480;
assign v5160 = ~(w16225 | w16481);
assign w16482 = v5160;
assign w16483 = w16199 & ~w16209;
assign v5161 = ~(w16210 | w16483);
assign w16484 = v5161;
assign w16485 = w16482 & w16484;
assign v5162 = ~(w16210 | w16485);
assign w16486 = v5162;
assign v5163 = ~(w16195 | w16486);
assign w16487 = v5163;
assign v5164 = ~(w16194 | w16487);
assign w16488 = v5164;
assign w16489 = w16179 & w16488;
assign v5165 = ~(w16177 | w16489);
assign w16490 = v5165;
assign v5166 = ~(w16153 | w16163);
assign w16491 = v5166;
assign v5167 = ~(w16164 | w16491);
assign w16492 = v5167;
assign w16493 = ~w16490 & w16492;
assign v5168 = ~(w16164 | w16493);
assign w16494 = v5168;
assign w16495 = w5765 & w12610;
assign w16496 = w6236 & ~w11683;
assign w16497 = w5983 & w11686;
assign w16498 = w5764 & w11689;
assign v5169 = ~(w16497 | w16498);
assign w16499 = v5169;
assign w16500 = ~w16496 & w16499;
assign w16501 = ~w16495 & w16500;
assign w16502 = ~pi17 & w16501;
assign w16503 = pi17 & ~w16501;
assign v5170 = ~(w16502 | w16503);
assign w16504 = v5170;
assign w16505 = w16494 & ~w16504;
assign w16506 = ~w16057 & w16067;
assign v5171 = ~(w16068 | w16506);
assign w16507 = v5171;
assign w16508 = ~w16494 & w16504;
assign v5172 = ~(w16505 | w16508);
assign w16509 = v5172;
assign w16510 = w16507 & w16509;
assign v5173 = ~(w16505 | w16510);
assign w16511 = v5173;
assign w16512 = w6389 & w11993;
assign w16513 = w7004 & w11984;
assign w16514 = w6388 & w11673;
assign w16515 = w6871 & w11671;
assign v5174 = ~(w16514 | w16515);
assign w16516 = v5174;
assign w16517 = ~w16513 & w16516;
assign w16518 = ~w16512 & w16517;
assign w16519 = ~pi14 & w16518;
assign w16520 = pi14 & ~w16518;
assign v5175 = ~(w16519 | w16520);
assign w16521 = v5175;
assign v5176 = ~(w16511 | w16521);
assign w16522 = v5176;
assign w16523 = w16082 & ~w16084;
assign v5177 = ~(w16085 | w16523);
assign w16524 = v5177;
assign w16525 = w16511 & w16521;
assign v5178 = ~(w16522 | w16525);
assign w16526 = v5178;
assign w16527 = ~w16524 & w16526;
assign v5179 = ~(w16522 | w16527);
assign w16528 = v5179;
assign w16529 = w7178 & ~w12277;
assign w16530 = w7765 & w12271;
assign w16531 = w7177 & w12155;
assign w16532 = w7466 & w12237;
assign v5180 = ~(w16531 | w16532);
assign w16533 = v5180;
assign w16534 = ~w16530 & w16533;
assign w16535 = ~w16529 & w16534;
assign w16536 = pi11 & w16535;
assign v5181 = ~(pi11 | w16535);
assign w16537 = v5181;
assign v5182 = ~(w16536 | w16537);
assign w16538 = v5182;
assign w16539 = w16528 & ~w16538;
assign w16540 = w16099 & ~w16101;
assign v5183 = ~(w16102 | w16540);
assign w16541 = v5183;
assign w16542 = ~w16528 & w16538;
assign v5184 = ~(w16539 | w16542);
assign w16543 = v5184;
assign w16544 = ~w16541 & w16543;
assign v5185 = ~(w16539 | w16544);
assign w16545 = v5185;
assign w16546 = ~w16140 & w16150;
assign v5186 = ~(w16151 | w16546);
assign w16547 = v5186;
assign w16548 = ~w16545 & w16547;
assign v5187 = ~(w16151 | w16548);
assign w16549 = v5187;
assign w16550 = pi08 & w12406;
assign w16551 = pi07 & ~w12406;
assign v5188 = ~(w16550 | w16551);
assign w16552 = v5188;
assign w16553 = w8139 & w16552;
assign v5189 = ~(w13299 | w16553);
assign w16554 = v5189;
assign w16555 = ~w16549 & w16554;
assign w16556 = w16549 & ~w16554;
assign v5190 = ~(w16555 | w16556);
assign w16557 = v5190;
assign v5191 = ~(w16120 | w16122);
assign w16558 = v5191;
assign v5192 = ~(w16123 | w16558);
assign w16559 = v5192;
assign w16560 = w16557 & w16559;
assign v5193 = ~(w16555 | w16560);
assign w16561 = v5193;
assign w16562 = ~w16138 & w16561;
assign w16563 = w16541 & ~w16543;
assign v5194 = ~(w16544 | w16563);
assign w16564 = v5194;
assign w16565 = w8141 & ~w12506;
assign w16566 = w8926 & ~w12406;
assign w16567 = w8140 & w12311;
assign w16568 = w8526 & w12381;
assign v5195 = ~(w16567 | w16568);
assign w16569 = v5195;
assign w16570 = ~w16566 & w16569;
assign w16571 = ~w16565 & w16570;
assign w16572 = pi08 & ~w16571;
assign w16573 = ~pi08 & w16571;
assign v5196 = ~(w16572 | w16573);
assign w16574 = v5196;
assign v5197 = ~(w16564 | w16574);
assign w16575 = v5197;
assign w16576 = w16524 & ~w16526;
assign v5198 = ~(w16527 | w16576);
assign w16577 = v5198;
assign w16578 = w16490 & ~w16492;
assign v5199 = ~(w16493 | w16578);
assign w16579 = v5199;
assign w16580 = w5765 & ~w12842;
assign w16581 = w6236 & w11686;
assign w16582 = w5983 & w11689;
assign w16583 = w5764 & ~w11695;
assign v5200 = ~(w16582 | w16583);
assign w16584 = v5200;
assign w16585 = ~w16581 & w16584;
assign w16586 = ~w16580 & w16585;
assign w16587 = pi17 & w16586;
assign v5201 = ~(pi17 | w16586);
assign w16588 = v5201;
assign v5202 = ~(w16587 | w16588);
assign w16589 = v5202;
assign w16590 = w16579 & ~w16589;
assign v5203 = ~(w16179 | w16488);
assign w16591 = v5203;
assign v5204 = ~(w16489 | w16591);
assign w16592 = v5204;
assign w16593 = w5765 & w12694;
assign w16594 = w6236 & w11689;
assign w16595 = w5764 & w11700;
assign w16596 = w5983 & ~w11695;
assign v5205 = ~(w16595 | w16596);
assign w16597 = v5205;
assign w16598 = ~w16594 & w16597;
assign w16599 = ~w16593 & w16598;
assign w16600 = pi17 & w16599;
assign v5206 = ~(pi17 | w16599);
assign w16601 = v5206;
assign v5207 = ~(w16600 | w16601);
assign w16602 = v5207;
assign w16603 = w16592 & ~w16602;
assign w16604 = ~w16592 & w16602;
assign v5208 = ~(w16603 | w16604);
assign w16605 = v5208;
assign w16606 = w5765 & ~w13008;
assign w16607 = w6236 & ~w11695;
assign w16608 = w5983 & w11700;
assign w16609 = w5764 & w11708;
assign v5209 = ~(w16608 | w16609);
assign w16610 = v5209;
assign w16611 = ~w16607 & w16610;
assign w16612 = ~w16606 & w16611;
assign w16613 = pi17 & w16612;
assign v5210 = ~(pi17 | w16612);
assign w16614 = v5210;
assign v5211 = ~(w16613 | w16614);
assign w16615 = v5211;
assign v5212 = ~(w16194 | w16195);
assign w16616 = v5212;
assign v5213 = ~(w16486 | w16616);
assign w16617 = v5213;
assign w16618 = w16486 & w16616;
assign v5214 = ~(w16617 | w16618);
assign w16619 = v5214;
assign w16620 = w16615 & ~w16619;
assign v5215 = ~(w16482 | w16484);
assign w16621 = v5215;
assign v5216 = ~(w16485 | w16621);
assign w16622 = v5216;
assign w16623 = w5765 & w12994;
assign w16624 = w6236 & w11700;
assign w16625 = w5764 & w11711;
assign w16626 = w5983 & w11708;
assign v5217 = ~(w16625 | w16626);
assign w16627 = v5217;
assign w16628 = ~w16624 & w16627;
assign w16629 = ~w16623 & w16628;
assign w16630 = ~pi17 & w16629;
assign w16631 = pi17 & ~w16629;
assign v5218 = ~(w16630 | w16631);
assign w16632 = v5218;
assign w16633 = w16622 & ~w16632;
assign w16634 = ~w16622 & w16632;
assign v5219 = ~(w16633 | w16634);
assign w16635 = v5219;
assign v5220 = ~(w16227 | w16480);
assign w16636 = v5220;
assign v5221 = ~(w16481 | w16636);
assign w16637 = v5221;
assign w16638 = w5765 & w13178;
assign w16639 = w6236 & w11708;
assign w16640 = w5764 & w11714;
assign w16641 = w5983 & w11711;
assign v5222 = ~(w16640 | w16641);
assign w16642 = v5222;
assign w16643 = ~w16639 & w16642;
assign w16644 = ~w16638 & w16643;
assign w16645 = pi17 & w16644;
assign v5223 = ~(pi17 | w16644);
assign w16646 = v5223;
assign v5224 = ~(w16645 | w16646);
assign w16647 = v5224;
assign w16648 = ~w16637 & w16647;
assign w16649 = w16637 & ~w16647;
assign w16650 = w5765 & w13194;
assign w16651 = w5764 & w11720;
assign w16652 = w6236 & w11711;
assign v5225 = ~(w16651 | w16652);
assign w16653 = v5225;
assign w16654 = w5983 & w11714;
assign w16655 = w16653 & ~w16654;
assign w16656 = ~w16650 & w16655;
assign w16657 = pi17 & w16656;
assign v5226 = ~(pi17 | w16656);
assign w16658 = v5226;
assign v5227 = ~(w16657 | w16658);
assign w16659 = v5227;
assign v5228 = ~(w16240 | w16241);
assign w16660 = v5228;
assign w16661 = w16478 & w16660;
assign v5229 = ~(w16478 | w16660);
assign w16662 = v5229;
assign v5230 = ~(w16661 | w16662);
assign w16663 = v5230;
assign v5231 = ~(w16659 | w16663);
assign w16664 = v5231;
assign w16665 = w16659 & w16663;
assign v5232 = ~(w16258 | w16476);
assign w16666 = v5232;
assign v5233 = ~(w16477 | w16666);
assign w16667 = v5233;
assign w16668 = w5765 & w13514;
assign w16669 = w6236 & w11714;
assign w16670 = w5764 & w11723;
assign w16671 = w5983 & w11720;
assign v5234 = ~(w16670 | w16671);
assign w16672 = v5234;
assign w16673 = ~w16669 & w16672;
assign w16674 = ~w16668 & w16673;
assign w16675 = ~pi17 & w16674;
assign w16676 = pi17 & ~w16674;
assign v5235 = ~(w16675 | w16676);
assign w16677 = v5235;
assign v5236 = ~(w16667 | w16677);
assign w16678 = v5236;
assign w16679 = w16667 & w16677;
assign w16680 = w5765 & ~w13310;
assign w16681 = w6236 & w11720;
assign w16682 = w5983 & w11723;
assign w16683 = w5764 & w11726;
assign v5237 = ~(w16682 | w16683);
assign w16684 = v5237;
assign w16685 = ~w16681 & w16684;
assign w16686 = ~w16680 & w16685;
assign w16687 = ~pi17 & w16686;
assign w16688 = pi17 & ~w16686;
assign v5238 = ~(w16687 | w16688);
assign w16689 = v5238;
assign v5239 = ~(w16271 | w16272);
assign w16690 = v5239;
assign w16691 = w16475 & w16690;
assign v5240 = ~(w16475 | w16690);
assign w16692 = v5240;
assign v5241 = ~(w16691 | w16692);
assign w16693 = v5241;
assign w16694 = ~w16689 & w16693;
assign w16695 = w16689 & ~w16693;
assign v5242 = ~(w16287 | w16473);
assign w16696 = v5242;
assign v5243 = ~(w16474 | w16696);
assign w16697 = v5243;
assign w16698 = w5765 & ~w13737;
assign w16699 = w5764 & w11729;
assign w16700 = w6236 & w11723;
assign v5244 = ~(w16699 | w16700);
assign w16701 = v5244;
assign w16702 = w5983 & w11726;
assign w16703 = w16701 & ~w16702;
assign w16704 = ~w16698 & w16703;
assign v5245 = ~(pi17 | w16704);
assign w16705 = v5245;
assign w16706 = pi17 & w16704;
assign v5246 = ~(w16705 | w16706);
assign w16707 = v5246;
assign w16708 = w16697 & ~w16707;
assign w16709 = ~w16697 & w16707;
assign w16710 = w5765 & w13864;
assign w16711 = w5983 & w11729;
assign w16712 = w6236 & w11726;
assign v5247 = ~(w16711 | w16712);
assign w16713 = v5247;
assign w16714 = w5764 & ~w11734;
assign w16715 = w16713 & ~w16714;
assign w16716 = ~w16710 & w16715;
assign v5248 = ~(pi17 | w16716);
assign w16717 = v5248;
assign w16718 = pi17 & w16716;
assign v5249 = ~(w16717 | w16718);
assign w16719 = v5249;
assign v5250 = ~(w16300 | w16301);
assign w16720 = v5250;
assign w16721 = w16472 & w16720;
assign v5251 = ~(w16472 | w16720);
assign w16722 = v5251;
assign v5252 = ~(w16721 | w16722);
assign w16723 = v5252;
assign v5253 = ~(w16719 | w16723);
assign w16724 = v5253;
assign w16725 = w16719 & w16723;
assign v5254 = ~(w16724 | w16725);
assign w16726 = v5254;
assign w16727 = w16468 & ~w16470;
assign v5255 = ~(w16471 | w16727);
assign w16728 = v5255;
assign w16729 = w5765 & ~w13703;
assign w16730 = w5983 & ~w11734;
assign w16731 = w6236 & w11729;
assign v5256 = ~(w16730 | w16731);
assign w16732 = v5256;
assign w16733 = w5764 & w11737;
assign w16734 = w16732 & ~w16733;
assign w16735 = ~w16729 & w16734;
assign w16736 = pi17 & w16735;
assign v5257 = ~(pi17 | w16735);
assign w16737 = v5257;
assign v5258 = ~(w16736 | w16737);
assign w16738 = v5258;
assign w16739 = ~w16728 & w16738;
assign w16740 = w16728 & ~w16738;
assign w16741 = w16464 & ~w16466;
assign v5259 = ~(w16467 | w16741);
assign w16742 = v5259;
assign w16743 = w5765 & w13882;
assign w16744 = w5983 & w11737;
assign w16745 = w6236 & ~w11734;
assign v5260 = ~(w16744 | w16745);
assign w16746 = v5260;
assign w16747 = w5764 & w11740;
assign w16748 = w16746 & ~w16747;
assign w16749 = ~w16743 & w16748;
assign w16750 = pi17 & w16749;
assign v5261 = ~(pi17 | w16749);
assign w16751 = v5261;
assign v5262 = ~(w16750 | w16751);
assign w16752 = v5262;
assign w16753 = w16742 & ~w16752;
assign w16754 = ~w16742 & w16752;
assign v5263 = ~(w16753 | w16754);
assign w16755 = v5263;
assign w16756 = w16460 & ~w16462;
assign v5264 = ~(w16463 | w16756);
assign w16757 = v5264;
assign w16758 = w5765 & w14288;
assign w16759 = w6236 & w11737;
assign w16760 = w5764 & ~w11745;
assign w16761 = w5983 & w11740;
assign v5265 = ~(w16760 | w16761);
assign w16762 = v5265;
assign w16763 = ~w16759 & w16762;
assign w16764 = ~w16758 & w16763;
assign w16765 = pi17 & ~w16764;
assign w16766 = ~pi17 & w16764;
assign v5266 = ~(w16765 | w16766);
assign w16767 = v5266;
assign v5267 = ~(w16757 | w16767);
assign w16768 = v5267;
assign w16769 = w16757 & w16767;
assign w16770 = w16456 & ~w16458;
assign v5268 = ~(w16459 | w16770);
assign w16771 = v5268;
assign w16772 = w6236 & w11740;
assign w16773 = w5983 & ~w11745;
assign w16774 = w5764 & w11748;
assign v5269 = ~(w16773 | w16774);
assign w16775 = v5269;
assign w16776 = ~w16772 & w16775;
assign w16777 = (w16776 & ~w14300) | (w16776 & w30364) | (~w14300 & w30364);
assign w16778 = pi17 & w16777;
assign v5270 = ~(pi17 | w16777);
assign w16779 = v5270;
assign v5271 = ~(w16778 | w16779);
assign w16780 = v5271;
assign w16781 = w16771 & ~w16780;
assign w16782 = w16452 & ~w16454;
assign v5272 = ~(w16455 | w16782);
assign w16783 = v5272;
assign w16784 = w5983 & w11748;
assign w16785 = w6236 & ~w11745;
assign v5273 = ~(w16784 | w16785);
assign w16786 = v5273;
assign w16787 = w5764 & w11759;
assign w16788 = w16786 & ~w16787;
assign w16789 = (w16788 & ~w13948) | (w16788 & w30183) | (~w13948 & w30183);
assign v5274 = ~(pi17 | w16789);
assign w16790 = v5274;
assign w16791 = pi17 & w16789;
assign v5275 = ~(w16790 | w16791);
assign w16792 = v5275;
assign w16793 = w16783 & ~w16792;
assign w16794 = w16448 & ~w16450;
assign v5276 = ~(w16451 | w16794);
assign w16795 = v5276;
assign w16796 = (w5765 & w11841) | (w5765 & w30045) | (w11841 & w30045);
assign w16797 = w6236 & w11748;
assign w16798 = w5983 & w11759;
assign w16799 = w5764 & w11761;
assign v5277 = ~(w16798 | w16799);
assign w16800 = v5277;
assign w16801 = ~w16797 & w16800;
assign w16802 = ~w16796 & w30184;
assign w16803 = (pi17 & w16796) | (pi17 & w30185) | (w16796 & w30185);
assign v5278 = ~(w16802 | w16803);
assign w16804 = v5278;
assign w16805 = w16795 & w16804;
assign w16806 = w16444 & ~w16446;
assign v5279 = ~(w16447 | w16806);
assign w16807 = v5279;
assign w16808 = w5764 & ~w11771;
assign w16809 = w6236 & w11759;
assign v5280 = ~(w16808 | w16809);
assign w16810 = v5280;
assign w16811 = w5983 & w11761;
assign w16812 = w16810 & ~w16811;
assign w16813 = (~w14356 & w30046) | (~w14356 & w30047) | (w30046 & w30047);
assign w16814 = (w14356 & w30048) | (w14356 & w30049) | (w30048 & w30049);
assign v5281 = ~(w16813 | w16814);
assign w16815 = v5281;
assign w16816 = w16807 & ~w16815;
assign w16817 = w16440 & ~w16442;
assign v5282 = ~(w16443 | w16817);
assign w16818 = v5282;
assign w16819 = w5764 & w11768;
assign w16820 = w5983 & ~w11771;
assign v5283 = ~(w16819 | w16820);
assign w16821 = v5283;
assign w16822 = w6236 & w11761;
assign w16823 = w16821 & ~w16822;
assign w16824 = (w14383 & w29722) | (w14383 & w29723) | (w29722 & w29723);
assign w16825 = (~w14383 & w29724) | (~w14383 & w29725) | (w29724 & w29725);
assign v5284 = ~(w16824 | w16825);
assign w16826 = v5284;
assign w16827 = w16818 & ~w16826;
assign w16828 = w16436 & ~w16438;
assign v5285 = ~(w16439 | w16828);
assign w16829 = v5285;
assign w16830 = w5765 & w14409;
assign w16831 = w5983 & w11768;
assign w16832 = (w6236 & ~w11766) | (w6236 & w29499) | (~w11766 & w29499);
assign w16833 = w5764 & w11776;
assign w16834 = ~w16832 & w29726;
assign w16835 = (~pi17 & w16830) | (~pi17 & w29727) | (w16830 & w29727);
assign w16836 = ~w16830 & w29728;
assign v5286 = ~(w16835 | w16836);
assign w16837 = v5286;
assign w16838 = w16829 & ~w16837;
assign v5287 = ~(w16425 | w16434);
assign w16839 = v5287;
assign v5288 = ~(w16435 | w16839);
assign w16840 = v5288;
assign w16841 = w5764 & w11784;
assign w16842 = w6236 & w11768;
assign w16843 = w5983 & w11776;
assign w16844 = (w29283 & ~w14461) | (w29283 & w30816) | (~w14461 & w30816);
assign w16845 = (w14461 & w30817) | (w14461 & w30818) | (w30817 & w30818);
assign v5289 = ~(w16844 | w16845);
assign w16846 = v5289;
assign w16847 = w16840 & ~w16846;
assign w16848 = pi20 & ~w16414;
assign v5290 = ~(w16420 | w16848);
assign w16849 = v5290;
assign w16850 = w16420 & w16848;
assign v5291 = ~(w16849 | w16850);
assign w16851 = v5291;
assign w16852 = w5983 & w11784;
assign w16853 = w6236 & w11776;
assign v5292 = ~(w16852 | w16853);
assign w16854 = v5292;
assign w16855 = w5764 & w11793;
assign w16856 = (w14504 & w29500) | (w14504 & w29501) | (w29500 & w29501);
assign w16857 = (~w14504 & w29502) | (~w14504 & w29503) | (w29502 & w29503);
assign v5293 = ~(w16856 | w16857);
assign w16858 = v5293;
assign v5294 = ~(w16851 | w16858);
assign w16859 = v5294;
assign w16860 = w16408 & ~w16413;
assign v5295 = ~(w16414 | w16860);
assign w16861 = v5295;
assign w16862 = w5765 & w14547;
assign w16863 = w5764 & w11803;
assign w16864 = w6236 & w11784;
assign w16865 = w5983 & w11793;
assign v5296 = ~(w16864 | w16865);
assign w16866 = v5296;
assign w16867 = (pi17 & w16862) | (pi17 & w29002) | (w16862 & w29002);
assign w16868 = ~w16862 & w29003;
assign v5297 = ~(w16867 | w16868);
assign w16869 = v5297;
assign w16870 = w16861 & w16869;
assign w16871 = w5756 & w11800;
assign w16872 = pi17 & w16871;
assign w16873 = w5765 & ~w14609;
assign w16874 = w6236 & w11798;
assign w16875 = w5983 & w11800;
assign v5298 = ~(w16874 | w16875);
assign w16876 = v5298;
assign w16877 = ~w16873 & w16876;
assign w16878 = ~w16872 & w16877;
assign w16879 = w5764 & w11800;
assign w16880 = (~w16879 & w14639) | (~w16879 & w29729) | (w14639 & w29729);
assign w16881 = w6236 & w11803;
assign w16882 = w5983 & w11798;
assign v5299 = ~(w16881 | w16882);
assign w16883 = v5299;
assign w16884 = w16880 & w16883;
assign w16885 = w16880 & w30520;
assign w16886 = w16878 & w16885;
assign w16887 = w16407 & w16886;
assign v5300 = ~(w16407 | w16886);
assign w16888 = v5300;
assign v5301 = ~(w16887 | w16888);
assign w16889 = v5301;
assign w16890 = w5765 & w14569;
assign w16891 = w5764 & w11798;
assign w16892 = w6236 & w11793;
assign w16893 = w5983 & w11803;
assign v5302 = ~(w16892 | w16893);
assign w16894 = v5302;
assign w16895 = ~w16891 & w16894;
assign w16896 = (pi17 & w16890) | (pi17 & w29504) | (w16890 & w29504);
assign w16897 = (w29505 & ~w14569) | (w29505 & w29730) | (~w14569 & w29730);
assign v5303 = ~(w16896 | w16897);
assign w16898 = v5303;
assign w16899 = w16889 & w16898;
assign w16900 = (~w16887 & ~w16898) | (~w16887 & w29731) | (~w16898 & w29731);
assign v5304 = ~(w16861 | w16869);
assign w16901 = v5304;
assign v5305 = ~(w16870 | w16901);
assign w16902 = v5305;
assign w16903 = ~w16900 & w16902;
assign w16904 = (~w16870 & ~w16902) | (~w16870 & w29506) | (~w16902 & w29506);
assign w16905 = w16851 & w16858;
assign v5306 = ~(w16859 | w16905);
assign w16906 = v5306;
assign w16907 = ~w16904 & w16906;
assign v5307 = ~(w16859 | w16907);
assign w16908 = v5307;
assign w16909 = ~w16840 & w16846;
assign v5308 = ~(w16847 | w16909);
assign w16910 = v5308;
assign w16911 = ~w16908 & w16910;
assign w16912 = (~w16847 & w16908) | (~w16847 & w31047) | (w16908 & w31047);
assign w16913 = ~w16829 & w16837;
assign v5309 = ~(w16838 | w16913);
assign w16914 = v5309;
assign w16915 = ~w16912 & w16914;
assign w16916 = (~w16838 & w16912) | (~w16838 & w29732) | (w16912 & w29732);
assign w16917 = ~w16818 & w16826;
assign v5310 = ~(w16827 | w16917);
assign w16918 = v5310;
assign w16919 = ~w16916 & w16918;
assign w16920 = (~w16827 & w16916) | (~w16827 & w29871) | (w16916 & w29871);
assign w16921 = ~w16807 & w16815;
assign v5311 = ~(w16816 | w16921);
assign w16922 = v5311;
assign w16923 = ~w16920 & w16922;
assign v5312 = ~(w16816 | w16923);
assign w16924 = v5312;
assign v5313 = ~(w16795 | w16804);
assign w16925 = v5313;
assign v5314 = ~(w16805 | w16925);
assign w16926 = v5314;
assign w16927 = ~w16924 & w16926;
assign w16928 = (~w16805 & w16924) | (~w16805 & w30050) | (w16924 & w30050);
assign w16929 = ~w16783 & w16792;
assign v5315 = ~(w16793 | w16929);
assign w16930 = v5315;
assign w16931 = ~w16928 & w16930;
assign w16932 = (~w16793 & w16928) | (~w16793 & w30819) | (w16928 & w30819);
assign w16933 = ~w16771 & w16780;
assign v5316 = ~(w16781 | w16933);
assign w16934 = v5316;
assign w16935 = ~w16932 & w16934;
assign w16936 = (~w16781 & w16932) | (~w16781 & w30186) | (w16932 & w30186);
assign w16937 = (~w16768 & ~w16936) | (~w16768 & w30365) | (~w16936 & w30365);
assign w16938 = w16755 & w16937;
assign w16939 = (~w16753 & ~w16755) | (~w16753 & w30820) | (~w16755 & w30820);
assign w16940 = (~w16739 & ~w16939) | (~w16739 & w30521) | (~w16939 & w30521);
assign w16941 = w16726 & w16940;
assign v5317 = ~(w16724 | w16941);
assign w16942 = v5317;
assign w16943 = (~w16709 & w16941) | (~w16709 & w30639) | (w16941 & w30639);
assign w16944 = (~w30639 & w30821) | (~w30639 & w30822) | (w30821 & w30822);
assign w16945 = (~w16694 & ~w16944) | (~w16694 & w31048) | (~w16944 & w31048);
assign w16946 = (~w16678 & w16945) | (~w16678 & w31194) | (w16945 & w31194);
assign w16947 = ~w16665 & w16946;
assign v5318 = ~(w16664 | w16947);
assign w16948 = v5318;
assign w16949 = (~w16648 & ~w16948) | (~w16648 & w31279) | (~w16948 & w31279);
assign w16950 = w16635 & ~w16949;
assign v5319 = ~(w16633 | w16950);
assign w16951 = v5319;
assign w16952 = ~w16615 & w16619;
assign v5320 = ~(w16620 | w16952);
assign w16953 = v5320;
assign w16954 = ~w16951 & w16953;
assign v5321 = ~(w16620 | w16954);
assign w16955 = v5321;
assign w16956 = w16605 & w16955;
assign v5322 = ~(w16603 | w16956);
assign w16957 = v5322;
assign w16958 = ~w16579 & w16589;
assign v5323 = ~(w16590 | w16958);
assign w16959 = v5323;
assign w16960 = ~w16957 & w16959;
assign v5324 = ~(w16590 | w16960);
assign w16961 = v5324;
assign w16962 = w6389 & w12469;
assign w16963 = w6871 & w11673;
assign w16964 = w7004 & w11671;
assign v5325 = ~(w16963 | w16964);
assign w16965 = v5325;
assign w16966 = w6388 & w11678;
assign w16967 = w16965 & ~w16966;
assign w16968 = ~w16962 & w16967;
assign v5326 = ~(pi14 | w16968);
assign w16969 = v5326;
assign w16970 = pi14 & w16968;
assign v5327 = ~(w16969 | w16970);
assign w16971 = v5327;
assign v5328 = ~(w16961 | w16971);
assign w16972 = v5328;
assign w16973 = w16961 & w16971;
assign v5329 = ~(w16972 | w16973);
assign w16974 = v5329;
assign v5330 = ~(w16507 | w16509);
assign w16975 = v5330;
assign v5331 = ~(w16510 | w16975);
assign w16976 = v5331;
assign w16977 = w16974 & ~w16976;
assign v5332 = ~(w16972 | w16977);
assign w16978 = v5332;
assign w16979 = w16577 & w16978;
assign v5333 = ~(w16577 | w16978);
assign w16980 = v5333;
assign v5334 = ~(w16979 | w16980);
assign w16981 = v5334;
assign w16982 = w7178 & ~w12351;
assign w16983 = w7466 & w12155;
assign w16984 = w7765 & w12237;
assign v5335 = ~(w16983 | w16984);
assign w16985 = v5335;
assign w16986 = w7177 & w12084;
assign w16987 = w16985 & ~w16986;
assign w16988 = ~w16982 & w16987;
assign w16989 = pi11 & w16988;
assign v5336 = ~(pi11 | w16988);
assign w16990 = v5336;
assign v5337 = ~(w16989 | w16990);
assign w16991 = v5337;
assign w16992 = w16981 & w16991;
assign v5338 = ~(w16979 | w16992);
assign w16993 = v5338;
assign w16994 = w16564 & w16574;
assign v5339 = ~(w16575 | w16994);
assign w16995 = v5339;
assign w16996 = ~w16993 & w16995;
assign v5340 = ~(w16575 | w16996);
assign w16997 = v5340;
assign w16998 = w8140 & w12381;
assign w16999 = w8141 & w12505;
assign v5341 = ~(w8526 | w16999);
assign w17000 = v5341;
assign v5342 = ~(w12406 | w17000);
assign w17001 = v5342;
assign v5343 = ~(w8926 | w17001);
assign w17002 = v5343;
assign w17003 = ~w16998 & w17002;
assign w17004 = ~pi08 & w17003;
assign w17005 = pi08 & ~w17003;
assign v5344 = ~(w17004 | w17005);
assign w17006 = v5344;
assign w17007 = w16997 & w17006;
assign w17008 = w16545 & ~w16547;
assign v5345 = ~(w16548 | w17008);
assign w17009 = v5345;
assign v5346 = ~(w16997 | w17006);
assign w17010 = v5346;
assign v5347 = ~(w17007 | w17010);
assign w17011 = v5347;
assign w17012 = w17009 & w17011;
assign v5348 = ~(w17007 | w17012);
assign w17013 = v5348;
assign v5349 = ~(w16557 | w16559);
assign w17014 = v5349;
assign v5350 = ~(w16560 | w17014);
assign w17015 = v5350;
assign w17016 = w17013 & ~w17015;
assign v5351 = ~(w16981 | w16991);
assign w17017 = v5351;
assign v5352 = ~(w16992 | w17017);
assign w17018 = v5352;
assign w17019 = ~w16974 & w16976;
assign v5353 = ~(w16977 | w17019);
assign w17020 = v5353;
assign w17021 = w16957 & ~w16959;
assign v5354 = ~(w16960 | w17021);
assign w17022 = v5354;
assign w17023 = w6389 & w12454;
assign w17024 = w6871 & w11678;
assign w17025 = w7004 & w11673;
assign v5355 = ~(w17024 | w17025);
assign w17026 = v5355;
assign w17027 = w6388 & ~w11683;
assign w17028 = w17026 & ~w17027;
assign w17029 = ~w17023 & w17028;
assign w17030 = pi14 & w17029;
assign v5356 = ~(pi14 | w17029);
assign w17031 = v5356;
assign v5357 = ~(w17030 | w17031);
assign w17032 = v5357;
assign w17033 = w17022 & ~w17032;
assign v5358 = ~(w16605 | w16955);
assign w17034 = v5358;
assign v5359 = ~(w16956 | w17034);
assign w17035 = v5359;
assign w17036 = w6389 & w12594;
assign w17037 = w7004 & w11678;
assign w17038 = w6871 & ~w11683;
assign w17039 = w6388 & w11686;
assign v5360 = ~(w17038 | w17039);
assign w17040 = v5360;
assign w17041 = ~w17037 & w17040;
assign w17042 = ~w17036 & w17041;
assign w17043 = pi14 & ~w17042;
assign w17044 = ~pi14 & w17042;
assign v5361 = ~(w17043 | w17044);
assign w17045 = v5361;
assign w17046 = w17035 & w17045;
assign v5362 = ~(w17035 | w17045);
assign w17047 = v5362;
assign v5363 = ~(w17046 | w17047);
assign w17048 = v5363;
assign w17049 = w16951 & ~w16953;
assign v5364 = ~(w16954 | w17049);
assign w17050 = v5364;
assign w17051 = w6389 & w12610;
assign w17052 = w7004 & ~w11683;
assign w17053 = w6871 & w11686;
assign w17054 = w6388 & w11689;
assign v5365 = ~(w17053 | w17054);
assign w17055 = v5365;
assign w17056 = ~w17052 & w17055;
assign w17057 = ~w17051 & w17056;
assign w17058 = pi14 & ~w17057;
assign w17059 = ~pi14 & w17057;
assign v5366 = ~(w17058 | w17059);
assign w17060 = v5366;
assign w17061 = ~w17050 & w17060;
assign w17062 = w17050 & ~w17060;
assign w17063 = ~w16635 & w16949;
assign v5367 = ~(w16950 | w17063);
assign w17064 = v5367;
assign w17065 = w6389 & ~w12842;
assign w17066 = w6871 & w11689;
assign w17067 = w7004 & w11686;
assign v5368 = ~(w17066 | w17067);
assign w17068 = v5368;
assign w17069 = w6388 & ~w11695;
assign w17070 = w17068 & ~w17069;
assign w17071 = ~w17065 & w17070;
assign v5369 = ~(pi14 | w17071);
assign w17072 = v5369;
assign w17073 = pi14 & w17071;
assign v5370 = ~(w17072 | w17073);
assign w17074 = v5370;
assign v5371 = ~(w17064 | w17074);
assign w17075 = v5371;
assign w17076 = w17064 & w17074;
assign w17077 = w6389 & w12694;
assign w17078 = w7004 & w11689;
assign w17079 = w6388 & w11700;
assign w17080 = w6871 & ~w11695;
assign v5372 = ~(w17079 | w17080);
assign w17081 = v5372;
assign w17082 = ~w17078 & w17081;
assign w17083 = ~w17077 & w17082;
assign w17084 = ~pi14 & w17083;
assign w17085 = pi14 & ~w17083;
assign v5373 = ~(w17084 | w17085);
assign w17086 = v5373;
assign v5374 = ~(w16648 | w16649);
assign w17087 = v5374;
assign w17088 = w16948 & ~w17087;
assign w17089 = ~w16948 & w17087;
assign v5375 = ~(w17088 | w17089);
assign w17090 = v5375;
assign v5376 = ~(w17086 | w17090);
assign w17091 = v5376;
assign w17092 = w17086 & w17090;
assign v5377 = ~(w17091 | w17092);
assign w17093 = v5377;
assign v5378 = ~(w16664 | w16665);
assign w17094 = v5378;
assign w17095 = ~w16946 & w17094;
assign w17096 = w16946 & ~w17094;
assign v5379 = ~(w17095 | w17096);
assign w17097 = v5379;
assign w17098 = w6389 & ~w13008;
assign w17099 = w6388 & w11708;
assign w17100 = w7004 & ~w11695;
assign v5380 = ~(w17099 | w17100);
assign w17101 = v5380;
assign w17102 = w6871 & w11700;
assign w17103 = w17101 & ~w17102;
assign w17104 = ~w17098 & w17103;
assign v5381 = ~(pi14 | w17104);
assign w17105 = v5381;
assign w17106 = pi14 & w17104;
assign v5382 = ~(w17105 | w17106);
assign w17107 = v5382;
assign w17108 = w17097 & w17107;
assign v5383 = ~(w17097 | w17107);
assign w17109 = v5383;
assign w17110 = w6389 & w12994;
assign w17111 = w7004 & w11700;
assign w17112 = w6871 & w11708;
assign w17113 = w6388 & w11711;
assign v5384 = ~(w17112 | w17113);
assign w17114 = v5384;
assign w17115 = ~w17111 & w17114;
assign w17116 = ~pi14 & w17115;
assign w17117 = ~w17110 & w17116;
assign w17118 = w6378 & w6383;
assign w17119 = w12994 & w17118;
assign w17120 = pi14 & ~w17115;
assign v5385 = ~(w17119 | w17120);
assign w17121 = v5385;
assign w17122 = ~w17117 & w17121;
assign v5386 = ~(w16678 | w16679);
assign w17123 = v5386;
assign v5387 = ~(w16945 | w17123);
assign w17124 = v5387;
assign w17125 = w16945 & w17123;
assign v5388 = ~(w17124 | w17125);
assign w17126 = v5388;
assign w17127 = w17122 & w17126;
assign v5389 = ~(w16694 | w16695);
assign w17128 = v5389;
assign v5390 = ~(w16944 | w17128);
assign w17129 = v5390;
assign w17130 = w16944 & w17128;
assign v5391 = ~(w17129 | w17130);
assign w17131 = v5391;
assign w17132 = w6389 & w13178;
assign w17133 = w7004 & w11708;
assign w17134 = w6388 & w11714;
assign w17135 = w6871 & w11711;
assign v5392 = ~(w17134 | w17135);
assign w17136 = v5392;
assign w17137 = ~w17133 & w17136;
assign w17138 = ~w17132 & w17137;
assign w17139 = pi14 & ~w17138;
assign w17140 = ~pi14 & w17138;
assign v5393 = ~(w17139 | w17140);
assign w17141 = v5393;
assign w17142 = ~w17131 & w17141;
assign w17143 = w6389 & w13194;
assign w17144 = w6388 & w11720;
assign w17145 = w7004 & w11711;
assign v5394 = ~(w17144 | w17145);
assign w17146 = v5394;
assign w17147 = w6871 & w11714;
assign w17148 = w17146 & ~w17147;
assign w17149 = ~w17143 & w17148;
assign w17150 = pi14 & w17149;
assign v5395 = ~(pi14 | w17149);
assign w17151 = v5395;
assign v5396 = ~(w17150 | w17151);
assign w17152 = v5396;
assign v5397 = ~(w16708 | w16709);
assign w17153 = v5397;
assign w17154 = w16942 & ~w17153;
assign w17155 = ~w16708 & w16943;
assign v5398 = ~(w17154 | w17155);
assign w17156 = v5398;
assign w17157 = ~w17152 & w17156;
assign w17158 = w17152 & ~w17156;
assign v5399 = ~(w17157 | w17158);
assign w17159 = v5399;
assign v5400 = ~(w16726 | w16940);
assign w17160 = v5400;
assign v5401 = ~(w16941 | w17160);
assign w17161 = v5401;
assign w17162 = w6389 & w13514;
assign w17163 = w7004 & w11714;
assign w17164 = w6388 & w11723;
assign w17165 = w6871 & w11720;
assign v5402 = ~(w17164 | w17165);
assign w17166 = v5402;
assign w17167 = ~w17163 & w17166;
assign w17168 = ~w17162 & w17167;
assign w17169 = pi14 & ~w17168;
assign w17170 = ~pi14 & w17168;
assign v5403 = ~(w17169 | w17170);
assign w17171 = v5403;
assign v5404 = ~(w17161 | w17171);
assign w17172 = v5404;
assign w17173 = w17161 & w17171;
assign w17174 = w6389 & ~w13310;
assign w17175 = w7004 & w11720;
assign w17176 = w6388 & w11726;
assign w17177 = w6871 & w11723;
assign v5405 = ~(w17176 | w17177);
assign w17178 = v5405;
assign w17179 = ~w17175 & w17178;
assign w17180 = ~w17174 & w17179;
assign w17181 = ~pi14 & w17180;
assign w17182 = pi14 & ~w17180;
assign v5406 = ~(w17181 | w17182);
assign w17183 = v5406;
assign v5407 = ~(w16739 | w16740);
assign w17184 = v5407;
assign w17185 = w16939 & w17184;
assign v5408 = ~(w16939 | w17184);
assign w17186 = v5408;
assign v5409 = ~(w17185 | w17186);
assign w17187 = v5409;
assign w17188 = w17183 & ~w17187;
assign v5410 = ~(w16755 | w16937);
assign w17189 = v5410;
assign v5411 = ~(w16938 | w17189);
assign w17190 = v5411;
assign w17191 = w6389 & ~w13737;
assign w17192 = w7004 & w11723;
assign w17193 = w6388 & w11729;
assign w17194 = w6871 & w11726;
assign v5412 = ~(w17193 | w17194);
assign w17195 = v5412;
assign w17196 = ~w17192 & w17195;
assign w17197 = ~w17191 & w17196;
assign w17198 = pi14 & ~w17197;
assign w17199 = ~pi14 & w17197;
assign v5413 = ~(w17198 | w17199);
assign w17200 = v5413;
assign v5414 = ~(w17190 | w17200);
assign w17201 = v5414;
assign w17202 = w6389 & w13864;
assign w17203 = w6871 & w11729;
assign w17204 = w7004 & w11726;
assign v5415 = ~(w17203 | w17204);
assign w17205 = v5415;
assign w17206 = w6388 & ~w11734;
assign w17207 = w17205 & ~w17206;
assign w17208 = ~w17202 & w17207;
assign v5416 = ~(pi14 | w17208);
assign w17209 = v5416;
assign w17210 = pi14 & w17208;
assign v5417 = ~(w17209 | w17210);
assign w17211 = v5417;
assign v5418 = ~(w16768 | w16769);
assign w17212 = v5418;
assign v5419 = ~(w16936 | w17212);
assign w17213 = v5419;
assign w17214 = w16936 & w17212;
assign v5420 = ~(w17213 | w17214);
assign w17215 = v5420;
assign v5421 = ~(w17211 | w17215);
assign w17216 = v5421;
assign w17217 = w17211 & w17215;
assign v5422 = ~(w17216 | w17217);
assign w17218 = v5422;
assign w17219 = w16932 & ~w16934;
assign v5423 = ~(w16935 | w17219);
assign w17220 = v5423;
assign w17221 = w6389 & ~w13703;
assign w17222 = w6871 & ~w11734;
assign w17223 = w7004 & w11729;
assign v5424 = ~(w17222 | w17223);
assign w17224 = v5424;
assign w17225 = w6388 & w11737;
assign w17226 = w17224 & ~w17225;
assign w17227 = ~w17221 & w17226;
assign w17228 = pi14 & w17227;
assign v5425 = ~(pi14 | w17227);
assign w17229 = v5425;
assign v5426 = ~(w17228 | w17229);
assign w17230 = v5426;
assign w17231 = ~w17220 & w17230;
assign w17232 = w17220 & ~w17230;
assign w17233 = w16928 & ~w16930;
assign v5427 = ~(w16931 | w17233);
assign w17234 = v5427;
assign w17235 = w6389 & w13882;
assign w17236 = w7004 & ~w11734;
assign w17237 = w6871 & w11737;
assign w17238 = w6388 & w11740;
assign v5428 = ~(w17237 | w17238);
assign w17239 = v5428;
assign w17240 = ~w17236 & w17239;
assign w17241 = ~w17235 & w17240;
assign w17242 = ~pi14 & w17241;
assign w17243 = pi14 & ~w17241;
assign v5429 = ~(w17242 | w17243);
assign w17244 = v5429;
assign w17245 = w17234 & w17244;
assign v5430 = ~(w17234 | w17244);
assign w17246 = v5430;
assign v5431 = ~(w17245 | w17246);
assign w17247 = v5431;
assign w17248 = w16924 & ~w16926;
assign v5432 = ~(w16927 | w17248);
assign w17249 = v5432;
assign w17250 = w6389 & w14288;
assign w17251 = w7004 & w11737;
assign w17252 = w6388 & ~w11745;
assign w17253 = w6871 & w11740;
assign v5433 = ~(w17252 | w17253);
assign w17254 = v5433;
assign w17255 = ~w17251 & w17254;
assign w17256 = ~w17250 & w17255;
assign w17257 = pi14 & ~w17256;
assign w17258 = ~pi14 & w17256;
assign v5434 = ~(w17257 | w17258);
assign w17259 = v5434;
assign v5435 = ~(w17249 | w17259);
assign w17260 = v5435;
assign w17261 = w17249 & w17259;
assign w17262 = w16920 & ~w16922;
assign v5436 = ~(w16923 | w17262);
assign w17263 = v5436;
assign w17264 = w7004 & w11740;
assign w17265 = w6871 & ~w11745;
assign w17266 = w6388 & w11748;
assign v5437 = ~(w17265 | w17266);
assign w17267 = v5437;
assign w17268 = ~w17264 & w17267;
assign w17269 = (w17268 & ~w14300) | (w17268 & w30051) | (~w14300 & w30051);
assign w17270 = pi14 & ~w17269;
assign w17271 = ~pi14 & w17269;
assign v5438 = ~(w17270 | w17271);
assign w17272 = v5438;
assign w17273 = w17263 & w17272;
assign w17274 = w16916 & ~w16918;
assign v5439 = ~(w16919 | w17274);
assign w17275 = v5439;
assign w17276 = w6871 & w11748;
assign w17277 = w7004 & ~w11745;
assign v5440 = ~(w17276 | w17277);
assign w17278 = v5440;
assign w17279 = w6388 & w11759;
assign w17280 = w17278 & ~w17279;
assign w17281 = (w17280 & ~w13948) | (w17280 & w30052) | (~w13948 & w30052);
assign v5441 = ~(pi14 | w17281);
assign w17282 = v5441;
assign w17283 = pi14 & w17281;
assign v5442 = ~(w17282 | w17283);
assign w17284 = v5442;
assign w17285 = w17275 & ~w17284;
assign w17286 = w16912 & ~w16914;
assign v5443 = ~(w16915 | w17286);
assign w17287 = v5443;
assign w17288 = (w6389 & w11841) | (w6389 & w29733) | (w11841 & w29733);
assign w17289 = w6871 & w11759;
assign w17290 = w7004 & w11748;
assign v5444 = ~(w17289 | w17290);
assign w17291 = v5444;
assign w17292 = w6388 & w11761;
assign w17293 = w17291 & ~w17292;
assign w17294 = ~w17288 & w17293;
assign v5445 = ~(pi14 | w17294);
assign w17295 = v5445;
assign w17296 = pi14 & w17294;
assign v5446 = ~(w17295 | w17296);
assign w17297 = v5446;
assign w17298 = w17287 & ~w17297;
assign w17299 = w16908 & ~w16910;
assign v5447 = ~(w16911 | w17299);
assign w17300 = v5447;
assign w17301 = w6388 & ~w11771;
assign w17302 = w7004 & w11759;
assign v5448 = ~(w17301 | w17302);
assign w17303 = v5448;
assign w17304 = w6871 & w11761;
assign w17305 = w17303 & ~w17304;
assign w17306 = (~w14356 & w29734) | (~w14356 & w29735) | (w29734 & w29735);
assign w17307 = (w14356 & w29736) | (w14356 & w29737) | (w29736 & w29737);
assign v5449 = ~(w17306 | w17307);
assign w17308 = v5449;
assign w17309 = w17300 & ~w17308;
assign w17310 = w16904 & ~w16906;
assign v5450 = ~(w16907 | w17310);
assign w17311 = v5450;
assign w17312 = w6871 & ~w11771;
assign w17313 = w6388 & w11768;
assign w17314 = w7004 & w11761;
assign v5451 = ~(w17313 | w17314);
assign w17315 = v5451;
assign w17316 = ~w17312 & w17315;
assign w17317 = (w14383 & w29508) | (w14383 & w29509) | (w29508 & w29509);
assign w17318 = (~w14383 & w29510) | (~w14383 & w29511) | (w29510 & w29511);
assign v5452 = ~(w17317 | w17318);
assign w17319 = v5452;
assign w17320 = w17311 & w17319;
assign w17321 = w16900 & ~w16902;
assign v5453 = ~(w16903 | w17321);
assign w17322 = v5453;
assign w17323 = w6871 & w11768;
assign w17324 = (w7004 & ~w11766) | (w7004 & w29285) | (~w11766 & w29285);
assign w17325 = w6388 & w11776;
assign w17326 = (w14409 & w29872) | (w14409 & w29873) | (w29872 & w29873);
assign w17327 = (w29287 & ~w14409) | (w29287 & w29874) | (~w14409 & w29874);
assign v5454 = ~(w17326 | w17327);
assign w17328 = v5454;
assign w17329 = w17322 & ~w17328;
assign v5455 = ~(w16889 | w16898);
assign w17330 = v5455;
assign v5456 = ~(w16899 | w17330);
assign w17331 = v5456;
assign w17332 = w11533 & w29288;
assign w17333 = w6388 & w11784;
assign w17334 = w6871 & w11776;
assign v5457 = ~(w17333 | w17334);
assign w17335 = v5457;
assign w17336 = ~w17332 & w17335;
assign w17337 = (~w14461 & w29289) | (~w14461 & w29290) | (w29289 & w29290);
assign w17338 = (w14461 & w29291) | (w14461 & w29292) | (w29291 & w29292);
assign v5458 = ~(w17337 | w17338);
assign w17339 = v5458;
assign w17340 = w17331 & w17339;
assign w17341 = pi17 & ~w16878;
assign v5459 = ~(w16884 | w17341);
assign w17342 = v5459;
assign w17343 = w16884 & w17341;
assign v5460 = ~(w17342 | w17343);
assign w17344 = v5460;
assign w17345 = w6871 & w11784;
assign w17346 = w7004 & w11776;
assign v5461 = ~(w17345 | w17346);
assign w17347 = v5461;
assign w17348 = w6388 & w11793;
assign w17349 = (w14504 & w29005) | (w14504 & w29006) | (w29005 & w29006);
assign w17350 = (~w14504 & w29007) | (~w14504 & w29008) | (w29007 & w29008);
assign v5462 = ~(w17349 | w17350);
assign w17351 = v5462;
assign v5463 = ~(w17344 | w17351);
assign w17352 = v5463;
assign w17353 = w16872 & ~w16877;
assign v5464 = ~(w16878 | w17353);
assign w17354 = v5464;
assign w17355 = w6389 & w14547;
assign w17356 = w6388 & w11803;
assign w17357 = w7004 & w11784;
assign w17358 = w6871 & w11793;
assign v5465 = ~(w17357 | w17358);
assign w17359 = v5465;
assign w17360 = (pi14 & w17355) | (pi14 & w28754) | (w17355 & w28754);
assign w17361 = ~w17355 & w28755;
assign v5466 = ~(w17360 | w17361);
assign w17362 = v5466;
assign w17363 = w17354 & w17362;
assign w17364 = w6383 & w11800;
assign w17365 = pi14 & w17364;
assign w17366 = w6389 & ~w14609;
assign w17367 = w7004 & w11798;
assign w17368 = w6871 & w11800;
assign v5467 = ~(w17367 | w17368);
assign w17369 = v5467;
assign w17370 = ~w17366 & w17369;
assign w17371 = ~w17365 & w17370;
assign w17372 = w6388 & w11800;
assign w17373 = (~w17372 & w14639) | (~w17372 & w29512) | (w14639 & w29512);
assign w17374 = w7004 & w11803;
assign w17375 = w6871 & w11798;
assign v5468 = ~(w17374 | w17375);
assign w17376 = v5468;
assign w17377 = w17373 & w17376;
assign w17378 = w17373 & w30522;
assign w17379 = w17371 & w17378;
assign w17380 = w16871 & w17379;
assign v5469 = ~(w16871 | w17379);
assign w17381 = v5469;
assign v5470 = ~(w17380 | w17381);
assign w17382 = v5470;
assign w17383 = w6389 & w14569;
assign w17384 = w6388 & w11798;
assign w17385 = w7004 & w11793;
assign w17386 = w6871 & w11803;
assign v5471 = ~(w17385 | w17386);
assign w17387 = v5471;
assign w17388 = (pi14 & w17383) | (pi14 & w29293) | (w17383 & w29293);
assign w17389 = ~w17383 & w29294;
assign v5472 = ~(w17388 | w17389);
assign w17390 = v5472;
assign w17391 = w17382 & w17390;
assign w17392 = (~w17380 & ~w17390) | (~w17380 & w29513) | (~w17390 & w29513);
assign v5473 = ~(w17354 | w17362);
assign w17393 = v5473;
assign v5474 = ~(w17363 | w17393);
assign w17394 = v5474;
assign w17395 = ~w17392 & w17394;
assign w17396 = (~w17363 & ~w17394) | (~w17363 & w29009) | (~w17394 & w29009);
assign w17397 = w17344 & w17351;
assign v5475 = ~(w17352 | w17397);
assign w17398 = v5475;
assign w17399 = ~w17396 & w17398;
assign v5476 = ~(w17352 | w17399);
assign w17400 = v5476;
assign v5477 = ~(w17331 | w17339);
assign w17401 = v5477;
assign v5478 = ~(w17340 | w17401);
assign w17402 = v5478;
assign w17403 = ~w17400 & w17402;
assign w17404 = (~w17340 & w17400) | (~w17340 & w29875) | (w17400 & w29875);
assign w17405 = ~w17322 & w17328;
assign v5479 = ~(w17329 | w17405);
assign w17406 = v5479;
assign w17407 = ~w17404 & w17406;
assign w17408 = (~w17329 & w17404) | (~w17329 & w29514) | (w17404 & w29514);
assign v5480 = ~(w17311 | w17319);
assign w17409 = v5480;
assign v5481 = ~(w17320 | w17409);
assign w17410 = v5481;
assign w17411 = ~w17408 & w17410;
assign w17412 = (~w17320 & w17408) | (~w17320 & w29876) | (w17408 & w29876);
assign w17413 = ~w17300 & w17308;
assign v5482 = ~(w17309 | w17413);
assign w17414 = v5482;
assign w17415 = ~w17412 & w17414;
assign v5483 = ~(w17309 | w17415);
assign w17416 = v5483;
assign w17417 = ~w17287 & w17297;
assign v5484 = ~(w17298 | w17417);
assign w17418 = v5484;
assign w17419 = ~w17416 & w17418;
assign w17420 = (~w17298 & w17416) | (~w17298 & w29738) | (w17416 & w29738);
assign w17421 = ~w17275 & w17284;
assign v5485 = ~(w17285 | w17421);
assign w17422 = v5485;
assign w17423 = ~w17420 & w17422;
assign w17424 = (~w17285 & w17420) | (~w17285 & w29877) | (w17420 & w29877);
assign v5486 = ~(w17263 | w17272);
assign w17425 = v5486;
assign v5487 = ~(w17273 | w17425);
assign w17426 = v5487;
assign w17427 = ~w17424 & w17426;
assign w17428 = (~w17273 & w17424) | (~w17273 & w29739) | (w17424 & w29739);
assign w17429 = (~w17260 & ~w17428) | (~w17260 & w30053) | (~w17428 & w30053);
assign w17430 = w17247 & w17429;
assign w17431 = (~w17245 & ~w17247) | (~w17245 & w30823) | (~w17247 & w30823);
assign w17432 = (~w17231 & ~w17431) | (~w17231 & w30187) | (~w17431 & w30187);
assign w17433 = w17218 & w17432;
assign v5488 = ~(w17216 | w17433);
assign w17434 = v5488;
assign w17435 = w17190 & w17200;
assign w17436 = (~w17201 & ~w30366) | (~w17201 & w30824) | (~w30366 & w30824);
assign w17437 = ~w17183 & w17187;
assign v5489 = ~(w17188 | w17437);
assign w17438 = v5489;
assign w17439 = w17436 & w17438;
assign v5490 = ~(w17188 | w17439);
assign w17440 = v5490;
assign w17441 = ~w17439 & w30523;
assign v5491 = ~(w17172 | w17441);
assign w17442 = v5491;
assign w17443 = w17159 & w17442;
assign w17444 = (~w17157 & ~w17159) | (~w17157 & w29740) | (~w17159 & w29740);
assign w17445 = w17131 & ~w17141;
assign v5492 = ~(w17142 | w17445);
assign w17446 = v5492;
assign w17447 = (~w17142 & w17444) | (~w17142 & w30640) | (w17444 & w30640);
assign v5493 = ~(w17122 | w17126);
assign w17448 = v5493;
assign v5494 = ~(w17127 | w17448);
assign w17449 = v5494;
assign w17450 = ~w17447 & w17449;
assign w17451 = (~w17127 & w17447) | (~w17127 & w31049) | (w17447 & w31049);
assign w17452 = (~w17108 & ~w17451) | (~w17108 & w31195) | (~w17451 & w31195);
assign w17453 = w17093 & ~w17452;
assign v5495 = ~(w17091 | w17453);
assign w17454 = v5495;
assign w17455 = ~w17076 & w17454;
assign v5496 = ~(w17075 | w17455);
assign w17456 = v5496;
assign v5497 = ~(w17062 | w17456);
assign w17457 = v5497;
assign v5498 = ~(w17061 | w17457);
assign w17458 = v5498;
assign w17459 = w17048 & ~w17458;
assign v5499 = ~(w17046 | w17459);
assign w17460 = v5499;
assign w17461 = ~w17022 & w17032;
assign v5500 = ~(w17033 | w17461);
assign w17462 = v5500;
assign w17463 = ~w17460 & w17462;
assign v5501 = ~(w17033 | w17463);
assign w17464 = v5501;
assign w17465 = w17020 & ~w17464;
assign w17466 = ~w17020 & w17464;
assign v5502 = ~(w17465 | w17466);
assign w17467 = v5502;
assign w17468 = w7178 & w12167;
assign w17469 = w7765 & w12155;
assign w17470 = w7177 & w11984;
assign w17471 = w7466 & w12084;
assign v5503 = ~(w17470 | w17471);
assign w17472 = v5503;
assign w17473 = ~w17469 & w17472;
assign w17474 = ~w17468 & w17473;
assign w17475 = ~pi11 & w17474;
assign w17476 = pi11 & ~w17474;
assign v5504 = ~(w17475 | w17476);
assign w17477 = v5504;
assign w17478 = w17467 & w17477;
assign v5505 = ~(w17465 | w17478);
assign w17479 = v5505;
assign v5506 = ~(w17018 | w17479);
assign w17480 = v5506;
assign w17481 = w17018 & w17479;
assign v5507 = ~(w17480 | w17481);
assign w17482 = v5507;
assign w17483 = w8141 & w12387;
assign w17484 = w8140 & w12271;
assign w17485 = w8926 & w12381;
assign v5508 = ~(w17484 | w17485);
assign w17486 = v5508;
assign w17487 = w8526 & w12311;
assign w17488 = w17486 & ~w17487;
assign w17489 = ~w17483 & w17488;
assign w17490 = pi08 & w17489;
assign v5509 = ~(pi08 | w17489);
assign w17491 = v5509;
assign v5510 = ~(w17490 | w17491);
assign w17492 = v5510;
assign w17493 = w17482 & ~w17492;
assign v5511 = ~(w17480 | w17493);
assign w17494 = v5511;
assign w17495 = w13697 & ~w17494;
assign w17496 = w16993 & ~w16995;
assign v5512 = ~(w16996 | w17496);
assign w17497 = v5512;
assign w17498 = ~w13697 & w17494;
assign v5513 = ~(w17495 | w17498);
assign w17499 = v5513;
assign w17500 = ~w17497 & w17499;
assign v5514 = ~(w17495 | w17500);
assign w17501 = v5514;
assign v5515 = ~(w17009 | w17011);
assign w17502 = v5515;
assign v5516 = ~(w17012 | w17502);
assign w17503 = v5516;
assign w17504 = ~w17501 & w17503;
assign w17505 = w17501 & ~w17503;
assign v5517 = ~(w17504 | w17505);
assign w17506 = v5517;
assign w17507 = w17497 & ~w17499;
assign v5518 = ~(w17500 | w17507);
assign w17508 = v5518;
assign w17509 = w17460 & ~w17462;
assign v5519 = ~(w17463 | w17509);
assign w17510 = v5519;
assign w17511 = w7178 & w12181;
assign w17512 = w7466 & w11984;
assign w17513 = w7765 & w12084;
assign v5520 = ~(w17512 | w17513);
assign w17514 = v5520;
assign w17515 = w7177 & w11671;
assign w17516 = w17514 & ~w17515;
assign w17517 = ~w17511 & w17516;
assign w17518 = pi11 & w17517;
assign v5521 = ~(pi11 | w17517);
assign w17519 = v5521;
assign v5522 = ~(w17518 | w17519);
assign w17520 = v5522;
assign w17521 = w17510 & ~w17520;
assign w17522 = ~w17510 & w17520;
assign v5523 = ~(w17521 | w17522);
assign w17523 = v5523;
assign w17524 = ~w17048 & w17458;
assign v5524 = ~(w17459 | w17524);
assign w17525 = v5524;
assign w17526 = w7178 & w11993;
assign w17527 = w7466 & w11671;
assign w17528 = w7765 & w11984;
assign v5525 = ~(w17527 | w17528);
assign w17529 = v5525;
assign w17530 = w7177 & w11673;
assign w17531 = w17529 & ~w17530;
assign w17532 = ~w17526 & w17531;
assign v5526 = ~(pi11 | w17532);
assign w17533 = v5526;
assign w17534 = pi11 & w17532;
assign v5527 = ~(w17533 | w17534);
assign w17535 = v5527;
assign w17536 = ~w17525 & w17535;
assign w17537 = w7178 & w12469;
assign w17538 = w7765 & w11671;
assign w17539 = w7466 & w11673;
assign w17540 = w7177 & w11678;
assign v5528 = ~(w17539 | w17540);
assign w17541 = v5528;
assign w17542 = ~w17538 & w17541;
assign w17543 = ~w17537 & w17542;
assign w17544 = pi11 & ~w17543;
assign w17545 = ~pi11 & w17543;
assign v5529 = ~(w17544 | w17545);
assign w17546 = v5529;
assign v5530 = ~(w17061 | w17062);
assign w17547 = v5530;
assign w17548 = w17456 & ~w17547;
assign w17549 = ~w17456 & w17547;
assign v5531 = ~(w17548 | w17549);
assign w17550 = v5531;
assign v5532 = ~(w17546 | w17550);
assign w17551 = v5532;
assign w17552 = w7178 & w12454;
assign w17553 = w7466 & w11678;
assign w17554 = w7765 & w11673;
assign v5533 = ~(w17553 | w17554);
assign w17555 = v5533;
assign w17556 = w7177 & ~w11683;
assign w17557 = w17555 & ~w17556;
assign w17558 = ~w17552 & w17557;
assign v5534 = ~(pi11 | w17558);
assign w17559 = v5534;
assign w17560 = pi11 & w17558;
assign v5535 = ~(w17559 | w17560);
assign w17561 = v5535;
assign v5536 = ~(w17075 | w17076);
assign w17562 = v5536;
assign v5537 = ~(w17454 | w17562);
assign w17563 = v5537;
assign w17564 = w17454 & w17562;
assign v5538 = ~(w17563 | w17564);
assign w17565 = v5538;
assign w17566 = w17561 & ~w17565;
assign w17567 = w9464 & w12594;
assign w17568 = w7765 & w11678;
assign w17569 = w7466 & ~w11683;
assign w17570 = w7177 & w11686;
assign v5539 = ~(w17569 | w17570);
assign w17571 = v5539;
assign w17572 = ~w17568 & w17571;
assign v5540 = ~(pi11 | w17572);
assign w17573 = v5540;
assign v5541 = ~(pi11 | w12594);
assign w17574 = v5541;
assign v5542 = ~(pi11 | w7178);
assign w17575 = v5542;
assign w17576 = w17572 & ~w17575;
assign w17577 = ~w17574 & w17576;
assign v5543 = ~(w17573 | w17577);
assign w17578 = v5543;
assign v5544 = ~(w17567 | w17578);
assign w17579 = v5544;
assign w17580 = ~w17093 & w17452;
assign v5545 = ~(w17453 | w17580);
assign w17581 = v5545;
assign w17582 = w17579 & ~w17581;
assign w17583 = w7765 & ~w11683;
assign w17584 = w7466 & w11686;
assign w17585 = w7177 & w11689;
assign v5546 = ~(w17584 | w17585);
assign w17586 = v5546;
assign w17587 = ~w17583 & w17586;
assign w17588 = pi11 & ~w17587;
assign w17589 = w7178 & w12610;
assign w17590 = ~pi11 & w17587;
assign w17591 = ~w17589 & w17590;
assign w17592 = w9464 & w12610;
assign v5547 = ~(w17591 | w17592);
assign w17593 = v5547;
assign w17594 = ~w17588 & w17593;
assign v5548 = ~(w17108 | w17109);
assign w17595 = v5548;
assign v5549 = ~(w17451 | w17595);
assign w17596 = v5549;
assign w17597 = w17451 & w17595;
assign v5550 = ~(w17596 | w17597);
assign w17598 = v5550;
assign w17599 = ~w17594 & w17598;
assign w17600 = w17594 & ~w17598;
assign v5551 = ~(w17599 | w17600);
assign w17601 = v5551;
assign w17602 = w17447 & ~w17449;
assign v5552 = ~(w17450 | w17602);
assign w17603 = v5552;
assign w17604 = w7178 & ~w12842;
assign w17605 = w7466 & w11689;
assign w17606 = w7765 & w11686;
assign v5553 = ~(w17605 | w17606);
assign w17607 = v5553;
assign w17608 = w7177 & ~w11695;
assign w17609 = w17607 & ~w17608;
assign w17610 = ~w17604 & w17609;
assign w17611 = pi11 & w17610;
assign v5554 = ~(pi11 | w17610);
assign w17612 = v5554;
assign v5555 = ~(w17611 | w17612);
assign w17613 = v5555;
assign w17614 = ~w17603 & w17613;
assign w17615 = w17603 & ~w17613;
assign w17616 = w7765 & w11689;
assign w17617 = w7177 & w11700;
assign w17618 = w7466 & ~w11695;
assign v5556 = ~(w17617 | w17618);
assign w17619 = v5556;
assign w17620 = ~w17616 & w17619;
assign w17621 = (w17620 & ~w12694) | (w17620 & w29741) | (~w12694 & w29741);
assign w17622 = ~pi11 & w17621;
assign w17623 = pi11 & ~w17621;
assign v5557 = ~(w17622 | w17623);
assign w17624 = v5557;
assign w17625 = w17446 & w17624;
assign v5558 = ~(w17446 | w17624);
assign w17626 = v5558;
assign v5559 = ~(w17625 | w17626);
assign w17627 = v5559;
assign w17628 = w17444 & w17627;
assign v5560 = ~(w17444 | w17627);
assign w17629 = v5560;
assign v5561 = ~(w17628 | w17629);
assign w17630 = v5561;
assign v5562 = ~(w17159 | w17442);
assign w17631 = v5562;
assign v5563 = ~(w17443 | w17631);
assign w17632 = v5563;
assign w17633 = w7178 & ~w13008;
assign w17634 = w7765 & ~w11695;
assign w17635 = w7466 & w11700;
assign w17636 = w7177 & w11708;
assign v5564 = ~(w17635 | w17636);
assign w17637 = v5564;
assign w17638 = ~w17634 & w17637;
assign w17639 = ~w17633 & w17638;
assign w17640 = pi11 & w17639;
assign v5565 = ~(pi11 | w17639);
assign w17641 = v5565;
assign v5566 = ~(w17640 | w17641);
assign w17642 = v5566;
assign w17643 = w17632 & ~w17642;
assign w17644 = ~w17632 & w17642;
assign w17645 = w7765 & w11700;
assign w17646 = w7466 & w11708;
assign w17647 = w7177 & w11711;
assign v5567 = ~(w17646 | w17647);
assign w17648 = v5567;
assign w17649 = ~w17645 & w17648;
assign w17650 = pi11 & ~w17649;
assign w17651 = w7178 & w12994;
assign w17652 = ~pi11 & w17649;
assign w17653 = ~w17651 & w17652;
assign w17654 = w9464 & w12994;
assign v5568 = ~(w17653 | w17654);
assign w17655 = v5568;
assign w17656 = ~w17650 & w17655;
assign v5569 = ~(w17172 | w17173);
assign w17657 = v5569;
assign v5570 = ~(w17440 | w17657);
assign w17658 = v5570;
assign w17659 = w17440 & w17657;
assign v5571 = ~(w17658 | w17659);
assign w17660 = v5571;
assign w17661 = w17656 & ~w17660;
assign w17662 = ~w17656 & w17660;
assign v5572 = ~(w17661 | w17662);
assign w17663 = v5572;
assign v5573 = ~(w17436 | w17438);
assign w17664 = v5573;
assign v5574 = ~(w17439 | w17664);
assign w17665 = v5574;
assign w17666 = w7178 & w13178;
assign w17667 = w7765 & w11708;
assign w17668 = w7177 & w11714;
assign w17669 = w7466 & w11711;
assign v5575 = ~(w17668 | w17669);
assign w17670 = v5575;
assign w17671 = ~w17667 & w17670;
assign w17672 = ~w17666 & w17671;
assign w17673 = ~pi11 & w17672;
assign w17674 = pi11 & ~w17672;
assign v5576 = ~(w17673 | w17674);
assign w17675 = v5576;
assign v5577 = ~(w17665 | w17675);
assign w17676 = v5577;
assign w17677 = w17665 & w17675;
assign w17678 = w7178 & w13194;
assign w17679 = w7765 & w11711;
assign w17680 = w7177 & w11720;
assign w17681 = w7466 & w11714;
assign v5578 = ~(w17680 | w17681);
assign w17682 = v5578;
assign w17683 = ~w17679 & w17682;
assign w17684 = ~w17678 & w17683;
assign w17685 = pi11 & ~w17684;
assign w17686 = ~pi11 & w17684;
assign v5579 = ~(w17685 | w17686);
assign w17687 = v5579;
assign v5580 = ~(w17201 | w17435);
assign w17688 = v5580;
assign w17689 = w17434 & ~w17688;
assign w17690 = ~w17434 & w17688;
assign v5581 = ~(w17689 | w17690);
assign w17691 = v5581;
assign w17692 = w17687 & w17691;
assign v5582 = ~(w17687 | w17691);
assign w17693 = v5582;
assign v5583 = ~(w17692 | w17693);
assign w17694 = v5583;
assign v5584 = ~(w17218 | w17432);
assign w17695 = v5584;
assign v5585 = ~(w17433 | w17695);
assign w17696 = v5585;
assign w17697 = w7178 & w13514;
assign w17698 = w7765 & w11714;
assign w17699 = w7177 & w11723;
assign w17700 = w7466 & w11720;
assign v5586 = ~(w17699 | w17700);
assign w17701 = v5586;
assign w17702 = ~w17698 & w17701;
assign w17703 = ~w17697 & w17702;
assign w17704 = pi11 & ~w17703;
assign w17705 = ~pi11 & w17703;
assign v5587 = ~(w17704 | w17705);
assign w17706 = v5587;
assign v5588 = ~(w17696 | w17706);
assign w17707 = v5588;
assign w17708 = w17696 & w17706;
assign w17709 = w7178 & ~w13310;
assign w17710 = w7765 & w11720;
assign w17711 = w7466 & w11723;
assign w17712 = w7177 & w11726;
assign v5589 = ~(w17711 | w17712);
assign w17713 = v5589;
assign w17714 = ~w17710 & w17713;
assign w17715 = ~w17709 & w17714;
assign w17716 = ~pi11 & w17715;
assign w17717 = pi11 & ~w17715;
assign v5590 = ~(w17716 | w17717);
assign w17718 = v5590;
assign v5591 = ~(w17231 | w17232);
assign w17719 = v5591;
assign w17720 = w17431 & w17719;
assign v5592 = ~(w17431 | w17719);
assign w17721 = v5592;
assign v5593 = ~(w17720 | w17721);
assign w17722 = v5593;
assign w17723 = w17718 & ~w17722;
assign w17724 = ~w17718 & w17722;
assign v5594 = ~(w17723 | w17724);
assign w17725 = v5594;
assign v5595 = ~(w17247 | w17429);
assign w17726 = v5595;
assign v5596 = ~(w17430 | w17726);
assign w17727 = v5596;
assign w17728 = w7178 & ~w13737;
assign w17729 = w7765 & w11723;
assign w17730 = w7177 & w11729;
assign w17731 = w7466 & w11726;
assign v5597 = ~(w17730 | w17731);
assign w17732 = v5597;
assign w17733 = ~w17729 & w17732;
assign w17734 = ~w17728 & w17733;
assign w17735 = pi11 & ~w17734;
assign w17736 = ~pi11 & w17734;
assign v5598 = ~(w17735 | w17736);
assign w17737 = v5598;
assign v5599 = ~(w17727 | w17737);
assign w17738 = v5599;
assign w17739 = w17727 & w17737;
assign v5600 = ~(w17260 | w17261);
assign w17740 = v5600;
assign w17741 = w17428 & w17740;
assign v5601 = ~(w17428 | w17740);
assign w17742 = v5601;
assign v5602 = ~(w17741 | w17742);
assign w17743 = v5602;
assign w17744 = w7178 & w13864;
assign w17745 = w7466 & w11729;
assign w17746 = w7765 & w11726;
assign v5603 = ~(w17745 | w17746);
assign w17747 = v5603;
assign w17748 = w7177 & ~w11734;
assign w17749 = w17747 & ~w17748;
assign w17750 = ~w17744 & w17749;
assign v5604 = ~(pi11 | w17750);
assign w17751 = v5604;
assign w17752 = pi11 & w17750;
assign v5605 = ~(w17751 | w17752);
assign w17753 = v5605;
assign v5606 = ~(w17743 | w17753);
assign w17754 = v5606;
assign w17755 = w17743 & w17753;
assign v5607 = ~(w17754 | w17755);
assign w17756 = v5607;
assign w17757 = w17424 & ~w17426;
assign v5608 = ~(w17427 | w17757);
assign w17758 = v5608;
assign w17759 = w7178 & ~w13703;
assign w17760 = w7765 & w11729;
assign w17761 = w7177 & w11737;
assign w17762 = w7466 & ~w11734;
assign v5609 = ~(w17761 | w17762);
assign w17763 = v5609;
assign w17764 = ~w17760 & w17763;
assign w17765 = ~w17759 & w17764;
assign w17766 = pi11 & w17765;
assign v5610 = ~(pi11 | w17765);
assign w17767 = v5610;
assign v5611 = ~(w17766 | w17767);
assign w17768 = v5611;
assign w17769 = ~w17758 & w17768;
assign w17770 = w17758 & ~w17768;
assign w17771 = w17420 & ~w17422;
assign v5612 = ~(w17423 | w17771);
assign w17772 = v5612;
assign w17773 = w7178 & w13882;
assign w17774 = w7466 & w11737;
assign w17775 = w7765 & ~w11734;
assign v5613 = ~(w17774 | w17775);
assign w17776 = v5613;
assign w17777 = w7177 & w11740;
assign w17778 = w17776 & ~w17777;
assign w17779 = ~w17773 & w17778;
assign w17780 = pi11 & w17779;
assign v5614 = ~(pi11 | w17779);
assign w17781 = v5614;
assign v5615 = ~(w17780 | w17781);
assign w17782 = v5615;
assign w17783 = w17772 & ~w17782;
assign w17784 = ~w17772 & w17782;
assign v5616 = ~(w17783 | w17784);
assign w17785 = v5616;
assign w17786 = w17416 & ~w17418;
assign v5617 = ~(w17419 | w17786);
assign w17787 = v5617;
assign w17788 = ~w14287 & w29742;
assign w17789 = w7765 & w11737;
assign w17790 = w7177 & ~w11745;
assign w17791 = w7466 & w11740;
assign v5618 = ~(w17790 | w17791);
assign w17792 = v5618;
assign w17793 = ~w17789 & w17792;
assign w17794 = ~w17788 & w17793;
assign w17795 = pi11 & ~w17794;
assign w17796 = ~pi11 & w17794;
assign v5619 = ~(w17795 | w17796);
assign w17797 = v5619;
assign v5620 = ~(w17787 | w17797);
assign w17798 = v5620;
assign w17799 = w17787 & w17797;
assign w17800 = w17412 & ~w17414;
assign v5621 = ~(w17415 | w17800);
assign w17801 = v5621;
assign w17802 = w7765 & w11740;
assign w17803 = w7466 & ~w11745;
assign w17804 = w7177 & w11748;
assign v5622 = ~(w17803 | w17804);
assign w17805 = v5622;
assign w17806 = ~w17802 & w17805;
assign w17807 = (w17806 & ~w14300) | (w17806 & w29743) | (~w14300 & w29743);
assign w17808 = pi11 & w17807;
assign v5623 = ~(pi11 | w17807);
assign w17809 = v5623;
assign v5624 = ~(w17808 | w17809);
assign w17810 = v5624;
assign w17811 = w17801 & ~w17810;
assign w17812 = w17408 & ~w17410;
assign v5625 = ~(w17411 | w17812);
assign w17813 = v5625;
assign w17814 = w7466 & w11748;
assign w17815 = w7765 & ~w11745;
assign v5626 = ~(w17814 | w17815);
assign w17816 = v5626;
assign w17817 = w7177 & w11759;
assign w17818 = w17816 & ~w17817;
assign w17819 = (w17818 & ~w13948) | (w17818 & w29744) | (~w13948 & w29744);
assign w17820 = pi11 & w17819;
assign v5627 = ~(pi11 | w17819);
assign w17821 = v5627;
assign v5628 = ~(w17820 | w17821);
assign w17822 = v5628;
assign w17823 = w17813 & ~w17822;
assign w17824 = w17404 & ~w17406;
assign v5629 = ~(w17407 | w17824);
assign w17825 = v5629;
assign w17826 = (w7178 & w11841) | (w7178 & w29515) | (w11841 & w29515);
assign w17827 = w7765 & w11748;
assign w17828 = w7466 & w11759;
assign w17829 = w7177 & w11761;
assign v5630 = ~(w17828 | w17829);
assign w17830 = v5630;
assign w17831 = ~w17827 & w17830;
assign w17832 = ~w17826 & w29745;
assign w17833 = (~pi11 & w17826) | (~pi11 & w29746) | (w17826 & w29746);
assign v5631 = ~(w17832 | w17833);
assign w17834 = v5631;
assign w17835 = w17825 & ~w17834;
assign w17836 = w17400 & ~w17402;
assign v5632 = ~(w17403 | w17836);
assign w17837 = v5632;
assign w17838 = w7177 & ~w11771;
assign w17839 = w7765 & w11759;
assign w17840 = w7466 & w11761;
assign v5633 = ~(w17839 | w17840);
assign w17841 = v5633;
assign w17842 = ~w17838 & w17841;
assign w17843 = (w14356 & w29516) | (w14356 & w29517) | (w29516 & w29517);
assign w17844 = (~w14356 & w29518) | (~w14356 & w29519) | (w29518 & w29519);
assign v5634 = ~(w17843 | w17844);
assign w17845 = v5634;
assign w17846 = w17837 & w17845;
assign w17847 = w17396 & ~w17398;
assign v5635 = ~(w17399 | w17847);
assign w17848 = v5635;
assign w17849 = w7466 & ~w11771;
assign w17850 = w7177 & w11768;
assign w17851 = (~w17850 & ~w11761) | (~w17850 & w29011) | (~w11761 & w29011);
assign w17852 = ~w17849 & w17851;
assign w17853 = (w14383 & w29012) | (w14383 & w29013) | (w29012 & w29013);
assign w17854 = (~w14383 & w29014) | (~w14383 & w29015) | (w29014 & w29015);
assign v5636 = ~(w17853 | w17854);
assign w17855 = v5636;
assign w17856 = w17848 & w17855;
assign w17857 = w17392 & ~w17394;
assign v5637 = ~(w17395 | w17857);
assign w17858 = v5637;
assign w17859 = w7466 & w11768;
assign w17860 = (w7765 & ~w11766) | (w7765 & w28756) | (~w11766 & w28756);
assign v5638 = ~(w17859 | w17860);
assign w17861 = v5638;
assign w17862 = w7177 & w11776;
assign w17863 = (w28757 & ~w14409) | (w28757 & w30367) | (~w14409 & w30367);
assign w17864 = (w14409 & w30368) | (w14409 & w30369) | (w30368 & w30369);
assign v5639 = ~(w17863 | w17864);
assign w17865 = v5639;
assign w17866 = w17858 & ~w17865;
assign v5640 = ~(w17382 | w17390);
assign w17867 = v5640;
assign v5641 = ~(w17391 | w17867);
assign w17868 = v5641;
assign w17869 = w11533 & w29016;
assign w17870 = w7177 & w11784;
assign w17871 = w7466 & w11776;
assign v5642 = ~(w17870 | w17871);
assign w17872 = v5642;
assign w17873 = (w14461 & w28508) | (w14461 & w28509) | (w28508 & w28509);
assign w17874 = (~w14461 & w28510) | (~w14461 & w28511) | (w28510 & w28511);
assign v5643 = ~(w17873 | w17874);
assign w17875 = v5643;
assign w17876 = w17868 & w17875;
assign w17877 = pi14 & ~w17371;
assign v5644 = ~(w17377 | w17877);
assign w17878 = v5644;
assign w17879 = w17377 & w17877;
assign v5645 = ~(w17878 | w17879);
assign w17880 = v5645;
assign w17881 = w7466 & w11784;
assign w17882 = w7765 & w11776;
assign v5646 = ~(w17881 | w17882);
assign w17883 = v5646;
assign w17884 = w7177 & w11793;
assign w17885 = (w14504 & w28512) | (w14504 & w28513) | (w28512 & w28513);
assign w17886 = (~w14504 & w28514) | (~w14504 & w28515) | (w28514 & w28515);
assign v5647 = ~(w17885 | w17886);
assign w17887 = v5647;
assign v5648 = ~(w17880 | w17887);
assign w17888 = v5648;
assign w17889 = w17365 & ~w17370;
assign v5649 = ~(w17371 | w17889);
assign w17890 = v5649;
assign w17891 = w7178 & w14547;
assign w17892 = w7177 & w11803;
assign w17893 = w7765 & w11784;
assign w17894 = w7466 & w11793;
assign v5650 = ~(w17893 | w17894);
assign w17895 = v5650;
assign w17896 = (pi11 & w17891) | (pi11 & w28328) | (w17891 & w28328);
assign w17897 = ~w17891 & w28329;
assign v5651 = ~(w17896 | w17897);
assign w17898 = v5651;
assign w17899 = w17890 & w17898;
assign w17900 = w7172 & w11800;
assign w17901 = pi11 & w17900;
assign w17902 = w7178 & ~w14609;
assign w17903 = w7765 & w11798;
assign w17904 = w7466 & w11800;
assign v5652 = ~(w17903 | w17904);
assign w17905 = v5652;
assign w17906 = ~w17902 & w17905;
assign w17907 = ~w17901 & w17906;
assign w17908 = pi11 & ~w17907;
assign w17909 = w7177 & w11800;
assign w17910 = (~w17909 & w14639) | (~w17909 & w28516) | (w14639 & w28516);
assign w17911 = w7765 & w11803;
assign w17912 = w7466 & w11798;
assign v5653 = ~(w17911 | w17912);
assign w17913 = v5653;
assign w17914 = w17910 & w17913;
assign w17915 = ~w17908 & w17914;
assign w17916 = pi11 & w17915;
assign w17917 = w17364 & w17916;
assign v5654 = ~(w17364 | w17916);
assign w17918 = v5654;
assign v5655 = ~(w17917 | w17918);
assign w17919 = v5655;
assign w17920 = w7178 & w14569;
assign w17921 = w7177 & w11798;
assign w17922 = w7765 & w11793;
assign w17923 = w7466 & w11803;
assign v5656 = ~(w17922 | w17923);
assign w17924 = v5656;
assign w17925 = (pi11 & w17920) | (pi11 & w28517) | (w17920 & w28517);
assign w17926 = ~w17920 & w28518;
assign v5657 = ~(w17925 | w17926);
assign w17927 = v5657;
assign w17928 = w17919 & w17927;
assign v5658 = ~(w17917 | w17928);
assign w17929 = v5658;
assign v5659 = ~(w17890 | w17898);
assign w17930 = v5659;
assign v5660 = ~(w17899 | w17930);
assign w17931 = v5660;
assign w17932 = ~w17929 & w17931;
assign w17933 = (~w17899 & ~w17931) | (~w17899 & w28519) | (~w17931 & w28519);
assign w17934 = w17880 & w17887;
assign v5661 = ~(w17888 | w17934);
assign w17935 = v5661;
assign w17936 = ~w17933 & w17935;
assign v5662 = ~(w17888 | w17936);
assign w17937 = v5662;
assign v5663 = ~(w17868 | w17875);
assign w17938 = v5663;
assign v5664 = ~(w17876 | w17938);
assign w17939 = v5664;
assign w17940 = ~w17937 & w17939;
assign w17941 = (~w17876 & w17937) | (~w17876 & w28759) | (w17937 & w28759);
assign w17942 = ~w17858 & w17865;
assign v5665 = ~(w17866 | w17942);
assign w17943 = v5665;
assign w17944 = ~w17941 & w17943;
assign w17945 = (~w17866 & w17941) | (~w17866 & w29520) | (w17941 & w29520);
assign v5666 = ~(w17848 | w17855);
assign w17946 = v5666;
assign v5667 = ~(w17856 | w17946);
assign w17947 = v5667;
assign w17948 = ~w17945 & w17947;
assign w17949 = (~w17856 & w17945) | (~w17856 & w29017) | (w17945 & w29017);
assign v5668 = ~(w17837 | w17845);
assign w17950 = v5668;
assign v5669 = ~(w17846 | w17950);
assign w17951 = v5669;
assign w17952 = ~w17949 & w17951;
assign w17953 = (~w17846 & w17949) | (~w17846 & w29521) | (w17949 & w29521);
assign w17954 = ~w17825 & w17834;
assign v5670 = ~(w17835 | w17954);
assign w17955 = v5670;
assign w17956 = ~w17953 & w17955;
assign w17957 = (~w17835 & w17953) | (~w17835 & w29878) | (w17953 & w29878);
assign w17958 = ~w17813 & w17822;
assign v5671 = ~(w17823 | w17958);
assign w17959 = v5671;
assign w17960 = ~w17957 & w17959;
assign w17961 = (~w17823 & w17957) | (~w17823 & w29747) | (w17957 & w29747);
assign w17962 = ~w17801 & w17810;
assign v5672 = ~(w17811 | w17962);
assign w17963 = v5672;
assign w17964 = ~w17961 & w17963;
assign w17965 = (~w17811 & w17961) | (~w17811 & w29522) | (w17961 & w29522);
assign w17966 = (~w17798 & ~w17965) | (~w17798 & w29018) | (~w17965 & w29018);
assign w17967 = w17785 & w17966;
assign w17968 = (~w17783 & ~w17785) | (~w17783 & w29019) | (~w17785 & w29019);
assign w17969 = (~w17769 & ~w17968) | (~w17769 & w29748) | (~w17968 & w29748);
assign w17970 = w17756 & w17969;
assign w17971 = (~w17754 & ~w17756) | (~w17754 & w29020) | (~w17756 & w29020);
assign w17972 = (w29020 & w30054) | (w29020 & w30055) | (w30054 & w30055);
assign v5673 = ~(w17738 | w17972);
assign w17973 = v5673;
assign w17974 = w17725 & w17973;
assign w17975 = (~w17723 & ~w17973) | (~w17723 & w30825) | (~w17973 & w30825);
assign w17976 = (~w29021 & w30826) | (~w29021 & w30827) | (w30826 & w30827);
assign w17977 = w17694 & w17976;
assign w17978 = (~w17692 & ~w17694) | (~w17692 & w29022) | (~w17694 & w29022);
assign w17979 = (w29022 & w30370) | (w29022 & w30371) | (w30370 & w30371);
assign v5674 = ~(w17676 | w17979);
assign w17980 = v5674;
assign w17981 = w17663 & w17980;
assign w17982 = (~w17661 & ~w17663) | (~w17661 & w29023) | (~w17663 & w29023);
assign w17983 = (~w17643 & w17982) | (~w17643 & w30524) | (w17982 & w30524);
assign v5675 = ~(w17630 | w17983);
assign w17984 = v5675;
assign w17985 = (w17624 & w17444) | (w17624 & w31050) | (w17444 & w31050);
assign w17986 = ~w17628 & w17985;
assign w17987 = (~w17986 & w17983) | (~w17986 & w30641) | (w17983 & w30641);
assign w17988 = (~w17614 & ~w17987) | (~w17614 & w29024) | (~w17987 & w29024);
assign w17989 = w17601 & ~w17988;
assign w17990 = (~w17599 & ~w17601) | (~w17599 & w29025) | (~w17601 & w29025);
assign w17991 = ~w17579 & w17581;
assign v5676 = ~(w17582 | w17991);
assign w17992 = v5676;
assign w17993 = w17990 & w17992;
assign w17994 = (~w17582 & ~w17990) | (~w17582 & w31196) | (~w17990 & w31196);
assign w17995 = ~w17561 & w17565;
assign v5677 = ~(w17566 | w17995);
assign w17996 = v5677;
assign w17997 = w17994 & w17996;
assign w17998 = (~w17566 & ~w17996) | (~w17566 & w29026) | (~w17996 & w29026);
assign w17999 = w17546 & w17550;
assign v5678 = ~(w17551 | w17999);
assign w18000 = v5678;
assign w18001 = ~w17998 & w18000;
assign w18002 = (~w17551 & ~w18000) | (~w17551 & w29027) | (~w18000 & w29027);
assign w18003 = w17525 & ~w17535;
assign v5679 = ~(w17536 | w18003);
assign w18004 = v5679;
assign w18005 = ~w18002 & w18004;
assign w18006 = (~w17536 & ~w18004) | (~w17536 & w29028) | (~w18004 & w29028);
assign w18007 = w17523 & w18006;
assign w18008 = w8526 & w12271;
assign w18009 = w8926 & w12311;
assign v5680 = ~(w18008 | w18009);
assign w18010 = v5680;
assign w18011 = w8140 & w12237;
assign w18012 = w18010 & ~w18011;
assign w18013 = (~w12318 & w29523) | (~w12318 & w29524) | (w29523 & w29524);
assign w18014 = (w12318 & w29525) | (w12318 & w29526) | (w29525 & w29526);
assign v5681 = ~(w18013 | w18014);
assign w18015 = v5681;
assign w18016 = (~w29029 & w31051) | (~w29029 & w31052) | (w31051 & w31052);
assign v5682 = ~(w17467 | w17477);
assign w18017 = v5682;
assign v5683 = ~(w17478 | w18017);
assign w18018 = v5683;
assign w18019 = (w29029 & w31053) | (w29029 & w31054) | (w31053 & w31054);
assign v5684 = ~(w18016 | w18019);
assign w18020 = v5684;
assign w18021 = w18018 & w18020;
assign w18022 = (~w18016 & ~w18020) | (~w18016 & w29527) | (~w18020 & w29527);
assign w18023 = pi05 & w12406;
assign w18024 = pi04 & ~w12406;
assign v5685 = ~(w18023 | w18024);
assign w18025 = v5685;
assign w18026 = w9400 & w18025;
assign v5686 = ~(w13695 | w18026);
assign w18027 = v5686;
assign w18028 = w18022 & ~w18027;
assign w18029 = ~w17482 & w17492;
assign v5687 = ~(w17493 | w18029);
assign w18030 = v5687;
assign w18031 = ~w18022 & w18027;
assign v5688 = ~(w18028 | w18031);
assign w18032 = v5688;
assign w18033 = ~w18030 & w18032;
assign v5689 = ~(w18028 | w18033);
assign w18034 = v5689;
assign w18035 = w17508 & w18034;
assign v5690 = ~(w18018 | w18020);
assign w18036 = v5690;
assign v5691 = ~(w18021 | w18036);
assign w18037 = v5691;
assign v5692 = ~(w17523 | w18006);
assign w18038 = v5692;
assign v5693 = ~(w18007 | w18038);
assign w18039 = v5693;
assign w18040 = w8141 & ~w12277;
assign w18041 = w8926 & w12271;
assign w18042 = w8140 & w12155;
assign w18043 = w8526 & w12237;
assign v5694 = ~(w18042 | w18043);
assign w18044 = v5694;
assign w18045 = ~w18041 & w18044;
assign w18046 = ~w18040 & w18045;
assign w18047 = pi08 & w18046;
assign v5695 = ~(pi08 | w18046);
assign w18048 = v5695;
assign v5696 = ~(w18047 | w18048);
assign w18049 = v5696;
assign w18050 = w18039 & ~w18049;
assign w18051 = w18002 & ~w18004;
assign v5697 = ~(w18005 | w18051);
assign w18052 = v5697;
assign w18053 = w8141 & ~w12351;
assign w18054 = w8926 & w12237;
assign w18055 = w8140 & w12084;
assign w18056 = w8526 & w12155;
assign v5698 = ~(w18055 | w18056);
assign w18057 = v5698;
assign w18058 = ~w18054 & w18057;
assign w18059 = ~w18053 & w18058;
assign w18060 = pi08 & ~w18059;
assign w18061 = ~pi08 & w18059;
assign v5699 = ~(w18060 | w18061);
assign w18062 = v5699;
assign w18063 = w18052 & ~w18062;
assign w18064 = w17998 & ~w18000;
assign v5700 = ~(w18001 | w18064);
assign w18065 = v5700;
assign w18066 = w8141 & w12167;
assign w18067 = w8140 & w11984;
assign w18068 = w8926 & w12155;
assign v5701 = ~(w18067 | w18068);
assign w18069 = v5701;
assign w18070 = w8526 & w12084;
assign w18071 = w18069 & ~w18070;
assign w18072 = ~w18066 & w18071;
assign w18073 = pi08 & w18072;
assign v5702 = ~(pi08 | w18072);
assign w18074 = v5702;
assign v5703 = ~(w18073 | w18074);
assign w18075 = v5703;
assign v5704 = ~(w18065 | w18075);
assign w18076 = v5704;
assign w18077 = w18065 & w18075;
assign v5705 = ~(w18076 | w18077);
assign w18078 = v5705;
assign v5706 = ~(w17994 | w17996);
assign w18079 = v5706;
assign v5707 = ~(w17997 | w18079);
assign w18080 = v5707;
assign w18081 = w8141 & w12181;
assign w18082 = w8526 & w11984;
assign w18083 = w8926 & w12084;
assign v5708 = ~(w18082 | w18083);
assign w18084 = v5708;
assign w18085 = w8140 & w11671;
assign w18086 = w18084 & ~w18085;
assign w18087 = ~w18081 & w18086;
assign v5709 = ~(pi08 | w18087);
assign w18088 = v5709;
assign w18089 = pi08 & w18087;
assign v5710 = ~(w18088 | w18089);
assign w18090 = v5710;
assign v5711 = ~(w18080 | w18090);
assign w18091 = v5711;
assign w18092 = w18080 & w18090;
assign v5712 = ~(w18091 | w18092);
assign w18093 = v5712;
assign v5713 = ~(w17990 | w17992);
assign w18094 = v5713;
assign v5714 = ~(w17993 | w18094);
assign w18095 = v5714;
assign w18096 = ~w11992 & w29528;
assign w18097 = w8926 & w11984;
assign w18098 = w8526 & w11671;
assign w18099 = w8140 & w11673;
assign v5715 = ~(w18098 | w18099);
assign w18100 = v5715;
assign w18101 = ~w18097 & w18100;
assign w18102 = ~w18096 & w18101;
assign w18103 = ~pi08 & w18102;
assign w18104 = pi08 & ~w18102;
assign v5716 = ~(w18103 | w18104);
assign w18105 = v5716;
assign w18106 = w18095 & w18105;
assign v5717 = ~(w18095 | w18105);
assign w18107 = v5717;
assign v5718 = ~(w18106 | w18107);
assign w18108 = v5718;
assign w18109 = w9920 & w12469;
assign w18110 = w8926 & w11671;
assign w18111 = w8526 & w11673;
assign w18112 = w8140 & w11678;
assign v5719 = ~(w18111 | w18112);
assign w18113 = v5719;
assign w18114 = ~w18110 & w18113;
assign w18115 = pi08 & ~w18114;
assign w18116 = ~pi08 & w18114;
assign w18117 = (w18116 & ~w12469) | (w18116 & w29529) | (~w12469 & w29529);
assign v5720 = ~(w18115 | w18117);
assign w18118 = v5720;
assign w18119 = ~w18109 & w18118;
assign w18120 = ~w17601 & w17988;
assign v5721 = ~(w17989 | w18120);
assign w18121 = v5721;
assign w18122 = ~w18119 & w18121;
assign w18123 = w18119 & ~w18121;
assign w18124 = w9920 & w12454;
assign w18125 = w8926 & w11673;
assign w18126 = w8526 & w11678;
assign w18127 = w8140 & ~w11683;
assign v5722 = ~(w18126 | w18127);
assign w18128 = v5722;
assign w18129 = ~w18125 & w18128;
assign w18130 = pi08 & ~w18129;
assign w18131 = ~pi08 & w18129;
assign w18132 = (w18131 & ~w12454) | (w18131 & w29530) | (~w12454 & w29530);
assign v5723 = ~(w18130 | w18132);
assign w18133 = v5723;
assign w18134 = ~w18124 & w18133;
assign v5724 = ~(w17614 | w17615);
assign w18135 = v5724;
assign w18136 = w17987 & w18135;
assign v5725 = ~(w17987 | w18135);
assign w18137 = v5725;
assign v5726 = ~(w18136 | w18137);
assign w18138 = v5726;
assign w18139 = w18134 & ~w18138;
assign w18140 = ~w18134 & w18138;
assign v5727 = ~(w18139 | w18140);
assign w18141 = v5727;
assign w18142 = w9920 & w12594;
assign w18143 = w8926 & w11678;
assign w18144 = w8526 & ~w11683;
assign w18145 = w8140 & w11686;
assign v5728 = ~(w18144 | w18145);
assign w18146 = v5728;
assign w18147 = ~w18143 & w18146;
assign w18148 = pi08 & ~w18147;
assign w18149 = ~pi08 & w18147;
assign w18150 = (w18149 & ~w12594) | (w18149 & w29531) | (~w12594 & w29531);
assign v5729 = ~(w18148 | w18150);
assign w18151 = v5729;
assign w18152 = ~w18142 & w18151;
assign w18153 = w17630 & w17983;
assign v5730 = ~(w17984 | w18153);
assign w18154 = v5730;
assign v5731 = ~(w18152 | w18154);
assign w18155 = v5731;
assign w18156 = w18152 & w18154;
assign w18157 = w9920 & w12610;
assign w18158 = w8926 & ~w11683;
assign w18159 = w8526 & w11686;
assign w18160 = w8140 & w11689;
assign v5732 = ~(w18159 | w18160);
assign w18161 = v5732;
assign w18162 = ~w18158 & w18161;
assign w18163 = pi08 & ~w18162;
assign w18164 = w8141 & w12610;
assign w18165 = ~pi08 & w18162;
assign w18166 = ~w18164 & w18165;
assign v5733 = ~(w18163 | w18166);
assign w18167 = v5733;
assign w18168 = ~w18157 & w18167;
assign v5734 = ~(w17643 | w17644);
assign w18169 = v5734;
assign w18170 = w17982 & ~w18169;
assign w18171 = ~w17982 & w18169;
assign v5735 = ~(w18170 | w18171);
assign w18172 = v5735;
assign w18173 = w18168 & w18172;
assign v5736 = ~(w18168 | w18172);
assign w18174 = v5736;
assign v5737 = ~(w18173 | w18174);
assign w18175 = v5737;
assign w18176 = w9920 & ~w12842;
assign w18177 = w8926 & w11686;
assign w18178 = w8526 & w11689;
assign w18179 = w8140 & ~w11695;
assign v5738 = ~(w18178 | w18179);
assign w18180 = v5738;
assign w18181 = ~w18177 & w18180;
assign w18182 = pi08 & ~w18181;
assign w18183 = w8141 & ~w12842;
assign w18184 = ~pi08 & w18181;
assign w18185 = ~w18183 & w18184;
assign v5739 = ~(w18182 | w18185);
assign w18186 = v5739;
assign w18187 = ~w18176 & w18186;
assign v5740 = ~(w17663 | w17980);
assign w18188 = v5740;
assign v5741 = ~(w17981 | w18188);
assign w18189 = v5741;
assign v5742 = ~(w18187 | w18189);
assign w18190 = v5742;
assign w18191 = w18187 & w18189;
assign w18192 = w8141 & w12694;
assign w18193 = w8926 & w11689;
assign w18194 = w8140 & w11700;
assign w18195 = w8526 & ~w11695;
assign v5743 = ~(w18194 | w18195);
assign w18196 = v5743;
assign w18197 = ~w18193 & w18196;
assign w18198 = ~w18192 & w18197;
assign w18199 = ~pi08 & w18198;
assign w18200 = pi08 & ~w18198;
assign v5744 = ~(w18199 | w18200);
assign w18201 = v5744;
assign v5745 = ~(w17676 | w17677);
assign w18202 = v5745;
assign v5746 = ~(w17978 | w18202);
assign w18203 = v5746;
assign w18204 = w17978 & w18202;
assign v5747 = ~(w18203 | w18204);
assign w18205 = v5747;
assign w18206 = w18201 & ~w18205;
assign w18207 = ~w18201 & w18205;
assign v5748 = ~(w18206 | w18207);
assign w18208 = v5748;
assign v5749 = ~(w17694 | w17976);
assign w18209 = v5749;
assign v5750 = ~(w17977 | w18209);
assign w18210 = v5750;
assign w18211 = w8141 & ~w13008;
assign w18212 = w8926 & ~w11695;
assign w18213 = w8526 & w11700;
assign w18214 = w8140 & w11708;
assign v5751 = ~(w18213 | w18214);
assign w18215 = v5751;
assign w18216 = ~w18212 & w18215;
assign w18217 = ~w18211 & w18216;
assign w18218 = pi08 & ~w18217;
assign w18219 = ~pi08 & w18217;
assign v5752 = ~(w18218 | w18219);
assign w18220 = v5752;
assign w18221 = w18210 & w18220;
assign v5753 = ~(w18210 | w18220);
assign w18222 = v5753;
assign w18223 = w8926 & w11700;
assign w18224 = w8526 & w11708;
assign w18225 = w8140 & w11711;
assign v5754 = ~(w18224 | w18225);
assign w18226 = v5754;
assign w18227 = ~w18223 & w18226;
assign w18228 = pi08 & ~w18227;
assign w18229 = w8141 & w12994;
assign w18230 = ~pi08 & w18227;
assign w18231 = ~w18229 & w18230;
assign w18232 = w9920 & w12994;
assign v5755 = ~(w18231 | w18232);
assign w18233 = v5755;
assign w18234 = ~w18228 & w18233;
assign v5756 = ~(w17707 | w17708);
assign w18235 = v5756;
assign w18236 = w17975 & w18235;
assign v5757 = ~(w17975 | w18235);
assign w18237 = v5757;
assign v5758 = ~(w18236 | w18237);
assign w18238 = v5758;
assign w18239 = w18234 & ~w18238;
assign w18240 = ~w18234 & w18238;
assign v5759 = ~(w18239 | w18240);
assign w18241 = v5759;
assign v5760 = ~(w17725 | w17973);
assign w18242 = v5760;
assign v5761 = ~(w17974 | w18242);
assign w18243 = v5761;
assign w18244 = w8141 & w13178;
assign w18245 = w8926 & w11708;
assign w18246 = w8140 & w11714;
assign w18247 = w8526 & w11711;
assign v5762 = ~(w18246 | w18247);
assign w18248 = v5762;
assign w18249 = ~w18245 & w18248;
assign w18250 = ~w18244 & w18249;
assign w18251 = ~pi08 & w18250;
assign w18252 = pi08 & ~w18250;
assign v5763 = ~(w18251 | w18252);
assign w18253 = v5763;
assign v5764 = ~(w18243 | w18253);
assign w18254 = v5764;
assign w18255 = w18243 & w18253;
assign w18256 = w8141 & w13194;
assign w18257 = w8140 & w11720;
assign w18258 = w8926 & w11711;
assign v5765 = ~(w18257 | w18258);
assign w18259 = v5765;
assign w18260 = w8526 & w11714;
assign w18261 = w18259 & ~w18260;
assign w18262 = ~w18256 & w18261;
assign v5766 = ~(pi08 | w18262);
assign w18263 = v5766;
assign w18264 = pi08 & w18262;
assign v5767 = ~(w18263 | w18264);
assign w18265 = v5767;
assign v5768 = ~(w17738 | w17739);
assign w18266 = v5768;
assign w18267 = w17971 & w18266;
assign v5769 = ~(w17971 | w18266);
assign w18268 = v5769;
assign v5770 = ~(w18267 | w18268);
assign w18269 = v5770;
assign v5771 = ~(w18265 | w18269);
assign w18270 = v5771;
assign w18271 = w18265 & w18269;
assign v5772 = ~(w18270 | w18271);
assign w18272 = v5772;
assign v5773 = ~(w17756 | w17969);
assign w18273 = v5773;
assign v5774 = ~(w17970 | w18273);
assign w18274 = v5774;
assign w18275 = w8141 & w13514;
assign w18276 = w8526 & w11720;
assign w18277 = w8926 & w11714;
assign v5775 = ~(w18276 | w18277);
assign w18278 = v5775;
assign w18279 = w8140 & w11723;
assign w18280 = w18278 & ~w18279;
assign w18281 = ~w18275 & w18280;
assign w18282 = pi08 & w18281;
assign v5776 = ~(pi08 | w18281);
assign w18283 = v5776;
assign v5777 = ~(w18282 | w18283);
assign w18284 = v5777;
assign w18285 = ~w18274 & w18284;
assign w18286 = w18274 & ~w18284;
assign w18287 = w8141 & ~w13310;
assign w18288 = w8926 & w11720;
assign w18289 = w8526 & w11723;
assign w18290 = w8140 & w11726;
assign v5778 = ~(w18289 | w18290);
assign w18291 = v5778;
assign w18292 = ~w18288 & w18291;
assign w18293 = ~w18287 & w18292;
assign w18294 = ~pi08 & w18293;
assign w18295 = pi08 & ~w18293;
assign v5779 = ~(w18294 | w18295);
assign w18296 = v5779;
assign v5780 = ~(w17769 | w17770);
assign w18297 = v5780;
assign w18298 = w17968 & w18297;
assign v5781 = ~(w17968 | w18297);
assign w18299 = v5781;
assign v5782 = ~(w18298 | w18299);
assign w18300 = v5782;
assign w18301 = w18296 & ~w18300;
assign w18302 = ~w18296 & w18300;
assign v5783 = ~(w18301 | w18302);
assign w18303 = v5783;
assign v5784 = ~(w17785 | w17966);
assign w18304 = v5784;
assign v5785 = ~(w17967 | w18304);
assign w18305 = v5785;
assign w18306 = w8141 & ~w13737;
assign w18307 = w8140 & w11729;
assign w18308 = w8926 & w11723;
assign v5786 = ~(w18307 | w18308);
assign w18309 = v5786;
assign w18310 = w8526 & w11726;
assign w18311 = w18309 & ~w18310;
assign w18312 = ~w18306 & w18311;
assign v5787 = ~(pi08 | w18312);
assign w18313 = v5787;
assign w18314 = pi08 & w18312;
assign v5788 = ~(w18313 | w18314);
assign w18315 = v5788;
assign w18316 = ~w18305 & w18315;
assign w18317 = w18305 & ~w18315;
assign w18318 = w8141 & w13864;
assign w18319 = w8526 & w11729;
assign w18320 = w8926 & w11726;
assign v5789 = ~(w18319 | w18320);
assign w18321 = v5789;
assign w18322 = w8140 & ~w11734;
assign w18323 = w18321 & ~w18322;
assign w18324 = ~w18318 & w18323;
assign v5790 = ~(pi08 | w18324);
assign w18325 = v5790;
assign w18326 = pi08 & w18324;
assign v5791 = ~(w18325 | w18326);
assign w18327 = v5791;
assign v5792 = ~(w17798 | w17799);
assign w18328 = v5792;
assign v5793 = ~(w17965 | w18328);
assign w18329 = v5793;
assign w18330 = w17965 & w18328;
assign v5794 = ~(w18329 | w18330);
assign w18331 = v5794;
assign v5795 = ~(w18327 | w18331);
assign w18332 = v5795;
assign w18333 = w17961 & ~w17963;
assign v5796 = ~(w17964 | w18333);
assign w18334 = v5796;
assign w18335 = w8141 & ~w13703;
assign w18336 = w8926 & w11729;
assign w18337 = w8526 & ~w11734;
assign w18338 = w8140 & w11737;
assign v5797 = ~(w18337 | w18338);
assign w18339 = v5797;
assign w18340 = ~w18336 & w18339;
assign w18341 = ~w18335 & w18340;
assign w18342 = pi08 & w18341;
assign v5798 = ~(pi08 | w18341);
assign w18343 = v5798;
assign v5799 = ~(w18342 | w18343);
assign w18344 = v5799;
assign w18345 = w18334 & ~w18344;
assign w18346 = w17957 & ~w17959;
assign v5800 = ~(w17960 | w18346);
assign w18347 = v5800;
assign w18348 = w8141 & w13882;
assign w18349 = w8926 & ~w11734;
assign w18350 = w8526 & w11737;
assign w18351 = w8140 & w11740;
assign v5801 = ~(w18350 | w18351);
assign w18352 = v5801;
assign w18353 = ~w18349 & w18352;
assign w18354 = ~w18348 & w18353;
assign w18355 = ~pi08 & w18354;
assign w18356 = pi08 & ~w18354;
assign v5802 = ~(w18355 | w18356);
assign w18357 = v5802;
assign w18358 = w18347 & w18357;
assign w18359 = w17953 & ~w17955;
assign v5803 = ~(w17956 | w18359);
assign w18360 = v5803;
assign w18361 = w8141 & w14288;
assign w18362 = w8926 & w11737;
assign w18363 = w8140 & ~w11745;
assign w18364 = w8526 & w11740;
assign v5804 = ~(w18363 | w18364);
assign w18365 = v5804;
assign w18366 = ~w18362 & w18365;
assign w18367 = ~w18361 & w18366;
assign w18368 = pi08 & ~w18367;
assign w18369 = ~pi08 & w18367;
assign v5805 = ~(w18368 | w18369);
assign w18370 = v5805;
assign w18371 = w18360 & w18370;
assign w18372 = w17949 & ~w17951;
assign v5806 = ~(w17952 | w18372);
assign w18373 = v5806;
assign w18374 = w8926 & w11740;
assign w18375 = w8526 & ~w11745;
assign w18376 = w8140 & w11748;
assign v5807 = ~(w18375 | w18376);
assign w18377 = v5807;
assign w18378 = ~w18374 & w18377;
assign w18379 = (w18378 & ~w14300) | (w18378 & w29532) | (~w14300 & w29532);
assign w18380 = pi08 & ~w18379;
assign w18381 = ~pi08 & w18379;
assign v5808 = ~(w18380 | w18381);
assign w18382 = v5808;
assign w18383 = w18373 & w18382;
assign w18384 = w17945 & ~w17947;
assign v5809 = ~(w17948 | w18384);
assign w18385 = v5809;
assign w18386 = w8926 & ~w11745;
assign w18387 = w8526 & w11748;
assign w18388 = w8140 & w11759;
assign v5810 = ~(w18387 | w18388);
assign w18389 = v5810;
assign w18390 = ~w18386 & w18389;
assign w18391 = (w18390 & ~w13948) | (w18390 & w29749) | (~w13948 & w29749);
assign w18392 = pi08 & w18391;
assign v5811 = ~(pi08 | w18391);
assign w18393 = v5811;
assign v5812 = ~(w18392 | w18393);
assign w18394 = v5812;
assign w18395 = w18385 & ~w18394;
assign w18396 = w17941 & ~w17943;
assign v5813 = ~(w17944 | w18396);
assign w18397 = v5813;
assign w18398 = w8926 & w11748;
assign w18399 = w8526 & w11759;
assign w18400 = w8140 & w11761;
assign v5814 = ~(w18399 | w18400);
assign w18401 = v5814;
assign w18402 = ~w18398 & w18401;
assign w18403 = (~w11841 & w29295) | (~w11841 & w29296) | (w29295 & w29296);
assign w18404 = pi08 & w18403;
assign v5815 = ~(pi08 | w18403);
assign w18405 = v5815;
assign v5816 = ~(w18404 | w18405);
assign w18406 = v5816;
assign w18407 = w18397 & ~w18406;
assign w18408 = w17937 & ~w17939;
assign v5817 = ~(w17940 | w18408);
assign w18409 = v5817;
assign w18410 = w8140 & ~w11771;
assign w18411 = w8926 & w11759;
assign v5818 = ~(w18410 | w18411);
assign w18412 = v5818;
assign w18413 = w8526 & w11761;
assign w18414 = w18412 & ~w18413;
assign w18415 = (w14356 & w29297) | (w14356 & w29298) | (w29297 & w29298);
assign w18416 = (~w14356 & w29299) | (~w14356 & w29300) | (w29299 & w29300);
assign v5819 = ~(w18415 | w18416);
assign w18417 = v5819;
assign w18418 = w18409 & ~w18417;
assign w18419 = w17933 & ~w17935;
assign v5820 = ~(w17936 | w18419);
assign w18420 = v5820;
assign w18421 = w8526 & ~w11771;
assign w18422 = w8926 & w11761;
assign w18423 = w8140 & w11768;
assign v5821 = ~(w18422 | w18423);
assign w18424 = v5821;
assign w18425 = ~w18421 & w18424;
assign w18426 = (w14383 & w28762) | (w14383 & w28763) | (w28762 & w28763);
assign w18427 = (~w14383 & w28764) | (~w14383 & w28765) | (w28764 & w28765);
assign v5822 = ~(w18426 | w18427);
assign w18428 = v5822;
assign w18429 = w18420 & w18428;
assign w18430 = w17929 & ~w17931;
assign v5823 = ~(w17932 | w18430);
assign w18431 = v5823;
assign w18432 = w8141 & w14409;
assign w18433 = w8526 & w11768;
assign w18434 = (w8926 & ~w11766) | (w8926 & w28520) | (~w11766 & w28520);
assign v5824 = ~(w18433 | w18434);
assign w18435 = v5824;
assign w18436 = w8140 & w11776;
assign w18437 = ~w18432 & w28521;
assign w18438 = (~pi08 & w18432) | (~pi08 & w28522) | (w18432 & w28522);
assign v5825 = ~(w18437 | w18438);
assign w18439 = v5825;
assign w18440 = w18431 & ~w18439;
assign v5826 = ~(w17919 | w17927);
assign w18441 = v5826;
assign v5827 = ~(w17928 | w18441);
assign w18442 = v5827;
assign w18443 = w8926 & w11768;
assign w18444 = w8140 & w11784;
assign w18445 = w8526 & w11776;
assign v5828 = ~(w18444 | w18445);
assign w18446 = v5828;
assign w18447 = ~w18443 & w18446;
assign w18448 = (w14461 & w28330) | (w14461 & w28331) | (w28330 & w28331);
assign w18449 = (~w14461 & w28332) | (~w14461 & w28333) | (w28332 & w28333);
assign v5829 = ~(w18448 | w18449);
assign w18450 = v5829;
assign w18451 = w18442 & w18450;
assign w18452 = w8141 & ~w14639;
assign w18453 = w8140 & w11800;
assign v5830 = ~(w18452 | w18453);
assign w18454 = v5830;
assign w18455 = w8926 & w11803;
assign w18456 = w8526 & w11798;
assign v5831 = ~(w18455 | w18456);
assign w18457 = v5831;
assign w18458 = w18454 & w18457;
assign w18459 = w8138 & w11800;
assign w18460 = pi08 & w18459;
assign w18461 = w8141 & ~w14609;
assign w18462 = w8926 & w11798;
assign w18463 = w8526 & w11800;
assign v5832 = ~(w18462 | w18463);
assign w18464 = v5832;
assign w18465 = ~w18461 & w18464;
assign w18466 = ~w18460 & w18465;
assign w18467 = pi08 & ~w18466;
assign w18468 = w18458 & ~w18467;
assign w18469 = pi08 & w18468;
assign v5833 = ~(w17900 | w18469);
assign w18470 = v5833;
assign w18471 = w8141 & w14569;
assign w18472 = w8526 & w11803;
assign w18473 = w8926 & w11793;
assign w18474 = w8140 & w11798;
assign v5834 = ~(w18473 | w18474);
assign w18475 = v5834;
assign w18476 = ~w18472 & w18475;
assign w18477 = (pi08 & w18471) | (pi08 & w28523) | (w18471 & w28523);
assign w18478 = ~w18471 & w28524;
assign v5835 = ~(w18477 | w18478);
assign w18479 = v5835;
assign w18480 = ~w18470 & w18479;
assign w18481 = w17901 & ~w17906;
assign v5836 = ~(w17907 | w18481);
assign w18482 = v5836;
assign v5837 = ~(pi08 | w18482);
assign w18483 = v5837;
assign w18484 = pi08 & w18482;
assign v5838 = ~(w18483 | w18484);
assign w18485 = v5838;
assign w18486 = w8141 & w14547;
assign w18487 = w8140 & w11803;
assign w18488 = w8526 & w11793;
assign w18489 = (~w18488 & ~w11784) | (~w18488 & w28766) | (~w11784 & w28766);
assign w18490 = ~w18487 & w18489;
assign w18491 = (w18485 & w18486) | (w18485 & w28525) | (w18486 & w28525);
assign w18492 = ~w18486 & w28526;
assign v5839 = ~(w18491 | w18492);
assign w18493 = v5839;
assign w18494 = w18480 & w18493;
assign w18495 = w18482 & ~w18493;
assign v5840 = ~(w18494 | w18495);
assign w18496 = v5840;
assign w18497 = w17908 & ~w17914;
assign v5841 = ~(w17915 | w18497);
assign w18498 = v5841;
assign v5842 = ~(pi08 | w18498);
assign w18499 = v5842;
assign w18500 = pi08 & w18498;
assign v5843 = ~(w18499 | w18500);
assign w18501 = v5843;
assign w18502 = w8526 & w11784;
assign w18503 = w8926 & w11776;
assign w18504 = w8140 & w11793;
assign v5844 = ~(w18503 | w18504);
assign w18505 = v5844;
assign w18506 = ~w18502 & w18505;
assign w18507 = (w14504 & w28767) | (w14504 & w28768) | (w28767 & w28768);
assign w18508 = (~w14504 & w28769) | (~w14504 & w28770) | (w28769 & w28770);
assign v5845 = ~(w18507 | w18508);
assign w18509 = v5845;
assign w18510 = ~w18496 & w18509;
assign w18511 = w18498 & ~w18509;
assign v5846 = ~(w18510 | w18511);
assign w18512 = v5846;
assign v5847 = ~(w18442 | w18450);
assign w18513 = v5847;
assign v5848 = ~(w18451 | w18513);
assign w18514 = v5848;
assign w18515 = ~w18512 & w18514;
assign w18516 = (~w18451 & ~w18514) | (~w18451 & w28528) | (~w18514 & w28528);
assign w18517 = ~w18431 & w18439;
assign v5849 = ~(w18440 | w18517);
assign w18518 = v5849;
assign w18519 = ~w18516 & w18518;
assign w18520 = (~w18440 & ~w18518) | (~w18440 & w29301) | (~w18518 & w29301);
assign v5850 = ~(w18420 | w18428);
assign w18521 = v5850;
assign v5851 = ~(w18429 | w18521);
assign w18522 = v5851;
assign w18523 = ~w18520 & w18522;
assign w18524 = (~w18429 & w18520) | (~w18429 & w28771) | (w18520 & w28771);
assign w18525 = ~w18409 & w18417;
assign v5852 = ~(w18418 | w18525);
assign w18526 = v5852;
assign w18527 = ~w18524 & w18526;
assign w18528 = (~w18418 & w18524) | (~w18418 & w29302) | (w18524 & w29302);
assign w18529 = ~w18397 & w18406;
assign v5853 = ~(w18407 | w18529);
assign w18530 = v5853;
assign w18531 = ~w18528 & w18530;
assign w18532 = (~w18407 & w18528) | (~w18407 & w28529) | (w18528 & w28529);
assign w18533 = ~w18385 & w18394;
assign v5854 = ~(w18395 | w18533);
assign w18534 = v5854;
assign w18535 = ~w18532 & w18534;
assign w18536 = (~w18395 & w18532) | (~w18395 & w29750) | (w18532 & w29750);
assign v5855 = ~(w18373 | w18382);
assign w18537 = v5855;
assign v5856 = ~(w18383 | w18537);
assign w18538 = v5856;
assign w18539 = ~w18536 & w18538;
assign w18540 = (~w18383 & w18536) | (~w18383 & w29303) | (w18536 & w29303);
assign v5857 = ~(w18360 | w18370);
assign w18541 = v5857;
assign v5858 = ~(w18371 | w18541);
assign w18542 = v5858;
assign w18543 = ~w18540 & w18542;
assign w18544 = (~w18371 & ~w18542) | (~w18371 & w28530) | (~w18542 & w28530);
assign v5859 = ~(w18347 | w18357);
assign w18545 = v5859;
assign v5860 = ~(w18358 | w18545);
assign w18546 = v5860;
assign w18547 = ~w18544 & w18546;
assign w18548 = (~w18358 & w18544) | (~w18358 & w29533) | (w18544 & w29533);
assign w18549 = ~w18334 & w18344;
assign v5861 = ~(w18345 | w18549);
assign w18550 = v5861;
assign w18551 = ~w18548 & w18550;
assign w18552 = (~w18345 & w18548) | (~w18345 & w29751) | (w18548 & w29751);
assign w18553 = w18327 & w18331;
assign v5862 = ~(w18332 | w18553);
assign w18554 = v5862;
assign w18555 = ~w18552 & w18554;
assign w18556 = (~w18332 & w18552) | (~w18332 & w29879) | (w18552 & w29879);
assign w18557 = (~w18316 & ~w18556) | (~w18316 & w29304) | (~w18556 & w29304);
assign w18558 = w18303 & w18557;
assign w18559 = (~w18301 & ~w18303) | (~w18301 & w28531) | (~w18303 & w28531);
assign w18560 = (~w18285 & ~w18559) | (~w18285 & w30056) | (~w18559 & w30056);
assign w18561 = w18272 & w18560;
assign w18562 = (~w18270 & ~w18272) | (~w18270 & w28532) | (~w18272 & w28532);
assign w18563 = (~w18254 & ~w18562) | (~w18254 & w30190) | (~w18562 & w30190);
assign w18564 = w18241 & w18563;
assign w18565 = (~w18239 & ~w18241) | (~w18239 & w28533) | (~w18241 & w28533);
assign w18566 = (~w28533 & w30191) | (~w28533 & w30192) | (w30191 & w30192);
assign w18567 = (~w18221 & w18565) | (~w18221 & w28772) | (w18565 & w28772);
assign w18568 = w18208 & ~w18567;
assign w18569 = (~w18206 & ~w18208) | (~w18206 & w28773) | (~w18208 & w28773);
assign w18570 = (~w18190 & ~w18569) | (~w18190 & w30193) | (~w18569 & w30193);
assign w18571 = w18175 & w18570;
assign w18572 = (~w18173 & ~w18175) | (~w18173 & w28534) | (~w18175 & w28534);
assign w18573 = (~w18155 & ~w18572) | (~w18155 & w28774) | (~w18572 & w28774);
assign w18574 = w18141 & w18573;
assign w18575 = (~w18139 & ~w18573) | (~w18139 & w30642) | (~w18573 & w30642);
assign w18576 = (~w18122 & ~w18575) | (~w18122 & w30525) | (~w18575 & w30525);
assign w18577 = w18108 & w18576;
assign w18578 = (~w18106 & ~w18108) | (~w18106 & w28775) | (~w18108 & w28775);
assign w18579 = w18093 & ~w18578;
assign w18580 = (~w18091 & w18578) | (~w18091 & w31197) | (w18578 & w31197);
assign w18581 = w18078 & ~w18580;
assign w18582 = (~w18076 & ~w18078) | (~w18076 & w28776) | (~w18078 & w28776);
assign w18583 = ~w18052 & w18062;
assign v5863 = ~(w18063 | w18583);
assign w18584 = v5863;
assign w18585 = w18582 & w18584;
assign w18586 = (~w18063 & ~w18584) | (~w18063 & w28777) | (~w18584 & w28777);
assign w18587 = ~w18039 & w18049;
assign v5864 = ~(w18050 | w18587);
assign w18588 = v5864;
assign w18589 = w18586 & w18588;
assign w18590 = (~w18050 & ~w18588) | (~w18050 & w28778) | (~w18588 & w28778);
assign w18591 = ~w18037 & w18590;
assign w18592 = w18037 & ~w18590;
assign v5865 = ~(w18591 | w18592);
assign w18593 = v5865;
assign w18594 = w9401 & w12381;
assign w18595 = (w28779 & ~w12502) | (w28779 & w29305) | (~w12502 & w29305);
assign v5866 = ~(w9891 | w18595);
assign w18596 = v5866;
assign v5867 = ~(w12406 | w18596);
assign w18597 = v5867;
assign v5868 = ~(w10419 | w18597);
assign w18598 = v5868;
assign w18599 = ~w18594 & w18598;
assign w18600 = ~pi05 & w18599;
assign w18601 = pi05 & ~w18599;
assign v5869 = ~(w18600 | w18601);
assign w18602 = v5869;
assign w18603 = w18593 & ~w18602;
assign w18604 = (~w18591 & ~w18593) | (~w18591 & w29306) | (~w18593 & w29306);
assign w18605 = w18030 & ~w18032;
assign v5870 = ~(w18033 | w18605);
assign w18606 = v5870;
assign w18607 = ~w18604 & w18606;
assign w18608 = w18604 & ~w18606;
assign v5871 = ~(w18607 | w18608);
assign w18609 = v5871;
assign w18610 = ~w18593 & w18602;
assign v5872 = ~(w18603 | w18610);
assign w18611 = v5872;
assign w18612 = (w10445 & ~w12505) | (w10445 & w30194) | (~w12505 & w30194);
assign w18613 = (w10419 & ~w12405) | (w10419 & w30195) | (~w12405 & w30195);
assign w18614 = w9401 & w12311;
assign w18615 = (~w18614 & ~w12381) | (~w18614 & w30196) | (~w12381 & w30196);
assign w18616 = ~w18613 & w18615;
assign w18617 = pi05 & ~w18616;
assign w18618 = ~pi05 & w18616;
assign w18619 = (w12505 & w28780) | (w12505 & w28781) | (w28780 & w28781);
assign v5873 = ~(w18617 | w18619);
assign w18620 = v5873;
assign w18621 = w18620 & w30197;
assign v5874 = ~(w18586 | w18588);
assign w18622 = v5874;
assign v5875 = ~(w18589 | w18622);
assign w18623 = v5875;
assign w18624 = (~w13657 & ~w18620) | (~w13657 & w30198) | (~w18620 & w30198);
assign v5876 = ~(w18621 | w18624);
assign w18625 = v5876;
assign w18626 = w18623 & w18625;
assign v5877 = ~(w18621 | w18626);
assign w18627 = v5877;
assign w18628 = w18611 & w18627;
assign v5878 = ~(w18582 | w18584);
assign w18629 = v5878;
assign v5879 = ~(w18585 | w18629);
assign w18630 = v5879;
assign w18631 = w10419 & w12381;
assign w18632 = w9401 & w12271;
assign w18633 = w9891 & w12311;
assign v5880 = ~(w18632 | w18633);
assign w18634 = v5880;
assign w18635 = ~w18631 & w18634;
assign w18636 = (w18635 & ~w12387) | (w18635 & w28782) | (~w12387 & w28782);
assign w18637 = ~pi05 & w18636;
assign w18638 = pi05 & ~w18636;
assign v5881 = ~(w18637 | w18638);
assign w18639 = v5881;
assign w18640 = ~w18630 & w18639;
assign w18641 = w18630 & ~w18639;
assign v5882 = ~(w18640 | w18641);
assign w18642 = v5882;
assign w18643 = ~w18078 & w18580;
assign v5883 = ~(w18581 | w18643);
assign w18644 = v5883;
assign w18645 = w10419 & w12311;
assign w18646 = w9891 & w12271;
assign w18647 = w9401 & w12237;
assign v5884 = ~(w18646 | w18647);
assign w18648 = v5884;
assign w18649 = ~w18645 & w18648;
assign w18650 = (w18649 & ~w12318) | (w18649 & w28783) | (~w12318 & w28783);
assign w18651 = pi05 & ~w18650;
assign w18652 = ~pi05 & w18650;
assign v5885 = ~(w18651 | w18652);
assign w18653 = v5885;
assign v5886 = ~(w18644 | w18653);
assign w18654 = v5886;
assign w18655 = ~w18093 & w18578;
assign v5887 = ~(w18579 | w18655);
assign w18656 = v5887;
assign w18657 = w10445 & ~w12277;
assign w18658 = w10419 & w12271;
assign w18659 = w9891 & w12237;
assign w18660 = w9401 & w12155;
assign v5888 = ~(w18659 | w18660);
assign w18661 = v5888;
assign w18662 = ~w18658 & w18661;
assign w18663 = pi05 & ~w18662;
assign w18664 = ~pi05 & w18662;
assign w18665 = (w18664 & w12277) | (w18664 & w30199) | (w12277 & w30199);
assign v5889 = ~(w18663 | w18665);
assign w18666 = v5889;
assign w18667 = ~w18657 & w18666;
assign w18668 = w18656 & w18667;
assign v5890 = ~(w18656 | w18667);
assign w18669 = v5890;
assign v5891 = ~(w18668 | w18669);
assign w18670 = v5891;
assign w18671 = w10419 & w12237;
assign w18672 = w9891 & w12155;
assign w18673 = w9401 & w12084;
assign v5892 = ~(w18672 | w18673);
assign w18674 = v5892;
assign w18675 = ~w18671 & w18674;
assign w18676 = pi05 & ~w18675;
assign w18677 = ~pi05 & w18675;
assign w18678 = (w18677 & w12351) | (w18677 & w28784) | (w12351 & w28784);
assign w18679 = w10445 & ~w12351;
assign v5893 = ~(w18678 | w18679);
assign w18680 = v5893;
assign w18681 = ~w18676 & w18680;
assign v5894 = ~(w18108 | w18576);
assign w18682 = v5894;
assign v5895 = ~(w18577 | w18682);
assign w18683 = v5895;
assign w18684 = w18681 & w18683;
assign w18685 = w10445 & w12167;
assign w18686 = w10447 & w12167;
assign w18687 = w10419 & w12155;
assign w18688 = w9891 & w12084;
assign w18689 = w9401 & w11984;
assign v5896 = ~(w18688 | w18689);
assign w18690 = v5896;
assign w18691 = ~w18687 & w18690;
assign w18692 = pi05 & w18691;
assign v5897 = ~(pi05 | w18691);
assign w18693 = v5897;
assign v5898 = ~(w18692 | w18693);
assign w18694 = v5898;
assign w18695 = ~w18686 & w18694;
assign v5899 = ~(w18685 | w18695);
assign w18696 = v5899;
assign v5900 = ~(w18122 | w18123);
assign w18697 = v5900;
assign w18698 = w18575 & ~w18697;
assign w18699 = ~w18575 & w18697;
assign v5901 = ~(w18698 | w18699);
assign w18700 = v5901;
assign w18701 = w18696 & w18700;
assign v5902 = ~(w18696 | w18700);
assign w18702 = v5902;
assign v5903 = ~(w18701 | w18702);
assign w18703 = v5903;
assign v5904 = ~(w18141 | w18573);
assign w18704 = v5904;
assign v5905 = ~(w18574 | w18704);
assign w18705 = v5905;
assign w18706 = w9891 & w11984;
assign w18707 = w10419 & w12084;
assign v5906 = ~(w18706 | w18707);
assign w18708 = v5906;
assign w18709 = w9401 & w11671;
assign w18710 = w18708 & ~w18709;
assign w18711 = (~w12181 & w30200) | (~w12181 & w30201) | (w30200 & w30201);
assign w18712 = (w12181 & w30202) | (w12181 & w30203) | (w30202 & w30203);
assign v5907 = ~(w18711 | w18712);
assign w18713 = v5907;
assign w18714 = w18705 & ~w18713;
assign w18715 = ~w18705 & w18713;
assign v5908 = ~(w18714 | w18715);
assign w18716 = v5908;
assign w18717 = w10445 & w11993;
assign w18718 = ~w11992 & w28786;
assign w18719 = w10419 & w11984;
assign w18720 = w9891 & w11671;
assign w18721 = w9401 & w11673;
assign v5909 = ~(w18720 | w18721);
assign w18722 = v5909;
assign w18723 = ~w18719 & w18722;
assign w18724 = pi05 & w18723;
assign v5910 = ~(pi05 | w18723);
assign w18725 = v5910;
assign v5911 = ~(w18724 | w18725);
assign w18726 = v5911;
assign w18727 = ~w18718 & w18726;
assign v5912 = ~(w18717 | w18727);
assign w18728 = v5912;
assign v5913 = ~(w18155 | w18156);
assign w18729 = v5913;
assign v5914 = ~(w18572 | w18729);
assign w18730 = v5914;
assign w18731 = w18572 & w18729;
assign v5915 = ~(w18730 | w18731);
assign w18732 = v5915;
assign w18733 = w18728 & ~w18732;
assign w18734 = ~w18728 & w18732;
assign v5916 = ~(w18175 | w18570);
assign w18735 = v5916;
assign v5917 = ~(w18571 | w18735);
assign w18736 = v5917;
assign w18737 = w9891 & w11673;
assign w18738 = w10419 & w11671;
assign v5918 = ~(w18737 | w18738);
assign w18739 = v5918;
assign w18740 = w9401 & w11678;
assign w18741 = w18739 & ~w18740;
assign w18742 = (w12469 & w30204) | (w12469 & w30205) | (w30204 & w30205);
assign w18743 = (~w12469 & w30206) | (~w12469 & w30207) | (w30206 & w30207);
assign v5919 = ~(w18742 | w18743);
assign w18744 = v5919;
assign w18745 = ~w18736 & w18744;
assign w18746 = w18736 & ~w18744;
assign w18747 = w10445 & w12454;
assign w18748 = w10447 & w12454;
assign w18749 = w10419 & w11673;
assign w18750 = w9891 & w11678;
assign w18751 = w9401 & ~w11683;
assign v5920 = ~(w18750 | w18751);
assign w18752 = v5920;
assign w18753 = ~w18749 & w18752;
assign w18754 = pi05 & w18753;
assign v5921 = ~(pi05 | w18753);
assign w18755 = v5921;
assign v5922 = ~(w18754 | w18755);
assign w18756 = v5922;
assign w18757 = ~w18748 & w18756;
assign v5923 = ~(w18747 | w18757);
assign w18758 = v5923;
assign v5924 = ~(w18190 | w18191);
assign w18759 = v5924;
assign v5925 = ~(w18569 | w18759);
assign w18760 = v5925;
assign w18761 = w18569 & w18759;
assign v5926 = ~(w18760 | w18761);
assign w18762 = v5926;
assign w18763 = w18758 & ~w18762;
assign w18764 = ~w18758 & w18762;
assign v5927 = ~(w18763 | w18764);
assign w18765 = v5927;
assign w18766 = w10445 & w12594;
assign w18767 = w10447 & w12594;
assign w18768 = w10419 & w11678;
assign w18769 = w9891 & ~w11683;
assign w18770 = w9401 & w11686;
assign v5928 = ~(w18769 | w18770);
assign w18771 = v5928;
assign w18772 = ~w18768 & w18771;
assign w18773 = pi05 & w18772;
assign v5929 = ~(pi05 | w18772);
assign w18774 = v5929;
assign v5930 = ~(w18773 | w18774);
assign w18775 = v5930;
assign w18776 = ~w18767 & w18775;
assign v5931 = ~(w18766 | w18776);
assign w18777 = v5931;
assign w18778 = ~w18208 & w18567;
assign v5932 = ~(w18568 | w18778);
assign w18779 = v5932;
assign v5933 = ~(w18777 | w18779);
assign w18780 = v5933;
assign w18781 = w18777 & w18779;
assign w18782 = w10445 & w12610;
assign w18783 = w10447 & w12610;
assign w18784 = w10419 & ~w11683;
assign w18785 = w9891 & w11686;
assign w18786 = w9401 & w11689;
assign v5934 = ~(w18785 | w18786);
assign w18787 = v5934;
assign w18788 = ~w18784 & w18787;
assign w18789 = pi05 & w18788;
assign v5935 = ~(pi05 | w18788);
assign w18790 = v5935;
assign v5936 = ~(w18789 | w18790);
assign w18791 = v5936;
assign w18792 = ~w18783 & w18791;
assign v5937 = ~(w18782 | w18792);
assign w18793 = v5937;
assign v5938 = ~(w18221 | w18222);
assign w18794 = v5938;
assign w18795 = w18565 & ~w18794;
assign w18796 = ~w18221 & w18566;
assign v5939 = ~(w18795 | w18796);
assign w18797 = v5939;
assign w18798 = w18793 & w18797;
assign v5940 = ~(w18793 | w18797);
assign w18799 = v5940;
assign v5941 = ~(w18798 | w18799);
assign w18800 = v5941;
assign v5942 = ~(w18241 | w18563);
assign w18801 = v5942;
assign v5943 = ~(w18564 | w18801);
assign w18802 = v5943;
assign w18803 = w10445 & ~w12842;
assign w18804 = w10447 & ~w12842;
assign w18805 = w10419 & w11686;
assign w18806 = w9891 & w11689;
assign w18807 = w9401 & ~w11695;
assign v5944 = ~(w18806 | w18807);
assign w18808 = v5944;
assign w18809 = ~w18805 & w18808;
assign w18810 = pi05 & w18809;
assign v5945 = ~(pi05 | w18809);
assign w18811 = v5945;
assign v5946 = ~(w18810 | w18811);
assign w18812 = v5946;
assign w18813 = ~w18804 & w18812;
assign v5947 = ~(w18803 | w18813);
assign w18814 = v5947;
assign w18815 = w18802 & w18814;
assign v5948 = ~(w18802 | w18814);
assign w18816 = v5948;
assign w18817 = w9402 & w12694;
assign w18818 = w10419 & w11689;
assign w18819 = w9401 & w11700;
assign w18820 = w9891 & ~w11695;
assign v5949 = ~(w18819 | w18820);
assign w18821 = v5949;
assign w18822 = ~w18818 & w18821;
assign w18823 = ~w18817 & w18822;
assign w18824 = pi05 & ~w18823;
assign w18825 = ~pi05 & w18823;
assign v5950 = ~(w18824 | w18825);
assign w18826 = v5950;
assign v5951 = ~(w18254 | w18255);
assign w18827 = v5951;
assign w18828 = w18562 & w18827;
assign v5952 = ~(w18562 | w18827);
assign w18829 = v5952;
assign v5953 = ~(w18828 | w18829);
assign w18830 = v5953;
assign w18831 = w18826 & ~w18830;
assign w18832 = ~w18826 & w18830;
assign v5954 = ~(w18831 | w18832);
assign w18833 = v5954;
assign v5955 = ~(w18272 | w18560);
assign w18834 = v5955;
assign v5956 = ~(w18561 | w18834);
assign w18835 = v5956;
assign w18836 = w9402 & ~w13008;
assign w18837 = w10419 & ~w11695;
assign w18838 = w9891 & w11700;
assign w18839 = w9401 & w11708;
assign v5957 = ~(w18838 | w18839);
assign w18840 = v5957;
assign w18841 = ~w18837 & w18840;
assign w18842 = ~w18836 & w18841;
assign w18843 = pi05 & w18842;
assign v5958 = ~(pi05 | w18842);
assign w18844 = v5958;
assign v5959 = ~(w18843 | w18844);
assign w18845 = v5959;
assign w18846 = ~w18835 & w18845;
assign w18847 = w18835 & ~w18845;
assign w18848 = ~w11884 & w28334;
assign w18849 = w10419 & w11700;
assign w18850 = w9401 & w11711;
assign w18851 = w9891 & w11708;
assign v5960 = ~(w18850 | w18851);
assign w18852 = v5960;
assign w18853 = ~w18849 & w18852;
assign w18854 = ~w18848 & w18853;
assign w18855 = ~pi05 & w18854;
assign w18856 = pi05 & ~w18854;
assign v5961 = ~(w18855 | w18856);
assign w18857 = v5961;
assign v5962 = ~(w18285 | w18286);
assign w18858 = v5962;
assign w18859 = w18559 & w18858;
assign v5963 = ~(w18559 | w18858);
assign w18860 = v5963;
assign v5964 = ~(w18859 | w18860);
assign w18861 = v5964;
assign w18862 = w18857 & ~w18861;
assign w18863 = ~w18857 & w18861;
assign v5965 = ~(w18862 | w18863);
assign w18864 = v5965;
assign v5966 = ~(w18303 | w18557);
assign w18865 = v5966;
assign v5967 = ~(w18558 | w18865);
assign w18866 = v5967;
assign w18867 = w9402 & w13178;
assign w18868 = w10419 & w11708;
assign w18869 = w9401 & w11714;
assign w18870 = w9891 & w11711;
assign v5968 = ~(w18869 | w18870);
assign w18871 = v5968;
assign w18872 = ~w18868 & w18871;
assign w18873 = ~w18867 & w18872;
assign w18874 = ~pi05 & w18873;
assign w18875 = pi05 & ~w18873;
assign v5969 = ~(w18874 | w18875);
assign w18876 = v5969;
assign v5970 = ~(w18866 | w18876);
assign w18877 = v5970;
assign w18878 = w18866 & w18876;
assign v5971 = ~(w18316 | w18317);
assign w18879 = v5971;
assign v5972 = ~(w18556 | w18879);
assign w18880 = v5972;
assign w18881 = w18556 & w18879;
assign v5973 = ~(w18880 | w18881);
assign w18882 = v5973;
assign w18883 = ~w11877 & w28030;
assign w18884 = w9891 & w11714;
assign w18885 = w10419 & w11711;
assign v5974 = ~(w18884 | w18885);
assign w18886 = v5974;
assign w18887 = w9401 & w11720;
assign w18888 = w18886 & ~w18887;
assign w18889 = ~w18883 & w18888;
assign v5975 = ~(pi05 | w18889);
assign w18890 = v5975;
assign w18891 = pi05 & w18889;
assign v5976 = ~(w18890 | w18891);
assign w18892 = v5976;
assign v5977 = ~(w18882 | w18892);
assign w18893 = v5977;
assign w18894 = w18552 & ~w18554;
assign v5978 = ~(w18555 | w18894);
assign w18895 = v5978;
assign w18896 = ~w11873 & w28031;
assign w18897 = w9891 & w11720;
assign w18898 = w10419 & w11714;
assign v5979 = ~(w18897 | w18898);
assign w18899 = v5979;
assign w18900 = w9401 & w11723;
assign w18901 = w18899 & ~w18900;
assign w18902 = ~w18896 & w18901;
assign v5980 = ~(pi05 | w18902);
assign w18903 = v5980;
assign w18904 = pi05 & w18902;
assign v5981 = ~(w18903 | w18904);
assign w18905 = v5981;
assign w18906 = w18895 & ~w18905;
assign w18907 = w18548 & ~w18550;
assign v5982 = ~(w18551 | w18907);
assign w18908 = v5982;
assign w18909 = (w9402 & w11869) | (w9402 & w28032) | (w11869 & w28032);
assign w18910 = w10419 & w11720;
assign w18911 = w9891 & w11723;
assign w18912 = w9401 & w11726;
assign v5983 = ~(w18911 | w18912);
assign w18913 = v5983;
assign w18914 = ~w18910 & w18913;
assign w18915 = ~w18909 & w18914;
assign w18916 = pi05 & w18915;
assign v5984 = ~(pi05 | w18915);
assign w18917 = v5984;
assign v5985 = ~(w18916 | w18917);
assign w18918 = v5985;
assign w18919 = w18908 & ~w18918;
assign w18920 = w18544 & ~w18546;
assign v5986 = ~(w18547 | w18920);
assign w18921 = v5986;
assign w18922 = (w9402 & w11865) | (w9402 & w28033) | (w11865 & w28033);
assign w18923 = w10419 & w11723;
assign w18924 = w9401 & w11729;
assign w18925 = w9891 & w11726;
assign v5987 = ~(w18924 | w18925);
assign w18926 = v5987;
assign w18927 = ~w18923 & w18926;
assign w18928 = ~w18922 & w18927;
assign w18929 = pi05 & w18928;
assign v5988 = ~(pi05 | w18928);
assign w18930 = v5988;
assign v5989 = ~(w18929 | w18930);
assign w18931 = v5989;
assign w18932 = w18921 & ~w18931;
assign w18933 = w18540 & ~w18542;
assign v5990 = ~(w18543 | w18933);
assign w18934 = v5990;
assign w18935 = ~w11861 & w28034;
assign w18936 = w9891 & w11729;
assign w18937 = w10419 & w11726;
assign v5991 = ~(w18936 | w18937);
assign w18938 = v5991;
assign w18939 = w9401 & ~w11734;
assign w18940 = w18938 & ~w18939;
assign w18941 = ~w18935 & w18940;
assign v5992 = ~(pi05 | w18941);
assign w18942 = v5992;
assign w18943 = pi05 & w18941;
assign v5993 = ~(w18942 | w18943);
assign w18944 = v5993;
assign w18945 = w18934 & ~w18944;
assign w18946 = w18536 & ~w18538;
assign v5994 = ~(w18539 | w18946);
assign w18947 = v5994;
assign w18948 = (w9402 & w11858) | (w9402 & w28035) | (w11858 & w28035);
assign w18949 = w10419 & w11729;
assign w18950 = w9891 & ~w11734;
assign w18951 = w9401 & w11737;
assign v5995 = ~(w18950 | w18951);
assign w18952 = v5995;
assign w18953 = ~w18949 & w18952;
assign w18954 = ~w18948 & w18953;
assign w18955 = pi05 & ~w18954;
assign w18956 = ~pi05 & w18954;
assign v5996 = ~(w18955 | w18956);
assign w18957 = v5996;
assign w18958 = w18947 & w18957;
assign w18959 = w18532 & ~w18534;
assign v5997 = ~(w18535 | w18959);
assign w18960 = v5997;
assign w18961 = ~w11854 & w28036;
assign w18962 = w10419 & ~w11734;
assign w18963 = w9891 & w11737;
assign w18964 = w9401 & w11740;
assign v5998 = ~(w18963 | w18964);
assign w18965 = v5998;
assign w18966 = ~w18962 & w18965;
assign w18967 = ~w18961 & w18966;
assign w18968 = ~pi05 & w18967;
assign w18969 = pi05 & ~w18967;
assign v5999 = ~(w18968 | w18969);
assign w18970 = v5999;
assign w18971 = w18960 & w18970;
assign w18972 = w18528 & ~w18530;
assign v6000 = ~(w18531 | w18972);
assign w18973 = v6000;
assign w18974 = ~w14287 & w29752;
assign w18975 = w10419 & w11737;
assign w18976 = w9401 & ~w11745;
assign w18977 = w9891 & w11740;
assign v6001 = ~(w18976 | w18977);
assign w18978 = v6001;
assign w18979 = ~w18975 & w18978;
assign w18980 = ~w18974 & w18979;
assign w18981 = pi05 & ~w18980;
assign w18982 = ~pi05 & w18980;
assign v6002 = ~(w18981 | w18982);
assign w18983 = v6002;
assign w18984 = w18973 & w18983;
assign w18985 = w18524 & ~w18526;
assign v6003 = ~(w18527 | w18985);
assign w18986 = v6003;
assign w18987 = w10419 & w11740;
assign w18988 = w9891 & ~w11745;
assign w18989 = w9401 & w11748;
assign v6004 = ~(w18988 | w18989);
assign w18990 = v6004;
assign w18991 = ~w18987 & w18990;
assign w18992 = (w18991 & ~w14300) | (w18991 & w29534) | (~w14300 & w29534);
assign w18993 = pi05 & w18992;
assign v6005 = ~(pi05 | w18992);
assign w18994 = v6005;
assign v6006 = ~(w18993 | w18994);
assign w18995 = v6006;
assign w18996 = w18986 & ~w18995;
assign w18997 = w18520 & ~w18522;
assign v6007 = ~(w18523 | w18997);
assign w18998 = v6007;
assign w18999 = w10419 & ~w11745;
assign w19000 = w9891 & w11748;
assign w19001 = w9401 & w11759;
assign v6008 = ~(w19000 | w19001);
assign w19002 = v6008;
assign w19003 = ~w18999 & w19002;
assign w19004 = (w19003 & ~w28037) | (w19003 & w29753) | (~w28037 & w29753);
assign w19005 = pi05 & w19004;
assign v6009 = ~(pi05 | w19004);
assign w19006 = v6009;
assign v6010 = ~(w19005 | w19006);
assign w19007 = v6010;
assign w19008 = w18998 & ~w19007;
assign w19009 = w18516 & ~w18518;
assign v6011 = ~(w18519 | w19009);
assign w19010 = v6011;
assign w19011 = w9891 & w11759;
assign w19012 = w10419 & w11748;
assign v6012 = ~(w19011 | w19012);
assign w19013 = v6012;
assign w19014 = w9401 & w11761;
assign w19015 = w19013 & ~w19014;
assign w19016 = (w14331 & w29307) | (w14331 & w29308) | (w29307 & w29308);
assign w19017 = (~w14331 & w29309) | (~w14331 & w29310) | (w29309 & w29310);
assign v6013 = ~(w19016 | w19017);
assign w19018 = v6013;
assign w19019 = w19010 & ~w19018;
assign w19020 = w18512 & ~w18514;
assign v6014 = ~(w18515 | w19020);
assign w19021 = v6014;
assign w19022 = w9401 & ~w11771;
assign w19023 = w10419 & w11759;
assign v6015 = ~(w19022 | w19023);
assign w19024 = v6015;
assign w19025 = w9891 & w11761;
assign w19026 = w19024 & ~w19025;
assign w19027 = (w14356 & w29311) | (w14356 & w29312) | (w29311 & w29312);
assign w19028 = (~w14356 & w29313) | (~w14356 & w29314) | (w29313 & w29314);
assign v6016 = ~(w19027 | w19028);
assign w19029 = v6016;
assign w19030 = w19021 & ~w19029;
assign w19031 = ~w19021 & w19029;
assign v6017 = ~(w19030 | w19031);
assign w19032 = v6017;
assign w19033 = w18496 & ~w18509;
assign v6018 = ~(w18510 | w19033);
assign w19034 = v6018;
assign w19035 = w10445 & ~w14383;
assign w19036 = w10447 & ~w14383;
assign w19037 = w9891 & ~w11771;
assign w19038 = w9401 & w11768;
assign w19039 = (~w19038 & ~w11761) | (~w19038 & w28790) | (~w11761 & w28790);
assign w19040 = ~w19037 & w19039;
assign w19041 = pi05 & w19040;
assign v6019 = ~(pi05 | w19040);
assign w19042 = v6019;
assign v6020 = ~(w19041 | w19042);
assign w19043 = v6020;
assign w19044 = ~w19036 & w19043;
assign w19045 = (~w19034 & w19044) | (~w19034 & w28791) | (w19044 & w28791);
assign w19046 = ~w19044 & w28792;
assign v6021 = ~(w19045 | w19046);
assign w19047 = v6021;
assign v6022 = ~(w18480 | w18493);
assign w19048 = v6022;
assign v6023 = ~(w18494 | w19048);
assign w19049 = v6023;
assign w19050 = w9402 & w14409;
assign w19051 = w9401 & w11776;
assign w19052 = (w10419 & ~w11766) | (w10419 & w28536) | (~w11766 & w28536);
assign w19053 = w9891 & w11768;
assign w19054 = ~w19052 & w29315;
assign w19055 = (pi05 & w19050) | (pi05 & w28537) | (w19050 & w28537);
assign w19056 = ~w19050 & w28538;
assign v6024 = ~(w19055 | w19056);
assign w19057 = v6024;
assign v6025 = ~(w19049 | w19057);
assign w19058 = v6025;
assign w19059 = w19049 & w19057;
assign w19060 = w18468 & w28539;
assign v6026 = ~(w18470 | w19060);
assign w19061 = v6026;
assign v6027 = ~(w18479 | w19061);
assign w19062 = v6027;
assign w19063 = w18479 & w19061;
assign v6028 = ~(w19062 | w19063);
assign w19064 = v6028;
assign w19065 = w10445 & w14461;
assign w19066 = w10447 & w14461;
assign w19067 = w11533 & w29316;
assign w19068 = w9891 & w11776;
assign w19069 = w9401 & w11784;
assign v6029 = ~(w19068 | w19069);
assign w19070 = v6029;
assign w19071 = ~w19067 & w19070;
assign w19072 = pi05 & w19071;
assign v6030 = ~(pi05 | w19071);
assign w19073 = v6030;
assign v6031 = ~(w19072 | w19073);
assign w19074 = v6031;
assign w19075 = ~w19066 & w19074;
assign w19076 = ~w19075 & w28335;
assign w19077 = w18460 & ~w18465;
assign v6032 = ~(w18466 | w19077);
assign w19078 = v6032;
assign w19079 = w9402 & w14547;
assign w19080 = w9891 & w11793;
assign w19081 = ~w11782 & w28038;
assign v6033 = ~(w19080 | w19081);
assign w19082 = v6033;
assign w19083 = w9401 & w11803;
assign w19084 = ~w19079 & w28039;
assign w19085 = (~pi05 & w19079) | (~pi05 & w28040) | (w19079 & w28040);
assign v6034 = ~(w19084 | w19085);
assign w19086 = v6034;
assign w19087 = w19078 & ~w19086;
assign w19088 = w9402 & ~w14639;
assign w19089 = w9401 & w11800;
assign v6035 = ~(w19088 | w19089);
assign w19090 = v6035;
assign w19091 = w10419 & w11803;
assign w19092 = w9891 & w11798;
assign v6036 = ~(w19091 | w19092);
assign w19093 = v6036;
assign w19094 = w19090 & w19093;
assign w19095 = w11394 & w11800;
assign w19096 = w9402 & ~w14609;
assign w19097 = w10419 & w11798;
assign w19098 = w9891 & w11800;
assign v6037 = ~(w19097 | w19098);
assign w19099 = v6037;
assign w19100 = ~w19096 & w19099;
assign w19101 = ~w19095 & w19100;
assign w19102 = pi05 & w19101;
assign w19103 = w19094 & w19102;
assign v6038 = ~(w18459 | w19103);
assign w19104 = v6038;
assign w19105 = w10445 & w14569;
assign w19106 = w10447 & w14569;
assign w19107 = w10419 & w11793;
assign w19108 = w9891 & w11803;
assign w19109 = w9401 & w11798;
assign v6039 = ~(w19108 | w19109);
assign w19110 = v6039;
assign w19111 = ~w19107 & w19110;
assign w19112 = pi05 & w19111;
assign v6040 = ~(pi05 | w19111);
assign w19113 = v6040;
assign v6041 = ~(w19112 | w19113);
assign w19114 = v6041;
assign w19115 = ~w19106 & w19114;
assign v6042 = ~(w19105 | w19115);
assign w19116 = v6042;
assign w19117 = ~w19104 & w19116;
assign w19118 = ~w19078 & w19086;
assign v6043 = ~(w19087 | w19118);
assign w19119 = v6043;
assign w19120 = w19117 & w19119;
assign w19121 = (~w19087 & ~w19119) | (~w19087 & w28336) | (~w19119 & w28336);
assign w19122 = w9401 & w11793;
assign w19123 = w10419 & w11776;
assign w19124 = w9891 & w11784;
assign v6044 = ~(w19123 | w19124);
assign w19125 = v6044;
assign w19126 = (~w14504 & w28042) | (~w14504 & w28043) | (w28042 & w28043);
assign w19127 = ~w18458 & w18467;
assign v6045 = ~(w18468 | w19127);
assign w19128 = v6045;
assign w19129 = ~pi05 & w19128;
assign w19130 = pi05 & ~w19128;
assign v6046 = ~(w19129 | w19130);
assign w19131 = v6046;
assign w19132 = w19126 & ~w19131;
assign w19133 = ~w19126 & w19131;
assign v6047 = ~(w19132 | w19133);
assign w19134 = v6047;
assign v6048 = ~(w19121 | w19134);
assign w19135 = v6048;
assign w19136 = w19128 & w19134;
assign v6049 = ~(w19135 | w19136);
assign w19137 = v6049;
assign w19138 = (~w19064 & w19075) | (~w19064 & w28044) | (w19075 & w28044);
assign v6050 = ~(w19076 | w19138);
assign w19139 = v6050;
assign w19140 = ~w19137 & w19139;
assign w19141 = (~w19076 & w19137) | (~w19076 & w28793) | (w19137 & w28793);
assign w19142 = (~w19058 & ~w19141) | (~w19058 & w28045) | (~w19141 & w28045);
assign w19143 = w19047 & ~w19142;
assign v6051 = ~(w19045 | w19143);
assign w19144 = v6051;
assign w19145 = w19032 & w19144;
assign w19146 = (~w19030 & ~w19032) | (~w19030 & w28046) | (~w19032 & w28046);
assign w19147 = ~w19010 & w19018;
assign v6052 = ~(w19019 | w19147);
assign w19148 = v6052;
assign w19149 = ~w19146 & w19148;
assign w19150 = (w28046 & w29535) | (w28046 & w29536) | (w29535 & w29536);
assign w19151 = ~w18998 & w19007;
assign v6053 = ~(w19008 | w19151);
assign w19152 = v6053;
assign w19153 = ~w19150 & w19152;
assign w19154 = (~w19008 & ~w19152) | (~w19008 & w28047) | (~w19152 & w28047);
assign w19155 = ~w18986 & w18995;
assign v6054 = ~(w18996 | w19155);
assign w19156 = v6054;
assign w19157 = ~w19154 & w19156;
assign w19158 = (~w18996 & w19154) | (~w18996 & w29317) | (w19154 & w29317);
assign v6055 = ~(w18973 | w18983);
assign w19159 = v6055;
assign v6056 = ~(w18984 | w19159);
assign w19160 = v6056;
assign w19161 = ~w19158 & w19160;
assign w19162 = (~w18984 & w19158) | (~w18984 & w29754) | (w19158 & w29754);
assign v6057 = ~(w18960 | w18970);
assign w19163 = v6057;
assign v6058 = ~(w18971 | w19163);
assign w19164 = v6058;
assign w19165 = ~w19162 & w19164;
assign w19166 = (~w18971 & w19162) | (~w18971 & w29537) | (w19162 & w29537);
assign v6059 = ~(w18947 | w18957);
assign w19167 = v6059;
assign v6060 = ~(w18958 | w19167);
assign w19168 = v6060;
assign w19169 = ~w19166 & w19168;
assign w19170 = (~w18958 & w19166) | (~w18958 & w29755) | (w19166 & w29755);
assign w19171 = ~w18934 & w18944;
assign v6061 = ~(w18945 | w19171);
assign w19172 = v6061;
assign w19173 = ~w19170 & w19172;
assign w19174 = (~w18945 & w19170) | (~w18945 & w29880) | (w19170 & w29880);
assign w19175 = ~w18921 & w18931;
assign v6062 = ~(w18932 | w19175);
assign w19176 = v6062;
assign w19177 = ~w19174 & w19176;
assign w19178 = (~w18932 & ~w19176) | (~w18932 & w28048) | (~w19176 & w28048);
assign w19179 = ~w18908 & w18918;
assign v6063 = ~(w18919 | w19179);
assign w19180 = v6063;
assign w19181 = ~w19178 & w19180;
assign w19182 = (~w18919 & ~w19180) | (~w18919 & w28049) | (~w19180 & w28049);
assign w19183 = ~w18895 & w18905;
assign v6064 = ~(w18906 | w19183);
assign w19184 = v6064;
assign w19185 = ~w19182 & w19184;
assign w19186 = (~w18906 & w19182) | (~w18906 & w30828) | (w19182 & w30828);
assign w19187 = w18882 & w18892;
assign v6065 = ~(w18893 | w19187);
assign w19188 = v6065;
assign w19189 = ~w19186 & w19188;
assign w19190 = (w28050 & w30829) | (w28050 & w30830) | (w30829 & w30830);
assign w19191 = (~w18877 & ~w19190) | (~w18877 & w30208) | (~w19190 & w30208);
assign w19192 = w18864 & w19191;
assign v6066 = ~(w18862 | w19192);
assign w19193 = v6066;
assign w19194 = (~w18846 & ~w19193) | (~w18846 & w28051) | (~w19193 & w28051);
assign w19195 = w18833 & w19194;
assign w19196 = (~w18831 & ~w18833) | (~w18831 & w28052) | (~w18833 & w28052);
assign w19197 = (~w18815 & w19196) | (~w18815 & w28337) | (w19196 & w28337);
assign w19198 = w18800 & ~w19197;
assign w19199 = (~w18798 & ~w18800) | (~w18798 & w28053) | (~w18800 & w28053);
assign w19200 = (~w18780 & ~w19199) | (~w18780 & w28338) | (~w19199 & w28338);
assign w19201 = w18765 & w19200;
assign w19202 = (~w18763 & ~w18765) | (~w18763 & w28339) | (~w18765 & w28339);
assign w19203 = (~w18745 & ~w19202) | (~w18745 & w30372) | (~w19202 & w30372);
assign w19204 = (~w18733 & ~w19203) | (~w18733 & w28340) | (~w19203 & w28340);
assign w19205 = w18716 & ~w19204;
assign w19206 = (~w18714 & ~w18716) | (~w18714 & w28341) | (~w18716 & w28341);
assign w19207 = w18703 & ~w19206;
assign w19208 = (~w18701 & w19206) | (~w18701 & w30643) | (w19206 & w30643);
assign v6067 = ~(w18681 | w18683);
assign w19209 = v6067;
assign v6068 = ~(w18684 | w19209);
assign w19210 = v6068;
assign w19211 = ~w19208 & w19210;
assign w19212 = (~w18684 & w19208) | (~w18684 & w31055) | (w19208 & w31055);
assign w19213 = w18670 & ~w19212;
assign w19214 = (~w18668 & ~w18670) | (~w18668 & w28342) | (~w18670 & w28342);
assign w19215 = w18644 & w18653;
assign v6069 = ~(w18654 | w19215);
assign w19216 = v6069;
assign w19217 = w19214 & w19216;
assign w19218 = (~w18654 & ~w19214) | (~w18654 & w31198) | (~w19214 & w31198);
assign w19219 = w18642 & w19218;
assign w19220 = (~w18640 & ~w18642) | (~w18640 & w30209) | (~w18642 & w30209);
assign v6070 = ~(w18623 | w18625);
assign w19221 = v6070;
assign v6071 = ~(w18626 | w19221);
assign w19222 = v6071;
assign w19223 = ~w19220 & w19222;
assign w19224 = w19220 & ~w19222;
assign v6072 = ~(w19223 | w19224);
assign w19225 = v6072;
assign w19226 = w10987 & w12406;
assign v6073 = ~(w13657 | w19226);
assign w19227 = v6073;
assign v6074 = ~(w18642 | w19218);
assign w19228 = v6074;
assign v6075 = ~(w19219 | w19228);
assign w19229 = v6075;
assign w19230 = w19227 & ~w19229;
assign v6076 = ~(w19214 | w19216);
assign w19231 = v6076;
assign v6077 = ~(w19217 | w19231);
assign w19232 = v6077;
assign w19233 = (w28343 & ~w12502) | (w28343 & w28794) | (~w12502 & w28794);
assign v6078 = ~(w11023 | w19233);
assign w19234 = v6078;
assign v6079 = ~(w12406 | w19234);
assign w19235 = v6079;
assign v6080 = ~(w11035 | w19235);
assign w19236 = v6080;
assign v6081 = ~(pi02 | w19236);
assign w19237 = v6081;
assign w19238 = w10986 & w12381;
assign w19239 = pi02 & ~w19238;
assign w19240 = w19236 & w19239;
assign v6082 = ~(w19237 | w19240);
assign w19241 = v6082;
assign w19242 = w19232 & w19241;
assign w19243 = ~w18670 & w19212;
assign v6083 = ~(w19213 | w19243);
assign w19244 = v6083;
assign w19245 = w11035 & ~w12406;
assign w19246 = w11023 & w12381;
assign v6084 = ~(w19245 | w19246);
assign w19247 = v6084;
assign w19248 = (w12505 & w28795) | (w12505 & w28796) | (w28795 & w28796);
assign v6085 = ~(pi02 | w19248);
assign w19249 = v6085;
assign w19250 = w10986 & w12311;
assign w19251 = pi02 & ~w19250;
assign w19252 = w19248 & w19251;
assign v6086 = ~(w19249 | w19252);
assign w19253 = v6086;
assign w19254 = w19244 & ~w19253;
assign w19255 = ~w19244 & w19253;
assign v6087 = ~(w19254 | w19255);
assign w19256 = v6087;
assign w19257 = w19208 & ~w19210;
assign v6088 = ~(w19211 | w19257);
assign w19258 = v6088;
assign w19259 = w11035 & w12381;
assign w19260 = w11023 & w12311;
assign v6089 = ~(w19259 | w19260);
assign w19261 = v6089;
assign w19262 = (w12387 & w28345) | (w12387 & w28346) | (w28345 & w28346);
assign w19263 = w10986 & w12271;
assign w19264 = pi02 & ~w19263;
assign w19265 = (~w12387 & w28347) | (~w12387 & w28348) | (w28347 & w28348);
assign v6090 = ~(w19262 | w19265);
assign w19266 = v6090;
assign w19267 = ~w19258 & w19266;
assign w19268 = w19258 & ~w19266;
assign v6091 = ~(w19267 | w19268);
assign w19269 = v6091;
assign w19270 = ~w18703 & w19206;
assign v6092 = ~(w19207 | w19270);
assign w19271 = v6092;
assign w19272 = w11035 & w12311;
assign w19273 = w11023 & w12271;
assign v6093 = ~(w19272 | w19273);
assign w19274 = v6093;
assign w19275 = (w12318 & w28797) | (w12318 & w28798) | (w28797 & w28798);
assign w19276 = w10986 & w12237;
assign w19277 = pi02 & ~w19276;
assign w19278 = (~w12318 & w28799) | (~w12318 & w28800) | (w28799 & w28800);
assign v6094 = ~(w19275 | w19278);
assign w19279 = v6094;
assign w19280 = ~w19271 & w19279;
assign w19281 = w19271 & ~w19279;
assign v6095 = ~(w19280 | w19281);
assign w19282 = v6095;
assign w19283 = ~w18716 & w19204;
assign v6096 = ~(w19205 | w19283);
assign w19284 = v6096;
assign w19285 = w11035 & w12271;
assign w19286 = w11023 & w12237;
assign v6097 = ~(w19285 | w19286);
assign w19287 = v6097;
assign w19288 = (~w12277 & w28801) | (~w12277 & w28802) | (w28801 & w28802);
assign w19289 = w10986 & w12155;
assign w19290 = pi02 & ~w19289;
assign w19291 = (w12277 & w28803) | (w12277 & w28804) | (w28803 & w28804);
assign v6098 = ~(w19288 | w19291);
assign w19292 = v6098;
assign w19293 = w19284 & ~w19292;
assign w19294 = ~w19284 & w19292;
assign v6099 = ~(w19293 | w19294);
assign w19295 = v6099;
assign w19296 = w11035 & w12237;
assign w19297 = w11023 & w12155;
assign v6100 = ~(w19296 | w19297);
assign w19298 = v6100;
assign w19299 = (~w12351 & w28805) | (~w12351 & w28806) | (w28805 & w28806);
assign w19300 = w10986 & w12084;
assign w19301 = pi02 & ~w19300;
assign w19302 = (w12351 & w28807) | (w12351 & w28808) | (w28807 & w28808);
assign v6101 = ~(w19299 | w19302);
assign w19303 = v6101;
assign v6102 = ~(w18733 | w18734);
assign w19304 = v6102;
assign v6103 = ~(w19203 | w19304);
assign w19305 = v6103;
assign w19306 = w19203 & w19304;
assign v6104 = ~(w19305 | w19306);
assign w19307 = v6104;
assign w19308 = ~w19303 & w19307;
assign w19309 = w19303 & ~w19307;
assign v6105 = ~(w19308 | w19309);
assign w19310 = v6105;
assign w19311 = w11035 & w12155;
assign w19312 = w11023 & w12084;
assign v6106 = ~(w19311 | w19312);
assign w19313 = v6106;
assign w19314 = (w12167 & w30210) | (w12167 & w30211) | (w30210 & w30211);
assign w19315 = w10986 & w11984;
assign w19316 = pi02 & ~w19315;
assign w19317 = (~w12167 & w30212) | (~w12167 & w30213) | (w30212 & w30213);
assign v6107 = ~(w19314 | w19317);
assign w19318 = v6107;
assign v6108 = ~(w18745 | w18746);
assign w19319 = v6108;
assign w19320 = w19202 & w19319;
assign v6109 = ~(w19202 | w19319);
assign w19321 = v6109;
assign v6110 = ~(w19320 | w19321);
assign w19322 = v6110;
assign w19323 = w19318 & w19322;
assign v6111 = ~(w19318 | w19322);
assign w19324 = v6111;
assign v6112 = ~(w18765 | w19200);
assign w19325 = v6112;
assign v6113 = ~(w19201 | w19325);
assign w19326 = v6113;
assign w19327 = w11035 & w12084;
assign w19328 = w11023 & w11984;
assign v6114 = ~(w19327 | w19328);
assign w19329 = v6114;
assign w19330 = (w12181 & w28809) | (w12181 & w28810) | (w28809 & w28810);
assign w19331 = w10986 & w11671;
assign w19332 = pi02 & ~w19331;
assign w19333 = (~w12181 & w28811) | (~w12181 & w28812) | (w28811 & w28812);
assign v6115 = ~(w19330 | w19333);
assign w19334 = v6115;
assign w19335 = w19326 & ~w19334;
assign w19336 = ~w19326 & w19334;
assign v6116 = ~(w19335 | w19336);
assign w19337 = v6116;
assign v6117 = ~(w18780 | w18781);
assign w19338 = v6117;
assign w19339 = w19199 & ~w19338;
assign w19340 = ~w19199 & w19338;
assign v6118 = ~(w19339 | w19340);
assign w19341 = v6118;
assign w19342 = ~w11992 & w28354;
assign w19343 = w11035 & w11984;
assign w19344 = w11023 & w11671;
assign v6119 = ~(w19343 | w19344);
assign w19345 = v6119;
assign w19346 = (~pi02 & w19342) | (~pi02 & w28813) | (w19342 & w28813);
assign w19347 = w10986 & w11673;
assign w19348 = pi02 & ~w19347;
assign w19349 = ~w19342 & w28814;
assign v6120 = ~(w19346 | w19349);
assign w19350 = v6120;
assign w19351 = w19341 & ~w19350;
assign w19352 = w11035 & w11673;
assign w19353 = w11023 & w11678;
assign v6121 = ~(w19352 | w19353);
assign w19354 = v6121;
assign w19355 = (w19354 & ~w12454) | (w19354 & w30214) | (~w12454 & w30214);
assign v6122 = ~(pi02 | w19355);
assign w19356 = v6122;
assign w19357 = w10986 & ~w11683;
assign w19358 = pi02 & ~w19357;
assign w19359 = w19355 & w19358;
assign v6123 = ~(w19356 | w19359);
assign w19360 = v6123;
assign v6124 = ~(w18815 | w18816);
assign w19361 = v6124;
assign w19362 = w19196 & ~w19361;
assign w19363 = ~w19196 & w19361;
assign v6125 = ~(w19362 | w19363);
assign w19364 = v6125;
assign w19365 = w19360 & ~w19364;
assign v6126 = ~(w18864 | w19191);
assign w19366 = v6126;
assign v6127 = ~(w19192 | w19366);
assign w19367 = v6127;
assign v6128 = ~(w18877 | w18878);
assign w19368 = v6128;
assign v6129 = ~(w19190 | w19368);
assign w19369 = v6129;
assign w19370 = w19190 & w19368;
assign v6130 = ~(w19369 | w19370);
assign w19371 = v6130;
assign w19372 = w19186 & ~w19188;
assign v6131 = ~(w19189 | w19372);
assign w19373 = v6131;
assign v6132 = ~(w4 | w13008);
assign w19374 = v6132;
assign w19375 = w11035 & ~w11695;
assign w19376 = w11023 & w11700;
assign v6133 = ~(w19375 | w19376);
assign w19377 = v6133;
assign w19378 = ~w19374 & w19377;
assign v6134 = ~(pi02 | w19378);
assign w19379 = v6134;
assign w19380 = w10986 & w11708;
assign w19381 = pi02 & ~w19380;
assign w19382 = w19378 & w19381;
assign v6135 = ~(w19379 | w19382);
assign w19383 = v6135;
assign w19384 = w19373 & ~w19383;
assign w19385 = ~w19373 & w19383;
assign w19386 = ~w4 & w12994;
assign w19387 = w11023 & w11708;
assign w19388 = w11035 & w11700;
assign v6136 = ~(w19387 | w19388);
assign w19389 = v6136;
assign w19390 = ~w19386 & w19389;
assign v6137 = ~(pi02 | w19390);
assign w19391 = v6137;
assign w19392 = w10986 & w11711;
assign w19393 = pi02 & ~w19392;
assign w19394 = w19390 & w19393;
assign v6138 = ~(w19391 | w19394);
assign w19395 = v6138;
assign w19396 = w19182 & ~w19184;
assign v6139 = ~(w19185 | w19396);
assign w19397 = v6139;
assign w19398 = ~w19395 & w19397;
assign w19399 = w19395 & ~w19397;
assign w19400 = ~w4 & w13178;
assign w19401 = w11035 & w11708;
assign w19402 = w11023 & w11711;
assign v6140 = ~(w19401 | w19402);
assign w19403 = v6140;
assign w19404 = ~w19400 & w19403;
assign v6141 = ~(pi02 | w19404);
assign w19405 = v6141;
assign w19406 = w10986 & w11714;
assign w19407 = pi02 & ~w19406;
assign w19408 = w19404 & w19407;
assign v6142 = ~(w19405 | w19408);
assign w19409 = v6142;
assign w19410 = w19178 & ~w19180;
assign v6143 = ~(w19181 | w19410);
assign w19411 = v6143;
assign w19412 = w19409 & ~w19411;
assign w19413 = w11035 & w11711;
assign w19414 = w11023 & w11714;
assign v6144 = ~(w19413 | w19414);
assign w19415 = v6144;
assign w19416 = pi02 & ~w19415;
assign w19417 = w1 & w13194;
assign w19418 = ~w4 & w13194;
assign w19419 = w10986 & w11720;
assign w19420 = pi02 & ~w19419;
assign w19421 = w19415 & ~w19420;
assign w19422 = ~w19418 & w19421;
assign v6145 = ~(w19417 | w19422);
assign w19423 = v6145;
assign w19424 = ~w19416 & w19423;
assign w19425 = w19174 & ~w19176;
assign v6146 = ~(w19177 | w19425);
assign w19426 = v6146;
assign v6147 = ~(w19424 | w19426);
assign w19427 = v6147;
assign w19428 = w19170 & ~w19172;
assign v6148 = ~(w19173 | w19428);
assign w19429 = v6148;
assign w19430 = ~w4 & w13514;
assign w19431 = w11035 & w11714;
assign w19432 = w11023 & w11720;
assign v6149 = ~(w19431 | w19432);
assign w19433 = v6149;
assign w19434 = ~w19430 & w19433;
assign v6150 = ~(pi02 | w19434);
assign w19435 = v6150;
assign w19436 = w10986 & w11723;
assign w19437 = pi02 & ~w19436;
assign w19438 = w19434 & w19437;
assign v6151 = ~(w19435 | w19438);
assign w19439 = v6151;
assign w19440 = w19429 & ~w19439;
assign w19441 = w19424 & w19426;
assign w19442 = ~w19429 & w19439;
assign w19443 = w19166 & ~w19168;
assign v6152 = ~(w19169 | w19443);
assign w19444 = v6152;
assign v6153 = ~(w4 | w13310);
assign w19445 = v6153;
assign w19446 = w11035 & w11720;
assign w19447 = w11023 & w11723;
assign v6154 = ~(w19446 | w19447);
assign w19448 = v6154;
assign w19449 = ~w19445 & w19448;
assign w19450 = pi02 & ~w19449;
assign w19451 = w10986 & w11726;
assign w19452 = pi02 & ~w19451;
assign w19453 = w19449 & ~w19452;
assign v6155 = ~(w19450 | w19453);
assign w19454 = v6155;
assign w19455 = w19444 & w19454;
assign w19456 = w19162 & ~w19164;
assign v6156 = ~(w19165 | w19456);
assign w19457 = v6156;
assign w19458 = w3 & w13864;
assign w19459 = w1 & w13864;
assign w19460 = w10987 & ~w11734;
assign w19461 = w11035 & w11726;
assign w19462 = w11023 & w11729;
assign v6157 = ~(w19461 | w19462);
assign w19463 = v6157;
assign w19464 = pi02 & w19463;
assign v6158 = ~(pi02 | w19463);
assign w19465 = v6158;
assign v6159 = ~(w19464 | w19465);
assign w19466 = v6159;
assign v6160 = ~(w19460 | w19466);
assign w19467 = v6160;
assign w19468 = ~w19459 & w19467;
assign v6161 = ~(w19458 | w19468);
assign w19469 = v6161;
assign w19470 = w19158 & ~w19160;
assign v6162 = ~(w19161 | w19470);
assign w19471 = v6162;
assign w19472 = w19469 & ~w19471;
assign w19473 = w19154 & ~w19156;
assign v6163 = ~(w19157 | w19473);
assign w19474 = v6163;
assign w19475 = w1 & ~w13703;
assign w19476 = w11023 & ~w11734;
assign w19477 = w11035 & w11729;
assign v6164 = ~(w19476 | w19477);
assign w19478 = v6164;
assign w19479 = w10987 & w11737;
assign w19480 = w19478 & ~w19479;
assign w19481 = ~w10988 & w19480;
assign w19482 = ~w13703 & w19481;
assign w19483 = ~pi02 & w19478;
assign w19484 = pi02 & ~w19480;
assign v6165 = ~(w19483 | w19484);
assign w19485 = v6165;
assign v6166 = ~(w19482 | w19485);
assign w19486 = v6166;
assign v6167 = ~(w19475 | w19486);
assign w19487 = v6167;
assign v6168 = ~(w19474 | w19487);
assign w19488 = v6168;
assign w19489 = w11023 & w11737;
assign w19490 = w11035 & ~w11734;
assign v6169 = ~(w19489 | w19490);
assign w19491 = v6169;
assign v6170 = ~(pi02 | w13882);
assign w19492 = v6170;
assign w19493 = w10987 & w11740;
assign v6171 = ~(w19492 | w19493);
assign w19494 = v6171;
assign w19495 = ~w10988 & w19494;
assign w19496 = w19491 & ~w19495;
assign w19497 = pi02 & ~w19491;
assign w19498 = w1 & w13882;
assign v6172 = ~(w19497 | w19498);
assign w19499 = v6172;
assign w19500 = ~w19496 & w19499;
assign w19501 = w19150 & ~w19152;
assign v6173 = ~(w19153 | w19501);
assign w19502 = v6173;
assign v6174 = ~(w19500 | w19502);
assign w19503 = v6174;
assign w19504 = ~w19047 & w19142;
assign v6175 = ~(w19143 | w19504);
assign w19505 = v6175;
assign w19506 = w3 & ~w14331;
assign w19507 = (w1 & w11841) | (w1 & w29318) | (w11841 & w29318);
assign w19508 = w11023 & w11759;
assign w19509 = w11035 & w11748;
assign v6176 = ~(w19508 | w19509);
assign w19510 = v6176;
assign w19511 = pi02 & ~w19510;
assign w19512 = w10986 & w11761;
assign w19513 = pi02 & ~w19512;
assign w19514 = w19510 & ~w19513;
assign v6177 = ~(w19511 | w19514);
assign w19515 = v6177;
assign w19516 = ~w19507 & w19515;
assign v6178 = ~(w19506 | w19516);
assign w19517 = v6178;
assign v6179 = ~(w19058 | w19059);
assign w19518 = v6179;
assign w19519 = w19141 & w19518;
assign v6180 = ~(w19141 | w19518);
assign w19520 = v6180;
assign v6181 = ~(w19519 | w19520);
assign w19521 = v6181;
assign v6182 = ~(w19517 | w19521);
assign w19522 = v6182;
assign w19523 = w19517 & w19521;
assign w19524 = w1 & w14356;
assign w19525 = w11023 & w11761;
assign w19526 = w11035 & w11759;
assign v6183 = ~(w19525 | w19526);
assign w19527 = v6183;
assign v6184 = ~(pi02 | w19527);
assign w19528 = v6184;
assign v6185 = ~(pi02 | w14356);
assign w19529 = v6185;
assign w19530 = w10987 & ~w11771;
assign w19531 = ~w19526 & w29031;
assign w19532 = ~w10988 & w19531;
assign w19533 = (~w19528 & w19529) | (~w19528 & w28355) | (w19529 & w28355);
assign v6186 = ~(w19524 | w19533);
assign w19534 = v6186;
assign w19535 = w19137 & ~w19139;
assign v6187 = ~(w19140 | w19535);
assign w19536 = v6187;
assign w19537 = w19534 & w19536;
assign w19538 = w11035 & w11761;
assign w19539 = (w11023 & ~w11766) | (w11023 & w29032) | (~w11766 & w29032);
assign v6188 = ~(w19538 | w19539);
assign w19540 = v6188;
assign w19541 = (~w14383 & w28540) | (~w14383 & w28541) | (w28540 & w28541);
assign w19542 = w10986 & w11768;
assign w19543 = pi02 & ~w19542;
assign w19544 = (w14383 & w28542) | (w14383 & w28543) | (w28542 & w28543);
assign v6189 = ~(w19541 | w19544);
assign w19545 = v6189;
assign w19546 = w19121 & w19134;
assign v6190 = ~(w19135 | w19546);
assign w19547 = v6190;
assign w19548 = ~w19545 & w19547;
assign w19549 = w19545 & ~w19547;
assign v6191 = ~(w19117 | w19119);
assign w19550 = v6191;
assign v6192 = ~(w19120 | w19550);
assign w19551 = v6192;
assign w19552 = ~w4 & w14409;
assign w19553 = w11023 & w11768;
assign w19554 = (w11035 & ~w11766) | (w11035 & w28544) | (~w11766 & w28544);
assign v6193 = ~(w19553 | w19554);
assign w19555 = v6193;
assign w19556 = w10986 & w11776;
assign w19557 = pi02 & ~w19556;
assign w19558 = ~w19552 & w28357;
assign w19559 = (pi02 & w19552) | (pi02 & w28358) | (w19552 & w28358);
assign v6194 = ~(w19558 | w19559);
assign w19560 = v6194;
assign w19561 = w19551 & w19560;
assign v6195 = ~(w19551 | w19560);
assign w19562 = v6195;
assign w19563 = w1 & w14461;
assign w19564 = w11533 & w28359;
assign w19565 = w11023 & w11776;
assign v6196 = ~(w19564 | w19565);
assign w19566 = v6196;
assign v6197 = ~(pi02 | w19566);
assign w19567 = v6197;
assign v6198 = ~(pi02 | w14461);
assign w19568 = v6198;
assign w19569 = w10987 & w11784;
assign w19570 = w19566 & ~w19569;
assign w19571 = ~w10988 & w19570;
assign w19572 = (~w19567 & w19568) | (~w19567 & w28190) | (w19568 & w28190);
assign w19573 = w18459 & w19103;
assign v6199 = ~(w19104 | w19573);
assign w19574 = v6199;
assign w19575 = w19116 & ~w19574;
assign w19576 = ~w19116 & w19574;
assign v6200 = ~(w19575 | w19576);
assign w19577 = v6200;
assign w19578 = ~w19572 & w28545;
assign w19579 = (w19577 & w19572) | (w19577 & w28360) | (w19572 & w28360);
assign w19580 = w19095 & ~w19100;
assign v6201 = ~(w19101 | w19580);
assign w19581 = v6201;
assign w19582 = w10987 & w11798;
assign w19583 = ~w11792 & w28546;
assign w19584 = w11023 & w11803;
assign v6202 = ~(w19583 | w19584);
assign w19585 = v6202;
assign w19586 = (~w14569 & w28361) | (~w14569 & w28362) | (w28361 & w28362);
assign w19587 = ~pi02 & pi03;
assign w19588 = w11800 & w19587;
assign w19589 = (w14569 & w28547) | (w14569 & w28548) | (w28547 & w28548);
assign w19590 = pi01 & w11798;
assign w19591 = pi00 & w11803;
assign v6203 = ~(w4 | w14609);
assign w19592 = v6203;
assign v6204 = ~(w19591 | w19592);
assign w19593 = v6204;
assign w19594 = w19593 & w28549;
assign w19595 = ~pi03 & w11800;
assign v6205 = ~(w19594 | w19595);
assign w19596 = v6205;
assign w19597 = pi02 & ~w19596;
assign w19598 = w19586 & w19597;
assign v6206 = ~(w19589 | w19598);
assign w19599 = v6206;
assign w19600 = w19581 & ~w19599;
assign w19601 = ~w19598 & w28550;
assign w19602 = ~w4 & w14547;
assign w19603 = w10987 & w11803;
assign w19604 = w11035 & w11784;
assign w19605 = w11023 & w11793;
assign w19606 = ~w19604 & w28551;
assign w19607 = ~w19602 & w28191;
assign w19608 = (pi02 & w19602) | (pi02 & w28192) | (w19602 & w28192);
assign v6207 = ~(w19607 | w19608);
assign w19609 = v6207;
assign w19610 = (~w19600 & ~w19609) | (~w19600 & w29033) | (~w19609 & w29033);
assign w19611 = w11035 & w11776;
assign w19612 = w11023 & w11784;
assign v6208 = ~(w19611 | w19612);
assign w19613 = v6208;
assign w19614 = (w14504 & w28193) | (w14504 & w28194) | (w28193 & w28194);
assign w19615 = w10986 & w11793;
assign w19616 = pi02 & ~w19615;
assign w19617 = (~w14504 & w28057) | (~w14504 & w28058) | (w28057 & w28058);
assign v6209 = ~(w19614 | w19617);
assign w19618 = v6209;
assign v6210 = ~(w19610 | w19618);
assign w19619 = v6210;
assign w19620 = pi05 & ~w19101;
assign w19621 = ~w19094 & w19620;
assign w19622 = w19094 & ~w19620;
assign v6211 = ~(w19621 | w19622);
assign w19623 = v6211;
assign w19624 = (w19623 & ~w19610) | (w19623 & w28195) | (~w19610 & w28195);
assign v6212 = ~(w19619 | w19624);
assign w19625 = v6212;
assign w19626 = (~w19578 & w19625) | (~w19578 & w29034) | (w19625 & w29034);
assign w19627 = (~w19561 & w19626) | (~w19561 & w28059) | (w19626 & w28059);
assign w19628 = (~w19548 & w19627) | (~w19548 & w28552) | (w19627 & w28552);
assign v6213 = ~(w19534 | w19536);
assign w19629 = v6213;
assign v6214 = ~(w19628 | w19629);
assign w19630 = v6214;
assign v6215 = ~(w19537 | w19630);
assign w19631 = v6215;
assign w19632 = (~w19522 & w19631) | (~w19522 & w28196) | (w19631 & w28196);
assign v6216 = ~(w19505 | w19632);
assign w19633 = v6216;
assign v6217 = ~(w19032 | w19144);
assign w19634 = v6217;
assign v6218 = ~(w19145 | w19634);
assign w19635 = v6218;
assign w19636 = w11035 & ~w11745;
assign w19637 = w11023 & w11748;
assign v6219 = ~(w19636 | w19637);
assign w19638 = v6219;
assign w19639 = (w19638 & ~w13948) | (w19638 & w28555) | (~w13948 & w28555);
assign w19640 = pi02 & ~w19639;
assign w19641 = w10986 & w11759;
assign w19642 = pi02 & ~w19641;
assign w19643 = w19639 & ~w19642;
assign v6220 = ~(w19640 | w19643);
assign w19644 = v6220;
assign w19645 = (~w28554 & w29035) | (~w28554 & w29036) | (w29035 & w29036);
assign v6221 = ~(w19635 | w19645);
assign w19646 = v6221;
assign w19647 = ~w19633 & w19646;
assign w19648 = ~w4 & w14300;
assign w19649 = w11035 & w11740;
assign w19650 = w11023 & ~w11745;
assign v6222 = ~(w19649 | w19650);
assign w19651 = v6222;
assign w19652 = ~w19648 & w19651;
assign v6223 = ~(pi02 | w19652);
assign w19653 = v6223;
assign w19654 = w10986 & w11748;
assign w19655 = pi02 & ~w19654;
assign w19656 = w19652 & w19655;
assign v6224 = ~(w19653 | w19656);
assign w19657 = v6224;
assign w19658 = (~w19657 & ~w19646) | (~w19657 & w29319) | (~w19646 & w29319);
assign w19659 = w19635 & w19645;
assign w19660 = w19633 & w19635;
assign v6225 = ~(w19659 | w19660);
assign w19661 = v6225;
assign w19662 = w19146 & ~w19148;
assign v6226 = ~(w19149 | w19662);
assign w19663 = v6226;
assign w19664 = w19661 & ~w19663;
assign w19665 = ~w4 & w14288;
assign w19666 = w11023 & w11740;
assign w19667 = w11035 & w11737;
assign v6227 = ~(w19666 | w19667);
assign w19668 = v6227;
assign w19669 = ~w19665 & w19668;
assign w19670 = pi02 & ~w19669;
assign w19671 = w10986 & ~w11745;
assign w19672 = pi02 & ~w19671;
assign w19673 = w19669 & ~w19672;
assign v6228 = ~(w19670 | w19673);
assign w19674 = v6228;
assign w19675 = (w19674 & ~w19664) | (w19674 & w29320) | (~w19664 & w29320);
assign w19676 = w19657 & w19661;
assign w19677 = ~w19647 & w19663;
assign w19678 = ~w19676 & w19677;
assign v6229 = ~(w19675 | w19678);
assign w19679 = v6229;
assign w19680 = w19502 & w19500;
assign w19681 = (~w19679 & w29756) | (~w19679 & w29757) | (w29756 & w29757);
assign w19682 = w19474 & w19487;
assign w19683 = (~w28197 & w28363) | (~w28197 & w28364) | (w28363 & w28364);
assign w19684 = ~w19681 & w19683;
assign w19685 = (w29758 & w29881) | (w29758 & w29882) | (w29881 & w29882);
assign v6230 = ~(w4 | w13737);
assign w19686 = v6230;
assign w19687 = w11035 & w11723;
assign w19688 = w11023 & w11726;
assign v6231 = ~(w19687 | w19688);
assign w19689 = v6231;
assign w19690 = ~w19686 & w19689;
assign w19691 = pi02 & ~w19690;
assign w19692 = w10986 & w11729;
assign w19693 = pi02 & ~w19692;
assign w19694 = w19690 & ~w19693;
assign v6232 = ~(w19691 | w19694);
assign w19695 = v6232;
assign w19696 = (~w19684 & w29759) | (~w19684 & w29760) | (w29759 & w29760);
assign v6233 = ~(w19685 | w19696);
assign w19697 = v6233;
assign v6234 = ~(w19444 | w19454);
assign w19698 = v6234;
assign w19699 = (~w19455 & w19697) | (~w19455 & w29883) | (w19697 & w29883);
assign w19700 = (~w19427 & ~w28198) | (~w19427 & w30057) | (~w28198 & w30057);
assign w19701 = ~w19409 & w19411;
assign w19702 = (~w19701 & ~w19700) | (~w19701 & w30215) | (~w19700 & w30215);
assign w19703 = (~w19398 & w19702) | (~w19398 & w29884) | (w19702 & w29884);
assign w19704 = ~w4 & w12694;
assign w19705 = w11035 & w11689;
assign w19706 = w11023 & ~w11695;
assign v6235 = ~(w19705 | w19706);
assign w19707 = v6235;
assign w19708 = ~w19704 & w19707;
assign w19709 = pi02 & ~w19708;
assign w19710 = w10986 & w11700;
assign w19711 = pi02 & ~w19710;
assign w19712 = w19708 & ~w19711;
assign v6236 = ~(w19709 | w19712);
assign w19713 = v6236;
assign w19714 = (~w29886 & w30831) | (~w29886 & w30832) | (w30831 & w30832);
assign v6237 = ~(w4 | w12842);
assign w19715 = v6237;
assign w19716 = w11035 & w11686;
assign w19717 = w11023 & w11689;
assign v6238 = ~(w19716 | w19717);
assign w19718 = v6238;
assign w19719 = ~w19715 & w19718;
assign w19720 = pi02 & ~w19719;
assign w19721 = w10986 & ~w11695;
assign w19722 = pi02 & ~w19721;
assign w19723 = w19719 & ~w19722;
assign v6239 = ~(w19720 | w19723);
assign w19724 = v6239;
assign w19725 = (~w30058 & w30833) | (~w30058 & w30834) | (w30833 & w30834);
assign w19726 = ~w19714 & w30059;
assign w19727 = w11035 & ~w11683;
assign w19728 = w11023 & w11686;
assign v6240 = ~(w19727 | w19728);
assign w19729 = v6240;
assign w19730 = (w19729 & ~w12610) | (w19729 & w29887) | (~w12610 & w29887);
assign v6241 = ~(pi02 | w19730);
assign w19731 = v6241;
assign w19732 = w10986 & w11689;
assign w19733 = pi02 & ~w19732;
assign w19734 = w19730 & w19733;
assign v6242 = ~(w19731 | w19734);
assign w19735 = v6242;
assign v6243 = ~(w18846 | w18847);
assign w19736 = v6243;
assign w19737 = (w19736 & w19192) | (w19736 & w30060) | (w19192 & w30060);
assign w19738 = ~w19192 & w30061;
assign v6244 = ~(w19737 | w19738);
assign w19739 = v6244;
assign w19740 = w19735 & ~w19739;
assign v6245 = ~(w19726 | w19740);
assign w19741 = v6245;
assign w19742 = ~w19735 & w19739;
assign w19743 = w11035 & w11678;
assign w19744 = w11023 & ~w11683;
assign v6246 = ~(w19743 | w19744);
assign w19745 = v6246;
assign w19746 = (~w29889 & w30062) | (~w29889 & w30063) | (w30062 & w30063);
assign w19747 = w10986 & w11686;
assign w19748 = pi02 & ~w19747;
assign w19749 = (w29889 & w30064) | (w29889 & w30065) | (w30064 & w30065);
assign v6247 = ~(w19746 | w19749);
assign w19750 = v6247;
assign v6248 = ~(w18833 | w19194);
assign w19751 = v6248;
assign v6249 = ~(w19195 | w19751);
assign w19752 = v6249;
assign w19753 = (~w19742 & ~w19752) | (~w19742 & w30066) | (~w19752 & w30066);
assign w19754 = w19750 & ~w19752;
assign w19755 = (~w30835 & w31056) | (~w30835 & w31057) | (w31056 & w31057);
assign w19756 = ~w19365 & w19755;
assign w19757 = ~w19360 & w19364;
assign w19758 = ~w18800 & w19197;
assign v6250 = ~(w19198 | w19758);
assign w19759 = v6250;
assign w19760 = w11035 & w11671;
assign w19761 = w11023 & w11673;
assign v6251 = ~(w19760 | w19761);
assign w19762 = v6251;
assign w19763 = (w12469 & w28559) | (w12469 & w28560) | (w28559 & w28560);
assign w19764 = w10986 & w11678;
assign w19765 = pi02 & ~w19764;
assign w19766 = (~w12469 & w28561) | (~w12469 & w28562) | (w28561 & w28562);
assign v6252 = ~(w19763 | w19766);
assign w19767 = v6252;
assign w19768 = w19759 & ~w19767;
assign v6253 = ~(w19757 | w19768);
assign w19769 = v6253;
assign w19770 = ~w19756 & w19769;
assign w19771 = ~w19759 & w19767;
assign w19772 = (w28144 & w29890) | (w28144 & w29891) | (w29890 & w29891);
assign w19773 = (~w19351 & ~w19772) | (~w19351 & w28815) | (~w19772 & w28815);
assign w19774 = w19337 & ~w19773;
assign v6254 = ~(w19335 | w19774);
assign w19775 = v6254;
assign w19776 = (~w19323 & ~w28200) | (~w19323 & w28365) | (~w28200 & w28365);
assign w19777 = w19310 & w19776;
assign w19778 = (~w19308 & ~w19310) | (~w19308 & w29892) | (~w19310 & w29892);
assign w19779 = w19295 & ~w19778;
assign w19780 = (~w19293 & w19778) | (~w19293 & w30526) | (w19778 & w30526);
assign w19781 = w19282 & w19780;
assign w19782 = w19269 & w19781;
assign w19783 = w19269 & w19280;
assign w19784 = (~w19267 & ~w19269) | (~w19267 & w28201) | (~w19269 & w28201);
assign w19785 = ~w19782 & w19784;
assign w19786 = w19256 & w19785;
assign v6255 = ~(w19232 | w19241);
assign w19787 = v6255;
assign v6256 = ~(w19242 | w19787);
assign w19788 = v6256;
assign w19789 = ~w19254 & w19788;
assign w19790 = w19788 & w29893;
assign w19791 = (~w19242 & ~w19789) | (~w19242 & w28202) | (~w19789 & w28202);
assign w19792 = ~w19227 & w19229;
assign v6257 = ~(w19230 | w19792);
assign w19793 = v6257;
assign w19794 = ~w19791 & w19793;
assign w19795 = (~w19230 & w19791) | (~w19230 & w31199) | (w19791 & w31199);
assign w19796 = ~w19794 & w29894;
assign w19797 = (~w19223 & ~w19795) | (~w19223 & w28366) | (~w19795 & w28366);
assign v6258 = ~(w18611 | w18627);
assign w19798 = v6258;
assign v6259 = ~(w18628 | w19798);
assign w19799 = v6259;
assign w19800 = (~w19795 & w29895) | (~w19795 & w29896) | (w29895 & w29896);
assign w19801 = (w19797 & w29037) | (w19797 & w29038) | (w29037 & w29038);
assign w19802 = (~w19797 & w29039) | (~w19797 & w29040) | (w29039 & w29040);
assign v6260 = ~(w17508 | w18034);
assign w19803 = v6260;
assign v6261 = ~(w18035 | w19803);
assign w19804 = v6261;
assign w19805 = (w29040 & w31280) | (w29040 & w31281) | (w31280 & w31281);
assign w19806 = (~w18035 & ~w19802) | (~w18035 & w31058) | (~w19802 & w31058);
assign w19807 = w17506 & ~w19806;
assign w19808 = (w17015 & w17012) | (w17015 & w29539) | (w17012 & w29539);
assign v6262 = ~(w17016 | w19808);
assign w19809 = v6262;
assign w19810 = ~w19807 & w29321;
assign w19811 = w16138 & ~w16561;
assign v6263 = ~(w16562 | w19811);
assign w19812 = v6263;
assign w19813 = (w19812 & w19810) | (w19812 & w29540) | (w19810 & w29540);
assign w19814 = (~w19810 & w29897) | (~w19810 & w29898) | (w29897 & w29898);
assign w19815 = ~w15394 & w15751;
assign v6264 = ~(w15752 | w19815);
assign w19816 = v6264;
assign w19817 = (~w19810 & w30218) | (~w19810 & w30219) | (w30218 & w30219);
assign w19818 = (w19810 & w30373) | (w19810 & w30374) | (w30373 & w30374);
assign w19819 = w15067 & ~w15391;
assign w19820 = (~w19810 & w31282) | (~w19810 & w31283) | (w31282 & w31283);
assign v6265 = ~(w15063 | w19820);
assign w19821 = v6265;
assign w19822 = ~w14778 & w14923;
assign v6266 = ~(w14924 | w19822);
assign w19823 = v6266;
assign w19824 = ~w19821 & w19823;
assign v6267 = ~(w14924 | w19824);
assign w19825 = v6267;
assign v6268 = ~(w14776 | w19825);
assign w19826 = v6268;
assign v6269 = ~(w14775 | w19826);
assign w19827 = v6269;
assign w19828 = w14219 & ~w19827;
assign v6270 = ~(w14217 | w19828);
assign w19829 = v6270;
assign w19830 = w14095 & ~w19829;
assign v6271 = ~(w14093 | w19830);
assign w19831 = v6271;
assign w19832 = w13620 & ~w13826;
assign w19833 = w19831 & ~w19832;
assign v6272 = ~(w13827 | w19833);
assign w19834 = v6272;
assign w19835 = w13618 & w19834;
assign v6273 = ~(w13616 | w19835);
assign w19836 = v6273;
assign w19837 = ~w13400 & w13494;
assign v6274 = ~(w13495 | w19837);
assign w19838 = v6274;
assign w19839 = ~w19836 & w19838;
assign v6275 = ~(w13495 | w19839);
assign w19840 = v6275;
assign w19841 = ~w13398 & w19840;
assign v6276 = ~(w13397 | w19841);
assign w19842 = v6276;
assign w19843 = w13082 & w19842;
assign v6277 = ~(w13080 | w19843);
assign w19844 = v6277;
assign w19845 = ~w12933 & w19844;
assign v6278 = ~(w12932 | w19845);
assign w19846 = v6278;
assign w19847 = ~w12834 & w19846;
assign v6279 = ~(w12833 | w19847);
assign w19848 = v6279;
assign w19849 = w12774 & ~w19848;
assign v6280 = ~(w12772 | w19849);
assign w19850 = v6280;
assign w19851 = w12537 & ~w19850;
assign w19852 = ~w12537 & w19850;
assign v6281 = ~(w19851 | w19852);
assign w19853 = v6281;
assign v6282 = ~(w12535 | w19851);
assign w19854 = v6282;
assign v6283 = ~(w12401 | w12413);
assign w19855 = v6283;
assign v6284 = ~(w12362 | w12398);
assign w19856 = v6284;
assign v6285 = ~(w12347 | w12359);
assign w19857 = v6285;
assign w19858 = ~w214 & w2429;
assign w19859 = w5843 & w19858;
assign w19860 = w12202 & w19859;
assign w19861 = w3895 & w19860;
assign w19862 = w3877 & w19861;
assign v6286 = ~(w564 | w674);
assign w19863 = v6286;
assign w19864 = w4044 & w19863;
assign w19865 = w2835 & w19864;
assign w19866 = w1597 & w1889;
assign w19867 = w4023 & w19866;
assign w19868 = w19865 & w19867;
assign w19869 = w19862 & w19868;
assign w19870 = ~w12346 & w19869;
assign w19871 = w12346 & ~w19869;
assign v6287 = ~(w19870 | w19871);
assign w19872 = v6287;
assign w19873 = w928 & ~w12277;
assign w19874 = w3406 & w12271;
assign w19875 = w3402 & w12237;
assign w19876 = w3399 & w12155;
assign v6288 = ~(w19875 | w19876);
assign w19877 = v6288;
assign w19878 = ~w19874 & w19877;
assign w19879 = ~w19873 & w19878;
assign w19880 = ~w19872 & w19879;
assign w19881 = w19872 & ~w19879;
assign v6289 = ~(w19880 | w19881);
assign w19882 = v6289;
assign w19883 = ~w19857 & w19882;
assign w19884 = w19857 & ~w19882;
assign v6290 = ~(w19883 | w19884);
assign w19885 = v6290;
assign w19886 = ~w19856 & w19885;
assign w19887 = w19856 & ~w19885;
assign v6291 = ~(w19886 | w19887);
assign w19888 = v6291;
assign v6292 = ~(pi26 | w38);
assign w19889 = v6292;
assign w19890 = w1563 & ~w19889;
assign w19891 = w3529 & ~w12506;
assign w19892 = w3760 & ~w12406;
assign w19893 = w3767 & w12311;
assign w19894 = w3763 & w12381;
assign v6293 = ~(w19893 | w19894);
assign w19895 = v6293;
assign w19896 = ~w19892 & w19895;
assign w19897 = ~w19891 & w19896;
assign w19898 = ~pi29 & w19897;
assign w19899 = pi29 & ~w19897;
assign v6294 = ~(w19898 | w19899);
assign w19900 = v6294;
assign w19901 = ~w19890 & w19900;
assign w19902 = w19890 & ~w19900;
assign v6295 = ~(w19901 | w19902);
assign w19903 = v6295;
assign w19904 = w19888 & w19903;
assign v6296 = ~(w19888 | w19903);
assign w19905 = v6296;
assign v6297 = ~(w19904 | w19905);
assign w19906 = v6297;
assign w19907 = w19855 & ~w19906;
assign w19908 = ~w19855 & w19906;
assign v6298 = ~(w19907 | w19908);
assign w19909 = v6298;
assign v6299 = ~(w19854 | w19909);
assign w19910 = v6299;
assign w19911 = w19854 & w19909;
assign v6300 = ~(w19910 | w19911);
assign w19912 = v6300;
assign w19913 = w19853 & ~w19912;
assign w19914 = ~w19853 & w19912;
assign v6301 = ~(w19913 | w19914);
assign w19915 = v6301;
assign w19916 = ~w12774 & w19848;
assign v6302 = ~(w19849 | w19916);
assign w19917 = v6302;
assign w19918 = w19853 & w19917;
assign v6303 = ~(w19853 | w19917);
assign w19919 = v6303;
assign v6304 = ~(w12833 | w12834);
assign w19920 = v6304;
assign w19921 = w19846 & ~w19920;
assign w19922 = ~w19846 & w19920;
assign v6305 = ~(w19921 | w19922);
assign w19923 = v6305;
assign w19924 = w19917 & ~w19923;
assign w19925 = ~w19917 & w19923;
assign v6306 = ~(w12932 | w12933);
assign w19926 = v6306;
assign w19927 = w19844 & w19926;
assign v6307 = ~(w19844 | w19926);
assign w19928 = v6307;
assign v6308 = ~(w19927 | w19928);
assign w19929 = v6308;
assign v6309 = ~(w19923 | w19929);
assign w19930 = v6309;
assign w19931 = w19923 & w19929;
assign v6310 = ~(w13082 | w19842);
assign w19932 = v6310;
assign v6311 = ~(w19843 | w19932);
assign w19933 = v6311;
assign w19934 = w19929 & ~w19933;
assign w19935 = ~w19929 & w19933;
assign v6312 = ~(w13397 | w13398);
assign w19936 = v6312;
assign v6313 = ~(w19840 | w19936);
assign w19937 = v6313;
assign w19938 = w19840 & w19936;
assign v6314 = ~(w19937 | w19938);
assign w19939 = v6314;
assign w19940 = w19933 & ~w19939;
assign w19941 = ~w19933 & w19939;
assign w19942 = w19836 & w19837;
assign w19943 = w13495 & ~w19836;
assign v6315 = ~(w19942 | w19943);
assign w19944 = v6315;
assign v6316 = ~(w19936 | w19944);
assign w19945 = v6316;
assign w19946 = w19936 & w19944;
assign v6317 = ~(w19945 | w19946);
assign w19947 = v6317;
assign v6318 = ~(w13827 | w19832);
assign w19948 = v6318;
assign w19949 = ~w19831 & w19948;
assign v6319 = ~(w19832 | w19949);
assign w19950 = v6319;
assign w19951 = ~w13618 & w19950;
assign v6320 = ~(w19835 | w19951);
assign w19952 = v6320;
assign w19953 = w19836 & ~w19838;
assign v6321 = ~(w19839 | w19953);
assign w19954 = v6321;
assign w19955 = w19952 & w19954;
assign v6322 = ~(w19952 | w19954);
assign w19956 = v6322;
assign w19957 = w19831 & ~w19948;
assign v6323 = ~(w19949 | w19957);
assign w19958 = v6323;
assign v6324 = ~(w19952 | w19958);
assign w19959 = v6324;
assign w19960 = ~w14095 & w19829;
assign v6325 = ~(w19830 | w19960);
assign w19961 = v6325;
assign w19962 = w19958 & w19961;
assign v6326 = ~(w19958 | w19961);
assign w19963 = v6326;
assign v6327 = ~(w19962 | w19963);
assign w19964 = v6327;
assign w19965 = ~w14219 & w19827;
assign v6328 = ~(w19828 | w19965);
assign w19966 = v6328;
assign v6329 = ~(w19961 | w19966);
assign w19967 = v6329;
assign v6330 = ~(w14775 | w14776);
assign w19968 = v6330;
assign v6331 = ~(w19825 | w19968);
assign w19969 = v6331;
assign w19970 = w19825 & w19968;
assign v6332 = ~(w19969 | w19970);
assign w19971 = v6332;
assign w19972 = w19966 & ~w19971;
assign w19973 = w19821 & ~w19823;
assign v6333 = ~(w19824 | w19973);
assign w19974 = v6333;
assign w19975 = ~w19971 & w19974;
assign v6334 = ~(w15392 | w19819);
assign w19976 = v6334;
assign w19977 = ~w19818 & w19976;
assign w19978 = (~w19819 & w19818) | (~w19819 & w30645) | (w19818 & w30645);
assign w19979 = ~w15065 & w19978;
assign v6335 = ~(w19820 | w19979);
assign w19980 = v6335;
assign w19981 = w19974 & w19980;
assign w19982 = w19818 & ~w19976;
assign v6336 = ~(w19977 | w19982);
assign w19983 = v6336;
assign w19984 = w19980 & w19983;
assign w19985 = (w19810 & w30646) | (w19810 & w30647) | (w30646 & w30647);
assign v6337 = ~(w19817 | w19985);
assign w19986 = v6337;
assign w19987 = w19983 & w19986;
assign w19988 = (w19810 & w30220) | (w19810 & w30221) | (w30220 & w30221);
assign v6338 = ~(w19814 | w19988);
assign w19989 = v6338;
assign w19990 = w19986 & w19989;
assign w19991 = ~w19810 & w29541;
assign v6339 = ~(w19813 | w19991);
assign w19992 = v6339;
assign w19993 = w19989 & ~w19992;
assign w19994 = ~w19989 & w19992;
assign v6340 = ~(w19993 | w19994);
assign w19995 = v6340;
assign w19996 = (~w19809 & w19807) | (~w19809 & w30069) | (w19807 & w30069);
assign v6341 = ~(w19810 | w19996);
assign w19997 = v6341;
assign v6342 = ~(w19992 | w19997);
assign w19998 = v6342;
assign w19999 = ~w17506 & w19806;
assign v6343 = ~(w19807 | w19999);
assign w20000 = v6343;
assign w20001 = ~w19997 & w20000;
assign w20002 = w19997 & ~w20000;
assign v6344 = ~(w20001 | w20002);
assign w20003 = v6344;
assign w20004 = (~w29040 & w31284) | (~w29040 & w31285) | (w31284 & w31285);
assign v6345 = ~(w19805 | w20004);
assign w20005 = v6345;
assign w20006 = w20000 & w20005;
assign w20007 = (~w19797 & w29041) | (~w19797 & w29042) | (w29041 & w29042);
assign v6346 = ~(w19801 | w20007);
assign w20008 = v6346;
assign w20009 = w20005 & ~w20008;
assign w20010 = (w19795 & w29899) | (w19795 & w29900) | (w29899 & w29900);
assign v6347 = ~(w19800 | w20010);
assign w20011 = v6347;
assign v6348 = ~(w20008 | w20011);
assign w20012 = v6348;
assign w20013 = (~w19225 & w19794) | (~w19225 & w29901) | (w19794 & w29901);
assign v6349 = ~(w19796 | w20013);
assign w20014 = v6349;
assign w20015 = ~w20011 & w20014;
assign w20016 = w20011 & ~w20014;
assign v6350 = ~(w20015 | w20016);
assign w20017 = v6350;
assign v6351 = ~(w19230 | w19791);
assign w20018 = v6351;
assign w20019 = w19791 & ~w19792;
assign v6352 = ~(w20018 | w20019);
assign w20020 = v6352;
assign w20021 = w19225 & w20020;
assign v6353 = ~(w19225 | w20020);
assign w20022 = v6353;
assign v6354 = ~(w20021 | w20022);
assign w20023 = v6354;
assign w20024 = w19786 & ~w19788;
assign w20025 = w19254 & ~w19788;
assign w20026 = ~w19790 & w28203;
assign w20027 = w19791 & ~w19793;
assign v6355 = ~(w19794 | w20027);
assign w20028 = v6355;
assign v6356 = ~(w20026 | w20028);
assign w20029 = v6356;
assign v6357 = ~(w19256 | w19785);
assign w20030 = v6357;
assign v6358 = ~(w19786 | w20030);
assign w20031 = v6358;
assign w20032 = w28203 & w30070;
assign w20033 = (~w20030 & w19790) | (~w20030 & w28204) | (w19790 & w28204);
assign v6359 = ~(w19282 | w19780);
assign w20034 = v6359;
assign v6360 = ~(w19269 | w19280);
assign w20035 = v6360;
assign v6361 = ~(w19783 | w20035);
assign w20036 = v6361;
assign w20037 = (~w19782 & w20036) | (~w19782 & w28205) | (w20036 & w28205);
assign v6362 = ~(w19781 | w20034);
assign w20038 = v6362;
assign w20039 = ~w19295 & w19778;
assign v6363 = ~(w19779 | w20039);
assign w20040 = v6363;
assign w20041 = ~w20038 & w20040;
assign v6364 = ~(w19310 | w19776);
assign w20042 = v6364;
assign v6365 = ~(w19777 | w20042);
assign w20043 = v6365;
assign v6366 = ~(w20040 | w20043);
assign w20044 = v6366;
assign w20045 = w20040 & w20043;
assign w20046 = ~w19337 & w19773;
assign v6367 = ~(w19774 | w20046);
assign w20047 = v6367;
assign v6368 = ~(w20043 | w20047);
assign w20048 = v6368;
assign v6369 = ~(w19323 | w19324);
assign w20049 = v6369;
assign w20050 = w19775 & w20049;
assign v6370 = ~(w19775 | w20049);
assign w20051 = v6370;
assign v6371 = ~(w20050 | w20051);
assign w20052 = v6371;
assign v6372 = ~(w20048 | w20052);
assign w20053 = v6372;
assign v6373 = ~(w20045 | w20053);
assign w20054 = v6373;
assign v6374 = ~(w20044 | w20054);
assign w20055 = v6374;
assign v6375 = ~(w20041 | w20055);
assign w20056 = v6375;
assign w20057 = w20037 & w20056;
assign w20058 = w20036 & w20038;
assign w20059 = w20038 & ~w20040;
assign w20060 = (~w20059 & ~w20036) | (~w20059 & w30071) | (~w20036 & w30071);
assign w20061 = ~w20057 & w20060;
assign v6376 = ~(w19781 | w20036);
assign w20062 = v6376;
assign w20063 = (~w19782 & w20036) | (~w19782 & w28206) | (w20036 & w28206);
assign w20064 = ~w19785 & w20063;
assign w20065 = ~w20064 & w28060;
assign w20066 = (~w19256 & w20064) | (~w19256 & w28061) | (w20064 & w28061);
assign v6377 = ~(w20065 | w20066);
assign w20067 = v6377;
assign w20068 = w20061 & w20067;
assign w20069 = w20031 & ~w20063;
assign w20070 = (~w20069 & ~w20067) | (~w20069 & w28062) | (~w20067 & w28062);
assign w20071 = (w28062 & w30648) | (w28062 & w30649) | (w30648 & w30649);
assign v6378 = ~(w20032 | w20071);
assign w20072 = v6378;
assign w20073 = w20026 & w20028;
assign w20074 = (~w20029 & ~w20072) | (~w20029 & w28207) | (~w20072 & w28207);
assign v6379 = ~(w20023 | w20074);
assign w20075 = v6379;
assign w20076 = w20014 & ~w20028;
assign w20077 = (~w20076 & w20074) | (~w20076 & w29902) | (w20074 & w29902);
assign w20078 = w20017 & ~w20077;
assign w20079 = (~w20015 & ~w20017) | (~w20015 & w28063) | (~w20017 & w28063);
assign w20080 = w20008 & w20011;
assign v6380 = ~(w20012 | w20080);
assign w20081 = v6380;
assign w20082 = (~w28063 & w31200) | (~w28063 & w31201) | (w31200 & w31201);
assign w20083 = (~w20012 & w20079) | (~w20012 & w28564) | (w20079 & w28564);
assign w20084 = ~w20005 & w20008;
assign v6381 = ~(w20009 | w20084);
assign w20085 = v6381;
assign w20086 = (~w20079 & w31286) | (~w20079 & w31287) | (w31286 & w31287);
assign w20087 = (~w20009 & w20083) | (~w20009 & w28817) | (w20083 & w28817);
assign v6382 = ~(w20000 | w20005);
assign w20088 = v6382;
assign v6383 = ~(w20006 | w20088);
assign w20089 = v6383;
assign w20090 = ~w20087 & w20089;
assign w20091 = (~w20006 & w20087) | (~w20006 & w29043) | (w20087 & w29043);
assign w20092 = w20003 & ~w20091;
assign w20093 = (~w20001 & w20091) | (~w20001 & w30072) | (w20091 & w30072);
assign w20094 = w19992 & w19997;
assign v6384 = ~(w19998 | w20094);
assign w20095 = v6384;
assign w20096 = ~w20093 & w20095;
assign w20097 = (~w19998 & w20093) | (~w19998 & w29322) | (w20093 & w29322);
assign w20098 = w19995 & ~w20097;
assign w20099 = (~w19993 & w20097) | (~w19993 & w29542) | (w20097 & w29542);
assign v6385 = ~(w19986 | w19989);
assign w20100 = v6385;
assign v6386 = ~(w19990 | w20100);
assign w20101 = v6386;
assign w20102 = (~w20097 & w30222) | (~w20097 & w30223) | (w30222 & w30223);
assign v6387 = ~(w19983 | w19986);
assign w20103 = v6387;
assign v6388 = ~(w19987 | w20103);
assign w20104 = v6388;
assign w20105 = (~w20099 & w30224) | (~w20099 & w30225) | (w30224 & w30225);
assign w20106 = (w20099 & w30375) | (w20099 & w30376) | (w30375 & w30376);
assign v6389 = ~(w19980 | w19983);
assign w20107 = v6389;
assign v6390 = ~(w19984 | w20107);
assign w20108 = v6390;
assign w20109 = ~w20106 & w20108;
assign w20110 = (~w19984 & w20106) | (~w19984 & w30226) | (w20106 & w30226);
assign v6391 = ~(w19974 | w19980);
assign w20111 = v6391;
assign v6392 = ~(w19981 | w20111);
assign w20112 = v6392;
assign w20113 = ~w20110 & w20112;
assign w20114 = (~w19981 & w20110) | (~w19981 & w30650) | (w20110 & w30650);
assign w20115 = w19971 & ~w19974;
assign v6393 = ~(w19975 | w20115);
assign w20116 = v6393;
assign w20117 = ~w20114 & w20116;
assign w20118 = (~w19975 & w20114) | (~w19975 & w30838) | (w20114 & w30838);
assign w20119 = ~w19966 & w19971;
assign v6394 = ~(w19972 | w20119);
assign w20120 = v6394;
assign w20121 = ~w20118 & w20120;
assign w20122 = (~w19972 & ~w20120) | (~w19972 & w28065) | (~w20120 & w28065);
assign w20123 = w19961 & w19966;
assign w20124 = (~w19967 & ~w20122) | (~w19967 & w28367) | (~w20122 & w28367);
assign w20125 = w19964 & w20124;
assign w20126 = (~w19962 & ~w19964) | (~w19962 & w28066) | (~w19964 & w28066);
assign w20127 = w19952 & w19958;
assign v6395 = ~(w19959 | w20127);
assign w20128 = v6395;
assign w20129 = w20126 & w20128;
assign w20130 = (~w19959 & ~w20128) | (~w19959 & w28067) | (~w20128 & w28067);
assign w20131 = ~w19956 & w20130;
assign v6396 = ~(w19955 | w20131);
assign w20132 = v6396;
assign w20133 = w19947 & ~w20132;
assign w20134 = ~w19939 & w19954;
assign v6397 = ~(w20133 | w20134);
assign w20135 = v6397;
assign v6398 = ~(w19941 | w20135);
assign w20136 = v6398;
assign v6399 = ~(w19940 | w20136);
assign w20137 = v6399;
assign w20138 = ~w19935 & w20137;
assign v6400 = ~(w19934 | w20138);
assign w20139 = v6400;
assign w20140 = ~w19931 & w20139;
assign v6401 = ~(w19930 | w20140);
assign w20141 = v6401;
assign v6402 = ~(w19925 | w20141);
assign w20142 = v6402;
assign v6403 = ~(w19924 | w20142);
assign w20143 = v6403;
assign v6404 = ~(w19919 | w20143);
assign w20144 = v6404;
assign v6405 = ~(w19918 | w20144);
assign w20145 = v6405;
assign w20146 = w19915 & ~w20145;
assign w20147 = (~w19913 & ~w19915) | (~w19913 & w28068) | (~w19915 & w28068);
assign v6406 = ~(w19883 | w19886);
assign w20148 = v6406;
assign w20149 = w4078 & w4188;
assign w20150 = w3304 & w20149;
assign w20151 = ~w267 & w20150;
assign w20152 = w3981 & w20151;
assign w20153 = ~w172 & w20152;
assign v6407 = ~(w12346 | w20153);
assign w20154 = v6407;
assign w20155 = w12346 & w20153;
assign v6408 = ~(w20154 | w20155);
assign w20156 = v6408;
assign w20157 = w19890 & w20156;
assign v6409 = ~(w19890 | w20156);
assign w20158 = v6409;
assign v6410 = ~(w20157 | w20158);
assign w20159 = v6410;
assign v6411 = ~(w19870 | w19879);
assign w20160 = v6411;
assign v6412 = ~(w19871 | w20160);
assign w20161 = v6412;
assign w20162 = ~w20159 & w20161;
assign w20163 = w20159 & ~w20161;
assign v6413 = ~(w20162 | w20163);
assign w20164 = v6413;
assign w20165 = w928 & w12318;
assign w20166 = w3406 & w12311;
assign w20167 = w3402 & w12271;
assign w20168 = w3399 & w12237;
assign v6414 = ~(w20167 | w20168);
assign w20169 = v6414;
assign w20170 = ~w20166 & w20169;
assign w20171 = ~w20165 & w20170;
assign w20172 = w20164 & ~w20171;
assign w20173 = ~w20164 & w20171;
assign v6415 = ~(w20172 | w20173);
assign w20174 = v6415;
assign w20175 = w3529 & w12505;
assign v6416 = ~(w3760 | w3763);
assign w20176 = v6416;
assign w20177 = w3766 & w12381;
assign w20178 = w20176 & ~w20177;
assign w20179 = ~w20175 & w20178;
assign w20180 = pi29 & w20179;
assign v6417 = ~(pi29 | w20179);
assign w20181 = v6417;
assign v6418 = ~(w20180 | w20181);
assign w20182 = v6418;
assign w20183 = w20174 & ~w20182;
assign w20184 = ~w20174 & w20182;
assign v6419 = ~(w20183 | w20184);
assign w20185 = v6419;
assign w20186 = w20148 & ~w20185;
assign w20187 = ~w20148 & w20185;
assign v6420 = ~(w20186 | w20187);
assign w20188 = v6420;
assign v6421 = ~(w19901 | w19904);
assign w20189 = v6421;
assign w20190 = ~w20188 & w20189;
assign w20191 = w20188 & ~w20189;
assign v6422 = ~(w20190 | w20191);
assign w20192 = v6422;
assign w20193 = (~w19850 & w29044) | (~w19850 & w29045) | (w29044 & w29045);
assign v6423 = ~(w19908 | w20193);
assign w20194 = v6423;
assign w20195 = w20192 & ~w20194;
assign w20196 = ~w20192 & w20194;
assign v6424 = ~(w20195 | w20196);
assign w20197 = v6424;
assign w20198 = ~w19912 & w20197;
assign w20199 = w19912 & ~w20197;
assign v6425 = ~(w20198 | w20199);
assign w20200 = v6425;
assign w20201 = ~w20147 & w20200;
assign w20202 = w20147 & ~w20200;
assign v6426 = ~(w20201 | w20202);
assign w20203 = v6426;
assign w20204 = w11035 & w20197;
assign w20205 = w11023 & ~w19912;
assign v6427 = ~(w20204 | w20205);
assign w20206 = v6427;
assign w20207 = (w20206 & ~w20203) | (w20206 & w29046) | (~w20203 & w29046);
assign v6428 = ~(pi02 | w20207);
assign w20208 = v6428;
assign w20209 = w10986 & w19853;
assign w20210 = pi02 & ~w20209;
assign w20211 = w20207 & w20210;
assign v6429 = ~(w20208 | w20211);
assign w20212 = v6429;
assign w20213 = ~w19947 & w20132;
assign v6430 = ~(w20133 | w20213);
assign w20214 = v6430;
assign w20215 = w8141 & w20214;
assign w20216 = w8926 & ~w19939;
assign w20217 = w8140 & w19952;
assign w20218 = w8526 & w19954;
assign v6431 = ~(w20217 | w20218);
assign w20219 = v6431;
assign w20220 = ~w20216 & w20219;
assign w20221 = ~w20215 & w20220;
assign w20222 = ~pi08 & w20221;
assign w20223 = pi08 & ~w20221;
assign v6432 = ~(w20222 | w20223);
assign w20224 = v6432;
assign w20225 = w7765 & w19961;
assign w20226 = w7466 & w19966;
assign w20227 = w7177 & ~w19971;
assign v6433 = ~(w20226 | w20227);
assign w20228 = v6433;
assign w20229 = ~w20225 & w20228;
assign w20230 = pi11 & ~w20229;
assign v6434 = ~(w19967 | w20123);
assign w20231 = v6434;
assign w20232 = ~w20122 & w20231;
assign w20233 = w20122 & ~w20231;
assign v6435 = ~(w20232 | w20233);
assign w20234 = v6435;
assign w20235 = w9464 & w20234;
assign v6436 = ~(w20230 | w20235);
assign w20236 = v6436;
assign w20237 = w7178 & w20234;
assign w20238 = ~pi11 & w20229;
assign w20239 = ~w20237 & w20238;
assign w20240 = w20236 & ~w20239;
assign w20241 = w3525 & w20047;
assign w20242 = w4152 & w20047;
assign w20243 = pi26 & w20242;
assign w20244 = ~w20047 & w20052;
assign w20245 = w20047 & ~w20052;
assign v6437 = ~(w20244 | w20245);
assign w20246 = v6437;
assign w20247 = w4153 & w20246;
assign w20248 = w4155 & ~w20052;
assign w20249 = w4158 & w20047;
assign v6438 = ~(w20248 | w20249);
assign w20250 = v6438;
assign w20251 = ~w20247 & w20250;
assign w20252 = ~w20247 & w30839;
assign w20253 = (pi26 & w20247) | (pi26 & w31059) | (w20247 & w31059);
assign v6439 = ~(w20047 | w20052);
assign w20254 = v6439;
assign v6440 = ~(w20043 | w20254);
assign w20255 = v6440;
assign w20256 = w20043 & w20254;
assign v6441 = ~(w20255 | w20256);
assign w20257 = v6441;
assign w20258 = ~w2873 & w20047;
assign w20259 = (~w20258 & ~w20257) | (~w20258 & w30840) | (~w20257 & w30840);
assign w20260 = w4155 & w20043;
assign w20261 = w4158 & ~w20052;
assign v6442 = ~(w20260 | w20261);
assign w20262 = v6442;
assign w20263 = w20259 & w20262;
assign w20264 = ~w20253 & w20263;
assign w20265 = w20263 & w31060;
assign w20266 = w20241 & w20265;
assign v6443 = ~(w20241 | w20265);
assign w20267 = v6443;
assign v6444 = ~(w20266 | w20267);
assign w20268 = v6444;
assign v6445 = ~(w20044 | w20045);
assign w20269 = v6445;
assign w20270 = w20053 & ~w20269;
assign w20271 = ~w20053 & w20269;
assign v6446 = ~(w20270 | w20271);
assign w20272 = v6446;
assign w20273 = w4158 & w20043;
assign w20274 = w4155 & w20040;
assign v6447 = ~(w2873 | w20052);
assign w20275 = v6447;
assign v6448 = ~(w20274 | w20275);
assign w20276 = v6448;
assign w20277 = (w20272 & w30841) | (w20272 & w30842) | (w30841 & w30842);
assign w20278 = (~w20272 & w30843) | (~w20272 & w30844) | (w30843 & w30844);
assign v6449 = ~(w20277 | w20278);
assign w20279 = v6449;
assign w20280 = w20268 & w20279;
assign w20281 = (~w20266 & ~w20279) | (~w20266 & w31061) | (~w20279 & w31061);
assign w20282 = pi29 & w20241;
assign w20283 = w3529 & w20246;
assign w20284 = w3760 & ~w20052;
assign w20285 = w3763 & w20047;
assign v6450 = ~(w20284 | w20285);
assign w20286 = v6450;
assign w20287 = ~w20283 & w20286;
assign w20288 = ~w20283 & w31062;
assign w20289 = w20282 & ~w20287;
assign v6451 = ~(w20288 | w20289);
assign w20290 = v6451;
assign v6452 = ~(w20041 | w20059);
assign w20291 = v6452;
assign w20292 = w20055 & ~w20291;
assign w20293 = ~w20055 & w20291;
assign v6453 = ~(w20292 | w20293);
assign w20294 = v6453;
assign w20295 = w4155 & ~w20038;
assign w20296 = ~w2873 & w20043;
assign w20297 = w4158 & w20040;
assign v6454 = ~(w20296 | w20297);
assign w20298 = v6454;
assign w20299 = ~w20295 & w20298;
assign w20300 = (w20294 & w30845) | (w20294 & w30846) | (w30845 & w30846);
assign w20301 = (~w20294 & w30847) | (~w20294 & w30848) | (w30847 & w30848);
assign v6455 = ~(w20300 | w20301);
assign w20302 = v6455;
assign w20303 = w20290 & w20302;
assign v6456 = ~(w20290 | w20302);
assign w20304 = v6456;
assign v6457 = ~(w20303 | w20304);
assign w20305 = v6457;
assign w20306 = ~w20281 & w20305;
assign w20307 = w20281 & ~w20305;
assign v6458 = ~(w20306 | w20307);
assign w20308 = v6458;
assign w20309 = (~w20070 & w20032) | (~w20070 & w28070) | (w20032 & w28070);
assign w20310 = ~w20032 & w20071;
assign v6459 = ~(w20309 | w20310);
assign w20311 = v6459;
assign w20312 = (w4764 & w20309) | (w4764 & w30652) | (w20309 & w30652);
assign w20313 = w4763 & ~w20063;
assign w20314 = w4913 & ~w20026;
assign w20315 = w4836 & w20031;
assign w20316 = ~w20312 & w30227;
assign w20317 = (~pi23 & w20312) | (~pi23 & w30228) | (w20312 & w30228);
assign v6460 = ~(w20316 | w20317);
assign w20318 = v6460;
assign w20319 = w20308 & ~w20318;
assign v6461 = ~(w20268 | w20279);
assign w20320 = v6461;
assign v6462 = ~(w20280 | w20320);
assign w20321 = v6462;
assign v6463 = ~(w20061 | w20067);
assign w20322 = v6463;
assign v6464 = ~(w20068 | w20322);
assign w20323 = v6464;
assign w20324 = w4913 & w20031;
assign w20325 = w4763 & ~w20038;
assign w20326 = w4836 & ~w20063;
assign v6465 = ~(w20325 | w20326);
assign w20327 = v6465;
assign w20328 = ~w20324 & w20327;
assign w20329 = (~w20323 & w30377) | (~w20323 & w30378) | (w30377 & w30378);
assign w20330 = (w20323 & w30379) | (w20323 & w30380) | (w30379 & w30380);
assign v6466 = ~(w20329 | w20330);
assign w20331 = v6466;
assign w20332 = w20321 & w20331;
assign w20333 = w20253 & ~w20263;
assign v6467 = ~(w20264 | w20333);
assign w20334 = v6467;
assign w20335 = w20037 & ~w20058;
assign w20336 = (~w20059 & w20055) | (~w20059 & w30653) | (w20055 & w30653);
assign w20337 = ~w20335 & w20336;
assign w20338 = w20335 & ~w20336;
assign v6468 = ~(w20337 | w20338);
assign w20339 = v6468;
assign w20340 = w4913 & ~w20063;
assign w20341 = w4763 & w20040;
assign w20342 = w4836 & ~w20038;
assign v6469 = ~(w20341 | w20342);
assign w20343 = v6469;
assign w20344 = (w20339 & w30381) | (w20339 & w30382) | (w30381 & w30382);
assign w20345 = (~w20339 & w30383) | (~w20339 & w30384) | (w30383 & w30384);
assign v6470 = ~(w20344 | w20345);
assign w20346 = v6470;
assign w20347 = w20334 & w20346;
assign w20348 = w20243 & ~w20251;
assign v6471 = ~(w20252 | w20348);
assign w20349 = v6471;
assign w20350 = w4913 & ~w20038;
assign w20351 = w4763 & w20043;
assign w20352 = (~w20351 & ~w20040) | (~w20351 & w30654) | (~w20040 & w30654);
assign w20353 = ~w20350 & w20352;
assign w20354 = (w20294 & w30385) | (w20294 & w30386) | (w30385 & w30386);
assign w20355 = (~w20294 & w30387) | (~w20294 & w30388) | (w30387 & w30388);
assign v6472 = ~(w20354 | w20355);
assign w20356 = v6472;
assign w20357 = w20349 & w20356;
assign w20358 = w10 & w20047;
assign w20359 = pi23 & w20358;
assign w20360 = w4764 & w20246;
assign w20361 = w4836 & w20047;
assign w20362 = w4913 & ~w20052;
assign v6473 = ~(w20361 | w20362);
assign w20363 = v6473;
assign w20364 = ~w20360 & w20363;
assign w20365 = ~w20360 & w30655;
assign w20366 = (pi23 & w20360) | (pi23 & w30849) | (w20360 & w30849);
assign w20367 = w4763 & w20047;
assign w20368 = (~w20367 & ~w20257) | (~w20367 & w30656) | (~w20257 & w30656);
assign w20369 = w4913 & w20043;
assign w20370 = w4836 & ~w20052;
assign v6474 = ~(w20369 | w20370);
assign w20371 = v6474;
assign w20372 = w20368 & w20371;
assign w20373 = ~w20366 & w20372;
assign w20374 = w20372 & w30850;
assign w20375 = w20242 & w20374;
assign v6475 = ~(w20242 | w20374);
assign w20376 = v6475;
assign v6476 = ~(w20375 | w20376);
assign w20377 = v6476;
assign w20378 = w4836 & w20043;
assign w20379 = w4763 & ~w20052;
assign w20380 = (~w20379 & ~w20040) | (~w20379 & w30657) | (~w20040 & w30657);
assign w20381 = ~w20378 & w20380;
assign w20382 = (w20272 & w30658) | (w20272 & w30659) | (w30658 & w30659);
assign w20383 = (~w20272 & w30660) | (~w20272 & w30661) | (w30660 & w30661);
assign v6477 = ~(w20382 | w20383);
assign w20384 = v6477;
assign w20385 = w20377 & w20384;
assign w20386 = (~w20375 & ~w20384) | (~w20375 & w30851) | (~w20384 & w30851);
assign v6478 = ~(w20349 | w20356);
assign w20387 = v6478;
assign v6479 = ~(w20357 | w20387);
assign w20388 = v6479;
assign w20389 = ~w20386 & w20388;
assign w20390 = (~w20357 & ~w20388) | (~w20357 & w30662) | (~w20388 & w30662);
assign v6480 = ~(w20334 | w20346);
assign w20391 = v6480;
assign v6481 = ~(w20347 | w20391);
assign w20392 = v6481;
assign w20393 = ~w20390 & w20392;
assign v6482 = ~(w20347 | w20393);
assign w20394 = v6482;
assign v6483 = ~(w20321 | w20331);
assign w20395 = v6483;
assign v6484 = ~(w20332 | w20395);
assign w20396 = v6484;
assign w20397 = ~w20394 & w20396;
assign v6485 = ~(w20332 | w20397);
assign w20398 = v6485;
assign w20399 = ~w20308 & w20318;
assign v6486 = ~(w20319 | w20399);
assign w20400 = v6486;
assign w20401 = ~w20398 & w20400;
assign w20402 = (~w20319 & ~w20400) | (~w20319 & w30389) | (~w20400 & w30389);
assign w20403 = (~w20303 & ~w20305) | (~w20303 & w30528) | (~w20305 & w30528);
assign w20404 = (pi29 & w20283) | (pi29 & w31202) | (w20283 & w31202);
assign w20405 = w3767 & w20047;
assign w20406 = (~w20405 & ~w20257) | (~w20405 & w31063) | (~w20257 & w31063);
assign w20407 = w3760 & w20043;
assign w20408 = w3763 & ~w20052;
assign v6487 = ~(w20407 | w20408);
assign w20409 = v6487;
assign w20410 = w20406 & w20409;
assign w20411 = ~w20404 & w20410;
assign w20412 = w20404 & ~w20410;
assign v6488 = ~(w20411 | w20412);
assign w20413 = v6488;
assign w20414 = (~w20036 & w31064) | (~w20036 & w31065) | (w31064 & w31065);
assign w20415 = w4158 & ~w20038;
assign w20416 = ~w2873 & w20040;
assign v6489 = ~(w20415 | w20416);
assign w20417 = v6489;
assign w20418 = ~w20414 & w20417;
assign w20419 = (w20339 & w30852) | (w20339 & w30853) | (w30852 & w30853);
assign w20420 = (~w20339 & w30854) | (~w20339 & w30855) | (w30854 & w30855);
assign v6490 = ~(w20419 | w20420);
assign w20421 = v6490;
assign w20422 = w20413 & w20421;
assign v6491 = ~(w20413 | w20421);
assign w20423 = v6491;
assign v6492 = ~(w20422 | w20423);
assign w20424 = v6492;
assign w20425 = w20403 & ~w20424;
assign w20426 = ~w20403 & w20424;
assign v6493 = ~(w20425 | w20426);
assign w20427 = v6493;
assign v6494 = ~(w20029 | w20073);
assign w20428 = v6494;
assign w20429 = w20072 & w20428;
assign v6495 = ~(w20072 | w20428);
assign w20430 = v6495;
assign v6496 = ~(w20429 | w20430);
assign w20431 = v6496;
assign w20432 = w4763 & w20031;
assign w20433 = (~w20432 & w20028) | (~w20432 & w30529) | (w20028 & w30529);
assign w20434 = w4836 & ~w20026;
assign w20435 = w20433 & ~w20434;
assign w20436 = (~w20431 & w30390) | (~w20431 & w30391) | (w30390 & w30391);
assign w20437 = (w20431 & w30392) | (w20431 & w30393) | (w30392 & w30393);
assign v6497 = ~(w20436 | w20437);
assign w20438 = v6497;
assign w20439 = w20427 & ~w20438;
assign w20440 = ~w20427 & w20438;
assign v6498 = ~(w20439 | w20440);
assign w20441 = v6498;
assign w20442 = ~w20402 & w20441;
assign w20443 = w20402 & ~w20441;
assign v6499 = ~(w20442 | w20443);
assign w20444 = v6499;
assign w20445 = (w28063 & w29047) | (w28063 & w29048) | (w29047 & w29048);
assign v6500 = ~(w20082 | w20445);
assign w20446 = v6500;
assign w20447 = w5531 & ~w20011;
assign w20448 = w5610 & ~w20008;
assign v6501 = ~(w20447 | w20448);
assign w20449 = v6501;
assign w20450 = w5113 & w20014;
assign w20451 = w20449 & ~w20450;
assign w20452 = (~w20446 & w30394) | (~w20446 & w30395) | (w30394 & w30395);
assign w20453 = (w20446 & w30396) | (w20446 & w30397) | (w30396 & w30397);
assign v6502 = ~(w20452 | w20453);
assign w20454 = v6502;
assign w20455 = w20444 & ~w20454;
assign w20456 = w20398 & ~w20400;
assign v6503 = ~(w20401 | w20456);
assign w20457 = v6503;
assign w20458 = ~w20017 & w20077;
assign v6504 = ~(w20078 | w20458);
assign w20459 = v6504;
assign w20460 = w5610 & ~w20011;
assign w20461 = w5531 & w20014;
assign w20462 = w5113 & ~w20028;
assign v6505 = ~(w20461 | w20462);
assign w20463 = v6505;
assign w20464 = ~w20460 & w20463;
assign w20465 = (~w20459 & w30398) | (~w20459 & w30399) | (w30398 & w30399);
assign w20466 = (w20459 & w30400) | (w20459 & w30401) | (w30400 & w30401);
assign v6506 = ~(w20465 | w20466);
assign w20467 = v6506;
assign w20468 = w20457 & w20467;
assign w20469 = w20394 & ~w20396;
assign v6507 = ~(w20397 | w20469);
assign w20470 = v6507;
assign w20471 = w20023 & w20074;
assign v6508 = ~(w20075 | w20471);
assign w20472 = v6508;
assign w20473 = w5531 & ~w20028;
assign w20474 = w5610 & w20014;
assign v6509 = ~(w20473 | w20474);
assign w20475 = v6509;
assign w20476 = w5113 & ~w20026;
assign w20477 = (~w20472 & w30231) | (~w20472 & w30232) | (w30231 & w30232);
assign w20478 = (w20472 & w30233) | (w20472 & w30234) | (w30233 & w30234);
assign v6510 = ~(w20477 | w20478);
assign w20479 = v6510;
assign w20480 = w20470 & ~w20479;
assign w20481 = w20390 & ~w20392;
assign v6511 = ~(w20393 | w20481);
assign w20482 = v6511;
assign w20483 = w5610 & ~w20028;
assign w20484 = w5113 & w20031;
assign w20485 = w5531 & ~w20026;
assign v6512 = ~(w20484 | w20485);
assign w20486 = v6512;
assign w20487 = ~w20483 & w20486;
assign w20488 = (w20431 & w29905) | (w20431 & w29906) | (w29905 & w29906);
assign w20489 = (~w20431 & w29907) | (~w20431 & w29908) | (w29907 & w29908);
assign v6513 = ~(w20488 | w20489);
assign w20490 = v6513;
assign w20491 = w20482 & w20490;
assign w20492 = w20386 & ~w20388;
assign v6514 = ~(w20389 | w20492);
assign w20493 = v6514;
assign w20494 = (w5610 & ~w28203) | (w5610 & w29909) | (~w28203 & w29909);
assign w20495 = w5113 & ~w20063;
assign w20496 = w5531 & w20031;
assign v6515 = ~(w20495 | w20496);
assign w20497 = v6515;
assign w20498 = (~w20309 & w30663) | (~w20309 & w30664) | (w30663 & w30664);
assign w20499 = (w20309 & w30665) | (w20309 & w30666) | (w30665 & w30666);
assign v6516 = ~(w20498 | w20499);
assign w20500 = v6516;
assign w20501 = w20493 & w20500;
assign v6517 = ~(w20377 | w20384);
assign w20502 = v6517;
assign v6518 = ~(w20385 | w20502);
assign w20503 = v6518;
assign w20504 = w5610 & w20031;
assign w20505 = w5113 & ~w20038;
assign w20506 = w5531 & ~w20063;
assign v6519 = ~(w20505 | w20506);
assign w20507 = v6519;
assign w20508 = ~w20504 & w20507;
assign w20509 = (~w20323 & w29768) | (~w20323 & w29769) | (w29768 & w29769);
assign w20510 = (w20323 & w29770) | (w20323 & w29771) | (w29770 & w29771);
assign v6520 = ~(w20509 | w20510);
assign w20511 = v6520;
assign w20512 = w20503 & w20511;
assign w20513 = w20366 & ~w20372;
assign v6521 = ~(w20373 | w20513);
assign w20514 = v6521;
assign w20515 = w5113 & w20040;
assign w20516 = w5531 & ~w20038;
assign v6522 = ~(w20515 | w20516);
assign w20517 = v6522;
assign w20518 = (w20517 & w20063) | (w20517 & w29772) | (w20063 & w29772);
assign w20519 = (~w20339 & w29773) | (~w20339 & w29774) | (w29773 & w29774);
assign w20520 = (w20339 & w29775) | (w20339 & w29776) | (w29775 & w29776);
assign v6523 = ~(w20519 | w20520);
assign w20521 = v6523;
assign w20522 = w20514 & w20521;
assign w20523 = w20359 & ~w20364;
assign v6524 = ~(w20365 | w20523);
assign w20524 = v6524;
assign w20525 = w5610 & ~w20038;
assign w20526 = w5113 & w20043;
assign w20527 = (~w20526 & ~w20040) | (~w20526 & w30530) | (~w20040 & w30530);
assign w20528 = ~w20525 & w20527;
assign w20529 = (~w20294 & w29777) | (~w20294 & w29778) | (w29777 & w29778);
assign w20530 = (w20294 & w29779) | (w20294 & w29780) | (w29779 & w29780);
assign v6525 = ~(w20529 | w20530);
assign w20531 = v6525;
assign w20532 = w20524 & w20531;
assign w20533 = w912 & w20047;
assign w20534 = pi20 & w20533;
assign w20535 = w5114 & w20246;
assign w20536 = w5531 & w20047;
assign w20537 = w5610 & ~w20052;
assign v6526 = ~(w20536 | w20537);
assign w20538 = v6526;
assign w20539 = ~w20535 & w20538;
assign w20540 = ~w20534 & w20539;
assign w20541 = w5113 & w20047;
assign w20542 = (~w20541 & ~w20257) | (~w20541 & w30402) | (~w20257 & w30402);
assign w20543 = w5610 & w20043;
assign w20544 = w5531 & ~w20052;
assign v6527 = ~(w20543 | w20544);
assign w20545 = v6527;
assign w20546 = w20542 & w20545;
assign w20547 = w20542 & w30531;
assign w20548 = w20540 & w20547;
assign w20549 = w20358 & w20548;
assign v6528 = ~(w20358 | w20548);
assign w20550 = v6528;
assign v6529 = ~(w20549 | w20550);
assign w20551 = v6529;
assign w20552 = w5610 & w20040;
assign w20553 = w5113 & ~w20052;
assign w20554 = w5531 & w20043;
assign v6530 = ~(w20553 | w20554);
assign w20555 = v6530;
assign w20556 = ~w20552 & w20555;
assign w20557 = (w20272 & w30403) | (w20272 & w30404) | (w30403 & w30404);
assign w20558 = (~w20272 & w30405) | (~w20272 & w30406) | (w30405 & w30406);
assign v6531 = ~(w20557 | w20558);
assign w20559 = v6531;
assign w20560 = w20551 & w20559;
assign w20561 = (~w20549 & ~w20559) | (~w20549 & w30532) | (~w20559 & w30532);
assign v6532 = ~(w20524 | w20531);
assign w20562 = v6532;
assign v6533 = ~(w20532 | w20562);
assign w20563 = v6533;
assign w20564 = ~w20561 & w20563;
assign w20565 = (~w20532 & ~w20563) | (~w20532 & w30236) | (~w20563 & w30236);
assign v6534 = ~(w20514 | w20521);
assign w20566 = v6534;
assign v6535 = ~(w20522 | w20566);
assign w20567 = v6535;
assign w20568 = ~w20565 & w20567;
assign w20569 = (~w20522 & ~w20567) | (~w20522 & w30237) | (~w20567 & w30237);
assign v6536 = ~(w20503 | w20511);
assign w20570 = v6536;
assign v6537 = ~(w20512 | w20570);
assign w20571 = v6537;
assign w20572 = ~w20569 & w20571;
assign w20573 = (~w20512 & ~w20571) | (~w20512 & w30238) | (~w20571 & w30238);
assign v6538 = ~(w20493 | w20500);
assign w20574 = v6538;
assign v6539 = ~(w20501 | w20574);
assign w20575 = v6539;
assign w20576 = ~w20573 & w20575;
assign w20577 = (~w20501 & ~w20575) | (~w20501 & w30239) | (~w20575 & w30239);
assign v6540 = ~(w20482 | w20490);
assign w20578 = v6540;
assign v6541 = ~(w20491 | w20578);
assign w20579 = v6541;
assign w20580 = ~w20577 & w20579;
assign w20581 = (~w20491 & w20577) | (~w20491 & w31066) | (w20577 & w31066);
assign w20582 = ~w20470 & w20479;
assign v6542 = ~(w20480 | w20582);
assign w20583 = v6542;
assign w20584 = ~w20581 & w20583;
assign w20585 = (~w20480 & w20581) | (~w20480 & w30667) | (w20581 & w30667);
assign v6543 = ~(w20457 | w20467);
assign w20586 = v6543;
assign v6544 = ~(w20468 | w20586);
assign w20587 = v6544;
assign w20588 = ~w20585 & w20587;
assign w20589 = (~w20468 & w20585) | (~w20468 & w30856) | (w20585 & w30856);
assign w20590 = ~w20444 & w20454;
assign v6545 = ~(w20455 | w20590);
assign w20591 = v6545;
assign w20592 = ~w20589 & w20591;
assign w20593 = (~w20455 & w20589) | (~w20455 & w30407) | (w20589 & w30407);
assign w20594 = (~w20439 & w20402) | (~w20439 & w31067) | (w20402 & w31067);
assign v6546 = ~(w20422 | w20426);
assign w20595 = v6546;
assign w20596 = ~w3405 & w20047;
assign w20597 = w20410 & w31203;
assign w20598 = w20596 & w20597;
assign v6547 = ~(w20596 | w20597);
assign w20599 = v6547;
assign v6548 = ~(w20598 | w20599);
assign w20600 = v6548;
assign w20601 = w3763 & w20043;
assign w20602 = w3760 & w20040;
assign w20603 = w3767 & ~w20052;
assign v6549 = ~(w20602 | w20603);
assign w20604 = v6549;
assign w20605 = (w20272 & w31068) | (w20272 & w31069) | (w31068 & w31069);
assign w20606 = (~w20272 & w31070) | (~w20272 & w31071) | (w31070 & w31071);
assign v6550 = ~(w20605 | w20606);
assign w20607 = v6550;
assign w20608 = w20600 & ~w20607;
assign w20609 = ~w20600 & w20607;
assign v6551 = ~(w20608 | w20609);
assign w20610 = v6551;
assign w20611 = w4155 & w20031;
assign v6552 = ~(w2873 | w20038);
assign w20612 = v6552;
assign w20613 = w4158 & ~w20063;
assign v6553 = ~(w20612 | w20613);
assign w20614 = v6553;
assign w20615 = ~w20611 & w20614;
assign w20616 = (~w20323 & w30858) | (~w20323 & w30859) | (w30858 & w30859);
assign w20617 = (w20323 & w30860) | (w20323 & w30861) | (w30860 & w30861);
assign v6554 = ~(w20616 | w20617);
assign w20618 = v6554;
assign v6555 = ~(w20610 | w20618);
assign w20619 = v6555;
assign w20620 = w20610 & w20618;
assign v6556 = ~(w20619 | w20620);
assign w20621 = v6556;
assign w20622 = ~w20595 & w20621;
assign w20623 = w20595 & ~w20621;
assign v6557 = ~(w20622 | w20623);
assign w20624 = v6557;
assign w20625 = w4836 & ~w20028;
assign w20626 = w4913 & w20014;
assign v6558 = ~(w20625 | w20626);
assign w20627 = v6558;
assign w20628 = w4763 & ~w20026;
assign w20629 = (~w20472 & w30533) | (~w20472 & w30534) | (w30533 & w30534);
assign w20630 = (w20472 & w30535) | (w20472 & w30536) | (w30535 & w30536);
assign v6559 = ~(w20629 | w20630);
assign w20631 = v6559;
assign w20632 = ~w20624 & w20631;
assign w20633 = w20624 & ~w20631;
assign v6560 = ~(w20632 | w20633);
assign w20634 = v6560;
assign w20635 = ~w20594 & w20634;
assign w20636 = w20594 & ~w20634;
assign v6561 = ~(w20635 | w20636);
assign w20637 = v6561;
assign w20638 = (w20079 & w29049) | (w20079 & w29050) | (w29049 & w29050);
assign v6562 = ~(w20086 | w20638);
assign w20639 = v6562;
assign w20640 = w5610 & w20005;
assign w20641 = w5113 & ~w20011;
assign w20642 = w5531 & ~w20008;
assign v6563 = ~(w20641 | w20642);
assign w20643 = v6563;
assign w20644 = ~w20640 & w20643;
assign w20645 = (~w20639 & w30537) | (~w20639 & w30538) | (w30537 & w30538);
assign w20646 = (w20639 & w30539) | (w20639 & w30540) | (w30539 & w30540);
assign v6564 = ~(w20645 | w20646);
assign w20647 = v6564;
assign v6565 = ~(w20637 | w20647);
assign w20648 = v6565;
assign w20649 = w20637 & w20647;
assign v6566 = ~(w20648 | w20649);
assign w20650 = v6566;
assign w20651 = ~w20593 & w20650;
assign w20652 = w20593 & ~w20650;
assign v6567 = ~(w20651 | w20652);
assign w20653 = v6567;
assign w20654 = (w28064 & w29544) | (w28064 & w29545) | (w29544 & w29545);
assign v6568 = ~(w20096 | w20654);
assign w20655 = v6568;
assign w20656 = w5983 & ~w19997;
assign w20657 = w6236 & ~w19992;
assign v6569 = ~(w20656 | w20657);
assign w20658 = v6569;
assign w20659 = w5764 & w20000;
assign w20660 = w20658 & ~w20659;
assign w20661 = (~w20655 & w30541) | (~w20655 & w30542) | (w30541 & w30542);
assign w20662 = (w20655 & w30543) | (w20655 & w30544) | (w30543 & w30544);
assign v6570 = ~(w20661 | w20662);
assign w20663 = v6570;
assign w20664 = w20653 & ~w20663;
assign w20665 = w20589 & ~w20591;
assign v6571 = ~(w20592 | w20665);
assign w20666 = v6571;
assign w20667 = ~w20003 & w20091;
assign v6572 = ~(w20092 | w20667);
assign w20668 = v6572;
assign w20669 = w6236 & ~w19997;
assign w20670 = w5764 & w20005;
assign w20671 = w5983 & w20000;
assign v6573 = ~(w20670 | w20671);
assign w20672 = v6573;
assign w20673 = ~w20669 & w20672;
assign w20674 = (~w20668 & w30411) | (~w20668 & w30412) | (w30411 & w30412);
assign w20675 = (w20668 & w30413) | (w20668 & w30414) | (w30413 & w30414);
assign v6574 = ~(w20674 | w20675);
assign w20676 = v6574;
assign w20677 = w20666 & w20676;
assign w20678 = w20585 & ~w20587;
assign v6575 = ~(w20588 | w20678);
assign w20679 = v6575;
assign w20680 = w20087 & ~w20089;
assign v6576 = ~(w20090 | w20680);
assign w20681 = v6576;
assign w20682 = w6236 & w20000;
assign w20683 = w5764 & ~w20008;
assign w20684 = w5983 & w20005;
assign v6577 = ~(w20683 | w20684);
assign w20685 = v6577;
assign w20686 = ~w20682 & w20685;
assign w20687 = (~w20681 & w30415) | (~w20681 & w30416) | (w30415 & w30416);
assign w20688 = (w20681 & w30417) | (w20681 & w30418) | (w30417 & w30418);
assign v6578 = ~(w20687 | w20688);
assign w20689 = v6578;
assign w20690 = w20679 & w20689;
assign w20691 = w20581 & ~w20583;
assign v6579 = ~(w20584 | w20691);
assign w20692 = v6579;
assign w20693 = w6236 & w20005;
assign w20694 = w5764 & ~w20011;
assign w20695 = w5983 & ~w20008;
assign v6580 = ~(w20694 | w20695);
assign w20696 = v6580;
assign w20697 = ~w20693 & w20696;
assign w20698 = (~w29546 & w30242) | (~w29546 & w30243) | (w30242 & w30243);
assign w20699 = (w29546 & w30244) | (w29546 & w30245) | (w30244 & w30245);
assign v6581 = ~(w20698 | w20699);
assign w20700 = v6581;
assign w20701 = w20692 & w20700;
assign w20702 = w20577 & ~w20579;
assign v6582 = ~(w20580 | w20702);
assign w20703 = v6582;
assign w20704 = w6236 & ~w20008;
assign w20705 = w5983 & ~w20011;
assign w20706 = w5764 & w20014;
assign v6583 = ~(w20705 | w20706);
assign w20707 = v6583;
assign w20708 = ~w20704 & w20707;
assign w20709 = (w29547 & ~w29323) | (w29547 & w29910) | (~w29323 & w29910);
assign w20710 = (w29323 & w29911) | (w29323 & w29912) | (w29911 & w29912);
assign v6584 = ~(w20709 | w20710);
assign w20711 = v6584;
assign w20712 = w20703 & w20711;
assign w20713 = w20573 & ~w20575;
assign v6585 = ~(w20576 | w20713);
assign w20714 = v6585;
assign w20715 = w6236 & ~w20011;
assign w20716 = w5983 & w20014;
assign w20717 = w5764 & ~w20028;
assign v6586 = ~(w20716 | w20717);
assign w20718 = v6586;
assign w20719 = ~w20715 & w20718;
assign w20720 = (~w20459 & w29549) | (~w20459 & w29550) | (w29549 & w29550);
assign w20721 = (w20459 & w29551) | (w20459 & w29552) | (w29551 & w29552);
assign v6587 = ~(w20720 | w20721);
assign w20722 = v6587;
assign w20723 = w20714 & w20722;
assign w20724 = w20569 & ~w20571;
assign v6588 = ~(w20572 | w20724);
assign w20725 = v6588;
assign w20726 = w5765 & w20472;
assign w20727 = w5983 & ~w20028;
assign w20728 = (~w20727 & ~w20014) | (~w20727 & w29553) | (~w20014 & w29553);
assign w20729 = w5764 & ~w20026;
assign w20730 = w20728 & ~w20729;
assign w20731 = ~w20726 & w29324;
assign w20732 = (~pi17 & w20726) | (~pi17 & w29325) | (w20726 & w29325);
assign v6589 = ~(w20731 | w20732);
assign w20733 = v6589;
assign w20734 = w20725 & ~w20733;
assign w20735 = w20565 & ~w20567;
assign v6590 = ~(w20568 | w20735);
assign w20736 = v6590;
assign w20737 = w6236 & ~w20028;
assign w20738 = w5764 & w20031;
assign w20739 = (~w20738 & w20026) | (~w20738 & w29554) | (w20026 & w29554);
assign w20740 = ~w20737 & w20739;
assign w20741 = (w20431 & w29326) | (w20431 & w29327) | (w29326 & w29327);
assign w20742 = (~w20431 & w29328) | (~w20431 & w29329) | (w29328 & w29329);
assign v6591 = ~(w20741 | w20742);
assign w20743 = v6591;
assign w20744 = w20736 & w20743;
assign w20745 = w20561 & ~w20563;
assign v6592 = ~(w20564 | w20745);
assign w20746 = v6592;
assign w20747 = w5764 & ~w20063;
assign w20748 = w5983 & w20031;
assign v6593 = ~(w20747 | w20748);
assign w20749 = v6593;
assign w20750 = (w20749 & w20026) | (w20749 & w29330) | (w20026 & w29330);
assign w20751 = (~w20309 & w30668) | (~w20309 & w30669) | (w30668 & w30669);
assign w20752 = (w20309 & w30670) | (w20309 & w30671) | (w30670 & w30671);
assign v6594 = ~(w20751 | w20752);
assign w20753 = v6594;
assign w20754 = w20746 & ~w20753;
assign v6595 = ~(w20551 | w20559);
assign w20755 = v6595;
assign v6596 = ~(w20560 | w20755);
assign w20756 = v6596;
assign w20757 = w6236 & w20031;
assign w20758 = w5764 & ~w20038;
assign w20759 = (~w20758 & w20063) | (~w20758 & w29555) | (w20063 & w29555);
assign w20760 = ~w20757 & w20759;
assign w20761 = (w20323 & w29335) | (w20323 & w29336) | (w29335 & w29336);
assign w20762 = (~w20323 & w29337) | (~w20323 & w29338) | (w29337 & w29338);
assign v6597 = ~(w20761 | w20762);
assign w20763 = v6597;
assign w20764 = w20756 & w20763;
assign w20765 = pi20 & ~w20540;
assign v6598 = ~(w20546 | w20765);
assign w20766 = v6598;
assign w20767 = w20546 & w20765;
assign v6599 = ~(w20766 | w20767);
assign w20768 = v6599;
assign w20769 = w5764 & w20040;
assign w20770 = (~w20769 & w20038) | (~w20769 & w29556) | (w20038 & w29556);
assign w20771 = (w20770 & w20063) | (w20770 & w29339) | (w20063 & w29339);
assign w20772 = (~w20339 & w29340) | (~w20339 & w29341) | (w29340 & w29341);
assign w20773 = (w20339 & w29342) | (w20339 & w29343) | (w29342 & w29343);
assign v6600 = ~(w20772 | w20773);
assign w20774 = v6600;
assign w20775 = ~w20768 & w20774;
assign w20776 = w20534 & ~w20539;
assign v6601 = ~(w20540 | w20776);
assign w20777 = v6601;
assign w20778 = w6236 & ~w20038;
assign w20779 = w5764 & w20043;
assign w20780 = (~w20779 & ~w20040) | (~w20779 & w30545) | (~w20040 & w30545);
assign w20781 = ~w20778 & w20780;
assign w20782 = (w20294 & w29344) | (w20294 & w29345) | (w29344 & w29345);
assign w20783 = (~w20294 & w29346) | (~w20294 & w29347) | (w29346 & w29347);
assign v6602 = ~(w20782 | w20783);
assign w20784 = v6602;
assign w20785 = w20777 & w20784;
assign w20786 = w5756 & w20047;
assign w20787 = pi17 & w20786;
assign w20788 = w5765 & w20246;
assign w20789 = w6236 & ~w20052;
assign w20790 = w5983 & w20047;
assign v6603 = ~(w20789 | w20790);
assign w20791 = v6603;
assign w20792 = ~w20788 & w20791;
assign w20793 = ~w20787 & w20792;
assign w20794 = w5764 & w20047;
assign w20795 = (~w20794 & ~w20257) | (~w20794 & w29781) | (~w20257 & w29781);
assign w20796 = w6236 & w20043;
assign w20797 = w5983 & ~w20052;
assign v6604 = ~(w20796 | w20797);
assign w20798 = v6604;
assign w20799 = w20795 & w20798;
assign w20800 = w20795 & w30546;
assign w20801 = w20793 & w20800;
assign w20802 = w20533 & w20801;
assign v6605 = ~(w20533 | w20801);
assign w20803 = v6605;
assign v6606 = ~(w20802 | w20803);
assign w20804 = v6606;
assign w20805 = w6236 & w20040;
assign w20806 = w5764 & ~w20052;
assign w20807 = w5983 & w20043;
assign v6607 = ~(w20806 | w20807);
assign w20808 = v6607;
assign w20809 = ~w20805 & w20808;
assign w20810 = (~w20272 & w29782) | (~w20272 & w29783) | (w29782 & w29783);
assign w20811 = (w20272 & w29784) | (w20272 & w29785) | (w29784 & w29785);
assign v6608 = ~(w20810 | w20811);
assign w20812 = v6608;
assign w20813 = w20804 & w20812;
assign w20814 = (~w20802 & ~w20812) | (~w20802 & w30547) | (~w20812 & w30547);
assign v6609 = ~(w20777 | w20784);
assign w20815 = v6609;
assign v6610 = ~(w20785 | w20815);
assign w20816 = v6610;
assign w20817 = ~w20814 & w20816;
assign w20818 = (~w20785 & ~w20816) | (~w20785 & w29558) | (~w20816 & w29558);
assign w20819 = w20768 & ~w20774;
assign v6611 = ~(w20775 | w20819);
assign w20820 = v6611;
assign w20821 = ~w20818 & w20820;
assign w20822 = (~w20775 & ~w20820) | (~w20775 & w29559) | (~w20820 & w29559);
assign v6612 = ~(w20756 | w20763);
assign w20823 = v6612;
assign v6613 = ~(w20764 | w20823);
assign w20824 = v6613;
assign w20825 = ~w20822 & w20824;
assign w20826 = (~w20764 & ~w20824) | (~w20764 & w29560) | (~w20824 & w29560);
assign w20827 = ~w20746 & w20753;
assign v6614 = ~(w20754 | w20827);
assign w20828 = v6614;
assign w20829 = ~w20826 & w20828;
assign w20830 = (~w20754 & ~w20828) | (~w20754 & w29561) | (~w20828 & w29561);
assign v6615 = ~(w20736 | w20743);
assign w20831 = v6615;
assign v6616 = ~(w20744 | w20831);
assign w20832 = v6616;
assign w20833 = ~w20830 & w20832;
assign w20834 = (~w20744 & w20830) | (~w20744 & w31072) | (w20830 & w31072);
assign w20835 = ~w20725 & w20733;
assign v6617 = ~(w20734 | w20835);
assign w20836 = v6617;
assign w20837 = ~w20834 & w20836;
assign w20838 = (~w20734 & ~w20836) | (~w20734 & w29562) | (~w20836 & w29562);
assign v6618 = ~(w20714 | w20722);
assign w20839 = v6618;
assign v6619 = ~(w20723 | w20839);
assign w20840 = v6619;
assign w20841 = (~w29562 & w30672) | (~w29562 & w30673) | (w30672 & w30673);
assign w20842 = (~w20723 & w20838) | (~w20723 & w29786) | (w20838 & w29786);
assign v6620 = ~(w20703 | w20711);
assign w20843 = v6620;
assign v6621 = ~(w20712 | w20843);
assign w20844 = v6621;
assign w20845 = ~w20842 & w20844;
assign w20846 = (~w20712 & w20842) | (~w20712 & w30674) | (w20842 & w30674);
assign v6622 = ~(w20692 | w20700);
assign w20847 = v6622;
assign v6623 = ~(w20701 | w20847);
assign w20848 = v6623;
assign w20849 = ~w20846 & w20848;
assign w20850 = (~w20701 & w20846) | (~w20701 & w30246) | (w20846 & w30246);
assign v6624 = ~(w20679 | w20689);
assign w20851 = v6624;
assign v6625 = ~(w20690 | w20851);
assign w20852 = v6625;
assign w20853 = ~w20850 & w20852;
assign w20854 = (~w20690 & w20850) | (~w20690 & w30675) | (w20850 & w30675);
assign v6626 = ~(w20666 | w20676);
assign w20855 = v6626;
assign v6627 = ~(w20677 | w20855);
assign w20856 = v6627;
assign w20857 = ~w20854 & w20856;
assign w20858 = (~w20677 & w20854) | (~w20677 & w30862) | (w20854 & w30862);
assign w20859 = ~w20653 & w20663;
assign v6628 = ~(w20664 | w20859);
assign w20860 = v6628;
assign w20861 = ~w20858 & w20860;
assign w20862 = (~w20664 & w20858) | (~w20664 & w30419) | (w20858 & w30419);
assign w20863 = (~w20649 & w20593) | (~w20649 & w31073) | (w20593 & w31073);
assign w20864 = (~w20633 & w20594) | (~w20633 & w30548) | (w20594 & w30548);
assign v6629 = ~(w20620 | w20622);
assign w20865 = v6629;
assign w20866 = (~w20598 & w20607) | (~w20598 & w31204) | (w20607 & w31204);
assign w20867 = w3278 & w4071;
assign w20868 = w4452 & w20867;
assign w20869 = ~w215 & w20868;
assign w20870 = ~w63 & w526;
assign w20871 = w580 & w1154;
assign w20872 = w1559 & w20871;
assign w20873 = w20870 & w20872;
assign w20874 = w1600 & w6710;
assign w20875 = w1041 & w12959;
assign w20876 = w20874 & w20875;
assign w20877 = w20873 & w20876;
assign w20878 = w20869 & w20877;
assign w20879 = ~w666 & w2750;
assign w20880 = w2455 & w6665;
assign w20881 = ~w201 & w20880;
assign w20882 = w20879 & w20881;
assign w20883 = w1574 & w5375;
assign w20884 = w1546 & w4987;
assign w20885 = w1370 & w1840;
assign w20886 = w20884 & w20885;
assign w20887 = ~w77 & w2256;
assign w20888 = ~w425 & w20887;
assign w20889 = w20886 & w20888;
assign w20890 = w20883 & w20889;
assign w20891 = w20882 & w20890;
assign w20892 = w20878 & w20891;
assign w20893 = ~w388 & w5000;
assign w20894 = w1128 & w20893;
assign w20895 = w442 & w20894;
assign w20896 = w2240 & w20895;
assign w20897 = w1937 & w14539;
assign w20898 = w20896 & w20897;
assign w20899 = w14434 & w20898;
assign w20900 = w20892 & w20899;
assign w20901 = w928 & w20246;
assign w20902 = w3406 & ~w20052;
assign w20903 = w3402 & w20047;
assign v6630 = ~(w20902 | w20903);
assign w20904 = v6630;
assign w20905 = ~w20901 & w20904;
assign v6631 = ~(w20900 | w20905);
assign w20906 = v6631;
assign w20907 = w20900 & w20905;
assign v6632 = ~(w20906 | w20907);
assign w20908 = v6632;
assign w20909 = w3760 & ~w20038;
assign w20910 = w3763 & w20040;
assign w20911 = w3767 & w20043;
assign v6633 = ~(w20910 | w20911);
assign w20912 = v6633;
assign w20913 = ~w20909 & w20912;
assign w20914 = (w20294 & w30863) | (w20294 & w30864) | (w30863 & w30864);
assign w20915 = (~w20294 & w30865) | (~w20294 & w30866) | (w30865 & w30866);
assign v6634 = ~(w20914 | w20915);
assign w20916 = v6634;
assign w20917 = w20908 & ~w20916;
assign w20918 = ~w20908 & w20916;
assign v6635 = ~(w20917 | w20918);
assign w20919 = v6635;
assign w20920 = ~w20866 & w20919;
assign w20921 = w20866 & ~w20919;
assign v6636 = ~(w20920 | w20921);
assign w20922 = v6636;
assign w20923 = (w4153 & w20309) | (w4153 & w30676) | (w20309 & w30676);
assign v6637 = ~(w2873 | w20063);
assign w20924 = v6637;
assign w20925 = w4155 & ~w20026;
assign w20926 = w4158 & w20031;
assign w20927 = ~w20923 & w30549;
assign w20928 = (~pi26 & w20923) | (~pi26 & w30550) | (w20923 & w30550);
assign v6638 = ~(w20927 | w20928);
assign w20929 = v6638;
assign w20930 = w20922 & ~w20929;
assign w20931 = ~w20922 & w20929;
assign v6639 = ~(w20930 | w20931);
assign w20932 = v6639;
assign w20933 = ~w20865 & w20932;
assign w20934 = w20865 & ~w20932;
assign v6640 = ~(w20933 | w20934);
assign w20935 = v6640;
assign w20936 = w4913 & ~w20011;
assign w20937 = w4836 & w20014;
assign w20938 = w4763 & ~w20028;
assign v6641 = ~(w20937 | w20938);
assign w20939 = v6641;
assign w20940 = ~w20936 & w20939;
assign w20941 = (~w20459 & w30867) | (~w20459 & w30868) | (w30867 & w30868);
assign w20942 = (w20459 & w30869) | (w20459 & w30870) | (w30869 & w30870);
assign v6642 = ~(w20941 | w20942);
assign w20943 = v6642;
assign v6643 = ~(w20935 | w20943);
assign w20944 = v6643;
assign w20945 = w20935 & w20943;
assign v6644 = ~(w20944 | w20945);
assign w20946 = v6644;
assign w20947 = ~w20864 & w20946;
assign w20948 = w20864 & ~w20946;
assign v6645 = ~(w20947 | w20948);
assign w20949 = v6645;
assign w20950 = w5610 & w20000;
assign w20951 = w5113 & ~w20008;
assign w20952 = w5531 & w20005;
assign v6646 = ~(w20951 | w20952);
assign w20953 = v6646;
assign w20954 = ~w20950 & w20953;
assign w20955 = (~w20681 & w30871) | (~w20681 & w30872) | (w30871 & w30872);
assign w20956 = (w20681 & w30873) | (w20681 & w30874) | (w30873 & w30874);
assign v6647 = ~(w20955 | w20956);
assign w20957 = v6647;
assign w20958 = w20949 & w20957;
assign v6648 = ~(w20949 | w20957);
assign w20959 = v6648;
assign v6649 = ~(w20958 | w20959);
assign w20960 = v6649;
assign w20961 = ~w20863 & w20960;
assign w20962 = w20863 & ~w20960;
assign v6650 = ~(w20961 | w20962);
assign w20963 = v6650;
assign w20964 = (w20093 & w29787) | (w20093 & w29788) | (w29787 & w29788);
assign v6651 = ~(w20098 | w20964);
assign w20965 = v6651;
assign w20966 = w5983 & ~w19992;
assign w20967 = w6236 & w19989;
assign v6652 = ~(w20966 | w20967);
assign w20968 = v6652;
assign w20969 = w5764 & ~w19997;
assign w20970 = w20968 & ~w20969;
assign w20971 = (w20970 & ~w20965) | (w20970 & w30552) | (~w20965 & w30552);
assign w20972 = pi17 & w20971;
assign v6653 = ~(pi17 | w20971);
assign w20973 = v6653;
assign v6654 = ~(w20972 | w20973);
assign w20974 = v6654;
assign w20975 = w20963 & ~w20974;
assign w20976 = ~w20963 & w20974;
assign v6655 = ~(w20975 | w20976);
assign w20977 = v6655;
assign w20978 = ~w20862 & w20977;
assign w20979 = w20862 & ~w20977;
assign v6656 = ~(w20978 | w20979);
assign w20980 = v6656;
assign w20981 = w20106 & ~w20108;
assign v6657 = ~(w20109 | w20981);
assign w20982 = v6657;
assign w20983 = w6389 & w20982;
assign w20984 = w6871 & w19983;
assign w20985 = w7004 & w19980;
assign v6658 = ~(w20984 | w20985);
assign w20986 = v6658;
assign w20987 = w6388 & w19986;
assign w20988 = w20986 & ~w20987;
assign w20989 = ~w20983 & w20988;
assign w20990 = pi14 & w20989;
assign v6659 = ~(pi14 | w20989);
assign w20991 = v6659;
assign v6660 = ~(w20990 | w20991);
assign w20992 = v6660;
assign w20993 = w20980 & ~w20992;
assign w20994 = w20858 & ~w20860;
assign v6661 = ~(w20861 | w20994);
assign w20995 = v6661;
assign w20996 = (w20099 & w30247) | (w20099 & w30248) | (w30247 & w30248);
assign v6662 = ~(w20105 | w20996);
assign w20997 = v6662;
assign w20998 = w6389 & w20997;
assign w20999 = w7004 & w19983;
assign w21000 = w6388 & w19989;
assign w21001 = w6871 & w19986;
assign v6663 = ~(w21000 | w21001);
assign w21002 = v6663;
assign w21003 = ~w20999 & w21002;
assign w21004 = ~w20998 & w21003;
assign w21005 = ~pi14 & w21004;
assign w21006 = pi14 & ~w21004;
assign v6664 = ~(w21005 | w21006);
assign w21007 = v6664;
assign w21008 = w20995 & w21007;
assign w21009 = w20854 & ~w20856;
assign v6665 = ~(w20857 | w21009);
assign w21010 = v6665;
assign w21011 = (w20097 & w30249) | (w20097 & w30250) | (w30249 & w30250);
assign v6666 = ~(w20102 | w21011);
assign w21012 = v6666;
assign w21013 = w6389 & w21012;
assign w21014 = w7004 & w19986;
assign w21015 = w6388 & ~w19992;
assign w21016 = w6871 & w19989;
assign v6667 = ~(w21015 | w21016);
assign w21017 = v6667;
assign w21018 = ~w21014 & w21017;
assign w21019 = ~w21013 & w21018;
assign w21020 = ~pi14 & w21019;
assign w21021 = pi14 & ~w21019;
assign v6668 = ~(w21020 | w21021);
assign w21022 = v6668;
assign w21023 = w21010 & w21022;
assign w21024 = w20850 & ~w20852;
assign v6669 = ~(w20853 | w21024);
assign w21025 = v6669;
assign w21026 = w7004 & w19989;
assign w21027 = w6388 & ~w19997;
assign w21028 = w6871 & ~w19992;
assign v6670 = ~(w21027 | w21028);
assign w21029 = v6670;
assign w21030 = ~w21026 & w21029;
assign w21031 = (w21030 & ~w20965) | (w21030 & w30553) | (~w20965 & w30553);
assign w21032 = ~pi14 & w21031;
assign w21033 = pi14 & ~w21031;
assign v6671 = ~(w21032 | w21033);
assign w21034 = v6671;
assign w21035 = w21025 & w21034;
assign w21036 = w20846 & ~w20848;
assign v6672 = ~(w20849 | w21036);
assign w21037 = v6672;
assign w21038 = w7004 & ~w19992;
assign w21039 = w6871 & ~w19997;
assign w21040 = w6388 & w20000;
assign v6673 = ~(w21039 | w21040);
assign w21041 = v6673;
assign w21042 = ~w21038 & w21041;
assign w21043 = (~w20655 & w30554) | (~w20655 & w30555) | (w30554 & w30555);
assign w21044 = (w20655 & w30556) | (w20655 & w30557) | (w30556 & w30557);
assign v6674 = ~(w21043 | w21044);
assign w21045 = v6674;
assign w21046 = w21037 & w21045;
assign w21047 = w20842 & ~w20844;
assign v6675 = ~(w20845 | w21047);
assign w21048 = v6675;
assign w21049 = w6388 & w20005;
assign w21050 = w7004 & ~w19997;
assign v6676 = ~(w21049 | w21050);
assign w21051 = v6676;
assign w21052 = w6871 & w20000;
assign w21053 = w21051 & ~w21052;
assign w21054 = (~w20668 & w30421) | (~w20668 & w30422) | (w30421 & w30422);
assign w21055 = (w20668 & w30423) | (w20668 & w30424) | (w30423 & w30424);
assign v6677 = ~(w21054 | w21055);
assign w21056 = v6677;
assign w21057 = w21048 & ~w21056;
assign w21058 = (w29562 & w30677) | (w29562 & w30678) | (w30677 & w30678);
assign v6678 = ~(w20841 | w21058);
assign w21059 = v6678;
assign w21060 = w7004 & w20000;
assign w21061 = w6388 & ~w20008;
assign w21062 = w6871 & w20005;
assign v6679 = ~(w21061 | w21062);
assign w21063 = v6679;
assign w21064 = ~w21060 & w21063;
assign w21065 = (~w20681 & w30425) | (~w20681 & w30426) | (w30425 & w30426);
assign w21066 = (w20681 & w30427) | (w20681 & w30428) | (w30427 & w30428);
assign v6680 = ~(w21065 | w21066);
assign w21067 = v6680;
assign w21068 = w21059 & w21067;
assign w21069 = w20834 & ~w20836;
assign v6681 = ~(w20837 | w21069);
assign w21070 = v6681;
assign w21071 = w6871 & ~w20008;
assign w21072 = w7004 & w20005;
assign v6682 = ~(w21071 | w21072);
assign w21073 = v6682;
assign w21074 = w6388 & ~w20011;
assign w21075 = w21073 & ~w21074;
assign w21076 = (~w29563 & w31074) | (~w29563 & w31075) | (w31074 & w31075);
assign w21077 = (w29563 & w31076) | (w29563 & w31077) | (w31076 & w31077);
assign v6683 = ~(w21076 | w21077);
assign w21078 = v6683;
assign w21079 = w21070 & ~w21078;
assign w21080 = w20830 & ~w20832;
assign v6684 = ~(w20833 | w21080);
assign w21081 = v6684;
assign w21082 = w6871 & ~w20011;
assign w21083 = w7004 & ~w20008;
assign v6685 = ~(w21082 | w21083);
assign w21084 = v6685;
assign w21085 = w6388 & w20014;
assign w21086 = (w29564 & ~w29348) | (w29564 & w29913) | (~w29348 & w29913);
assign w21087 = (w29348 & w29914) | (w29348 & w29915) | (w29914 & w29915);
assign v6686 = ~(w21086 | w21087);
assign w21088 = v6686;
assign w21089 = w21081 & ~w21088;
assign w21090 = w20826 & ~w20828;
assign v6687 = ~(w20829 | w21090);
assign w21091 = v6687;
assign w21092 = w6871 & w20014;
assign w21093 = w7004 & ~w20011;
assign w21094 = w6388 & ~w20028;
assign w21095 = ~w21093 & w29566;
assign w21096 = (~w20459 & w29567) | (~w20459 & w29568) | (w29567 & w29568);
assign w21097 = (w20459 & w29569) | (w20459 & w29570) | (w29569 & w29570);
assign v6688 = ~(w21096 | w21097);
assign w21098 = v6688;
assign w21099 = w21091 & ~w21098;
assign w21100 = w20822 & ~w20824;
assign v6689 = ~(w20825 | w21100);
assign w21101 = v6689;
assign w21102 = w6389 & w20472;
assign w21103 = w6871 & ~w20028;
assign w21104 = (~w21103 & ~w20014) | (~w21103 & w29571) | (~w20014 & w29571);
assign w21105 = w6388 & ~w20026;
assign w21106 = w21104 & ~w21105;
assign w21107 = ~w21102 & w29349;
assign w21108 = (~pi14 & w21102) | (~pi14 & w29350) | (w21102 & w29350);
assign v6690 = ~(w21107 | w21108);
assign w21109 = v6690;
assign w21110 = w21101 & ~w21109;
assign w21111 = w20818 & ~w20820;
assign v6691 = ~(w20821 | w21111);
assign w21112 = v6691;
assign w21113 = w7004 & ~w20028;
assign w21114 = w6388 & w20031;
assign w21115 = (~w21114 & w20026) | (~w21114 & w29572) | (w20026 & w29572);
assign w21116 = ~w21113 & w21115;
assign w21117 = (w20431 & w29351) | (w20431 & w29352) | (w29351 & w29352);
assign w21118 = (~w20431 & w29353) | (~w20431 & w29354) | (w29353 & w29354);
assign v6692 = ~(w21117 | w21118);
assign w21119 = v6692;
assign w21120 = w21112 & w21119;
assign w21121 = w20814 & ~w20816;
assign v6693 = ~(w20817 | w21121);
assign w21122 = v6693;
assign w21123 = w6388 & ~w20063;
assign w21124 = (w28203 & w29916) | (w28203 & w29917) | (w29916 & w29917);
assign w21125 = w6871 & w20031;
assign w21126 = (~w20309 & w30679) | (~w20309 & w30680) | (w30679 & w30680);
assign w21127 = (w20309 & w30681) | (w20309 & w30682) | (w30681 & w30682);
assign v6694 = ~(w21126 | w21127);
assign w21128 = v6694;
assign w21129 = w21122 & ~w21128;
assign v6695 = ~(w20804 | w20812);
assign w21130 = v6695;
assign v6696 = ~(w20813 | w21130);
assign w21131 = v6696;
assign w21132 = w7004 & w20031;
assign w21133 = w6388 & ~w20038;
assign w21134 = (~w21133 & w20063) | (~w21133 & w29573) | (w20063 & w29573);
assign w21135 = ~w21132 & w21134;
assign w21136 = (w20323 & w29356) | (w20323 & w29357) | (w29356 & w29357);
assign w21137 = (~w20323 & w29358) | (~w20323 & w29359) | (w29358 & w29359);
assign v6697 = ~(w21136 | w21137);
assign w21138 = v6697;
assign w21139 = w21131 & w21138;
assign w21140 = pi17 & ~w20793;
assign v6698 = ~(w20799 | w21140);
assign w21141 = v6698;
assign w21142 = w20799 & w21140;
assign v6699 = ~(w21141 | w21142);
assign w21143 = v6699;
assign w21144 = w6388 & w20040;
assign w21145 = (~w21144 & w20038) | (~w21144 & w29574) | (w20038 & w29574);
assign w21146 = (w21145 & w20063) | (w21145 & w29360) | (w20063 & w29360);
assign w21147 = (~w20339 & w29361) | (~w20339 & w29362) | (w29361 & w29362);
assign w21148 = (w20339 & w29363) | (w20339 & w29364) | (w29363 & w29364);
assign v6700 = ~(w21147 | w21148);
assign w21149 = v6700;
assign w21150 = ~w21143 & w21149;
assign w21151 = w20787 & ~w20792;
assign v6701 = ~(w20793 | w21151);
assign w21152 = v6701;
assign w21153 = w7004 & ~w20038;
assign w21154 = w6388 & w20043;
assign w21155 = (~w21154 & ~w20040) | (~w21154 & w30558) | (~w20040 & w30558);
assign w21156 = ~w21153 & w21155;
assign w21157 = (~w20294 & w29365) | (~w20294 & w29366) | (w29365 & w29366);
assign w21158 = (w20294 & w29367) | (w20294 & w29368) | (w29367 & w29368);
assign v6702 = ~(w21157 | w21158);
assign w21159 = v6702;
assign w21160 = w21152 & w21159;
assign w21161 = w6383 & w20047;
assign w21162 = pi14 & w21161;
assign w21163 = w6389 & w20246;
assign w21164 = w7004 & ~w20052;
assign w21165 = w6871 & w20047;
assign v6703 = ~(w21164 | w21165);
assign w21166 = v6703;
assign w21167 = ~w21163 & w21166;
assign w21168 = ~w21162 & w21167;
assign w21169 = w6388 & w20047;
assign w21170 = (~w21169 & ~w20257) | (~w21169 & w29918) | (~w20257 & w29918);
assign w21171 = w7004 & w20043;
assign w21172 = w6871 & ~w20052;
assign v6704 = ~(w21171 | w21172);
assign w21173 = v6704;
assign w21174 = w21170 & w21173;
assign w21175 = w21170 & w30559;
assign w21176 = w21168 & w21175;
assign w21177 = w20786 & w21176;
assign v6705 = ~(w20786 | w21176);
assign w21178 = v6705;
assign v6706 = ~(w21177 | w21178);
assign w21179 = v6706;
assign w21180 = w7004 & w20040;
assign w21181 = w6388 & ~w20052;
assign w21182 = w6871 & w20043;
assign v6707 = ~(w21181 | w21182);
assign w21183 = v6707;
assign w21184 = ~w21180 & w21183;
assign w21185 = (w20272 & w30253) | (w20272 & w30254) | (w30253 & w30254);
assign w21186 = (~w20272 & w30255) | (~w20272 & w30256) | (w30255 & w30256);
assign v6708 = ~(w21185 | w21186);
assign w21187 = v6708;
assign w21188 = w21179 & w21187;
assign w21189 = (~w21177 & ~w21187) | (~w21177 & w30560) | (~w21187 & w30560);
assign v6709 = ~(w21152 | w21159);
assign w21190 = v6709;
assign v6710 = ~(w21160 | w21190);
assign w21191 = v6710;
assign w21192 = ~w21189 & w21191;
assign w21193 = (~w21160 & ~w21191) | (~w21160 & w29576) | (~w21191 & w29576);
assign w21194 = w21143 & ~w21149;
assign v6711 = ~(w21150 | w21194);
assign w21195 = v6711;
assign w21196 = ~w21193 & w21195;
assign w21197 = (~w21150 & ~w21195) | (~w21150 & w29577) | (~w21195 & w29577);
assign v6712 = ~(w21131 | w21138);
assign w21198 = v6712;
assign v6713 = ~(w21139 | w21198);
assign w21199 = v6713;
assign w21200 = ~w21197 & w21199;
assign w21201 = (~w21139 & ~w21199) | (~w21139 & w29578) | (~w21199 & w29578);
assign w21202 = ~w21122 & w21128;
assign v6714 = ~(w21129 | w21202);
assign w21203 = v6714;
assign w21204 = ~w21201 & w21203;
assign w21205 = (~w21129 & ~w21203) | (~w21129 & w29369) | (~w21203 & w29369);
assign v6715 = ~(w21112 | w21119);
assign w21206 = v6715;
assign v6716 = ~(w21120 | w21206);
assign w21207 = v6716;
assign w21208 = ~w21205 & w21207;
assign w21209 = (~w21120 & w21205) | (~w21120 & w31078) | (w21205 & w31078);
assign w21210 = ~w21101 & w21109;
assign v6717 = ~(w21110 | w21210);
assign w21211 = v6717;
assign w21212 = ~w21209 & w21211;
assign w21213 = (~w21110 & ~w21211) | (~w21110 & w29919) | (~w21211 & w29919);
assign w21214 = ~w21091 & w21098;
assign v6718 = ~(w21099 | w21214);
assign w21215 = v6718;
assign w21216 = (~w29919 & w30683) | (~w29919 & w30684) | (w30683 & w30684);
assign w21217 = (~w21099 & w21213) | (~w21099 & w29579) | (w21213 & w29579);
assign w21218 = ~w21081 & w21088;
assign v6719 = ~(w21089 | w21218);
assign w21219 = v6719;
assign w21220 = ~w21217 & w21219;
assign w21221 = (~w21089 & w21217) | (~w21089 & w30685) | (w21217 & w30685);
assign w21222 = ~w21070 & w21078;
assign v6720 = ~(w21079 | w21222);
assign w21223 = v6720;
assign w21224 = ~w21221 & w21223;
assign w21225 = (~w21079 & w21221) | (~w21079 & w31079) | (w21221 & w31079);
assign v6721 = ~(w21059 | w21067);
assign w21226 = v6721;
assign v6722 = ~(w21068 | w21226);
assign w21227 = v6722;
assign w21228 = ~w21225 & w21227;
assign w21229 = (~w21068 & w21225) | (~w21068 & w30257) | (w21225 & w30257);
assign w21230 = ~w21048 & w21056;
assign v6723 = ~(w21057 | w21230);
assign w21231 = v6723;
assign w21232 = ~w21229 & w21231;
assign w21233 = (~w21057 & w21229) | (~w21057 & w30429) | (w21229 & w30429);
assign v6724 = ~(w21037 | w21045);
assign w21234 = v6724;
assign v6725 = ~(w21046 | w21234);
assign w21235 = v6725;
assign w21236 = ~w21233 & w21235;
assign w21237 = (~w21046 & w21233) | (~w21046 & w30686) | (w21233 & w30686);
assign v6726 = ~(w21025 | w21034);
assign w21238 = v6726;
assign v6727 = ~(w21035 | w21238);
assign w21239 = v6727;
assign w21240 = ~w21237 & w21239;
assign w21241 = (~w21035 & w21237) | (~w21035 & w30561) | (w21237 & w30561);
assign v6728 = ~(w21010 | w21022);
assign w21242 = v6728;
assign v6729 = ~(w21023 | w21242);
assign w21243 = v6729;
assign w21244 = ~w21241 & w21243;
assign w21245 = (~w21023 & w21241) | (~w21023 & w30687) | (w21241 & w30687);
assign v6730 = ~(w20995 | w21007);
assign w21246 = v6730;
assign v6731 = ~(w21008 | w21246);
assign w21247 = v6731;
assign w21248 = ~w21245 & w21247;
assign w21249 = (~w21008 & w21245) | (~w21008 & w30875) | (w21245 & w30875);
assign w21250 = ~w20980 & w20992;
assign v6732 = ~(w20993 | w21250);
assign w21251 = v6732;
assign w21252 = ~w21249 & w21251;
assign v6733 = ~(w20993 | w21252);
assign w21253 = v6733;
assign w21254 = (~w20975 & w20862) | (~w20975 & w31080) | (w20862 & w31080);
assign w21255 = (~w20958 & w20863) | (~w20958 & w30562) | (w20863 & w30562);
assign w21256 = (~w20945 & w20864) | (~w20945 & w30876) | (w20864 & w30876);
assign v6734 = ~(w20930 | w20933);
assign w21257 = v6734;
assign w21258 = (~w20917 & ~w20919) | (~w20917 & w31081) | (~w20919 & w31081);
assign w21259 = w371 & w3431;
assign w21260 = w3205 & w4268;
assign w21261 = w478 & w21260;
assign w21262 = w21259 & w21261;
assign v6735 = ~(w108 | w673);
assign w21263 = v6735;
assign w21264 = w2188 & w21263;
assign w21265 = w675 & w2027;
assign w21266 = w21264 & w21265;
assign w21267 = ~w997 & w2371;
assign v6736 = ~(w221 | w303);
assign w21268 = v6736;
assign w21269 = w2053 & w21268;
assign w21270 = w21267 & w21269;
assign w21271 = w5330 & w21270;
assign w21272 = w21266 & w21271;
assign w21273 = w21262 & w21272;
assign w21274 = w1898 & w6589;
assign w21275 = w14434 & w21274;
assign w21276 = w21273 & w21275;
assign w21277 = ~w20906 & w21276;
assign w21278 = w20906 & ~w21276;
assign v6737 = ~(w21277 | w21278);
assign w21279 = v6737;
assign w21280 = w928 & w20257;
assign w21281 = w3399 & w20047;
assign v6738 = ~(w21280 | w21281);
assign w21282 = v6738;
assign w21283 = w3406 & w20043;
assign w21284 = w3402 & ~w20052;
assign v6739 = ~(w21283 | w21284);
assign w21285 = v6739;
assign w21286 = w21282 & w21285;
assign w21287 = ~w21279 & w21286;
assign w21288 = w21279 & ~w21286;
assign v6740 = ~(w21287 | w21288);
assign w21289 = v6740;
assign w21290 = w3529 & ~w20339;
assign w21291 = w3763 & ~w20038;
assign w21292 = w3760 & ~w20063;
assign v6741 = ~(w21291 | w21292);
assign w21293 = v6741;
assign w21294 = w3767 & w20040;
assign w21295 = (~pi29 & w21290) | (~pi29 & w30877) | (w21290 & w30877);
assign w21296 = ~w21290 & w30878;
assign v6742 = ~(w21295 | w21296);
assign w21297 = v6742;
assign w21298 = w21289 & ~w21297;
assign w21299 = ~w21289 & w21297;
assign v6743 = ~(w21298 | w21299);
assign w21300 = v6743;
assign w21301 = w21258 & ~w21300;
assign w21302 = ~w21258 & w21300;
assign v6744 = ~(w21301 | w21302);
assign w21303 = v6744;
assign w21304 = ~w2873 & w20031;
assign w21305 = w4155 & ~w20028;
assign v6745 = ~(w21304 | w21305);
assign w21306 = v6745;
assign w21307 = w4158 & ~w20026;
assign w21308 = (w20431 & w30879) | (w20431 & w30880) | (w30879 & w30880);
assign w21309 = (~w20431 & w30881) | (~w20431 & w30882) | (w30881 & w30882);
assign v6746 = ~(w21308 | w21309);
assign w21310 = v6746;
assign w21311 = w21303 & ~w21310;
assign w21312 = ~w21303 & w21310;
assign v6747 = ~(w21311 | w21312);
assign w21313 = v6747;
assign w21314 = ~w21257 & w21313;
assign w21315 = w21257 & ~w21313;
assign v6748 = ~(w21314 | w21315);
assign w21316 = v6748;
assign w21317 = w4836 & ~w20011;
assign w21318 = w4913 & ~w20008;
assign v6749 = ~(w21317 | w21318);
assign w21319 = v6749;
assign w21320 = w4763 & w20014;
assign w21321 = w21319 & ~w21320;
assign w21322 = (~w20446 & w30883) | (~w20446 & w30884) | (w30883 & w30884);
assign w21323 = (w20446 & w30885) | (w20446 & w30886) | (w30885 & w30886);
assign v6750 = ~(w21322 | w21323);
assign w21324 = v6750;
assign w21325 = ~w21316 & w21324;
assign w21326 = w21316 & ~w21324;
assign v6751 = ~(w21325 | w21326);
assign w21327 = v6751;
assign w21328 = ~w21256 & w21327;
assign w21329 = w21256 & ~w21327;
assign v6752 = ~(w21328 | w21329);
assign w21330 = v6752;
assign w21331 = w5610 & ~w19997;
assign w21332 = w5113 & w20005;
assign w21333 = w5531 & w20000;
assign v6753 = ~(w21332 | w21333);
assign w21334 = v6753;
assign w21335 = ~w21331 & w21334;
assign w21336 = (~w20668 & w30887) | (~w20668 & w30888) | (w30887 & w30888);
assign w21337 = (w20668 & w30889) | (w20668 & w30890) | (w30889 & w30890);
assign v6754 = ~(w21336 | w21337);
assign w21338 = v6754;
assign w21339 = ~w21330 & w21338;
assign w21340 = w21330 & ~w21338;
assign v6755 = ~(w21339 | w21340);
assign w21341 = v6755;
assign w21342 = ~w21255 & w21341;
assign w21343 = w21255 & ~w21341;
assign v6756 = ~(w21342 | w21343);
assign w21344 = v6756;
assign w21345 = w5765 & w21012;
assign w21346 = w6236 & w19986;
assign w21347 = w5983 & w19989;
assign w21348 = w5764 & ~w19992;
assign v6757 = ~(w21347 | w21348);
assign w21349 = v6757;
assign w21350 = ~w21346 & w21349;
assign w21351 = ~w21345 & w21350;
assign w21352 = ~pi17 & w21351;
assign w21353 = pi17 & ~w21351;
assign v6758 = ~(w21352 | w21353);
assign w21354 = v6758;
assign w21355 = w21344 & w21354;
assign v6759 = ~(w21344 | w21354);
assign w21356 = v6759;
assign v6760 = ~(w21355 | w21356);
assign w21357 = v6760;
assign w21358 = w21254 & ~w21357;
assign w21359 = ~w21254 & w21357;
assign v6761 = ~(w21358 | w21359);
assign w21360 = v6761;
assign w21361 = w20110 & ~w20112;
assign v6762 = ~(w20113 | w21361);
assign w21362 = v6762;
assign w21363 = w6389 & w21362;
assign w21364 = w7004 & w19974;
assign w21365 = w6871 & w19980;
assign w21366 = w6388 & w19983;
assign v6763 = ~(w21365 | w21366);
assign w21367 = v6763;
assign w21368 = ~w21364 & w21367;
assign w21369 = ~w21363 & w21368;
assign w21370 = ~pi14 & w21369;
assign w21371 = pi14 & ~w21369;
assign v6764 = ~(w21370 | w21371);
assign w21372 = v6764;
assign w21373 = w21360 & w21372;
assign v6765 = ~(w21360 | w21372);
assign w21374 = v6765;
assign v6766 = ~(w21373 | w21374);
assign w21375 = v6766;
assign w21376 = ~w21253 & w21375;
assign w21377 = w21253 & ~w21375;
assign v6767 = ~(w21376 | w21377);
assign w21378 = v6767;
assign w21379 = w20240 & w21378;
assign v6768 = ~(w20240 | w21378);
assign w21380 = v6768;
assign v6769 = ~(w21379 | w21380);
assign w21381 = v6769;
assign w21382 = w21249 & ~w21251;
assign v6770 = ~(w21252 | w21382);
assign w21383 = v6770;
assign w21384 = w20118 & ~w20120;
assign v6771 = ~(w20121 | w21384);
assign w21385 = v6771;
assign w21386 = w7178 & w21385;
assign w21387 = w7765 & w19966;
assign w21388 = w7177 & w19974;
assign w21389 = w7466 & ~w19971;
assign v6772 = ~(w21388 | w21389);
assign w21390 = v6772;
assign w21391 = ~w21387 & w21390;
assign w21392 = ~w21386 & w21391;
assign w21393 = ~pi11 & w21392;
assign w21394 = pi11 & ~w21392;
assign v6773 = ~(w21393 | w21394);
assign w21395 = v6773;
assign w21396 = w21383 & w21395;
assign v6774 = ~(w21383 | w21395);
assign w21397 = v6774;
assign w21398 = w21245 & ~w21247;
assign v6775 = ~(w21248 | w21398);
assign w21399 = v6775;
assign w21400 = w20114 & ~w20116;
assign v6776 = ~(w20117 | w21400);
assign w21401 = v6776;
assign w21402 = w7178 & w21401;
assign w21403 = w7765 & ~w19971;
assign w21404 = w7177 & w19980;
assign w21405 = w7466 & w19974;
assign v6777 = ~(w21404 | w21405);
assign w21406 = v6777;
assign w21407 = ~w21403 & w21406;
assign w21408 = ~w21402 & w21407;
assign w21409 = pi11 & w21408;
assign v6778 = ~(pi11 | w21408);
assign w21410 = v6778;
assign v6779 = ~(w21409 | w21410);
assign w21411 = v6779;
assign w21412 = w21399 & ~w21411;
assign w21413 = w21241 & ~w21243;
assign v6780 = ~(w21244 | w21413);
assign w21414 = v6780;
assign w21415 = w7178 & w21362;
assign w21416 = w7466 & w19980;
assign w21417 = w7765 & w19974;
assign v6781 = ~(w21416 | w21417);
assign w21418 = v6781;
assign w21419 = w7177 & w19983;
assign w21420 = w21418 & ~w21419;
assign w21421 = ~w21415 & w21420;
assign w21422 = pi11 & w21421;
assign v6782 = ~(pi11 | w21421);
assign w21423 = v6782;
assign v6783 = ~(w21422 | w21423);
assign w21424 = v6783;
assign w21425 = w21414 & ~w21424;
assign w21426 = w21237 & ~w21239;
assign v6784 = ~(w21240 | w21426);
assign w21427 = v6784;
assign w21428 = w7178 & w20982;
assign w21429 = w7765 & w19980;
assign w21430 = w7466 & w19983;
assign w21431 = w7177 & w19986;
assign v6785 = ~(w21430 | w21431);
assign w21432 = v6785;
assign w21433 = ~w21429 & w21432;
assign w21434 = ~w21428 & w21433;
assign w21435 = ~pi11 & w21434;
assign w21436 = pi11 & ~w21434;
assign v6786 = ~(w21435 | w21436);
assign w21437 = v6786;
assign w21438 = w21427 & w21437;
assign w21439 = w21233 & ~w21235;
assign v6787 = ~(w21236 | w21439);
assign w21440 = v6787;
assign w21441 = w7178 & w20997;
assign w21442 = w7765 & w19983;
assign w21443 = w7177 & w19989;
assign w21444 = w7466 & w19986;
assign v6788 = ~(w21443 | w21444);
assign w21445 = v6788;
assign w21446 = ~w21442 & w21445;
assign w21447 = ~w21441 & w21446;
assign w21448 = ~pi11 & w21447;
assign w21449 = pi11 & ~w21447;
assign v6789 = ~(w21448 | w21449);
assign w21450 = v6789;
assign w21451 = w21440 & w21450;
assign w21452 = w21229 & ~w21231;
assign v6790 = ~(w21232 | w21452);
assign w21453 = v6790;
assign w21454 = w7178 & w21012;
assign w21455 = w7765 & w19986;
assign w21456 = w7177 & ~w19992;
assign w21457 = w7466 & w19989;
assign v6791 = ~(w21456 | w21457);
assign w21458 = v6791;
assign w21459 = ~w21455 & w21458;
assign w21460 = ~w21454 & w21459;
assign w21461 = ~pi11 & w21460;
assign w21462 = pi11 & ~w21460;
assign v6792 = ~(w21461 | w21462);
assign w21463 = v6792;
assign w21464 = w21453 & w21463;
assign w21465 = w21225 & ~w21227;
assign v6793 = ~(w21228 | w21465);
assign w21466 = v6793;
assign w21467 = w7765 & w19989;
assign w21468 = w7177 & ~w19997;
assign w21469 = w7466 & ~w19992;
assign v6794 = ~(w21468 | w21469);
assign w21470 = v6794;
assign w21471 = ~w21467 & w21470;
assign w21472 = (w21471 & ~w20965) | (w21471 & w30430) | (~w20965 & w30430);
assign w21473 = ~pi11 & w21472;
assign w21474 = pi11 & ~w21472;
assign v6795 = ~(w21473 | w21474);
assign w21475 = v6795;
assign w21476 = w21466 & w21475;
assign w21477 = w21221 & ~w21223;
assign v6796 = ~(w21224 | w21477);
assign w21478 = v6796;
assign w21479 = w7466 & ~w19997;
assign w21480 = w7765 & ~w19992;
assign v6797 = ~(w21479 | w21480);
assign w21481 = v6797;
assign w21482 = w7177 & w20000;
assign w21483 = w21481 & ~w21482;
assign w21484 = (~w20655 & w30431) | (~w20655 & w30432) | (w30431 & w30432);
assign w21485 = (w20655 & w30433) | (w20655 & w30434) | (w30433 & w30434);
assign v6798 = ~(w21484 | w21485);
assign w21486 = v6798;
assign w21487 = w21478 & ~w21486;
assign w21488 = w21217 & ~w21219;
assign v6799 = ~(w21220 | w21488);
assign w21489 = v6799;
assign w21490 = w7765 & ~w19997;
assign w21491 = w7177 & w20005;
assign w21492 = w7466 & w20000;
assign v6800 = ~(w21491 | w21492);
assign w21493 = v6800;
assign w21494 = ~w21490 & w21493;
assign w21495 = (~w20668 & w30259) | (~w20668 & w30260) | (w30259 & w30260);
assign w21496 = (w20668 & w30261) | (w20668 & w30262) | (w30261 & w30262);
assign v6801 = ~(w21495 | w21496);
assign w21497 = v6801;
assign w21498 = w21489 & ~w21497;
assign w21499 = (w29919 & w30688) | (w29919 & w30689) | (w30688 & w30689);
assign v6802 = ~(w21216 | w21499);
assign w21500 = v6802;
assign w21501 = w7765 & w20000;
assign w21502 = w7177 & ~w20008;
assign w21503 = w7466 & w20005;
assign v6803 = ~(w21502 | w21503);
assign w21504 = v6803;
assign w21505 = ~w21501 & w21504;
assign w21506 = (~w20681 & w30263) | (~w20681 & w30264) | (w30263 & w30264);
assign w21507 = (w20681 & w30265) | (w20681 & w30266) | (w30265 & w30266);
assign v6804 = ~(w21506 | w21507);
assign w21508 = v6804;
assign w21509 = w21500 & w21508;
assign w21510 = w21209 & ~w21211;
assign v6805 = ~(w21212 | w21510);
assign w21511 = v6805;
assign w21512 = w7466 & ~w20008;
assign w21513 = w7765 & w20005;
assign v6806 = ~(w21512 | w21513);
assign w21514 = v6806;
assign w21515 = w7177 & ~w20011;
assign w21516 = w21514 & ~w21515;
assign w21517 = (~w29580 & w31082) | (~w29580 & w31083) | (w31082 & w31083);
assign w21518 = (w29580 & w31084) | (w29580 & w31085) | (w31084 & w31085);
assign v6807 = ~(w21517 | w21518);
assign w21519 = v6807;
assign w21520 = w21511 & ~w21519;
assign w21521 = w21205 & ~w21207;
assign v6808 = ~(w21208 | w21521);
assign w21522 = v6808;
assign w21523 = w7466 & ~w20011;
assign w21524 = w7765 & ~w20008;
assign v6809 = ~(w21523 | w21524);
assign w21525 = v6809;
assign w21526 = w7177 & w20014;
assign w21527 = (w29581 & ~w29370) | (w29581 & w29920) | (~w29370 & w29920);
assign w21528 = (w29370 & w29921) | (w29370 & w29922) | (w29921 & w29922);
assign v6810 = ~(w21527 | w21528);
assign w21529 = v6810;
assign w21530 = w21522 & ~w21529;
assign w21531 = w21201 & ~w21203;
assign v6811 = ~(w21204 | w21531);
assign w21532 = v6811;
assign w21533 = w7765 & ~w20011;
assign w21534 = w7466 & w20014;
assign w21535 = w7177 & ~w20028;
assign v6812 = ~(w21534 | w21535);
assign w21536 = v6812;
assign w21537 = ~w21533 & w21536;
assign w21538 = (~w20459 & w29583) | (~w20459 & w29584) | (w29583 & w29584);
assign w21539 = (w20459 & w29585) | (w20459 & w29586) | (w29585 & w29586);
assign v6813 = ~(w21538 | w21539);
assign w21540 = v6813;
assign w21541 = w21532 & w21540;
assign w21542 = w21197 & ~w21199;
assign v6814 = ~(w21200 | w21542);
assign w21543 = v6814;
assign w21544 = w7178 & w20472;
assign w21545 = w7466 & ~w20028;
assign w21546 = (~w21545 & ~w20014) | (~w21545 & w29587) | (~w20014 & w29587);
assign w21547 = w7177 & ~w20026;
assign w21548 = w21546 & ~w21547;
assign w21549 = ~w21544 & w29371;
assign w21550 = (~pi11 & w21544) | (~pi11 & w29372) | (w21544 & w29372);
assign v6815 = ~(w21549 | w21550);
assign w21551 = v6815;
assign w21552 = w21543 & ~w21551;
assign w21553 = w21193 & ~w21195;
assign v6816 = ~(w21196 | w21553);
assign w21554 = v6816;
assign w21555 = w7765 & ~w20028;
assign w21556 = w7177 & w20031;
assign w21557 = (~w21556 & w20026) | (~w21556 & w29588) | (w20026 & w29588);
assign w21558 = ~w21555 & w21557;
assign w21559 = (~w20431 & w29373) | (~w20431 & w29374) | (w29373 & w29374);
assign w21560 = (w20431 & w29375) | (w20431 & w29376) | (w29375 & w29376);
assign v6817 = ~(w21559 | w21560);
assign w21561 = v6817;
assign w21562 = w21554 & ~w21561;
assign w21563 = w21189 & ~w21191;
assign v6818 = ~(w21192 | w21563);
assign w21564 = v6818;
assign w21565 = w7177 & ~w20063;
assign w21566 = w7466 & w20031;
assign v6819 = ~(w21565 | w21566);
assign w21567 = v6819;
assign w21568 = (w21567 & w20026) | (w21567 & w29377) | (w20026 & w29377);
assign w21569 = (~w20309 & w30690) | (~w20309 & w30691) | (w30690 & w30691);
assign w21570 = (w20309 & w30692) | (w20309 & w30693) | (w30692 & w30693);
assign v6820 = ~(w21569 | w21570);
assign w21571 = v6820;
assign w21572 = w21564 & w21571;
assign v6821 = ~(w21179 | w21187);
assign w21573 = v6821;
assign v6822 = ~(w21188 | w21573);
assign w21574 = v6822;
assign w21575 = w7466 & ~w20063;
assign w21576 = w7765 & w20031;
assign w21577 = w7177 & ~w20038;
assign w21578 = ~w21576 & w29382;
assign w21579 = (~w20323 & w29383) | (~w20323 & w29384) | (w29383 & w29384);
assign w21580 = (w20323 & w29385) | (w20323 & w29386) | (w29385 & w29386);
assign v6823 = ~(w21579 | w21580);
assign w21581 = v6823;
assign w21582 = w21574 & ~w21581;
assign w21583 = pi14 & ~w21168;
assign v6824 = ~(w21174 | w21583);
assign w21584 = v6824;
assign w21585 = w21174 & w21583;
assign v6825 = ~(w21584 | w21585);
assign w21586 = v6825;
assign w21587 = w7177 & w20040;
assign w21588 = (~w21587 & w20038) | (~w21587 & w29589) | (w20038 & w29589);
assign w21589 = (w21588 & w20063) | (w21588 & w29387) | (w20063 & w29387);
assign w21590 = (w20339 & w29388) | (w20339 & w29389) | (w29388 & w29389);
assign w21591 = (~w20339 & w29390) | (~w20339 & w29391) | (w29390 & w29391);
assign v6826 = ~(w21590 | w21591);
assign w21592 = v6826;
assign w21593 = ~w21586 & w21592;
assign w21594 = w21162 & ~w21167;
assign v6827 = ~(w21168 | w21594);
assign w21595 = v6827;
assign w21596 = w7765 & ~w20038;
assign w21597 = w7177 & w20043;
assign w21598 = (~w21597 & ~w20040) | (~w21597 & w30565) | (~w20040 & w30565);
assign w21599 = ~w21596 & w21598;
assign w21600 = (w20294 & w29392) | (w20294 & w29393) | (w29392 & w29393);
assign w21601 = (~w20294 & w29394) | (~w20294 & w29395) | (w29394 & w29395);
assign v6828 = ~(w21600 | w21601);
assign w21602 = v6828;
assign w21603 = w21595 & w21602;
assign w21604 = w7172 & w20047;
assign w21605 = pi11 & w21604;
assign w21606 = w7178 & w20246;
assign w21607 = w7765 & ~w20052;
assign w21608 = w7466 & w20047;
assign v6829 = ~(w21607 | w21608);
assign w21609 = v6829;
assign w21610 = ~w21606 & w21609;
assign w21611 = ~w21605 & w21610;
assign w21612 = w7177 & w20047;
assign w21613 = (~w21612 & ~w20257) | (~w21612 & w29794) | (~w20257 & w29794);
assign w21614 = w7765 & w20043;
assign w21615 = w7466 & ~w20052;
assign v6830 = ~(w21614 | w21615);
assign w21616 = v6830;
assign w21617 = w21613 & w21616;
assign w21618 = w21613 & w30075;
assign w21619 = w21611 & w21618;
assign w21620 = w21161 & w21619;
assign v6831 = ~(w21161 | w21619);
assign w21621 = v6831;
assign v6832 = ~(w21620 | w21621);
assign w21622 = v6832;
assign w21623 = w7765 & w20040;
assign w21624 = w7177 & ~w20052;
assign w21625 = w7466 & w20043;
assign v6833 = ~(w21624 | w21625);
assign w21626 = v6833;
assign w21627 = ~w21623 & w21626;
assign w21628 = (w20272 & w29795) | (w20272 & w29796) | (w29795 & w29796);
assign w21629 = (~w20272 & w29797) | (~w20272 & w29798) | (w29797 & w29798);
assign v6834 = ~(w21628 | w21629);
assign w21630 = v6834;
assign w21631 = w21622 & ~w21630;
assign w21632 = (~w21620 & w21630) | (~w21620 & w30566) | (w21630 & w30566);
assign v6835 = ~(w21595 | w21602);
assign w21633 = v6835;
assign v6836 = ~(w21603 | w21633);
assign w21634 = v6836;
assign w21635 = ~w21632 & w21634;
assign w21636 = (~w21603 & ~w21634) | (~w21603 & w29591) | (~w21634 & w29591);
assign w21637 = w21586 & ~w21592;
assign v6837 = ~(w21593 | w21637);
assign w21638 = v6837;
assign w21639 = ~w21636 & w21638;
assign w21640 = (~w21593 & ~w21638) | (~w21593 & w29592) | (~w21638 & w29592);
assign w21641 = ~w21574 & w21581;
assign v6838 = ~(w21582 | w21641);
assign w21642 = v6838;
assign w21643 = ~w21640 & w21642;
assign w21644 = (~w21582 & ~w21642) | (~w21582 & w29593) | (~w21642 & w29593);
assign v6839 = ~(w21564 | w21571);
assign w21645 = v6839;
assign v6840 = ~(w21572 | w21645);
assign w21646 = v6840;
assign w21647 = ~w21644 & w21646;
assign w21648 = (~w21572 & ~w21646) | (~w21572 & w29594) | (~w21646 & w29594);
assign w21649 = ~w21554 & w21561;
assign v6841 = ~(w21562 | w21649);
assign w21650 = v6841;
assign w21651 = ~w21648 & w21650;
assign w21652 = (~w21562 & w21648) | (~w21562 & w31086) | (w21648 & w31086);
assign w21653 = ~w21543 & w21551;
assign v6842 = ~(w21552 | w21653);
assign w21654 = v6842;
assign w21655 = ~w21652 & w21654;
assign w21656 = (~w21552 & ~w21654) | (~w21552 & w29595) | (~w21654 & w29595);
assign v6843 = ~(w21532 | w21540);
assign w21657 = v6843;
assign v6844 = ~(w21541 | w21657);
assign w21658 = v6844;
assign w21659 = (~w29595 & w30694) | (~w29595 & w30695) | (w30694 & w30695);
assign w21660 = (~w21541 & w21656) | (~w21541 & w29799) | (w21656 & w29799);
assign w21661 = ~w21522 & w21529;
assign v6845 = ~(w21530 | w21661);
assign w21662 = v6845;
assign w21663 = ~w21660 & w21662;
assign w21664 = (~w21530 & w21660) | (~w21530 & w30696) | (w21660 & w30696);
assign w21665 = ~w21511 & w21519;
assign v6846 = ~(w21520 | w21665);
assign w21666 = v6846;
assign w21667 = ~w21664 & w21666;
assign w21668 = (~w21520 & w21664) | (~w21520 & w31087) | (w21664 & w31087);
assign v6847 = ~(w21500 | w21508);
assign w21669 = v6847;
assign v6848 = ~(w21509 | w21669);
assign w21670 = v6848;
assign w21671 = ~w21668 & w21670;
assign w21672 = (~w21509 & w21668) | (~w21509 & w30076) | (w21668 & w30076);
assign w21673 = ~w21489 & w21497;
assign v6849 = ~(w21498 | w21673);
assign w21674 = v6849;
assign w21675 = ~w21672 & w21674;
assign w21676 = (~w21498 & w21672) | (~w21498 & w30267) | (w21672 & w30267);
assign w21677 = ~w21478 & w21486;
assign v6850 = ~(w21487 | w21677);
assign w21678 = v6850;
assign w21679 = ~w21676 & w21678;
assign w21680 = (~w21487 & w21676) | (~w21487 & w30697) | (w21676 & w30697);
assign v6851 = ~(w21466 | w21475);
assign w21681 = v6851;
assign v6852 = ~(w21476 | w21681);
assign w21682 = v6852;
assign w21683 = ~w21680 & w21682;
assign w21684 = (~w21476 & w21680) | (~w21476 & w31088) | (w21680 & w31088);
assign v6853 = ~(w21453 | w21463);
assign w21685 = v6853;
assign v6854 = ~(w21464 | w21685);
assign w21686 = v6854;
assign w21687 = ~w21684 & w21686;
assign w21688 = (~w21464 & w21684) | (~w21464 & w30435) | (w21684 & w30435);
assign v6855 = ~(w21440 | w21450);
assign w21689 = v6855;
assign v6856 = ~(w21451 | w21689);
assign w21690 = v6856;
assign w21691 = ~w21688 & w21690;
assign w21692 = (~w21451 & w21688) | (~w21451 & w30567) | (w21688 & w30567);
assign v6857 = ~(w21427 | w21437);
assign w21693 = v6857;
assign v6858 = ~(w21438 | w21693);
assign w21694 = v6858;
assign w21695 = ~w21692 & w21694;
assign w21696 = (~w21438 & w21692) | (~w21438 & w30698) | (w21692 & w30698);
assign w21697 = ~w21414 & w21424;
assign v6859 = ~(w21425 | w21697);
assign w21698 = v6859;
assign w21699 = ~w21696 & w21698;
assign w21700 = (~w21425 & w21696) | (~w21425 & w31089) | (w21696 & w31089);
assign w21701 = ~w21399 & w21411;
assign v6860 = ~(w21412 | w21701);
assign w21702 = v6860;
assign w21703 = ~w21700 & w21702;
assign w21704 = (~w21412 & w21700) | (~w21412 & w30891) | (w21700 & w30891);
assign w21705 = (~w21396 & w21704) | (~w21396 & w31205) | (w21704 & w31205);
assign w21706 = w21381 & ~w21705;
assign w21707 = (~w21379 & ~w21381) | (~w21379 & w31206) | (~w21381 & w31206);
assign w21708 = w7765 & w19958;
assign w21709 = w7177 & w19966;
assign w21710 = w7466 & w19961;
assign v6861 = ~(w21709 | w21710);
assign w21711 = v6861;
assign w21712 = ~w21708 & w21711;
assign w21713 = ~pi11 & w21712;
assign v6862 = ~(w20123 | w20232);
assign w21714 = v6862;
assign w21715 = ~w19964 & w21714;
assign v6863 = ~(w20125 | w21715);
assign w21716 = v6863;
assign w21717 = w7178 & w21716;
assign w21718 = w21713 & ~w21717;
assign w21719 = w9464 & w21716;
assign w21720 = pi11 & ~w21712;
assign v6864 = ~(w21719 | w21720);
assign w21721 = v6864;
assign w21722 = ~w21718 & w21721;
assign w21723 = (~w21355 & w21254) | (~w21355 & w30568) | (w21254 & w30568);
assign w21724 = (~w21340 & w21255) | (~w21340 & w30892) | (w21255 & w30892);
assign v6865 = ~(w21326 | w21328);
assign w21725 = v6865;
assign w21726 = (~w21311 & w21257) | (~w21311 & w31090) | (w21257 & w31090);
assign w21727 = (~w21298 & ~w21300) | (~w21298 & w31091) | (~w21300 & w31091);
assign v6866 = ~(w21278 | w21288);
assign w21728 = v6866;
assign w21729 = w2418 & w5435;
assign v6867 = ~(w168 | w643);
assign w21730 = v6867;
assign w21731 = w1409 & w21730;
assign w21732 = w1462 & w21731;
assign w21733 = w4625 & w21732;
assign w21734 = ~w353 & w1066;
assign w21735 = w990 & w1535;
assign w21736 = w21734 & w21735;
assign w21737 = w21733 & w21736;
assign w21738 = w4571 & w6590;
assign w21739 = w3463 & w21738;
assign w21740 = w21737 & w21739;
assign w21741 = w789 & w21740;
assign w21742 = w21729 & w21741;
assign w21743 = w2599 & w21742;
assign w21744 = w1847 & w21743;
assign w21745 = w3406 & w20040;
assign w21746 = w3399 & ~w20052;
assign w21747 = w3402 & w20043;
assign v6868 = ~(w21746 | w21747);
assign w21748 = v6868;
assign w21749 = ~w21745 & w21748;
assign w21750 = (~w20272 & w31288) | (~w20272 & w31289) | (w31288 & w31289);
assign w21751 = (w20272 & w31290) | (w20272 & w31291) | (w31290 & w31291);
assign v6869 = ~(w21750 | w21751);
assign w21752 = v6869;
assign w21753 = ~w21728 & w21752;
assign w21754 = w21728 & ~w21752;
assign v6870 = ~(w21753 | w21754);
assign w21755 = v6870;
assign w21756 = w3760 & w20031;
assign w21757 = w3767 & ~w20038;
assign w21758 = w3763 & ~w20063;
assign v6871 = ~(w21757 | w21758);
assign w21759 = v6871;
assign w21760 = ~w21756 & w21759;
assign w21761 = (~w20323 & w31092) | (~w20323 & w31093) | (w31092 & w31093);
assign w21762 = (w20323 & w31094) | (w20323 & w31095) | (w31094 & w31095);
assign v6872 = ~(w21761 | w21762);
assign w21763 = v6872;
assign v6873 = ~(w21755 | w21763);
assign w21764 = v6873;
assign w21765 = w21755 & w21763;
assign v6874 = ~(w21764 | w21765);
assign w21766 = v6874;
assign w21767 = w21727 & ~w21766;
assign w21768 = ~w21727 & w21766;
assign v6875 = ~(w21767 | w21768);
assign w21769 = v6875;
assign v6876 = ~(w2873 | w20026);
assign w21770 = v6876;
assign w21771 = (~w21770 & ~w20014) | (~w21770 & w31292) | (~w20014 & w31292);
assign w21772 = w4158 & ~w20028;
assign w21773 = w21771 & ~w21772;
assign w21774 = (~w20472 & w31207) | (~w20472 & w31208) | (w31207 & w31208);
assign w21775 = (w20472 & w31209) | (w20472 & w31210) | (w31209 & w31210);
assign v6877 = ~(w21774 | w21775);
assign w21776 = v6877;
assign w21777 = w21769 & ~w21776;
assign w21778 = ~w21769 & w21776;
assign v6878 = ~(w21777 | w21778);
assign w21779 = v6878;
assign w21780 = ~w21726 & w21779;
assign w21781 = w21726 & ~w21779;
assign v6879 = ~(w21780 | w21781);
assign w21782 = v6879;
assign w21783 = w4913 & w20005;
assign w21784 = w4763 & ~w20011;
assign w21785 = w4836 & ~w20008;
assign v6880 = ~(w21784 | w21785);
assign w21786 = v6880;
assign w21787 = ~w21783 & w21786;
assign w21788 = (w31097 & w31211) | (w31097 & w31212) | (w31211 & w31212);
assign w21789 = (~w31097 & w31213) | (~w31097 & w31214) | (w31213 & w31214);
assign v6881 = ~(w21788 | w21789);
assign w21790 = v6881;
assign w21791 = w21782 & w21790;
assign v6882 = ~(w21782 | w21790);
assign w21792 = v6882;
assign v6883 = ~(w21791 | w21792);
assign w21793 = v6883;
assign w21794 = ~w21725 & w21793;
assign w21795 = w21725 & ~w21793;
assign v6884 = ~(w21794 | w21795);
assign w21796 = v6884;
assign w21797 = w5610 & ~w19992;
assign w21798 = w5531 & ~w19997;
assign w21799 = w5113 & w20000;
assign v6885 = ~(w21798 | w21799);
assign w21800 = v6885;
assign w21801 = ~w21797 & w21800;
assign w21802 = (w21801 & ~w20655) | (w21801 & w30894) | (~w20655 & w30894);
assign w21803 = pi20 & w21802;
assign v6886 = ~(pi20 | w21802);
assign w21804 = v6886;
assign v6887 = ~(w21803 | w21804);
assign w21805 = v6887;
assign w21806 = w21796 & ~w21805;
assign w21807 = ~w21796 & w21805;
assign v6888 = ~(w21806 | w21807);
assign w21808 = v6888;
assign w21809 = ~w21724 & w21808;
assign w21810 = w21724 & ~w21808;
assign v6889 = ~(w21809 | w21810);
assign w21811 = v6889;
assign w21812 = w5765 & w20997;
assign w21813 = w6236 & w19983;
assign w21814 = w5764 & w19989;
assign w21815 = w5983 & w19986;
assign v6890 = ~(w21814 | w21815);
assign w21816 = v6890;
assign w21817 = ~w21813 & w21816;
assign w21818 = ~w21812 & w21817;
assign w21819 = ~pi17 & w21818;
assign w21820 = pi17 & ~w21818;
assign v6891 = ~(w21819 | w21820);
assign w21821 = v6891;
assign w21822 = w21811 & w21821;
assign v6892 = ~(w21811 | w21821);
assign w21823 = v6892;
assign v6893 = ~(w21822 | w21823);
assign w21824 = v6893;
assign w21825 = ~w21723 & w21824;
assign w21826 = w21723 & ~w21824;
assign v6894 = ~(w21825 | w21826);
assign w21827 = v6894;
assign w21828 = w6389 & w21401;
assign w21829 = w6871 & w19974;
assign w21830 = w7004 & ~w19971;
assign v6895 = ~(w21829 | w21830);
assign w21831 = v6895;
assign w21832 = w6388 & w19980;
assign w21833 = w21831 & ~w21832;
assign w21834 = ~w21828 & w21833;
assign w21835 = pi14 & w21834;
assign v6896 = ~(pi14 | w21834);
assign w21836 = v6896;
assign v6897 = ~(w21835 | w21836);
assign w21837 = v6897;
assign w21838 = w21827 & ~w21837;
assign w21839 = ~w21827 & w21837;
assign v6898 = ~(w21838 | w21839);
assign w21840 = v6898;
assign w21841 = ~w21252 & w31098;
assign v6899 = ~(w21374 | w21841);
assign w21842 = v6899;
assign w21843 = w21840 & w21842;
assign v6900 = ~(w21840 | w21842);
assign w21844 = v6900;
assign v6901 = ~(w21843 | w21844);
assign w21845 = v6901;
assign w21846 = w21722 & w21845;
assign v6902 = ~(w21722 | w21845);
assign w21847 = v6902;
assign v6903 = ~(w21846 | w21847);
assign w21848 = v6903;
assign v6904 = ~(w21707 | w21848);
assign w21849 = v6904;
assign w21850 = w21707 & w21848;
assign v6905 = ~(w21849 | w21850);
assign w21851 = v6905;
assign w21852 = ~w20224 & w21851;
assign w21853 = w20224 & ~w21851;
assign v6906 = ~(w21852 | w21853);
assign w21854 = v6906;
assign w21855 = ~w21381 & w21705;
assign v6907 = ~(w21706 | w21855);
assign w21856 = v6907;
assign w21857 = w8926 & w19954;
assign w21858 = w8140 & w19958;
assign w21859 = w8526 & w19952;
assign v6908 = ~(w21858 | w21859);
assign w21860 = v6908;
assign w21861 = ~w21857 & w21860;
assign w21862 = pi08 & ~w21861;
assign v6909 = ~(w19955 | w19956);
assign w21863 = v6909;
assign w21864 = w20130 & ~w21863;
assign w21865 = ~w20130 & w21863;
assign v6910 = ~(w21864 | w21865);
assign w21866 = v6910;
assign w21867 = w8141 & ~w21866;
assign w21868 = ~pi08 & w21861;
assign w21869 = ~w21867 & w21868;
assign w21870 = w9920 & ~w21866;
assign v6911 = ~(w21869 | w21870);
assign w21871 = v6911;
assign w21872 = ~w21862 & w21871;
assign v6912 = ~(w21856 | w21872);
assign w21873 = v6912;
assign w21874 = w21856 & w21872;
assign w21875 = w8926 & w19952;
assign w21876 = w8526 & w19958;
assign w21877 = w8140 & w19961;
assign v6913 = ~(w21876 | w21877);
assign w21878 = v6913;
assign w21879 = ~w21875 & w21878;
assign w21880 = ~pi08 & w21879;
assign v6914 = ~(w20126 | w20128);
assign w21881 = v6914;
assign v6915 = ~(w20129 | w21881);
assign w21882 = v6915;
assign w21883 = w8141 & ~w21882;
assign w21884 = w21880 & ~w21883;
assign w21885 = w9920 & ~w21882;
assign w21886 = pi08 & ~w21879;
assign v6916 = ~(w21885 | w21886);
assign w21887 = v6916;
assign w21888 = ~w21884 & w21887;
assign v6917 = ~(w21396 | w21397);
assign w21889 = v6917;
assign w21890 = ~w21704 & w21889;
assign w21891 = w21704 & ~w21889;
assign v6918 = ~(w21890 | w21891);
assign w21892 = v6918;
assign w21893 = w21888 & w21892;
assign v6919 = ~(w21888 | w21892);
assign w21894 = v6919;
assign v6920 = ~(w21893 | w21894);
assign w21895 = v6920;
assign w21896 = w8141 & w21716;
assign w21897 = w8926 & w19958;
assign w21898 = w8526 & w19961;
assign w21899 = w8140 & w19966;
assign v6921 = ~(w21898 | w21899);
assign w21900 = v6921;
assign w21901 = ~w21897 & w21900;
assign w21902 = ~pi08 & w21901;
assign w21903 = ~w21896 & w21902;
assign w21904 = w9920 & w21716;
assign w21905 = pi08 & ~w21901;
assign v6922 = ~(w21904 | w21905);
assign w21906 = v6922;
assign w21907 = ~w21903 & w21906;
assign w21908 = w21700 & ~w21702;
assign v6923 = ~(w21703 | w21908);
assign w21909 = v6923;
assign v6924 = ~(w21907 | w21909);
assign w21910 = v6924;
assign w21911 = w21907 & w21909;
assign w21912 = w21696 & ~w21698;
assign v6925 = ~(w21699 | w21912);
assign w21913 = v6925;
assign w21914 = w9920 & w20234;
assign w21915 = w8926 & w19961;
assign w21916 = w8526 & w19966;
assign w21917 = w8140 & ~w19971;
assign v6926 = ~(w21916 | w21917);
assign w21918 = v6926;
assign w21919 = ~w21915 & w21918;
assign w21920 = pi08 & ~w21919;
assign w21921 = w8141 & w20234;
assign w21922 = ~pi08 & w21919;
assign w21923 = ~w21921 & w21922;
assign v6927 = ~(w21920 | w21923);
assign w21924 = v6927;
assign w21925 = ~w21914 & w21924;
assign w21926 = w21913 & w21925;
assign v6928 = ~(w21913 | w21925);
assign w21927 = v6928;
assign v6929 = ~(w21926 | w21927);
assign w21928 = v6929;
assign w21929 = w21692 & ~w21694;
assign v6930 = ~(w21695 | w21929);
assign w21930 = v6930;
assign w21931 = w8141 & w21385;
assign w21932 = w8526 & ~w19971;
assign w21933 = w8926 & w19966;
assign v6931 = ~(w21932 | w21933);
assign w21934 = v6931;
assign w21935 = w8140 & w19974;
assign w21936 = w21934 & ~w21935;
assign w21937 = ~w21931 & w21936;
assign w21938 = pi08 & w21937;
assign v6932 = ~(pi08 | w21937);
assign w21939 = v6932;
assign v6933 = ~(w21938 | w21939);
assign w21940 = v6933;
assign w21941 = ~w21930 & w21940;
assign w21942 = w21930 & ~w21940;
assign w21943 = w21688 & ~w21690;
assign v6934 = ~(w21691 | w21943);
assign w21944 = v6934;
assign w21945 = w8141 & w21401;
assign w21946 = w8926 & ~w19971;
assign w21947 = w8526 & w19974;
assign w21948 = w8140 & w19980;
assign v6935 = ~(w21947 | w21948);
assign w21949 = v6935;
assign w21950 = ~w21946 & w21949;
assign w21951 = ~w21945 & w21950;
assign w21952 = ~pi08 & w21951;
assign w21953 = pi08 & ~w21951;
assign v6936 = ~(w21952 | w21953);
assign w21954 = v6936;
assign w21955 = w21944 & w21954;
assign v6937 = ~(w21944 | w21954);
assign w21956 = v6937;
assign v6938 = ~(w21955 | w21956);
assign w21957 = v6938;
assign w21958 = w21684 & ~w21686;
assign v6939 = ~(w21687 | w21958);
assign w21959 = v6939;
assign w21960 = w8141 & w21362;
assign w21961 = w8926 & w19974;
assign w21962 = w8526 & w19980;
assign w21963 = w8140 & w19983;
assign v6940 = ~(w21962 | w21963);
assign w21964 = v6940;
assign w21965 = ~w21961 & w21964;
assign w21966 = ~w21960 & w21965;
assign w21967 = pi08 & ~w21966;
assign w21968 = ~pi08 & w21966;
assign v6941 = ~(w21967 | w21968);
assign w21969 = v6941;
assign v6942 = ~(w21959 | w21969);
assign w21970 = v6942;
assign w21971 = w21680 & ~w21682;
assign v6943 = ~(w21683 | w21971);
assign w21972 = v6943;
assign w21973 = w8141 & w20982;
assign w21974 = w8526 & w19983;
assign w21975 = w8926 & w19980;
assign v6944 = ~(w21974 | w21975);
assign w21976 = v6944;
assign w21977 = w8140 & w19986;
assign w21978 = w21976 & ~w21977;
assign w21979 = ~w21973 & w21978;
assign w21980 = pi08 & w21979;
assign v6945 = ~(pi08 | w21979);
assign w21981 = v6945;
assign v6946 = ~(w21980 | w21981);
assign w21982 = v6946;
assign w21983 = w21972 & ~w21982;
assign w21984 = w21676 & ~w21678;
assign v6947 = ~(w21679 | w21984);
assign w21985 = v6947;
assign w21986 = w8141 & w20997;
assign w21987 = w8926 & w19983;
assign w21988 = w8140 & w19989;
assign w21989 = w8526 & w19986;
assign v6948 = ~(w21988 | w21989);
assign w21990 = v6948;
assign w21991 = ~w21987 & w21990;
assign w21992 = ~w21986 & w21991;
assign w21993 = ~pi08 & w21992;
assign w21994 = pi08 & ~w21992;
assign v6949 = ~(w21993 | w21994);
assign w21995 = v6949;
assign w21996 = w21985 & w21995;
assign w21997 = w21672 & ~w21674;
assign v6950 = ~(w21675 | w21997);
assign w21998 = v6950;
assign w21999 = w8141 & w21012;
assign w22000 = w8140 & ~w19992;
assign w22001 = w8926 & w19986;
assign v6951 = ~(w22000 | w22001);
assign w22002 = v6951;
assign w22003 = w8526 & w19989;
assign w22004 = w22002 & ~w22003;
assign w22005 = ~w21999 & w22004;
assign w22006 = pi08 & w22005;
assign v6952 = ~(pi08 | w22005);
assign w22007 = v6952;
assign v6953 = ~(w22006 | w22007);
assign w22008 = v6953;
assign w22009 = w21998 & ~w22008;
assign w22010 = w21668 & ~w21670;
assign v6954 = ~(w21671 | w22010);
assign w22011 = v6954;
assign w22012 = w8926 & w19989;
assign w22013 = w8140 & ~w19997;
assign w22014 = w8526 & ~w19992;
assign v6955 = ~(w22013 | w22014);
assign w22015 = v6955;
assign w22016 = ~w22012 & w22015;
assign w22017 = (w22016 & ~w20965) | (w22016 & w30268) | (~w20965 & w30268);
assign w22018 = ~pi08 & w22017;
assign w22019 = pi08 & ~w22017;
assign v6956 = ~(w22018 | w22019);
assign w22020 = v6956;
assign w22021 = w22011 & w22020;
assign w22022 = w21664 & ~w21666;
assign v6957 = ~(w21667 | w22022);
assign w22023 = v6957;
assign w22024 = w8926 & ~w19992;
assign w22025 = w8526 & ~w19997;
assign w22026 = w8140 & w20000;
assign v6958 = ~(w22025 | w22026);
assign w22027 = v6958;
assign w22028 = ~w22024 & w22027;
assign w22029 = (~w29800 & w30269) | (~w29800 & w30270) | (w30269 & w30270);
assign w22030 = (w29800 & w30271) | (w29800 & w30272) | (w30271 & w30272);
assign v6959 = ~(w22029 | w22030);
assign w22031 = v6959;
assign w22032 = w22023 & ~w22031;
assign w22033 = w21660 & ~w21662;
assign v6960 = ~(w21663 | w22033);
assign w22034 = v6960;
assign w22035 = w8140 & w20005;
assign w22036 = w8926 & ~w19997;
assign v6961 = ~(w22035 | w22036);
assign w22037 = v6961;
assign w22038 = w8526 & w20000;
assign w22039 = w22037 & ~w22038;
assign w22040 = (~w20668 & w30078) | (~w20668 & w30079) | (w30078 & w30079);
assign w22041 = (w20668 & w30080) | (w20668 & w30081) | (w30080 & w30081);
assign v6962 = ~(w22040 | w22041);
assign w22042 = v6962;
assign w22043 = w22034 & ~w22042;
assign w22044 = (w29595 & w30700) | (w29595 & w30701) | (w30700 & w30701);
assign v6963 = ~(w21659 | w22044);
assign w22045 = v6963;
assign w22046 = w8926 & w20000;
assign w22047 = w8140 & ~w20008;
assign w22048 = w8526 & w20005;
assign v6964 = ~(w22047 | w22048);
assign w22049 = v6964;
assign w22050 = ~w22046 & w22049;
assign w22051 = (w20681 & w30082) | (w20681 & w30083) | (w30082 & w30083);
assign w22052 = (~w20681 & w30084) | (~w20681 & w30085) | (w30084 & w30085);
assign v6965 = ~(w22051 | w22052);
assign w22053 = v6965;
assign w22054 = w22045 & w22053;
assign w22055 = w21652 & ~w21654;
assign v6966 = ~(w21655 | w22055);
assign w22056 = v6966;
assign w22057 = w8926 & w20005;
assign w22058 = w8140 & ~w20011;
assign w22059 = w8526 & ~w20008;
assign v6967 = ~(w22058 | w22059);
assign w22060 = v6967;
assign w22061 = ~w22057 & w22060;
assign w22062 = (w29597 & ~w29396) | (w29597 & w29802) | (~w29396 & w29802);
assign w22063 = (w29396 & w29803) | (w29396 & w29804) | (w29803 & w29804);
assign v6968 = ~(w22062 | w22063);
assign w22064 = v6968;
assign w22065 = w22056 & w22064;
assign w22066 = w21648 & ~w21650;
assign v6969 = ~(w21651 | w22066);
assign w22067 = v6969;
assign w22068 = w8526 & ~w20011;
assign w22069 = w8926 & ~w20008;
assign v6970 = ~(w22068 | w22069);
assign w22070 = v6970;
assign w22071 = w8140 & w20014;
assign w22072 = w22070 & ~w22071;
assign w22073 = (w29397 & ~w29063) | (w29397 & w29923) | (~w29063 & w29923);
assign w22074 = (w29063 & w29924) | (w29063 & w29925) | (w29924 & w29925);
assign v6971 = ~(w22073 | w22074);
assign w22075 = v6971;
assign w22076 = w22067 & ~w22075;
assign w22077 = w21644 & ~w21646;
assign v6972 = ~(w21647 | w22077);
assign w22078 = v6972;
assign w22079 = w8926 & ~w20011;
assign w22080 = w8140 & ~w20028;
assign w22081 = (~w22080 & ~w20014) | (~w22080 & w29599) | (~w20014 & w29599);
assign w22082 = ~w22079 & w22081;
assign w22083 = (~w20459 & w29399) | (~w20459 & w29400) | (w29399 & w29400);
assign w22084 = (w20459 & w29401) | (w20459 & w29402) | (w29401 & w29402);
assign v6973 = ~(w22083 | w22084);
assign w22085 = v6973;
assign w22086 = w22078 & w22085;
assign w22087 = w21640 & ~w21642;
assign v6974 = ~(w21643 | w22087);
assign w22088 = v6974;
assign w22089 = w8141 & w20472;
assign w22090 = w8526 & ~w20028;
assign w22091 = (~w22090 & ~w20014) | (~w22090 & w29403) | (~w20014 & w29403);
assign w22092 = w8140 & ~w20026;
assign w22093 = w22091 & ~w22092;
assign w22094 = ~w22089 & w29065;
assign w22095 = (~pi08 & w22089) | (~pi08 & w29066) | (w22089 & w29066);
assign v6975 = ~(w22094 | w22095);
assign w22096 = v6975;
assign w22097 = w22088 & ~w22096;
assign w22098 = w21636 & ~w21638;
assign v6976 = ~(w21639 | w22098);
assign w22099 = v6976;
assign w22100 = w8926 & ~w20028;
assign w22101 = w8140 & w20031;
assign w22102 = (~w22101 & w20026) | (~w22101 & w29404) | (w20026 & w29404);
assign w22103 = ~w22100 & w22102;
assign w22104 = (w20431 & w29067) | (w20431 & w29068) | (w29067 & w29068);
assign w22105 = (~w20431 & w29069) | (~w20431 & w29070) | (w29069 & w29070);
assign v6977 = ~(w22104 | w22105);
assign w22106 = v6977;
assign w22107 = w22099 & w22106;
assign w22108 = w21632 & ~w21634;
assign v6978 = ~(w21635 | w22108);
assign w22109 = v6978;
assign w22110 = w8140 & ~w20063;
assign w22111 = (~w22110 & w20026) | (~w22110 & w29071) | (w20026 & w29071);
assign w22112 = w8526 & w20031;
assign w22113 = (w20026 & w29405) | (w20026 & w29406) | (w29405 & w29406);
assign w22114 = (w20311 & w29072) | (w20311 & w29073) | (w29072 & w29073);
assign w22115 = (~w20311 & w29074) | (~w20311 & w29075) | (w29074 & w29075);
assign v6979 = ~(w22114 | w22115);
assign w22116 = v6979;
assign w22117 = w22109 & ~w22116;
assign w22118 = ~w21622 & w21630;
assign v6980 = ~(w21631 | w22118);
assign w22119 = v6980;
assign w22120 = w8526 & ~w20063;
assign w22121 = w8926 & w20031;
assign v6981 = ~(w22120 | w22121);
assign w22122 = v6981;
assign w22123 = w8140 & ~w20038;
assign w22124 = ~w22121 & w29407;
assign w22125 = (~w20323 & w29076) | (~w20323 & w29077) | (w29076 & w29077);
assign w22126 = (w20323 & w29078) | (w20323 & w29079) | (w29078 & w29079);
assign v6982 = ~(w22125 | w22126);
assign w22127 = v6982;
assign w22128 = w22119 & ~w22127;
assign w22129 = pi11 & ~w21611;
assign v6983 = ~(w21617 | w22129);
assign w22130 = v6983;
assign w22131 = w21617 & w22129;
assign v6984 = ~(w22130 | w22131);
assign w22132 = v6984;
assign w22133 = w8140 & w20040;
assign w22134 = (~w22133 & w20038) | (~w22133 & w29408) | (w20038 & w29408);
assign w22135 = (w22134 & w20063) | (w22134 & w29080) | (w20063 & w29080);
assign w22136 = (w20339 & w29081) | (w20339 & w29082) | (w29081 & w29082);
assign w22137 = (~w20339 & w29083) | (~w20339 & w29084) | (w29083 & w29084);
assign v6985 = ~(w22136 | w22137);
assign w22138 = v6985;
assign w22139 = ~w22132 & w22138;
assign w22140 = w21605 & ~w21610;
assign v6986 = ~(w21611 | w22140);
assign w22141 = v6986;
assign w22142 = w8926 & ~w20038;
assign w22143 = w8140 & w20043;
assign w22144 = (~w22143 & ~w20040) | (~w22143 & w30702) | (~w20040 & w30702);
assign w22145 = ~w22142 & w22144;
assign w22146 = (~w20294 & w29085) | (~w20294 & w29086) | (w29085 & w29086);
assign w22147 = (w20294 & w29087) | (w20294 & w29088) | (w29087 & w29088);
assign v6987 = ~(w22146 | w22147);
assign w22148 = v6987;
assign w22149 = w22141 & w22148;
assign w22150 = w8141 & w20246;
assign w22151 = w8526 & w20047;
assign w22152 = w8926 & ~w20052;
assign v6988 = ~(w22151 | w22152);
assign w22153 = v6988;
assign w22154 = ~w22150 & w22153;
assign w22155 = w8138 & w20047;
assign w22156 = pi08 & w22155;
assign w22157 = w22154 & ~w22156;
assign w22158 = w8140 & w20047;
assign w22159 = (~w22158 & ~w20257) | (~w22158 & w29600) | (~w20257 & w29600);
assign w22160 = w8926 & w20043;
assign w22161 = w8526 & ~w20052;
assign v6989 = ~(w22160 | w22161);
assign w22162 = v6989;
assign w22163 = w22159 & w22162;
assign w22164 = w22159 & w30703;
assign w22165 = w22157 & w22164;
assign w22166 = w21604 & w22165;
assign v6990 = ~(w21604 | w22165);
assign w22167 = v6990;
assign v6991 = ~(w22166 | w22167);
assign w22168 = v6991;
assign w22169 = w8526 & w20043;
assign w22170 = w8140 & ~w20052;
assign w22171 = (~w20040 & w30704) | (~w20040 & w30705) | (w30704 & w30705);
assign w22172 = (w20272 & w29602) | (w20272 & w29603) | (w29602 & w29603);
assign w22173 = (~w20272 & w29604) | (~w20272 & w29605) | (w29604 & w29605);
assign v6992 = ~(w22172 | w22173);
assign w22174 = v6992;
assign w22175 = w22168 & w22174;
assign w22176 = (~w22166 & ~w22174) | (~w22166 & w30706) | (~w22174 & w30706);
assign v6993 = ~(w22141 | w22148);
assign w22177 = v6993;
assign v6994 = ~(w22149 | w22177);
assign w22178 = v6994;
assign w22179 = ~w22176 & w22178;
assign w22180 = (~w22149 & ~w22178) | (~w22149 & w29410) | (~w22178 & w29410);
assign w22181 = w22132 & ~w22138;
assign v6995 = ~(w22139 | w22181);
assign w22182 = v6995;
assign w22183 = ~w22180 & w22182;
assign w22184 = (~w22139 & ~w22182) | (~w22139 & w29411) | (~w22182 & w29411);
assign w22185 = ~w22119 & w22127;
assign v6996 = ~(w22128 | w22185);
assign w22186 = v6996;
assign w22187 = ~w22184 & w22186;
assign w22188 = (~w22128 & ~w22186) | (~w22128 & w29412) | (~w22186 & w29412);
assign w22189 = ~w22109 & w22116;
assign v6997 = ~(w22117 | w22189);
assign w22190 = v6997;
assign w22191 = ~w22188 & w22190;
assign w22192 = (~w22117 & ~w22190) | (~w22117 & w29413) | (~w22190 & w29413);
assign v6998 = ~(w22099 | w22106);
assign w22193 = v6998;
assign v6999 = ~(w22107 | w22193);
assign w22194 = v6999;
assign w22195 = ~w22192 & w22194;
assign w22196 = (~w22107 & w22192) | (~w22107 & w31099) | (w22192 & w31099);
assign w22197 = ~w22088 & w22096;
assign v7000 = ~(w22097 | w22197);
assign w22198 = v7000;
assign w22199 = ~w22196 & w22198;
assign w22200 = (~w22097 & ~w22198) | (~w22097 & w29414) | (~w22198 & w29414);
assign v7001 = ~(w22078 | w22085);
assign w22201 = v7001;
assign v7002 = ~(w22086 | w22201);
assign w22202 = v7002;
assign w22203 = (~w29414 & w30707) | (~w29414 & w30708) | (w30707 & w30708);
assign w22204 = (~w22086 & w22200) | (~w22086 & w29805) | (w22200 & w29805);
assign w22205 = ~w22067 & w22075;
assign v7003 = ~(w22076 | w22205);
assign w22206 = v7003;
assign w22207 = ~w22204 & w22206;
assign v7004 = ~(w22076 | w22207);
assign w22208 = v7004;
assign v7005 = ~(w22056 | w22064);
assign w22209 = v7005;
assign v7006 = ~(w22065 | w22209);
assign w22210 = v7006;
assign w22211 = ~w22208 & w22210;
assign w22212 = (~w22065 & w22208) | (~w22065 & w29606) | (w22208 & w29606);
assign v7007 = ~(w22045 | w22053);
assign w22213 = v7007;
assign v7008 = ~(w22054 | w22213);
assign w22214 = v7008;
assign w22215 = ~w22212 & w22214;
assign w22216 = (~w22054 & w22212) | (~w22054 & w29926) | (w22212 & w29926);
assign w22217 = ~w22034 & w22042;
assign v7009 = ~(w22043 | w22217);
assign w22218 = v7009;
assign w22219 = ~w22216 & w22218;
assign w22220 = (~w22043 & w22216) | (~w22043 & w30086) | (w22216 & w30086);
assign w22221 = ~w22023 & w22031;
assign v7010 = ~(w22032 | w22221);
assign w22222 = v7010;
assign w22223 = ~w22220 & w22222;
assign w22224 = (~w22032 & w22220) | (~w22032 & w30709) | (w22220 & w30709);
assign v7011 = ~(w22011 | w22020);
assign w22225 = v7011;
assign v7012 = ~(w22021 | w22225);
assign w22226 = v7012;
assign w22227 = ~w22224 & w22226;
assign w22228 = (~w22021 & w22224) | (~w22021 & w31100) | (w22224 & w31100);
assign w22229 = ~w21998 & w22008;
assign v7013 = ~(w22009 | w22229);
assign w22230 = v7013;
assign w22231 = ~w22228 & w22230;
assign w22232 = (~w22009 & w22228) | (~w22009 & w30273) | (w22228 & w30273);
assign v7014 = ~(w21985 | w21995);
assign w22233 = v7014;
assign v7015 = ~(w21996 | w22233);
assign w22234 = v7015;
assign w22235 = ~w22232 & w22234;
assign w22236 = (~w21996 & w22232) | (~w21996 & w30436) | (w22232 & w30436);
assign w22237 = ~w21972 & w21982;
assign v7016 = ~(w21983 | w22237);
assign w22238 = v7016;
assign w22239 = ~w22236 & w22238;
assign w22240 = (~w21983 & w22236) | (~w21983 & w30710) | (w22236 & w30710);
assign w22241 = w21959 & w21969;
assign v7017 = ~(w21970 | w22241);
assign w22242 = v7017;
assign w22243 = w22240 & w22242;
assign w22244 = (~w21970 & ~w22240) | (~w21970 & w31101) | (~w22240 & w31101);
assign w22245 = w21957 & w22244;
assign w22246 = (~w21955 & ~w22244) | (~w21955 & w30569) | (~w22244 & w30569);
assign w22247 = (~w21941 & ~w22246) | (~w21941 & w30895) | (~w22246 & w30895);
assign w22248 = w21928 & w22247;
assign v7018 = ~(w21926 | w22248);
assign w22249 = v7018;
assign w22250 = ~w22248 & w31102;
assign v7019 = ~(w21910 | w22250);
assign w22251 = v7019;
assign w22252 = w21895 & w22251;
assign w22253 = (~w21893 & ~w22251) | (~w21893 & w31215) | (~w22251 & w31215);
assign w22254 = ~w21874 & w22253;
assign v7020 = ~(w21873 | w22254);
assign w22255 = v7020;
assign w22256 = w21854 & ~w22255;
assign w22257 = ~w21854 & w22255;
assign v7021 = ~(w22256 | w22257);
assign w22258 = v7021;
assign v7022 = ~(w19930 | w19931);
assign w22259 = v7022;
assign v7023 = ~(w20139 | w22259);
assign w22260 = v7023;
assign w22261 = w20139 & w22259;
assign v7024 = ~(w22260 | w22261);
assign w22262 = v7024;
assign w22263 = w10445 & w22262;
assign w22264 = w10447 & w22262;
assign w22265 = w10419 & ~w19923;
assign w22266 = w9401 & w19933;
assign w22267 = w9891 & ~w19929;
assign v7025 = ~(w22266 | w22267);
assign w22268 = v7025;
assign w22269 = ~w22265 & w22268;
assign w22270 = pi05 & w22269;
assign v7026 = ~(pi05 | w22269);
assign w22271 = v7026;
assign v7027 = ~(w22270 | w22271);
assign w22272 = v7027;
assign w22273 = ~w22264 & w22272;
assign v7028 = ~(w22263 | w22273);
assign w22274 = v7028;
assign w22275 = ~w22258 & w22274;
assign w22276 = w22258 & ~w22274;
assign v7029 = ~(w22275 | w22276);
assign w22277 = v7029;
assign v7030 = ~(w21873 | w21874);
assign w22278 = v7030;
assign v7031 = ~(w22253 | w22278);
assign w22279 = v7031;
assign w22280 = w22253 & w22278;
assign v7032 = ~(w22279 | w22280);
assign w22281 = v7032;
assign v7033 = ~(w19934 | w19935);
assign w22282 = v7033;
assign v7034 = ~(w20137 | w22282);
assign w22283 = v7034;
assign w22284 = w20137 & w22282;
assign v7035 = ~(w22283 | w22284);
assign w22285 = v7035;
assign w22286 = w9402 & ~w22285;
assign w22287 = w10419 & ~w19929;
assign w22288 = w9401 & ~w19939;
assign w22289 = w9891 & w19933;
assign v7036 = ~(w22288 | w22289);
assign w22290 = v7036;
assign w22291 = ~w22287 & w22290;
assign w22292 = ~w22286 & w22291;
assign w22293 = ~pi05 & w22292;
assign w22294 = pi05 & ~w22292;
assign v7037 = ~(w22293 | w22294);
assign w22295 = v7037;
assign w22296 = w22281 & ~w22295;
assign w22297 = ~w22281 & w22295;
assign v7038 = ~(w22296 | w22297);
assign w22298 = v7038;
assign v7039 = ~(w21895 | w22251);
assign w22299 = v7039;
assign v7040 = ~(w22252 | w22299);
assign w22300 = v7040;
assign v7041 = ~(w19940 | w19941);
assign w22301 = v7041;
assign w22302 = w20135 & w22301;
assign v7042 = ~(w20135 | w22301);
assign w22303 = v7042;
assign v7043 = ~(w22302 | w22303);
assign w22304 = v7043;
assign w22305 = w9402 & ~w22304;
assign w22306 = w10419 & w19933;
assign w22307 = w9401 & w19954;
assign w22308 = w9891 & ~w19939;
assign v7044 = ~(w22307 | w22308);
assign w22309 = v7044;
assign w22310 = ~w22306 & w22309;
assign w22311 = ~w22305 & w22310;
assign w22312 = ~pi05 & w22311;
assign w22313 = pi05 & ~w22311;
assign v7045 = ~(w22312 | w22313);
assign w22314 = v7045;
assign v7046 = ~(w22300 | w22314);
assign w22315 = v7046;
assign w22316 = w22300 & w22314;
assign w22317 = w9402 & w20214;
assign w22318 = w9891 & w19954;
assign w22319 = w10419 & ~w19939;
assign v7047 = ~(w22318 | w22319);
assign w22320 = v7047;
assign w22321 = w9401 & w19952;
assign w22322 = w22320 & ~w22321;
assign w22323 = ~w22317 & w22322;
assign v7048 = ~(pi05 | w22323);
assign w22324 = v7048;
assign w22325 = pi05 & w22323;
assign v7049 = ~(w22324 | w22325);
assign w22326 = v7049;
assign v7050 = ~(w21910 | w21911);
assign w22327 = v7050;
assign w22328 = w22249 & w22327;
assign v7051 = ~(w22249 | w22327);
assign w22329 = v7051;
assign v7052 = ~(w22328 | w22329);
assign w22330 = v7052;
assign v7053 = ~(w22326 | w22330);
assign w22331 = v7053;
assign w22332 = w22326 & w22330;
assign v7054 = ~(w22331 | w22332);
assign w22333 = v7054;
assign v7055 = ~(w21928 | w22247);
assign w22334 = v7055;
assign v7056 = ~(w22248 | w22334);
assign w22335 = v7056;
assign w22336 = w9402 & ~w21866;
assign w22337 = w9891 & w19952;
assign w22338 = w10419 & w19954;
assign v7057 = ~(w22337 | w22338);
assign w22339 = v7057;
assign w22340 = w9401 & w19958;
assign w22341 = w22339 & ~w22340;
assign w22342 = ~w22336 & w22341;
assign w22343 = pi05 & w22342;
assign v7058 = ~(pi05 | w22342);
assign w22344 = v7058;
assign v7059 = ~(w22343 | w22344);
assign w22345 = v7059;
assign w22346 = ~w22335 & w22345;
assign w22347 = w22335 & ~w22345;
assign w22348 = w9402 & ~w21882;
assign w22349 = w10419 & w19952;
assign w22350 = w9891 & w19958;
assign w22351 = w9401 & w19961;
assign v7060 = ~(w22350 | w22351);
assign w22352 = v7060;
assign w22353 = ~w22349 & w22352;
assign w22354 = ~w22348 & w22353;
assign w22355 = pi05 & ~w22354;
assign w22356 = ~pi05 & w22354;
assign v7061 = ~(w22355 | w22356);
assign w22357 = v7061;
assign v7062 = ~(w21941 | w21942);
assign w22358 = v7062;
assign w22359 = w22246 & w22358;
assign v7063 = ~(w22246 | w22358);
assign w22360 = v7063;
assign v7064 = ~(w22359 | w22360);
assign w22361 = v7064;
assign w22362 = w22357 & ~w22361;
assign v7065 = ~(w21957 | w22244);
assign w22363 = v7065;
assign v7066 = ~(w22245 | w22363);
assign w22364 = v7066;
assign w22365 = w9402 & w21716;
assign w22366 = w9891 & w19961;
assign w22367 = w10419 & w19958;
assign v7067 = ~(w22366 | w22367);
assign w22368 = v7067;
assign w22369 = w9401 & w19966;
assign w22370 = w22368 & ~w22369;
assign w22371 = ~w22365 & w22370;
assign v7068 = ~(pi05 | w22371);
assign w22372 = v7068;
assign w22373 = pi05 & w22371;
assign v7069 = ~(w22372 | w22373);
assign w22374 = v7069;
assign w22375 = w22364 & ~w22374;
assign v7070 = ~(w22240 | w22242);
assign w22376 = v7070;
assign v7071 = ~(w22243 | w22376);
assign w22377 = v7071;
assign w22378 = w9402 & w20234;
assign w22379 = w9891 & w19966;
assign w22380 = w10419 & w19961;
assign v7072 = ~(w22379 | w22380);
assign w22381 = v7072;
assign w22382 = w9401 & ~w19971;
assign w22383 = w22381 & ~w22382;
assign w22384 = ~w22378 & w22383;
assign v7073 = ~(pi05 | w22384);
assign w22385 = v7073;
assign w22386 = pi05 & w22384;
assign v7074 = ~(w22385 | w22386);
assign w22387 = v7074;
assign v7075 = ~(w22377 | w22387);
assign w22388 = v7075;
assign w22389 = w22236 & ~w22238;
assign v7076 = ~(w22239 | w22389);
assign w22390 = v7076;
assign w22391 = w9402 & w21385;
assign w22392 = w9891 & ~w19971;
assign w22393 = w10419 & w19966;
assign v7077 = ~(w22392 | w22393);
assign w22394 = v7077;
assign w22395 = w9401 & w19974;
assign w22396 = w22394 & ~w22395;
assign w22397 = ~w22391 & w22396;
assign v7078 = ~(pi05 | w22397);
assign w22398 = v7078;
assign w22399 = pi05 & w22397;
assign v7079 = ~(w22398 | w22399);
assign w22400 = v7079;
assign w22401 = w22390 & ~w22400;
assign w22402 = w22232 & ~w22234;
assign v7080 = ~(w22235 | w22402);
assign w22403 = v7080;
assign w22404 = w9402 & w21401;
assign w22405 = w10419 & ~w19971;
assign w22406 = w9401 & w19980;
assign w22407 = w9891 & w19974;
assign v7081 = ~(w22406 | w22407);
assign w22408 = v7081;
assign w22409 = ~w22405 & w22408;
assign w22410 = ~w22404 & w22409;
assign w22411 = pi05 & w22410;
assign v7082 = ~(pi05 | w22410);
assign w22412 = v7082;
assign v7083 = ~(w22411 | w22412);
assign w22413 = v7083;
assign w22414 = w22403 & ~w22413;
assign w22415 = w22228 & ~w22230;
assign v7084 = ~(w22231 | w22415);
assign w22416 = v7084;
assign w22417 = w9402 & w21362;
assign w22418 = w9891 & w19980;
assign w22419 = w10419 & w19974;
assign v7085 = ~(w22418 | w22419);
assign w22420 = v7085;
assign w22421 = w9401 & w19983;
assign w22422 = w22420 & ~w22421;
assign w22423 = ~w22417 & w22422;
assign w22424 = pi05 & w22423;
assign v7086 = ~(pi05 | w22423);
assign w22425 = v7086;
assign v7087 = ~(w22424 | w22425);
assign w22426 = v7087;
assign w22427 = w22416 & ~w22426;
assign w22428 = w22224 & ~w22226;
assign v7088 = ~(w22227 | w22428);
assign w22429 = v7088;
assign w22430 = w9402 & w20982;
assign w22431 = w9891 & w19983;
assign w22432 = w10419 & w19980;
assign v7089 = ~(w22431 | w22432);
assign w22433 = v7089;
assign w22434 = w9401 & w19986;
assign w22435 = w22433 & ~w22434;
assign w22436 = ~w22430 & w22435;
assign v7090 = ~(pi05 | w22436);
assign w22437 = v7090;
assign w22438 = pi05 & w22436;
assign v7091 = ~(w22437 | w22438);
assign w22439 = v7091;
assign w22440 = w22429 & ~w22439;
assign w22441 = w22220 & ~w22222;
assign v7092 = ~(w22223 | w22441);
assign w22442 = v7092;
assign w22443 = w9402 & w20997;
assign w22444 = w10419 & w19983;
assign w22445 = w9401 & w19989;
assign w22446 = w9891 & w19986;
assign v7093 = ~(w22445 | w22446);
assign w22447 = v7093;
assign w22448 = ~w22444 & w22447;
assign w22449 = ~w22443 & w22448;
assign w22450 = ~pi05 & w22449;
assign w22451 = pi05 & ~w22449;
assign v7094 = ~(w22450 | w22451);
assign w22452 = v7094;
assign w22453 = w22442 & w22452;
assign w22454 = w22216 & ~w22218;
assign v7095 = ~(w22219 | w22454);
assign w22455 = v7095;
assign w22456 = w9402 & w21012;
assign w22457 = w9401 & ~w19992;
assign w22458 = w10419 & w19986;
assign v7096 = ~(w22457 | w22458);
assign w22459 = v7096;
assign w22460 = w9891 & w19989;
assign w22461 = w22459 & ~w22460;
assign w22462 = ~w22456 & w22461;
assign v7097 = ~(pi05 | w22462);
assign w22463 = v7097;
assign w22464 = pi05 & w22462;
assign v7098 = ~(w22463 | w22464);
assign w22465 = v7098;
assign w22466 = w22455 & ~w22465;
assign w22467 = w22212 & ~w22214;
assign v7099 = ~(w22215 | w22467);
assign w22468 = v7099;
assign w22469 = w10419 & w19989;
assign w22470 = w9401 & ~w19997;
assign w22471 = w9891 & ~w19992;
assign v7100 = ~(w22470 | w22471);
assign w22472 = v7100;
assign w22473 = ~w22469 & w22472;
assign w22474 = (w20098 & w29806) | (w20098 & w29807) | (w29806 & w29807);
assign w22475 = pi05 & ~w22474;
assign w22476 = ~pi05 & w22474;
assign v7101 = ~(w22475 | w22476);
assign w22477 = v7101;
assign w22478 = w22468 & w22477;
assign w22479 = w22208 & ~w22210;
assign v7102 = ~(w22211 | w22479);
assign w22480 = v7102;
assign w22481 = ~w20096 & w29808;
assign w22482 = w10419 & ~w19992;
assign w22483 = w9891 & ~w19997;
assign w22484 = w9401 & w20000;
assign v7103 = ~(w22483 | w22484);
assign w22485 = v7103;
assign w22486 = ~w22482 & w22485;
assign w22487 = ~w22481 & w22486;
assign w22488 = ~pi05 & w22487;
assign w22489 = pi05 & ~w22487;
assign v7104 = ~(w22488 | w22489);
assign w22490 = v7104;
assign w22491 = w22480 & w22490;
assign w22492 = w22204 & ~w22206;
assign v7105 = ~(w22207 | w22492);
assign w22493 = v7105;
assign w22494 = w10419 & ~w19997;
assign w22495 = w9401 & w20005;
assign w22496 = w9891 & w20000;
assign v7106 = ~(w22495 | w22496);
assign w22497 = v7106;
assign w22498 = ~w22494 & w22497;
assign w22499 = (~w20668 & w29809) | (~w20668 & w29810) | (w29809 & w29810);
assign w22500 = (w20668 & w29811) | (w20668 & w29812) | (w29811 & w29812);
assign v7107 = ~(w22499 | w22500);
assign w22501 = v7107;
assign w22502 = w22493 & w22501;
assign w22503 = (w29414 & w30711) | (w29414 & w30712) | (w30711 & w30712);
assign v7108 = ~(w22203 | w22503);
assign w22504 = v7108;
assign w22505 = w10419 & w20000;
assign w22506 = w9401 & ~w20008;
assign w22507 = w9891 & w20005;
assign v7109 = ~(w22506 | w22507);
assign w22508 = v7109;
assign w22509 = ~w22505 & w22508;
assign w22510 = (w22509 & ~w20681) | (w22509 & w29608) | (~w20681 & w29608);
assign w22511 = pi05 & ~w22510;
assign w22512 = ~pi05 & w22510;
assign v7110 = ~(w22511 | w22512);
assign w22513 = v7110;
assign w22514 = w22504 & w22513;
assign w22515 = w22196 & ~w22198;
assign v7111 = ~(w22199 | w22515);
assign w22516 = v7111;
assign w22517 = w10419 & w20005;
assign w22518 = w9401 & ~w20011;
assign w22519 = w9891 & ~w20008;
assign v7112 = ~(w22518 | w22519);
assign w22520 = v7112;
assign w22521 = ~w22517 & w22520;
assign w22522 = (w29089 & w29813) | (w29089 & w29814) | (w29813 & w29814);
assign w22523 = (w29610 & ~w29089) | (w29610 & w29815) | (~w29089 & w29815);
assign v7113 = ~(w22522 | w22523);
assign w22524 = v7113;
assign w22525 = w22516 & w22524;
assign w22526 = w22192 & ~w22194;
assign v7114 = ~(w22195 | w22526);
assign w22527 = v7114;
assign w22528 = w9891 & ~w20011;
assign w22529 = w10419 & ~w20008;
assign w22530 = w9401 & w20014;
assign w22531 = ~w22529 & w29927;
assign w22532 = (~w29091 & w29928) | (~w29091 & w29929) | (w29928 & w29929);
assign w22533 = (w29091 & w29930) | (w29091 & w29931) | (w29930 & w29931);
assign v7115 = ~(w22532 | w22533);
assign w22534 = v7115;
assign w22535 = w22527 & ~w22534;
assign w22536 = w22188 & ~w22190;
assign v7116 = ~(w22191 | w22536);
assign w22537 = v7116;
assign w22538 = w9891 & w20014;
assign w22539 = w10419 & ~w20011;
assign w22540 = w9401 & ~w20028;
assign w22541 = ~w22539 & w29092;
assign w22542 = (~w20459 & w29093) | (~w20459 & w29094) | (w29093 & w29094);
assign w22543 = (w20459 & w29095) | (w20459 & w29096) | (w29095 & w29096);
assign v7117 = ~(w22542 | w22543);
assign w22544 = v7117;
assign w22545 = w22537 & ~w22544;
assign w22546 = w22184 & ~w22186;
assign v7118 = ~(w22187 | w22546);
assign w22547 = v7118;
assign w22548 = w9402 & w20472;
assign w22549 = w9891 & ~w20028;
assign w22550 = w10419 & w20014;
assign v7119 = ~(w22549 | w22550);
assign w22551 = v7119;
assign w22552 = w9401 & ~w20026;
assign w22553 = ~w22548 & w28370;
assign w22554 = (~pi05 & w22548) | (~pi05 & w28371) | (w22548 & w28371);
assign v7120 = ~(w22553 | w22554);
assign w22555 = v7120;
assign w22556 = w22547 & ~w22555;
assign w22557 = w22180 & ~w22182;
assign v7121 = ~(w22183 | w22557);
assign w22558 = v7121;
assign w22559 = w10419 & ~w20028;
assign w22560 = w9401 & w20031;
assign w22561 = (~w22560 & w20026) | (~w22560 & w29097) | (w20026 & w29097);
assign w22562 = ~w22559 & w22561;
assign w22563 = (~w20431 & w28822) | (~w20431 & w28823) | (w28822 & w28823);
assign w22564 = (w20431 & w28824) | (w20431 & w28825) | (w28824 & w28825);
assign v7122 = ~(w22563 | w22564);
assign w22565 = v7122;
assign w22566 = w22558 & w22565;
assign w22567 = w22176 & ~w22178;
assign v7123 = ~(w22179 | w22567);
assign w22568 = v7123;
assign w22569 = w9401 & ~w20063;
assign w22570 = w10419 & ~w20026;
assign w22571 = (~w22569 & w20026) | (~w22569 & w29098) | (w20026 & w29098);
assign w22572 = w9891 & w20031;
assign w22573 = (~w20311 & w28373) | (~w20311 & w28374) | (w28373 & w28374);
assign w22574 = (w20311 & w28375) | (w20311 & w28376) | (w28375 & w28376);
assign v7124 = ~(w22573 | w22574);
assign w22575 = v7124;
assign w22576 = w22568 & ~w22575;
assign w22577 = ~w22568 & w22575;
assign v7125 = ~(w22576 | w22577);
assign w22578 = v7125;
assign v7126 = ~(w22168 | w22174);
assign w22579 = v7126;
assign v7127 = ~(w22175 | w22579);
assign w22580 = v7127;
assign w22581 = w10419 & w20031;
assign w22582 = w9401 & ~w20038;
assign w22583 = (~w22582 & w20063) | (~w22582 & w29099) | (w20063 & w29099);
assign w22584 = ~w22581 & w22583;
assign w22585 = (w20323 & w28377) | (w20323 & w28378) | (w28377 & w28378);
assign w22586 = (~w20323 & w28379) | (~w20323 & w28380) | (w28379 & w28380);
assign v7128 = ~(w22585 | w22586);
assign w22587 = v7128;
assign v7129 = ~(w22580 | w22587);
assign w22588 = v7129;
assign w22589 = w22580 & w22587;
assign w22590 = ~w22154 & w22156;
assign v7130 = ~(w22157 | w22590);
assign w22591 = v7130;
assign w22592 = w10419 & ~w20038;
assign w22593 = w9401 & w20043;
assign w22594 = w9891 & w20040;
assign v7131 = ~(w22593 | w22594);
assign w22595 = v7131;
assign w22596 = ~w22592 & w22595;
assign w22597 = pi05 & ~w22596;
assign w22598 = ~pi05 & w22596;
assign w22599 = (w22598 & w20294) | (w22598 & w28071) | (w20294 & w28071);
assign w22600 = w10445 & ~w20294;
assign v7132 = ~(w22599 | w22600);
assign w22601 = v7132;
assign w22602 = w22601 & w28210;
assign w22603 = w11394 & w20047;
assign w22604 = w9402 & w20246;
assign w22605 = w10419 & ~w20052;
assign w22606 = w9891 & w20047;
assign v7133 = ~(w22605 | w22606);
assign w22607 = v7133;
assign w22608 = ~w22604 & w22607;
assign w22609 = ~w22603 & w22608;
assign w22610 = pi05 & ~w22609;
assign w22611 = w9402 & w20257;
assign w22612 = w9401 & w20047;
assign v7134 = ~(w22611 | w22612);
assign w22613 = v7134;
assign w22614 = w10419 & w20043;
assign w22615 = w9891 & ~w20052;
assign v7135 = ~(w22614 | w22615);
assign w22616 = v7135;
assign w22617 = w22613 & w22616;
assign w22618 = ~w22610 & w22617;
assign w22619 = pi05 & w22618;
assign v7136 = ~(w22155 | w22619);
assign w22620 = v7136;
assign w22621 = w10419 & w20040;
assign w22622 = w9401 & ~w20052;
assign w22623 = w9891 & w20043;
assign v7137 = ~(w22622 | w22623);
assign w22624 = v7137;
assign w22625 = ~w22621 & w22624;
assign w22626 = (w22625 & w20272) | (w22625 & w29100) | (w20272 & w29100);
assign w22627 = pi05 & w22626;
assign v7138 = ~(pi05 | w22626);
assign w22628 = v7138;
assign v7139 = ~(w22627 | w22628);
assign w22629 = v7139;
assign v7140 = ~(w22620 | w22629);
assign w22630 = v7140;
assign w22631 = (~w22591 & ~w22601) | (~w22591 & w28211) | (~w22601 & w28211);
assign v7141 = ~(w22602 | w22631);
assign w22632 = v7141;
assign w22633 = w22630 & w22632;
assign w22634 = (~w22602 & ~w22632) | (~w22602 & w28567) | (~w22632 & w28567);
assign w22635 = pi08 & ~w22157;
assign v7142 = ~(w22163 | w22635);
assign w22636 = v7142;
assign w22637 = w22163 & w22635;
assign v7143 = ~(w22636 | w22637);
assign w22638 = v7143;
assign w22639 = w10419 & ~w20063;
assign w22640 = w9891 & ~w20038;
assign w22641 = w9401 & w20040;
assign v7144 = ~(w22640 | w22641);
assign w22642 = v7144;
assign w22643 = (w22642 & w20063) | (w22642 & w28826) | (w20063 & w28826);
assign w22644 = (~w20339 & w28381) | (~w20339 & w28382) | (w28381 & w28382);
assign w22645 = (w20339 & w28383) | (w20339 & w28384) | (w28383 & w28384);
assign v7145 = ~(w22644 | w22645);
assign w22646 = v7145;
assign w22647 = w22638 & w22646;
assign v7146 = ~(w22638 | w22646);
assign w22648 = v7146;
assign v7147 = ~(w22647 | w22648);
assign w22649 = v7147;
assign v7148 = ~(w22634 | w22649);
assign w22650 = v7148;
assign w22651 = ~w22638 & w22646;
assign w22652 = (~w22651 & w22649) | (~w22651 & w28827) | (w22649 & w28827);
assign w22653 = ~w22589 & w22652;
assign v7149 = ~(w22588 | w22653);
assign w22654 = v7149;
assign w22655 = w22578 & w22654;
assign w22656 = (~w22576 & ~w22578) | (~w22576 & w28212) | (~w22578 & w28212);
assign v7150 = ~(w22558 | w22565);
assign w22657 = v7150;
assign v7151 = ~(w22566 | w22657);
assign w22658 = v7151;
assign w22659 = ~w22656 & w22658;
assign w22660 = (~w22566 & ~w22658) | (~w22566 & w28213) | (~w22658 & w28213);
assign w22661 = ~w22547 & w22555;
assign v7152 = ~(w22556 | w22661);
assign w22662 = v7152;
assign w22663 = ~w22660 & w22662;
assign w22664 = (~w22556 & ~w22662) | (~w22556 & w28828) | (~w22662 & w28828);
assign w22665 = ~w22537 & w22544;
assign v7153 = ~(w22545 | w22665);
assign w22666 = v7153;
assign w22667 = ~w22664 & w22666;
assign w22668 = (~w22545 & w22664) | (~w22545 & w29816) | (w22664 & w29816);
assign w22669 = ~w22527 & w22534;
assign v7154 = ~(w22535 | w22669);
assign w22670 = v7154;
assign w22671 = ~w22668 & w22670;
assign w22672 = (~w22535 & ~w22670) | (~w22535 & w28214) | (~w22670 & w28214);
assign v7155 = ~(w22516 | w22524);
assign w22673 = v7155;
assign v7156 = ~(w22525 | w22673);
assign w22674 = v7156;
assign w22675 = ~w22672 & w22674;
assign w22676 = (~w22525 & w22672) | (~w22525 & w29611) | (w22672 & w29611);
assign v7157 = ~(w22504 | w22513);
assign w22677 = v7157;
assign v7158 = ~(w22514 | w22677);
assign w22678 = v7158;
assign w22679 = ~w22676 & w22678;
assign w22680 = (~w22514 & w22676) | (~w22514 & w29932) | (w22676 & w29932);
assign v7159 = ~(w22493 | w22501);
assign w22681 = v7159;
assign v7160 = ~(w22502 | w22681);
assign w22682 = v7160;
assign w22683 = ~w22680 & w22682;
assign w22684 = (~w22502 & w22680) | (~w22502 & w29101) | (w22680 & w29101);
assign v7161 = ~(w22480 | w22490);
assign w22685 = v7161;
assign v7162 = ~(w22491 | w22685);
assign w22686 = v7162;
assign w22687 = ~w22684 & w22686;
assign w22688 = (~w22491 & ~w22686) | (~w22491 & w28215) | (~w22686 & w28215);
assign v7163 = ~(w22468 | w22477);
assign w22689 = v7163;
assign v7164 = ~(w22478 | w22689);
assign w22690 = v7164;
assign w22691 = ~w22688 & w22690;
assign w22692 = (~w22478 & w22688) | (~w22478 & w29416) | (w22688 & w29416);
assign w22693 = ~w22455 & w22465;
assign v7165 = ~(w22466 | w22693);
assign w22694 = v7165;
assign w22695 = ~w22692 & w22694;
assign w22696 = (~w22466 & w22692) | (~w22466 & w30087) | (w22692 & w30087);
assign v7166 = ~(w22442 | w22452);
assign w22697 = v7166;
assign v7167 = ~(w22453 | w22697);
assign w22698 = v7167;
assign w22699 = ~w22696 & w22698;
assign w22700 = (~w22453 & w22696) | (~w22453 & w29933) | (w22696 & w29933);
assign w22701 = ~w22429 & w22439;
assign v7168 = ~(w22440 | w22701);
assign w22702 = v7168;
assign w22703 = ~w22700 & w22702;
assign w22704 = (~w22440 & w22700) | (~w22440 & w30713) | (w22700 & w30713);
assign w22705 = ~w22416 & w22426;
assign v7169 = ~(w22427 | w22705);
assign w22706 = v7169;
assign w22707 = ~w22704 & w22706;
assign w22708 = (~w22427 & ~w22706) | (~w22427 & w28216) | (~w22706 & w28216);
assign w22709 = ~w22403 & w22413;
assign v7170 = ~(w22414 | w22709);
assign w22710 = v7170;
assign w22711 = ~w22708 & w22710;
assign w22712 = (~w22414 & w22708) | (~w22414 & w30274) | (w22708 & w30274);
assign w22713 = ~w22390 & w22400;
assign v7171 = ~(w22401 | w22713);
assign w22714 = v7171;
assign w22715 = ~w22712 & w22714;
assign w22716 = (~w22401 & w22712) | (~w22401 & w30437) | (w22712 & w30437);
assign w22717 = w22377 & w22387;
assign v7172 = ~(w22388 | w22717);
assign w22718 = v7172;
assign w22719 = ~w22716 & w22718;
assign w22720 = (~w22388 & w22716) | (~w22388 & w30714) | (w22716 & w30714);
assign w22721 = ~w22364 & w22374;
assign v7173 = ~(w22375 | w22721);
assign w22722 = v7173;
assign w22723 = ~w22720 & w22722;
assign w22724 = (~w22375 & w22720) | (~w22375 & w31103) | (w22720 & w31103);
assign w22725 = ~w22357 & w22361;
assign v7174 = ~(w22362 | w22725);
assign w22726 = v7174;
assign w22727 = ~w22724 & w22726;
assign w22728 = (~w22362 & w22724) | (~w22362 & w30570) | (w22724 & w30570);
assign w22729 = (~w22346 & ~w22728) | (~w22346 & w28829) | (~w22728 & w28829);
assign w22730 = w22333 & w22729;
assign w22731 = (~w22331 & ~w22333) | (~w22331 & w28830) | (~w22333 & w28830);
assign w22732 = (~w22315 & ~w22731) | (~w22315 & w30896) | (~w22731 & w30896);
assign w22733 = w22298 & ~w22732;
assign w22734 = (~w22296 & w22732) | (~w22296 & w31216) | (w22732 & w31216);
assign w22735 = w22277 & w22734;
assign w22736 = (~w22275 & ~w22277) | (~w22275 & w28831) | (~w22277 & w28831);
assign w22737 = (~w21852 & w22255) | (~w21852 & w28385) | (w22255 & w28385);
assign w22738 = (~w21847 & w21706) | (~w21847 & w28832) | (w21706 & w28832);
assign w22739 = w7765 & w19952;
assign w22740 = w7466 & w19958;
assign w22741 = w7177 & w19961;
assign v7175 = ~(w22740 | w22741);
assign w22742 = v7175;
assign w22743 = ~w22739 & w22742;
assign w22744 = ~pi11 & w22743;
assign w22745 = w7178 & ~w21882;
assign w22746 = w22744 & ~w22745;
assign w22747 = w9464 & ~w21882;
assign w22748 = pi11 & ~w22743;
assign v7176 = ~(w22747 | w22748);
assign w22749 = v7176;
assign w22750 = ~w22746 & w22749;
assign w22751 = (~w21838 & ~w21842) | (~w21838 & w28386) | (~w21842 & w28386);
assign w22752 = (~w21822 & w21723) | (~w21822 & w30897) | (w21723 & w30897);
assign v7177 = ~(w21806 | w21809);
assign w22753 = v7177;
assign w22754 = (~w21791 & w21725) | (~w21791 & w30088) | (w21725 & w30088);
assign w22755 = (~w21777 & w21726) | (~w21777 & w30275) | (w21726 & w30275);
assign v7178 = ~(w21765 | w21768);
assign w22756 = v7178;
assign v7179 = ~(w21750 | w21753);
assign w22757 = v7179;
assign w22758 = w1641 & w14482;
assign w22759 = ~w465 & w1457;
assign w22760 = ~w49 & w5838;
assign w22761 = w22759 & w22760;
assign w22762 = w766 & w2752;
assign w22763 = w22761 & w22762;
assign w22764 = w207 & w22763;
assign w22765 = w688 & w3722;
assign w22766 = w257 & w22765;
assign v7180 = ~(w131 | w388);
assign w22767 = v7180;
assign w22768 = w22766 & w22767;
assign w22769 = w22764 & w22768;
assign w22770 = w22758 & w22769;
assign w22771 = w3406 & ~w20038;
assign w22772 = w3402 & w20040;
assign w22773 = w3399 & w20043;
assign v7181 = ~(w22772 | w22773);
assign w22774 = v7181;
assign w22775 = ~w22771 & w22774;
assign w22776 = (w22775 & w20294) | (w22775 & w31293) | (w20294 & w31293);
assign v7182 = ~(w22770 | w22776);
assign w22777 = v7182;
assign w22778 = w22770 & w22776;
assign v7183 = ~(w22777 | w22778);
assign w22779 = v7183;
assign w22780 = ~w22757 & w22779;
assign w22781 = w22757 & ~w22779;
assign v7184 = ~(w22780 | w22781);
assign w22782 = v7184;
assign w22783 = (w3529 & w20309) | (w3529 & w30715) | (w20309 & w30715);
assign w22784 = w3767 & ~w20063;
assign w22785 = w3760 & ~w20026;
assign v7185 = ~(w22784 | w22785);
assign w22786 = v7185;
assign w22787 = w3763 & w20031;
assign w22788 = ~w22783 & w31104;
assign w22789 = (~pi29 & w22783) | (~pi29 & w31105) | (w22783 & w31105);
assign v7186 = ~(w22788 | w22789);
assign w22790 = v7186;
assign w22791 = w22782 & ~w22790;
assign w22792 = ~w22782 & w22790;
assign v7187 = ~(w22791 | w22792);
assign w22793 = v7187;
assign w22794 = ~w22756 & w22793;
assign w22795 = w22756 & ~w22793;
assign v7188 = ~(w22794 | w22795);
assign w22796 = v7188;
assign v7189 = ~(w2873 | w20028);
assign w22797 = v7189;
assign w22798 = w4155 & ~w20011;
assign v7190 = ~(w22797 | w22798);
assign w22799 = v7190;
assign w22800 = w4158 & w20014;
assign w22801 = (w20459 & w31106) | (w20459 & w31107) | (w31106 & w31107);
assign w22802 = (~w20459 & w31108) | (~w20459 & w31109) | (w31108 & w31109);
assign v7191 = ~(w22801 | w22802);
assign w22803 = v7191;
assign w22804 = ~w22796 & w22803;
assign w22805 = w22796 & ~w22803;
assign v7192 = ~(w22804 | w22805);
assign w22806 = v7192;
assign w22807 = ~w22755 & w22806;
assign w22808 = w22755 & ~w22806;
assign v7193 = ~(w22807 | w22808);
assign w22809 = v7193;
assign w22810 = w4913 & w20000;
assign w22811 = w4763 & ~w20008;
assign w22812 = w4836 & w20005;
assign v7194 = ~(w22811 | w22812);
assign w22813 = v7194;
assign w22814 = ~w22810 & w22813;
assign w22815 = (~w20681 & w31294) | (~w20681 & w31295) | (w31294 & w31295);
assign w22816 = (w20681 & w31296) | (w20681 & w31297) | (w31296 & w31297);
assign v7195 = ~(w22815 | w22816);
assign w22817 = v7195;
assign w22818 = w22809 & w22817;
assign v7196 = ~(w22809 | w22817);
assign w22819 = v7196;
assign v7197 = ~(w22818 | w22819);
assign w22820 = v7197;
assign w22821 = ~w22754 & w22820;
assign w22822 = w22754 & ~w22820;
assign v7198 = ~(w22821 | w22822);
assign w22823 = v7198;
assign w22824 = w5114 & w20965;
assign w22825 = w5610 & w19989;
assign w22826 = w5113 & ~w19997;
assign w22827 = w5531 & ~w19992;
assign v7199 = ~(w22826 | w22827);
assign w22828 = v7199;
assign w22829 = ~w22825 & w22828;
assign w22830 = ~w22824 & w22829;
assign w22831 = ~pi20 & w22830;
assign w22832 = pi20 & ~w22830;
assign v7200 = ~(w22831 | w22832);
assign w22833 = v7200;
assign w22834 = w22823 & w22833;
assign v7201 = ~(w22823 | w22833);
assign w22835 = v7201;
assign v7202 = ~(w22834 | w22835);
assign w22836 = v7202;
assign w22837 = ~w22753 & w22836;
assign w22838 = w22753 & ~w22836;
assign v7203 = ~(w22837 | w22838);
assign w22839 = v7203;
assign w22840 = w5765 & w20982;
assign w22841 = w5983 & w19983;
assign w22842 = w6236 & w19980;
assign v7204 = ~(w22841 | w22842);
assign w22843 = v7204;
assign w22844 = w5764 & w19986;
assign w22845 = w22843 & ~w22844;
assign w22846 = ~w22840 & w22845;
assign w22847 = pi17 & w22846;
assign v7205 = ~(pi17 | w22846);
assign w22848 = v7205;
assign v7206 = ~(w22847 | w22848);
assign w22849 = v7206;
assign w22850 = w22839 & ~w22849;
assign w22851 = ~w22839 & w22849;
assign v7207 = ~(w22850 | w22851);
assign w22852 = v7207;
assign w22853 = w22752 & ~w22852;
assign w22854 = ~w22752 & w22852;
assign v7208 = ~(w22853 | w22854);
assign w22855 = v7208;
assign w22856 = w6389 & w21385;
assign w22857 = w7004 & w19966;
assign w22858 = w6871 & ~w19971;
assign w22859 = w6388 & w19974;
assign v7209 = ~(w22858 | w22859);
assign w22860 = v7209;
assign w22861 = ~w22857 & w22860;
assign w22862 = ~w22856 & w22861;
assign w22863 = pi14 & ~w22862;
assign w22864 = ~pi14 & w22862;
assign v7210 = ~(w22863 | w22864);
assign w22865 = v7210;
assign w22866 = w22855 & w22865;
assign v7211 = ~(w22855 | w22865);
assign w22867 = v7211;
assign v7212 = ~(w22866 | w22867);
assign w22868 = v7212;
assign w22869 = w22751 & ~w22868;
assign w22870 = ~w22751 & w22868;
assign v7213 = ~(w22869 | w22870);
assign w22871 = v7213;
assign v7214 = ~(w22750 | w22871);
assign w22872 = v7214;
assign w22873 = w22750 & w22871;
assign v7215 = ~(w22872 | w22873);
assign w22874 = v7215;
assign w22875 = w8926 & w19933;
assign w22876 = w8140 & w19954;
assign w22877 = w8526 & ~w19939;
assign v7216 = ~(w22876 | w22877);
assign w22878 = v7216;
assign w22879 = ~w22875 & w22878;
assign w22880 = (~w22304 & w28387) | (~w22304 & w28388) | (w28387 & w28388);
assign w22881 = (w22304 & w28389) | (w22304 & w28390) | (w28389 & w28390);
assign v7217 = ~(w22880 | w22881);
assign w22882 = v7217;
assign v7218 = ~(w22874 | w22882);
assign w22883 = v7218;
assign w22884 = w22874 & w22882;
assign v7219 = ~(w22883 | w22884);
assign w22885 = v7219;
assign w22886 = ~w22738 & w22885;
assign w22887 = w22738 & ~w22885;
assign v7220 = ~(w22886 | w22887);
assign w22888 = v7220;
assign w22889 = ~w22737 & w22888;
assign w22890 = w22737 & ~w22888;
assign v7221 = ~(w22889 | w22890);
assign w22891 = v7221;
assign v7222 = ~(w19924 | w19925);
assign w22892 = v7222;
assign w22893 = w20141 & w22892;
assign v7223 = ~(w20141 | w22892);
assign w22894 = v7223;
assign v7224 = ~(w22893 | w22894);
assign w22895 = v7224;
assign w22896 = w10445 & ~w22895;
assign w22897 = w10419 & w19917;
assign w22898 = w9401 & ~w19929;
assign w22899 = w9891 & ~w19923;
assign v7225 = ~(w22898 | w22899);
assign w22900 = v7225;
assign w22901 = ~w22897 & w22900;
assign w22902 = pi05 & ~w22901;
assign w22903 = ~pi05 & w22901;
assign w22904 = (w22903 & w22895) | (w22903 & w28391) | (w22895 & w28391);
assign v7226 = ~(w22902 | w22904);
assign w22905 = v7226;
assign w22906 = ~w22896 & w22905;
assign w22907 = w22891 & w22906;
assign v7227 = ~(w22891 | w22906);
assign w22908 = v7227;
assign v7228 = ~(w22907 | w22908);
assign w22909 = v7228;
assign w22910 = w22736 & ~w22909;
assign w22911 = ~w22736 & w22909;
assign v7229 = ~(w22910 | w22911);
assign w22912 = v7229;
assign w22913 = ~w20212 & w22912;
assign w22914 = w20212 & ~w22912;
assign v7230 = ~(w22913 | w22914);
assign w22915 = v7230;
assign w22916 = ~w19915 & w20145;
assign v7231 = ~(w20146 | w22916);
assign w22917 = v7231;
assign w22918 = w11035 & ~w19912;
assign w22919 = w11023 & w19853;
assign v7232 = ~(w22918 | w22919);
assign w22920 = v7232;
assign w22921 = (w22920 & ~w22917) | (w22920 & w28219) | (~w22917 & w28219);
assign v7233 = ~(pi02 | w22921);
assign w22922 = v7233;
assign w22923 = w10986 & w19917;
assign w22924 = pi02 & ~w22923;
assign w22925 = w22921 & w22924;
assign v7234 = ~(w22922 | w22925);
assign w22926 = v7234;
assign v7235 = ~(w22277 | w22734);
assign w22927 = v7235;
assign v7236 = ~(w22735 | w22927);
assign w22928 = v7236;
assign w22929 = ~w22926 & w22928;
assign w22930 = w22926 & ~w22928;
assign w22931 = ~w22298 & w22732;
assign v7237 = ~(w22733 | w22931);
assign w22932 = v7237;
assign v7238 = ~(w19918 | w19919);
assign w22933 = v7238;
assign w22934 = w20143 & ~w22933;
assign w22935 = ~w20143 & w22933;
assign v7239 = ~(w22934 | w22935);
assign w22936 = v7239;
assign w22937 = w11035 & w19853;
assign w22938 = w11023 & w19917;
assign v7240 = ~(w22937 | w22938);
assign w22939 = v7240;
assign w22940 = (w22939 & ~w22936) | (w22939 & w28072) | (~w22936 & w28072);
assign w22941 = w10986 & ~w19923;
assign w22942 = pi02 & ~w22941;
assign w22943 = w22940 & ~w22942;
assign w22944 = pi02 & ~w22940;
assign v7241 = ~(w22943 | w22944);
assign w22945 = v7241;
assign w22946 = ~w22932 & w22945;
assign v7242 = ~(w4 | w22895);
assign w22947 = v7242;
assign w22948 = w11035 & w19917;
assign w22949 = w11023 & ~w19923;
assign v7243 = ~(w22948 | w22949);
assign w22950 = v7243;
assign w22951 = ~w22947 & w22950;
assign v7244 = ~(pi02 | w22951);
assign w22952 = v7244;
assign w22953 = w10986 & ~w19929;
assign w22954 = pi02 & ~w22953;
assign w22955 = w22951 & w22954;
assign v7245 = ~(w22952 | w22955);
assign w22956 = v7245;
assign v7246 = ~(w22315 | w22316);
assign w22957 = v7246;
assign w22958 = w22731 & w22957;
assign v7247 = ~(w22731 | w22957);
assign w22959 = v7247;
assign v7248 = ~(w22958 | w22959);
assign w22960 = v7248;
assign v7249 = ~(w22956 | w22960);
assign w22961 = v7249;
assign v7250 = ~(w22333 | w22729);
assign w22962 = v7250;
assign v7251 = ~(w22730 | w22962);
assign w22963 = v7251;
assign w22964 = ~w4 & w22262;
assign w22965 = w11023 & ~w19929;
assign w22966 = w11035 & ~w19923;
assign v7252 = ~(w22965 | w22966);
assign w22967 = v7252;
assign w22968 = ~w22964 & w22967;
assign v7253 = ~(pi02 | w22968);
assign w22969 = v7253;
assign w22970 = w10986 & w19933;
assign w22971 = pi02 & ~w22970;
assign w22972 = w22968 & w22971;
assign v7254 = ~(w22969 | w22972);
assign w22973 = v7254;
assign w22974 = w22963 & ~w22973;
assign w22975 = ~w22963 & w22973;
assign v7255 = ~(w22346 | w22347);
assign w22976 = v7255;
assign v7256 = ~(w22728 | w22976);
assign w22977 = v7256;
assign w22978 = w22728 & w22976;
assign v7257 = ~(w22977 | w22978);
assign w22979 = v7257;
assign v7258 = ~(w4 | w22285);
assign w22980 = v7258;
assign w22981 = w11035 & ~w19929;
assign w22982 = w11023 & w19933;
assign v7259 = ~(w22981 | w22982);
assign w22983 = v7259;
assign w22984 = ~w22980 & w22983;
assign v7260 = ~(pi02 | w22984);
assign w22985 = v7260;
assign w22986 = w10986 & ~w19939;
assign w22987 = pi02 & ~w22986;
assign w22988 = w22984 & w22987;
assign v7261 = ~(w22985 | w22988);
assign w22989 = v7261;
assign v7262 = ~(w22979 | w22989);
assign w22990 = v7262;
assign w22991 = w22979 & w22989;
assign v7263 = ~(w4 | w22304);
assign w22992 = v7263;
assign w22993 = w11023 & ~w19939;
assign w22994 = w11035 & w19933;
assign v7264 = ~(w22993 | w22994);
assign w22995 = v7264;
assign w22996 = ~w22992 & w22995;
assign v7265 = ~(pi02 | w22996);
assign w22997 = v7265;
assign w22998 = w10986 & w19954;
assign w22999 = pi02 & ~w22998;
assign w23000 = w22996 & w22999;
assign v7266 = ~(w22997 | w23000);
assign w23001 = v7266;
assign w23002 = w22724 & ~w22726;
assign v7267 = ~(w22727 | w23002);
assign w23003 = v7267;
assign w23004 = ~w23001 & w23003;
assign w23005 = w23001 & ~w23003;
assign w23006 = ~w4 & w20214;
assign w23007 = w11035 & ~w19939;
assign w23008 = w11023 & w19954;
assign v7268 = ~(w23007 | w23008);
assign w23009 = v7268;
assign w23010 = ~w23006 & w23009;
assign v7269 = ~(pi02 | w23010);
assign w23011 = v7269;
assign w23012 = w10986 & w19952;
assign w23013 = pi02 & ~w23012;
assign w23014 = w23010 & w23013;
assign v7270 = ~(w23011 | w23014);
assign w23015 = v7270;
assign w23016 = w22720 & ~w22722;
assign v7271 = ~(w22723 | w23016);
assign w23017 = v7271;
assign w23018 = ~w23015 & w23017;
assign w23019 = w23015 & ~w23017;
assign w23020 = w1 & ~w21866;
assign w23021 = w11023 & w19952;
assign w23022 = w11035 & w19954;
assign v7272 = ~(w23021 | w23022);
assign w23023 = v7272;
assign v7273 = ~(pi02 | w23023);
assign w23024 = v7273;
assign w23025 = w10987 & w19958;
assign w23026 = (~w23025 & ~w21866) | (~w23025 & w28073) | (~w21866 & w28073);
assign w23027 = ~w10988 & w23023;
assign w23028 = w23026 & w23027;
assign v7274 = ~(w23024 | w23028);
assign w23029 = v7274;
assign v7275 = ~(w23020 | w23029);
assign w23030 = v7275;
assign w23031 = w22716 & ~w22718;
assign v7276 = ~(w22719 | w23031);
assign w23032 = v7276;
assign w23033 = w23030 & w23032;
assign w23034 = w22712 & ~w22714;
assign v7277 = ~(w22715 | w23034);
assign w23035 = v7277;
assign w23036 = w22708 & ~w22710;
assign v7278 = ~(w22711 | w23036);
assign w23037 = v7278;
assign w23038 = w22704 & ~w22706;
assign v7279 = ~(w22707 | w23038);
assign w23039 = v7279;
assign w23040 = w1 & w21385;
assign w23041 = w11023 & ~w19971;
assign w23042 = w11035 & w19966;
assign v7280 = ~(w23041 | w23042);
assign w23043 = v7280;
assign v7281 = ~(pi02 | w23043);
assign w23044 = v7281;
assign v7282 = ~(pi02 | w21385);
assign w23045 = v7282;
assign w23046 = w10987 & w19974;
assign w23047 = w23043 & ~w23046;
assign w23048 = ~w10988 & w23047;
assign w23049 = (~w23044 & w23045) | (~w23044 & w28074) | (w23045 & w28074);
assign v7283 = ~(w23040 | w23049);
assign w23050 = v7283;
assign w23051 = w22700 & ~w22702;
assign v7284 = ~(w22703 | w23051);
assign w23052 = v7284;
assign w23053 = w23050 & w23052;
assign v7285 = ~(w23050 | w23052);
assign w23054 = v7285;
assign w23055 = w3 & w21401;
assign w23056 = w1 & w21401;
assign w23057 = w10987 & w19980;
assign w23058 = w11023 & w19974;
assign w23059 = (~w23058 & w19971) | (~w23058 & w28075) | (w19971 & w28075);
assign w23060 = pi02 & w23059;
assign v7286 = ~(pi02 | w23059);
assign w23061 = v7286;
assign v7287 = ~(w23060 | w23061);
assign w23062 = v7287;
assign v7288 = ~(w23057 | w23062);
assign w23063 = v7288;
assign w23064 = ~w23056 & w23063;
assign v7289 = ~(w23055 | w23064);
assign w23065 = v7289;
assign w23066 = w22696 & ~w22698;
assign v7290 = ~(w22699 | w23066);
assign w23067 = v7290;
assign w23068 = w23065 & ~w23067;
assign w23069 = w11023 & w19980;
assign w23070 = w11035 & w19974;
assign v7291 = ~(w23069 | w23070);
assign w23071 = v7291;
assign w23072 = pi02 & ~w23071;
assign w23073 = w1 & w21362;
assign w23074 = w10987 & w19983;
assign v7292 = ~(w23073 | w23074);
assign w23075 = v7292;
assign w23076 = ~w23072 & w23075;
assign w23077 = w3 & w21362;
assign w23078 = w23071 & ~w23077;
assign w23079 = ~pi02 & w23078;
assign w23080 = w23076 & ~w23079;
assign w23081 = w22692 & ~w22694;
assign v7293 = ~(w22695 | w23081);
assign w23082 = v7293;
assign v7294 = ~(w23080 | w23082);
assign w23083 = v7294;
assign w23084 = w22688 & ~w22690;
assign v7295 = ~(w22691 | w23084);
assign w23085 = v7295;
assign w23086 = ~w4 & w20982;
assign w23087 = w11035 & w19980;
assign w23088 = w11023 & w19983;
assign v7296 = ~(w23087 | w23088);
assign w23089 = v7296;
assign w23090 = ~w23086 & w23089;
assign w23091 = pi02 & ~w23090;
assign w23092 = w10986 & w19986;
assign w23093 = pi02 & ~w23092;
assign w23094 = w23090 & ~w23093;
assign v7297 = ~(w23091 | w23094);
assign w23095 = v7297;
assign w23096 = w23085 & w23095;
assign w23097 = w22684 & ~w22686;
assign v7298 = ~(w22687 | w23097);
assign w23098 = v7298;
assign w23099 = ~w4 & w20997;
assign w23100 = w11035 & w19983;
assign w23101 = w11023 & w19986;
assign v7299 = ~(w23100 | w23101);
assign w23102 = v7299;
assign w23103 = ~w23099 & w23102;
assign v7300 = ~(pi02 | w23103);
assign w23104 = v7300;
assign w23105 = w10986 & w19989;
assign w23106 = pi02 & ~w23105;
assign w23107 = w23103 & w23106;
assign v7301 = ~(w23104 | w23107);
assign w23108 = v7301;
assign w23109 = w23098 & ~w23108;
assign w23110 = ~w23098 & w23108;
assign w23111 = w22680 & ~w22682;
assign v7302 = ~(w22683 | w23111);
assign w23112 = v7302;
assign w23113 = w11035 & w19986;
assign w23114 = w11023 & w19989;
assign v7303 = ~(w23113 | w23114);
assign w23115 = v7303;
assign w23116 = (w23115 & ~w21012) | (w23115 & w29817) | (~w21012 & w29817);
assign v7304 = ~(pi02 | w23116);
assign w23117 = v7304;
assign w23118 = w10986 & ~w19992;
assign w23119 = pi02 & ~w23118;
assign w23120 = w23116 & w23119;
assign v7305 = ~(w23117 | w23120);
assign w23121 = v7305;
assign w23122 = ~w23112 & w23121;
assign w23123 = w23112 & ~w23121;
assign w23124 = w1 & w20965;
assign w23125 = w11035 & w19989;
assign w23126 = w11023 & ~w19992;
assign v7306 = ~(w23125 | w23126);
assign w23127 = v7306;
assign v7307 = ~(pi02 | w23127);
assign w23128 = v7307;
assign w23129 = w10987 & ~w19997;
assign w23130 = ~w10988 & w23127;
assign w23131 = ~w23129 & w23130;
assign w23132 = (~w20965 & w29818) | (~w20965 & w29819) | (w29818 & w29819);
assign v7308 = ~(w23124 | w23132);
assign w23133 = v7308;
assign w23134 = w22676 & ~w22678;
assign v7309 = ~(w22679 | w23134);
assign w23135 = v7309;
assign v7310 = ~(w23133 | w23135);
assign w23136 = v7310;
assign w23137 = w23133 & w23135;
assign w23138 = w3 & w20655;
assign w23139 = ~w20096 & w29613;
assign w23140 = w10987 & w20000;
assign w23141 = w11035 & ~w19992;
assign w23142 = w11023 & ~w19997;
assign v7311 = ~(w23141 | w23142);
assign w23143 = v7311;
assign w23144 = pi02 & w23143;
assign v7312 = ~(pi02 | w23143);
assign w23145 = v7312;
assign v7313 = ~(w23144 | w23145);
assign w23146 = v7313;
assign v7314 = ~(w23140 | w23146);
assign w23147 = v7314;
assign w23148 = ~w23139 & w23147;
assign v7315 = ~(w23138 | w23148);
assign w23149 = v7315;
assign w23150 = w22672 & ~w22674;
assign v7316 = ~(w22675 | w23150);
assign w23151 = v7316;
assign w23152 = w23149 & ~w23151;
assign w23153 = ~w23149 & w23151;
assign w23154 = w11023 & w20000;
assign w23155 = w11035 & ~w19997;
assign v7317 = ~(w23154 | w23155);
assign w23156 = v7317;
assign w23157 = pi02 & ~w23156;
assign w23158 = (~w23157 & ~w20668) | (~w23157 & w29614) | (~w20668 & w29614);
assign w23159 = w10987 & w20005;
assign v7318 = ~(w10988 | w23159);
assign w23160 = v7318;
assign w23161 = (~w20668 & w29615) | (~w20668 & w29616) | (w29615 & w29616);
assign w23162 = w23158 & ~w23161;
assign w23163 = w22668 & ~w22670;
assign v7319 = ~(w22671 | w23163);
assign w23164 = v7319;
assign w23165 = w23162 & w23164;
assign v7320 = ~(w23162 | w23164);
assign w23166 = v7320;
assign w23167 = w22664 & ~w22666;
assign v7321 = ~(w22667 | w23167);
assign w23168 = v7321;
assign w23169 = w11035 & w20000;
assign w23170 = w11023 & w20005;
assign v7322 = ~(w23169 | w23170);
assign w23171 = v7322;
assign w23172 = (w20681 & w29418) | (w20681 & w29419) | (w29418 & w29419);
assign w23173 = w10986 & ~w20008;
assign w23174 = pi02 & ~w23173;
assign w23175 = (~w20681 & w29420) | (~w20681 & w29421) | (w29420 & w29421);
assign v7323 = ~(w23172 | w23175);
assign w23176 = v7323;
assign w23177 = ~w23168 & w23176;
assign w23178 = w23168 & ~w23176;
assign w23179 = w22660 & ~w22662;
assign v7324 = ~(w22663 | w23179);
assign w23180 = v7324;
assign w23181 = w11035 & w20005;
assign w23182 = w11023 & ~w20008;
assign v7325 = ~(w23181 | w23182);
assign w23183 = v7325;
assign w23184 = (~w29104 & w29820) | (~w29104 & w29821) | (w29820 & w29821);
assign w23185 = w10986 & ~w20011;
assign w23186 = pi02 & ~w23185;
assign w23187 = (w29104 & w29822) | (w29104 & w29823) | (w29822 & w29823);
assign v7326 = ~(w23184 | w23187);
assign w23188 = v7326;
assign w23189 = ~w23180 & w23188;
assign w23190 = w23180 & ~w23188;
assign w23191 = w22656 & ~w22658;
assign v7327 = ~(w22659 | w23191);
assign w23192 = v7327;
assign w23193 = w11035 & ~w20008;
assign w23194 = w11023 & ~w20011;
assign v7328 = ~(w23193 | w23194);
assign w23195 = v7328;
assign w23196 = (w20082 & w29105) | (w20082 & w29106) | (w29105 & w29106);
assign v7329 = ~(pi02 | w23196);
assign w23197 = v7329;
assign w23198 = w10986 & w20014;
assign w23199 = pi02 & ~w23198;
assign w23200 = w23196 & w23199;
assign v7330 = ~(w23197 | w23200);
assign w23201 = v7330;
assign w23202 = ~w23192 & w23201;
assign w23203 = w3 & w20459;
assign w23204 = w1 & w20459;
assign w23205 = w10987 & ~w20028;
assign w23206 = w11023 & w20014;
assign w23207 = w11035 & ~w20011;
assign w23208 = ~w23207 & w28835;
assign w23209 = (~pi02 & w23207) | (~pi02 & w28836) | (w23207 & w28836);
assign v7331 = ~(w23208 | w23209);
assign w23210 = v7331;
assign v7332 = ~(w23205 | w23210);
assign w23211 = v7332;
assign w23212 = ~w23204 & w23211;
assign v7333 = ~(w23203 | w23212);
assign w23213 = v7333;
assign v7334 = ~(w22578 | w22654);
assign w23214 = v7334;
assign v7335 = ~(w22655 | w23214);
assign w23215 = v7335;
assign w23216 = w23213 & ~w23215;
assign w23217 = w1 & w20472;
assign w23218 = w11023 & ~w20028;
assign w23219 = (~w23218 & ~w20014) | (~w23218 & w29107) | (~w20014 & w29107);
assign v7336 = ~(pi02 | w23219);
assign w23220 = v7336;
assign v7337 = ~(pi02 | w20472);
assign w23221 = v7337;
assign w23222 = w10987 & ~w20026;
assign w23223 = ~w10988 & w23219;
assign w23224 = ~w23222 & w23223;
assign w23225 = (~w23220 & w23221) | (~w23220 & w29108) | (w23221 & w29108);
assign v7338 = ~(w23217 | w23225);
assign w23226 = v7338;
assign v7339 = ~(w22588 | w22589);
assign w23227 = v7339;
assign w23228 = w22652 & w23227;
assign v7340 = ~(w22652 | w23227);
assign w23229 = v7340;
assign v7341 = ~(w23228 | w23229);
assign w23230 = v7341;
assign w23231 = ~w23226 & w23230;
assign w23232 = w22634 & w22649;
assign v7342 = ~(w22650 | w23232);
assign w23233 = v7342;
assign w23234 = w11023 & ~w20026;
assign w23235 = w11035 & ~w20028;
assign v7343 = ~(w23234 | w23235);
assign w23236 = v7343;
assign w23237 = (w20431 & w29109) | (w20431 & w29110) | (w29109 & w29110);
assign w23238 = w10986 & w20031;
assign w23239 = pi02 & ~w23238;
assign w23240 = (~w20431 & w29111) | (~w20431 & w29112) | (w29111 & w29112);
assign v7344 = ~(w23237 | w23240);
assign w23241 = v7344;
assign w23242 = w23233 & w23241;
assign v7345 = ~(w22630 | w22632);
assign w23243 = v7345;
assign v7346 = ~(w22633 | w23243);
assign w23244 = v7346;
assign w23245 = w11023 & w20031;
assign w23246 = (~w23245 & w20026) | (~w23245 & w29113) | (w20026 & w29113);
assign w23247 = (~w20311 & w29114) | (~w20311 & w29115) | (w29114 & w29115);
assign w23248 = w10986 & ~w20063;
assign w23249 = pi02 & ~w23248;
assign w23250 = (w20311 & w29116) | (w20311 & w29117) | (w29116 & w29117);
assign v7347 = ~(w23247 | w23250);
assign w23251 = v7347;
assign w23252 = w23244 & ~w23251;
assign w23253 = ~w23244 & w23251;
assign w23254 = w22155 & w22619;
assign v7348 = ~(w22620 | w23254);
assign w23255 = v7348;
assign w23256 = w22629 & ~w23255;
assign w23257 = ~w22629 & w23255;
assign v7349 = ~(w23256 | w23257);
assign w23258 = v7349;
assign w23259 = w11023 & ~w20063;
assign w23260 = w11035 & w20031;
assign v7350 = ~(w23259 | w23260);
assign w23261 = v7350;
assign w23262 = pi02 & ~w23261;
assign w23263 = (~w23262 & ~w20323) | (~w23262 & w29118) | (~w20323 & w29118);
assign w23264 = w10987 & ~w20038;
assign v7351 = ~(w10988 | w23264);
assign w23265 = v7351;
assign w23266 = (~w20323 & w29119) | (~w20323 & w29120) | (w29119 & w29120);
assign w23267 = w23263 & ~w23266;
assign w23268 = w22610 & ~w22617;
assign v7352 = ~(w22618 | w23268);
assign w23269 = v7352;
assign w23270 = w11023 & ~w20038;
assign w23271 = (~w23270 & w20063) | (~w23270 & w28838) | (w20063 & w28838);
assign w23272 = (~w20339 & w28839) | (~w20339 & w28840) | (w28839 & w28840);
assign w23273 = w10986 & w20040;
assign w23274 = pi02 & ~w23273;
assign w23275 = (w20339 & w28841) | (w20339 & w28842) | (w28841 & w28842);
assign v7353 = ~(w23272 | w23275);
assign w23276 = v7353;
assign w23277 = ~w23269 & w23276;
assign w23278 = w23269 & ~w23276;
assign v7354 = ~(w4 | w20272);
assign w23279 = v7354;
assign w23280 = w11023 & w20043;
assign w23281 = w11035 & w20040;
assign v7355 = ~(w23280 | w23281);
assign w23282 = v7355;
assign w23283 = ~w23279 & w23282;
assign w23284 = ~w10986 & w20047;
assign w23285 = ~pi00 & w20052;
assign v7356 = ~(w23284 | w23285);
assign w23286 = v7356;
assign v7357 = ~(pi03 | w23286);
assign w23287 = v7357;
assign w23288 = pi00 & w20043;
assign w23289 = w20244 & ~w23288;
assign v7358 = ~(w23287 | w23289);
assign w23290 = v7358;
assign w23291 = pi02 & ~w23290;
assign w23292 = w23283 & ~w23291;
assign w23293 = w19587 & w20047;
assign v7359 = ~(w23283 | w23293);
assign w23294 = v7359;
assign v7360 = ~(w23292 | w23294);
assign w23295 = v7360;
assign w23296 = w22603 & ~w22608;
assign v7361 = ~(w22609 | w23296);
assign w23297 = v7361;
assign w23298 = w11023 & w20040;
assign w23299 = (~w23298 & w20038) | (~w23298 & w28568) | (w20038 & w28568);
assign w23300 = w10986 & w20043;
assign w23301 = w23299 & ~w23300;
assign w23302 = (w20294 & w28569) | (w20294 & w28570) | (w28569 & w28570);
assign v7362 = ~(pi02 | w23299);
assign w23303 = v7362;
assign w23304 = (~w23303 & w20294) | (~w23303 & w28571) | (w20294 & w28571);
assign w23305 = ~w23302 & w23304;
assign w23306 = w23297 & ~w23305;
assign v7363 = ~(w23295 | w23306);
assign w23307 = v7363;
assign w23308 = ~w23297 & w23305;
assign v7364 = ~(w23307 | w23308);
assign w23309 = v7364;
assign v7365 = ~(w23278 | w23309);
assign w23310 = v7365;
assign v7366 = ~(w23277 | w23310);
assign w23311 = v7366;
assign w23312 = (~w23258 & ~w23311) | (~w23258 & w29121) | (~w23311 & w29121);
assign v7367 = ~(w23267 | w23311);
assign w23313 = v7367;
assign v7368 = ~(w23312 | w23313);
assign w23314 = v7368;
assign w23315 = ~w23253 & w23314;
assign v7369 = ~(w23252 | w23315);
assign w23316 = v7369;
assign v7370 = ~(w23233 | w23241);
assign w23317 = v7370;
assign v7371 = ~(w23316 | w23317);
assign w23318 = v7371;
assign v7372 = ~(w23242 | w23318);
assign w23319 = v7372;
assign v7373 = ~(w23231 | w23319);
assign w23320 = v7373;
assign w23321 = w23226 & ~w23230;
assign w23322 = (~w28843 & w29824) | (~w28843 & w29825) | (w29824 & w29825);
assign w23323 = ~w23320 & w23322;
assign v7374 = ~(w23216 | w23323);
assign w23324 = v7374;
assign w23325 = w23192 & ~w23201;
assign w23326 = (~w23202 & w23324) | (~w23202 & w29122) | (w23324 & w29122);
assign w23327 = (~w23189 & w23326) | (~w23189 & w28572) | (w23326 & w28572);
assign w23328 = (~w23177 & w23327) | (~w23177 & w29422) | (w23327 & w29422);
assign w23329 = (~w23165 & ~w23328) | (~w23165 & w29826) | (~w23328 & w29826);
assign w23330 = ~w23153 & w23329;
assign v7375 = ~(w23152 | w23330);
assign w23331 = v7375;
assign w23332 = (~w23136 & w23331) | (~w23136 & w29617) | (w23331 & w29617);
assign w23333 = (~w23122 & w23332) | (~w23122 & w29934) | (w23332 & w29934);
assign w23334 = ~w23110 & w23333;
assign v7376 = ~(w23109 | w23334);
assign w23335 = v7376;
assign v7377 = ~(w23085 | w23095);
assign w23336 = v7377;
assign w23337 = (~w23096 & w23335) | (~w23096 & w29935) | (w23335 & w29935);
assign v7378 = ~(w23083 | w23337);
assign w23338 = v7378;
assign w23339 = w23080 & w23082;
assign w23340 = (~w23339 & ~w23067) | (~w23339 & w29936) | (~w23067 & w29936);
assign w23341 = (~w23068 & ~w23340) | (~w23068 & w28077) | (~w23340 & w28077);
assign w23342 = ~w23054 & w23341;
assign w23343 = (~w23053 & ~w23341) | (~w23053 & w29937) | (~w23341 & w29937);
assign w23344 = w23039 & ~w23343;
assign w23345 = ~w4 & w20234;
assign w23346 = w11035 & w19961;
assign w23347 = w11023 & w19966;
assign v7379 = ~(w23346 | w23347);
assign w23348 = v7379;
assign w23349 = ~w23345 & w23348;
assign w23350 = pi02 & ~w23349;
assign w23351 = w10986 & ~w19971;
assign w23352 = pi02 & ~w23351;
assign w23353 = w23349 & ~w23352;
assign v7380 = ~(w23350 | w23353);
assign w23354 = v7380;
assign w23355 = (w23354 & w23342) | (w23354 & w30716) | (w23342 & w30716);
assign w23356 = ~w4 & w21716;
assign w23357 = w11035 & w19958;
assign w23358 = w11023 & w19961;
assign v7381 = ~(w23357 | w23358);
assign w23359 = v7381;
assign w23360 = ~w23356 & w23359;
assign w23361 = pi02 & ~w23360;
assign w23362 = w10986 & w19966;
assign w23363 = pi02 & ~w23362;
assign w23364 = w23360 & ~w23363;
assign v7382 = ~(w23361 | w23364);
assign w23365 = v7382;
assign w23366 = (w23365 & ~w29938) | (w23365 & w30717) | (~w29938 & w30717);
assign v7383 = ~(w4 | w21882);
assign w23367 = v7383;
assign w23368 = w11035 & w19952;
assign w23369 = w11023 & w19958;
assign v7384 = ~(w23368 | w23369);
assign w23370 = v7384;
assign w23371 = ~w23367 & w23370;
assign w23372 = pi02 & ~w23371;
assign w23373 = w10986 & w19961;
assign w23374 = pi02 & ~w23373;
assign w23375 = w23371 & ~w23374;
assign v7385 = ~(w23372 | w23375);
assign w23376 = v7385;
assign w23377 = (~w23032 & w23029) | (~w23032 & w28079) | (w23029 & w28079);
assign w23378 = ~w23366 & w30438;
assign v7386 = ~(w23377 | w23378);
assign w23379 = v7386;
assign w23380 = (~w30440 & w30720) | (~w30440 & w30721) | (w30720 & w30721);
assign w23381 = (~w23004 & w23380) | (~w23004 & w30722) | (w23380 & w30722);
assign w23382 = (~w22990 & w23381) | (~w22990 & w31111) | (w23381 & w31111);
assign w23383 = (~w22974 & w23382) | (~w22974 & w31298) | (w23382 & w31298);
assign w23384 = ~w22961 & w23383;
assign w23385 = w22956 & w22960;
assign w23386 = w22932 & ~w22945;
assign v7387 = ~(w23385 | w23386);
assign w23387 = v7387;
assign w23388 = (~w22946 & ~w23387) | (~w22946 & w28080) | (~w23387 & w28080);
assign v7388 = ~(w22930 | w23388);
assign w23389 = v7388;
assign v7389 = ~(w22929 | w23389);
assign w23390 = v7389;
assign w23391 = ~w22915 & w23390;
assign w23392 = (~w22908 & ~w22736) | (~w22908 & w28395) | (~w22736 & w28395);
assign w23393 = w10445 & w22936;
assign w23394 = w10447 & w22936;
assign w23395 = w10419 & w19853;
assign w23396 = w9891 & w19917;
assign w23397 = w9401 & ~w19923;
assign v7390 = ~(w23396 | w23397);
assign w23398 = v7390;
assign w23399 = ~w23395 & w23398;
assign w23400 = pi05 & w23399;
assign v7391 = ~(pi05 | w23399);
assign w23401 = v7391;
assign v7392 = ~(w23400 | w23401);
assign w23402 = v7392;
assign w23403 = ~w23394 & w23402;
assign v7393 = ~(w23393 | w23403);
assign w23404 = v7393;
assign w23405 = w22738 & w22874;
assign w23406 = w22882 & ~w23405;
assign w23407 = ~w22886 & w23406;
assign w23408 = w8926 & ~w19929;
assign w23409 = w8140 & ~w19939;
assign w23410 = w8526 & w19933;
assign v7394 = ~(w23409 | w23410);
assign w23411 = v7394;
assign w23412 = ~w23408 & w23411;
assign w23413 = (w23412 & w22285) | (w23412 & w28396) | (w22285 & w28396);
assign w23414 = ~pi08 & w23413;
assign w23415 = pi08 & ~w23413;
assign v7395 = ~(w23414 | w23415);
assign w23416 = v7395;
assign w23417 = (~w22873 & ~w22738) | (~w22873 & w28397) | (~w22738 & w28397);
assign v7396 = ~(w22850 | w22854);
assign w23418 = v7396;
assign w23419 = (~w22834 & w22753) | (~w22834 & w30089) | (w22753 & w30089);
assign w23420 = (~w22818 & w22754) | (~w22818 & w29940) | (w22754 & w29940);
assign w23421 = (~w22805 & w22755) | (~w22805 & w30441) | (w22755 & w30441);
assign v7397 = ~(w22791 | w22794);
assign w23422 = v7397;
assign v7398 = ~(w22777 | w22780);
assign w23423 = v7398;
assign w23424 = w622 & w6044;
assign w23425 = w682 & w23424;
assign w23426 = w4971 & w23425;
assign w23427 = w4255 & w23426;
assign w23428 = w12622 & w23427;
assign w23429 = w726 & w2575;
assign w23430 = w12552 & w23429;
assign w23431 = w1267 & w23430;
assign w23432 = w5187 & w23431;
assign w23433 = w809 & w4609;
assign w23434 = w23432 & w23433;
assign w23435 = w23428 & w23434;
assign w23436 = w928 & ~w20339;
assign w23437 = w3406 & ~w20063;
assign w23438 = w3399 & w20040;
assign w23439 = w3402 & ~w20038;
assign v7399 = ~(w23438 | w23439);
assign w23440 = v7399;
assign w23441 = ~w23437 & w23440;
assign w23442 = ~w23436 & w23441;
assign v7400 = ~(w23435 | w23442);
assign w23443 = v7400;
assign w23444 = w23435 & w23442;
assign v7401 = ~(w23443 | w23444);
assign w23445 = v7401;
assign w23446 = ~w23423 & w23445;
assign w23447 = w23423 & ~w23445;
assign v7402 = ~(w23446 | w23447);
assign w23448 = v7402;
assign w23449 = w3760 & ~w20028;
assign w23450 = w3767 & w20031;
assign w23451 = w3763 & ~w20026;
assign v7403 = ~(w23450 | w23451);
assign w23452 = v7403;
assign w23453 = ~w23449 & w23452;
assign w23454 = (w20431 & w31217) | (w20431 & w31218) | (w31217 & w31218);
assign w23455 = (~w20431 & w31219) | (~w20431 & w31220) | (w31219 & w31220);
assign v7404 = ~(w23454 | w23455);
assign w23456 = v7404;
assign w23457 = w23448 & w23456;
assign v7405 = ~(w23448 | w23456);
assign w23458 = v7405;
assign v7406 = ~(w23457 | w23458);
assign w23459 = v7406;
assign w23460 = ~w23422 & w23459;
assign w23461 = w23422 & ~w23459;
assign v7407 = ~(w23460 | w23461);
assign w23462 = v7407;
assign w23463 = w4158 & ~w20011;
assign w23464 = w4155 & ~w20008;
assign v7408 = ~(w23463 | w23464);
assign w23465 = v7408;
assign w23466 = ~w2873 & w20014;
assign w23467 = w23465 & ~w23466;
assign w23468 = (w23467 & ~w20446) | (w23467 & w30723) | (~w20446 & w30723);
assign w23469 = pi26 & w23468;
assign v7409 = ~(pi26 | w23468);
assign w23470 = v7409;
assign v7410 = ~(w23469 | w23470);
assign w23471 = v7410;
assign w23472 = w23462 & ~w23471;
assign w23473 = ~w23462 & w23471;
assign v7411 = ~(w23472 | w23473);
assign w23474 = v7411;
assign w23475 = ~w23421 & w23474;
assign w23476 = w23421 & ~w23474;
assign v7412 = ~(w23475 | w23476);
assign w23477 = v7412;
assign w23478 = w4913 & ~w19997;
assign w23479 = w4763 & w20005;
assign w23480 = w4836 & w20000;
assign v7413 = ~(w23479 | w23480);
assign w23481 = v7413;
assign w23482 = ~w23478 & w23481;
assign w23483 = (w23482 & ~w20668) | (w23482 & w30724) | (~w20668 & w30724);
assign w23484 = ~pi23 & w23483;
assign w23485 = pi23 & ~w23483;
assign v7414 = ~(w23484 | w23485);
assign w23486 = v7414;
assign w23487 = w23477 & w23486;
assign v7415 = ~(w23477 | w23486);
assign w23488 = v7415;
assign v7416 = ~(w23487 | w23488);
assign w23489 = v7416;
assign w23490 = ~w23420 & w23489;
assign w23491 = w23420 & ~w23489;
assign v7417 = ~(w23490 | w23491);
assign w23492 = v7417;
assign w23493 = w5114 & w21012;
assign w23494 = w5610 & w19986;
assign w23495 = w5113 & ~w19992;
assign w23496 = w5531 & w19989;
assign v7418 = ~(w23495 | w23496);
assign w23497 = v7418;
assign w23498 = ~w23494 & w23497;
assign w23499 = ~w23493 & w23498;
assign w23500 = ~pi20 & w23499;
assign w23501 = pi20 & ~w23499;
assign v7419 = ~(w23500 | w23501);
assign w23502 = v7419;
assign w23503 = w23492 & w23502;
assign v7420 = ~(w23492 | w23502);
assign w23504 = v7420;
assign v7421 = ~(w23503 | w23504);
assign w23505 = v7421;
assign w23506 = w23419 & ~w23505;
assign w23507 = ~w23419 & w23505;
assign v7422 = ~(w23506 | w23507);
assign w23508 = v7422;
assign w23509 = w5765 & w21362;
assign w23510 = w6236 & w19974;
assign w23511 = w5983 & w19980;
assign w23512 = w5764 & w19983;
assign v7423 = ~(w23511 | w23512);
assign w23513 = v7423;
assign w23514 = ~w23510 & w23513;
assign w23515 = ~w23509 & w23514;
assign w23516 = pi17 & w23515;
assign v7424 = ~(pi17 | w23515);
assign w23517 = v7424;
assign v7425 = ~(w23516 | w23517);
assign w23518 = v7425;
assign w23519 = w23508 & ~w23518;
assign w23520 = ~w23508 & w23518;
assign v7426 = ~(w23519 | w23520);
assign w23521 = v7426;
assign w23522 = w23418 & ~w23521;
assign w23523 = ~w23418 & w23521;
assign v7427 = ~(w23522 | w23523);
assign w23524 = v7427;
assign w23525 = w7004 & w19961;
assign w23526 = w6871 & w19966;
assign w23527 = w6388 & ~w19971;
assign v7428 = ~(w23526 | w23527);
assign w23528 = v7428;
assign w23529 = ~w23525 & w23528;
assign w23530 = pi14 & ~w23529;
assign w23531 = w17118 & w20234;
assign v7429 = ~(w23530 | w23531);
assign w23532 = v7429;
assign w23533 = w6389 & w20234;
assign w23534 = ~pi14 & w23529;
assign w23535 = ~w23533 & w23534;
assign w23536 = w23532 & ~w23535;
assign w23537 = w23524 & w23536;
assign v7430 = ~(w23524 | w23536);
assign w23538 = v7430;
assign v7431 = ~(w23537 | w23538);
assign w23539 = v7431;
assign w23540 = (~w28575 & w30899) | (~w28575 & w30900) | (w30899 & w30900);
assign w23541 = w23539 & w23540;
assign v7432 = ~(w23539 | w23540);
assign w23542 = v7432;
assign v7433 = ~(w23541 | w23542);
assign w23543 = v7433;
assign w23544 = w7765 & w19954;
assign w23545 = w7466 & w19952;
assign w23546 = w7177 & w19958;
assign v7434 = ~(w23545 | w23546);
assign w23547 = v7434;
assign w23548 = ~w23544 & w23547;
assign w23549 = pi11 & ~w23548;
assign w23550 = w7178 & ~w21866;
assign w23551 = ~pi11 & w23548;
assign w23552 = ~w23550 & w23551;
assign w23553 = w9464 & ~w21866;
assign v7435 = ~(w23552 | w23553);
assign w23554 = v7435;
assign w23555 = ~w23549 & w23554;
assign v7436 = ~(w23543 | w23555);
assign w23556 = v7436;
assign w23557 = w23543 & w23555;
assign v7437 = ~(w23556 | w23557);
assign w23558 = v7437;
assign w23559 = w23417 & ~w23558;
assign w23560 = ~w23417 & w23558;
assign v7438 = ~(w23559 | w23560);
assign w23561 = v7438;
assign w23562 = w23416 & w23561;
assign v7439 = ~(w23416 | w23561);
assign w23563 = v7439;
assign v7440 = ~(w23562 | w23563);
assign w23564 = v7440;
assign w23565 = (~w22737 & w29941) | (~w22737 & w29942) | (w29941 & w29942);
assign w23566 = (w22890 & w23564) | (w22890 & w28576) | (w23564 & w28576);
assign v7441 = ~(w23565 | w23566);
assign w23567 = v7441;
assign w23568 = w23404 & ~w23567;
assign w23569 = ~w23404 & w23567;
assign v7442 = ~(w23568 | w23569);
assign w23570 = v7442;
assign w23571 = ~w23392 & w23570;
assign w23572 = w23392 & ~w23570;
assign v7443 = ~(w23571 | w23572);
assign w23573 = v7443;
assign v7444 = ~(w20183 | w20187);
assign w23574 = v7444;
assign v7445 = ~(w20154 | w20157);
assign w23575 = v7445;
assign w23576 = ~w172 & w4186;
assign w23577 = w4008 & w23576;
assign w23578 = w20149 & w23577;
assign w23579 = ~w23575 & w23578;
assign w23580 = w23575 & ~w23578;
assign v7446 = ~(w23579 | w23580);
assign w23581 = v7446;
assign w23582 = w928 & w12387;
assign w23583 = w3406 & w12381;
assign w23584 = w3402 & w12311;
assign v7447 = ~(w20168 | w23584);
assign w23585 = v7447;
assign w23586 = ~w23583 & w23585;
assign w23587 = ~w23582 & w23586;
assign w23588 = ~w23581 & w23587;
assign w23589 = w23581 & ~w23587;
assign v7448 = ~(w23588 | w23589);
assign w23590 = v7448;
assign v7449 = ~(w20163 | w20172);
assign w23591 = v7449;
assign w23592 = ~w23590 & w23591;
assign w23593 = w23590 & ~w23591;
assign v7450 = ~(w23592 | w23593);
assign w23594 = v7450;
assign w23595 = pi28 & w20176;
assign v7451 = ~(pi29 | w20176);
assign w23596 = v7451;
assign v7452 = ~(w23595 | w23596);
assign w23597 = v7452;
assign w23598 = w23594 & ~w23597;
assign w23599 = ~w23594 & w23597;
assign v7453 = ~(w23598 | w23599);
assign w23600 = v7453;
assign w23601 = ~w23574 & w23600;
assign w23602 = w23574 & ~w23600;
assign v7454 = ~(w23601 | w23602);
assign w23603 = v7454;
assign w23604 = (w19850 & w28577) | (w19850 & w28578) | (w28577 & w28578);
assign w23605 = ~w23603 & w23604;
assign w23606 = w23603 & ~w23604;
assign v7455 = ~(w23605 | w23606);
assign w23607 = v7455;
assign w23608 = w20197 & w23607;
assign v7456 = ~(w20197 | w23607);
assign w23609 = v7456;
assign v7457 = ~(w23608 | w23609);
assign w23610 = v7457;
assign w23611 = (~w20198 & w20147) | (~w20198 & w29123) | (w20147 & w29123);
assign w23612 = ~w20201 & w28222;
assign w23613 = (w23610 & w20201) | (w23610 & w28223) | (w20201 & w28223);
assign v7458 = ~(w23612 | w23613);
assign w23614 = v7458;
assign w23615 = w11035 & w23607;
assign w23616 = w11023 & w20197;
assign v7459 = ~(w23615 | w23616);
assign w23617 = v7459;
assign w23618 = (w23614 & w28400) | (w23614 & w28401) | (w28400 & w28401);
assign w23619 = w10986 & ~w19912;
assign w23620 = pi02 & ~w23619;
assign w23621 = (~w23614 & w28402) | (~w23614 & w28403) | (w28402 & w28403);
assign v7460 = ~(w23618 | w23621);
assign w23622 = v7460;
assign w23623 = w23573 & ~w23622;
assign w23624 = ~w23573 & w23622;
assign v7461 = ~(w23623 | w23624);
assign w23625 = v7461;
assign v7462 = ~(w22913 | w23625);
assign w23626 = v7462;
assign w23627 = w22913 & w23625;
assign v7463 = ~(w23626 | w23627);
assign w23628 = v7463;
assign w23629 = ~w23391 & w23628;
assign w23630 = w23391 & ~w23628;
assign v7464 = ~(w23629 | w23630);
assign w23631 = v7464;
assign w23632 = w22915 & ~w23390;
assign w23633 = w23629 & ~w23632;
assign w23634 = (~w23608 & w23611) | (~w23608 & w28084) | (w23611 & w28084);
assign v7465 = ~(w23593 | w23598);
assign w23635 = v7465;
assign v7466 = ~(w23579 | w23589);
assign w23636 = v7466;
assign w23637 = w4061 & w4189;
assign w23638 = ~w23578 & w23637;
assign w23639 = w23578 & ~w23637;
assign v7467 = ~(w23638 | w23639);
assign w23640 = v7467;
assign w23641 = w23636 & w23640;
assign v7468 = ~(w23636 | w23640);
assign w23642 = v7468;
assign v7469 = ~(w23641 | w23642);
assign w23643 = v7469;
assign w23644 = pi31 & ~w12311;
assign w23645 = w18 & ~w23644;
assign w23646 = w928 & ~w12506;
assign v7470 = ~(w3406 | w23646);
assign w23647 = v7470;
assign w23648 = ~w23645 & w23647;
assign w23649 = ~w23597 & w23648;
assign w23650 = w23597 & ~w23648;
assign v7471 = ~(w23649 | w23650);
assign w23651 = v7471;
assign w23652 = w23643 & ~w23651;
assign w23653 = ~w23643 & w23651;
assign v7472 = ~(w23652 | w23653);
assign w23654 = v7472;
assign v7473 = ~(w23635 | w23654);
assign w23655 = v7473;
assign w23656 = w23635 & w23654;
assign v7474 = ~(w23655 | w23656);
assign w23657 = v7474;
assign v7475 = ~(w23601 | w23604);
assign w23658 = v7475;
assign w23659 = ~w23602 & w23604;
assign v7476 = ~(w23658 | w23659);
assign w23660 = v7476;
assign w23661 = w23657 & w23660;
assign v7477 = ~(w23657 | w23660);
assign w23662 = v7477;
assign v7478 = ~(w23661 | w23662);
assign w23663 = v7478;
assign w23664 = (~w23611 & w28224) | (~w23611 & w28225) | (w28224 & w28225);
assign w23665 = (w23611 & w28226) | (w23611 & w28227) | (w28226 & w28227);
assign v7479 = ~(w23664 | w23665);
assign w23666 = v7479;
assign v7480 = ~(w23601 | w23606);
assign w23667 = v7480;
assign w23668 = ~w23657 & w23667;
assign w23669 = w23657 & ~w23667;
assign v7481 = ~(w23668 | w23669);
assign w23670 = v7481;
assign w23671 = w11035 & w23670;
assign w23672 = w11023 & w23607;
assign v7482 = ~(w23671 | w23672);
assign w23673 = v7482;
assign w23674 = (w23673 & ~w23666) | (w23673 & w28404) | (~w23666 & w28404);
assign v7483 = ~(pi02 | w23674);
assign w23675 = v7483;
assign w23676 = w10986 & w20197;
assign w23677 = pi02 & ~w23676;
assign w23678 = w23674 & w23677;
assign v7484 = ~(w23675 | w23678);
assign w23679 = v7484;
assign w23680 = w23404 & w23567;
assign w23681 = (~w23680 & ~w23392) | (~w23680 & w31112) | (~w23392 & w31112);
assign w23682 = w10445 & w22917;
assign w23683 = w10447 & w22917;
assign w23684 = w10419 & ~w19912;
assign w23685 = w9891 & w19853;
assign w23686 = w9401 & w19917;
assign v7485 = ~(w23685 | w23686);
assign w23687 = v7485;
assign w23688 = ~w23684 & w23687;
assign w23689 = pi05 & w23688;
assign v7486 = ~(pi05 | w23688);
assign w23690 = v7486;
assign v7487 = ~(w23689 | w23690);
assign w23691 = v7487;
assign w23692 = ~w23683 & w23691;
assign v7488 = ~(w23682 | w23692);
assign w23693 = v7488;
assign w23694 = w7178 & w20214;
assign w23695 = w7765 & ~w19939;
assign w23696 = w7177 & w19952;
assign w23697 = w7466 & w19954;
assign v7489 = ~(w23696 | w23697);
assign w23698 = v7489;
assign w23699 = ~w23695 & w23698;
assign w23700 = ~w23694 & w23699;
assign w23701 = ~pi11 & w23700;
assign w23702 = pi11 & ~w23700;
assign v7490 = ~(w23701 | w23702);
assign w23703 = v7490;
assign w23704 = (~w23537 & ~w23539) | (~w23537 & w31113) | (~w23539 & w31113);
assign w23705 = w7004 & w19958;
assign w23706 = w6871 & w19961;
assign w23707 = w6388 & w19966;
assign v7491 = ~(w23706 | w23707);
assign w23708 = v7491;
assign w23709 = ~w23705 & w23708;
assign w23710 = pi14 & ~w23709;
assign w23711 = w6389 & w21716;
assign w23712 = ~pi14 & w23709;
assign w23713 = ~w23711 & w23712;
assign w23714 = w17118 & w21716;
assign v7492 = ~(w23713 | w23714);
assign w23715 = v7492;
assign w23716 = ~w23710 & w23715;
assign w23717 = (~w23519 & w23418) | (~w23519 & w30090) | (w23418 & w30090);
assign w23718 = (~w23503 & w23419) | (~w23503 & w29943) | (w23419 & w29943);
assign w23719 = (~w23487 & w23420) | (~w23487 & w30442) | (w23420 & w30442);
assign v7493 = ~(w23472 | w23475);
assign w23720 = v7493;
assign w23721 = (~w23457 & w23422) | (~w23457 & w30725) | (w23422 & w30725);
assign w23722 = (~w23443 & w23423) | (~w23443 & w30726) | (w23423 & w30726);
assign w23723 = w740 & w752;
assign w23724 = w2325 & w23723;
assign w23725 = w2363 & w2397;
assign w23726 = w23724 & w23725;
assign w23727 = w185 & w23726;
assign w23728 = w13251 & w23727;
assign w23729 = w6569 & w6664;
assign w23730 = w3019 & w23729;
assign w23731 = w23728 & w23730;
assign w23732 = ~w886 & w2673;
assign v7494 = ~(w214 | w978);
assign w23733 = v7494;
assign w23734 = w2119 & w23733;
assign w23735 = w2241 & w23734;
assign w23736 = w3633 & w23735;
assign w23737 = w23732 & w23736;
assign w23738 = w1377 & w23737;
assign w23739 = w23731 & w23738;
assign w23740 = w3406 & w20031;
assign w23741 = w3402 & ~w20063;
assign w23742 = w3399 & ~w20038;
assign v7495 = ~(w23741 | w23742);
assign w23743 = v7495;
assign w23744 = ~w23740 & w23743;
assign w23745 = (w23744 & ~w20323) | (w23744 & w30901) | (~w20323 & w30901);
assign v7496 = ~(w23739 | w23745);
assign w23746 = v7496;
assign w23747 = w23739 & w23745;
assign v7497 = ~(w23746 | w23747);
assign w23748 = v7497;
assign w23749 = ~w23722 & w23748;
assign w23750 = w23722 & ~w23748;
assign v7498 = ~(w23749 | w23750);
assign w23751 = v7498;
assign w23752 = w3763 & ~w20028;
assign w23753 = w3760 & w20014;
assign v7499 = ~(w23752 | w23753);
assign w23754 = v7499;
assign w23755 = w3767 & ~w20026;
assign w23756 = w23754 & ~w23755;
assign w23757 = (~w20472 & w31299) | (~w20472 & w31300) | (w31299 & w31300);
assign w23758 = (w20472 & w31301) | (w20472 & w31302) | (w31301 & w31302);
assign v7500 = ~(w23757 | w23758);
assign w23759 = v7500;
assign w23760 = ~w23751 & w23759;
assign w23761 = w23751 & ~w23759;
assign v7501 = ~(w23760 | w23761);
assign w23762 = v7501;
assign w23763 = ~w23721 & w23762;
assign w23764 = w23721 & ~w23762;
assign v7502 = ~(w23763 | w23764);
assign w23765 = v7502;
assign w23766 = w4155 & w20005;
assign w23767 = w4158 & ~w20008;
assign v7503 = ~(w2873 | w20011);
assign w23768 = v7503;
assign v7504 = ~(w23767 | w23768);
assign w23769 = v7504;
assign w23770 = ~w23766 & w23769;
assign w23771 = (w23770 & ~w20639) | (w23770 & w30903) | (~w20639 & w30903);
assign w23772 = ~pi26 & w23771;
assign w23773 = pi26 & ~w23771;
assign v7505 = ~(w23772 | w23773);
assign w23774 = v7505;
assign v7506 = ~(w23765 | w23774);
assign w23775 = v7506;
assign w23776 = w23765 & w23774;
assign v7507 = ~(w23775 | w23776);
assign w23777 = v7507;
assign w23778 = ~w23720 & w23777;
assign w23779 = w23720 & ~w23777;
assign v7508 = ~(w23778 | w23779);
assign w23780 = v7508;
assign w23781 = w4913 & ~w19992;
assign w23782 = w4836 & ~w19997;
assign w23783 = w4763 & w20000;
assign v7509 = ~(w23782 | w23783);
assign w23784 = v7509;
assign w23785 = ~w23781 & w23784;
assign w23786 = (w23785 & ~w20655) | (w23785 & w30904) | (~w20655 & w30904);
assign w23787 = ~pi23 & w23786;
assign w23788 = pi23 & ~w23786;
assign v7510 = ~(w23787 | w23788);
assign w23789 = v7510;
assign v7511 = ~(w23780 | w23789);
assign w23790 = v7511;
assign w23791 = w23780 & w23789;
assign v7512 = ~(w23790 | w23791);
assign w23792 = v7512;
assign w23793 = ~w23719 & w23792;
assign w23794 = w23719 & ~w23792;
assign v7513 = ~(w23793 | w23794);
assign w23795 = v7513;
assign w23796 = w5114 & w20997;
assign w23797 = w5610 & w19983;
assign w23798 = w5113 & w19989;
assign w23799 = w5531 & w19986;
assign v7514 = ~(w23798 | w23799);
assign w23800 = v7514;
assign w23801 = ~w23797 & w23800;
assign w23802 = ~w23796 & w23801;
assign w23803 = ~pi20 & w23802;
assign w23804 = pi20 & ~w23802;
assign v7515 = ~(w23803 | w23804);
assign w23805 = v7515;
assign w23806 = w23795 & w23805;
assign v7516 = ~(w23795 | w23805);
assign w23807 = v7516;
assign v7517 = ~(w23806 | w23807);
assign w23808 = v7517;
assign w23809 = ~w23718 & w23808;
assign w23810 = w23718 & ~w23808;
assign v7518 = ~(w23809 | w23810);
assign w23811 = v7518;
assign w23812 = w5765 & w21401;
assign w23813 = w5983 & w19974;
assign w23814 = w6236 & ~w19971;
assign v7519 = ~(w23813 | w23814);
assign w23815 = v7519;
assign w23816 = w5764 & w19980;
assign w23817 = w23815 & ~w23816;
assign w23818 = ~w23812 & w23817;
assign w23819 = pi17 & w23818;
assign v7520 = ~(pi17 | w23818);
assign w23820 = v7520;
assign v7521 = ~(w23819 | w23820);
assign w23821 = v7521;
assign w23822 = w23811 & ~w23821;
assign w23823 = ~w23811 & w23821;
assign v7522 = ~(w23822 | w23823);
assign w23824 = v7522;
assign w23825 = ~w23717 & w23824;
assign w23826 = w23717 & ~w23824;
assign v7523 = ~(w23825 | w23826);
assign w23827 = v7523;
assign w23828 = w23716 & w23827;
assign v7524 = ~(w23716 | w23827);
assign w23829 = v7524;
assign v7525 = ~(w23828 | w23829);
assign w23830 = v7525;
assign v7526 = ~(w23704 | w23830);
assign w23831 = v7526;
assign w23832 = w23704 & w23830;
assign v7527 = ~(w23831 | w23832);
assign w23833 = v7527;
assign w23834 = ~w23703 & w23833;
assign w23835 = w23703 & ~w23833;
assign v7528 = ~(w23834 | w23835);
assign w23836 = v7528;
assign w23837 = (~w23556 & ~w23417) | (~w23556 & w28579) | (~w23417 & w28579);
assign w23838 = w23836 & ~w23837;
assign w23839 = ~w23836 & w23837;
assign v7529 = ~(w23838 | w23839);
assign w23840 = v7529;
assign w23841 = w9920 & w22262;
assign w23842 = w8926 & ~w19923;
assign w23843 = w8526 & ~w19929;
assign w23844 = w8140 & w19933;
assign v7530 = ~(w23843 | w23844);
assign w23845 = v7530;
assign w23846 = ~w23842 & w23845;
assign w23847 = pi08 & ~w23846;
assign w23848 = ~pi08 & w23846;
assign w23849 = (w22262 & w28405) | (w22262 & w28406) | (w28405 & w28406);
assign w23850 = ~w23841 & w23849;
assign w23851 = ~w23840 & w23850;
assign w23852 = w23840 & ~w23850;
assign v7531 = ~(w23851 | w23852);
assign w23853 = v7531;
assign w23854 = (~w22890 & w28580) | (~w22890 & w28581) | (w28580 & w28581);
assign w23855 = (w22890 & w29944) | (w22890 & w29945) | (w29944 & w29945);
assign w23856 = (~w22890 & w29946) | (~w22890 & w29947) | (w29946 & w29947);
assign v7532 = ~(w23855 | w23856);
assign w23857 = v7532;
assign w23858 = (~w23857 & w23692) | (~w23857 & w28407) | (w23692 & w28407);
assign w23859 = ~w23692 & w28408;
assign v7533 = ~(w23858 | w23859);
assign w23860 = v7533;
assign w23861 = w23681 & ~w23860;
assign w23862 = ~w23681 & w23860;
assign v7534 = ~(w23861 | w23862);
assign w23863 = v7534;
assign w23864 = ~w23679 & w23863;
assign w23865 = w23679 & ~w23863;
assign w23866 = (~w23624 & w23632) | (~w23624 & w28229) | (w23632 & w28229);
assign w23867 = w23866 & w23868;
assign v7535 = ~(w23864 | w23865);
assign w23868 = v7535;
assign v7536 = ~(w23866 | w23868);
assign w23869 = v7536;
assign v7537 = ~(w23867 | w23869);
assign w23870 = v7537;
assign w23871 = w23633 & w23870;
assign v7538 = ~(w23633 | w23870);
assign w23872 = v7538;
assign v7539 = ~(w23871 | w23872);
assign w23873 = v7539;
assign w23874 = w10419 & w20197;
assign w23875 = w9891 & ~w19912;
assign w23876 = w9401 & w19853;
assign v7540 = ~(w23875 | w23876);
assign w23877 = v7540;
assign w23878 = ~w23874 & w23877;
assign w23879 = (~w20203 & w28409) | (~w20203 & w28410) | (w28409 & w28410);
assign w23880 = (w20203 & w28411) | (w20203 & w28412) | (w28411 & w28412);
assign v7541 = ~(w23879 | w23880);
assign w23881 = v7541;
assign w23882 = (~w23851 & w23854) | (~w23851 & w28086) | (w23854 & w28086);
assign v7542 = ~(w23834 | w23838);
assign w23883 = v7542;
assign w23884 = w7765 & w19933;
assign w23885 = w7177 & w19954;
assign w23886 = w7466 & ~w19939;
assign v7543 = ~(w23885 | w23886);
assign w23887 = v7543;
assign w23888 = ~w23884 & w23887;
assign w23889 = (w23888 & w22304) | (w23888 & w28413) | (w22304 & w28413);
assign w23890 = ~pi11 & w23889;
assign w23891 = pi11 & ~w23889;
assign v7544 = ~(w23890 | w23891);
assign w23892 = v7544;
assign w23893 = (~w23829 & ~w23704) | (~w23829 & w29948) | (~w23704 & w29948);
assign w23894 = w17118 & ~w21882;
assign w23895 = w7004 & w19952;
assign w23896 = w6871 & w19958;
assign w23897 = w6388 & w19961;
assign v7545 = ~(w23896 | w23897);
assign w23898 = v7545;
assign w23899 = ~w23895 & w23898;
assign w23900 = pi14 & ~w23899;
assign w23901 = w6389 & ~w21882;
assign w23902 = ~pi14 & w23899;
assign w23903 = ~w23901 & w23902;
assign v7546 = ~(w23900 | w23903);
assign w23904 = v7546;
assign w23905 = ~w23894 & w23904;
assign w23906 = (~w23822 & w23717) | (~w23822 & w29949) | (w23717 & w29949);
assign v7547 = ~(w23791 | w23793);
assign w23907 = v7547;
assign w23908 = (~w23776 & w23720) | (~w23776 & w30727) | (w23720 & w30727);
assign w23909 = (~w23761 & w23721) | (~w23761 & w30905) | (w23721 & w30905);
assign w23910 = (~w23746 & w23722) | (~w23746 & w30906) | (w23722 & w30906);
assign w23911 = ~w469 & w1237;
assign w23912 = w12661 & w13290;
assign w23913 = w12012 & w23912;
assign w23914 = w23911 & w23913;
assign w23915 = w442 & w2516;
assign w23916 = w565 & w23915;
assign w23917 = w3051 & w6686;
assign w23918 = w3552 & w23917;
assign w23919 = w23916 & w23918;
assign w23920 = w1620 & w1624;
assign w23921 = ~w711 & w23920;
assign w23922 = ~w437 & w23921;
assign w23923 = w23919 & w23922;
assign w23924 = w23914 & w23923;
assign w23925 = w1185 & w2392;
assign w23926 = w23924 & w23925;
assign w23927 = w3406 & ~w20026;
assign w23928 = w3399 & ~w20063;
assign w23929 = w3402 & w20031;
assign v7548 = ~(w23928 | w23929);
assign w23930 = v7548;
assign w23931 = ~w23927 & w23930;
assign w23932 = (~w30728 & w30907) | (~w30728 & w30908) | (w30907 & w30908);
assign v7549 = ~(w23926 | w23932);
assign w23933 = v7549;
assign w23934 = w23926 & w23932;
assign v7550 = ~(w23933 | w23934);
assign w23935 = v7550;
assign w23936 = ~w23910 & w23935;
assign w23937 = w23910 & ~w23935;
assign v7551 = ~(w23936 | w23937);
assign w23938 = v7551;
assign w23939 = w3763 & w20014;
assign w23940 = w3760 & ~w20011;
assign v7552 = ~(w23939 | w23940);
assign w23941 = v7552;
assign w23942 = w3767 & ~w20028;
assign w23943 = w23941 & ~w23942;
assign w23944 = (w23943 & ~w20459) | (w23943 & w31303) | (~w20459 & w31303);
assign v7553 = ~(pi29 | w23944);
assign w23945 = v7553;
assign w23946 = pi29 & w23944;
assign v7554 = ~(w23945 | w23946);
assign w23947 = v7554;
assign w23948 = w23938 & ~w23947;
assign w23949 = ~w23938 & w23947;
assign v7555 = ~(w23948 | w23949);
assign w23950 = v7555;
assign w23951 = ~w23909 & w23950;
assign w23952 = w23909 & ~w23950;
assign v7556 = ~(w23951 | w23952);
assign w23953 = v7556;
assign w23954 = w4155 & w20000;
assign v7557 = ~(w2873 | w20008);
assign w23955 = v7557;
assign w23956 = w4158 & w20005;
assign v7558 = ~(w23955 | w23956);
assign w23957 = v7558;
assign w23958 = ~w23954 & w23957;
assign w23959 = (w23958 & ~w20681) | (w23958 & w31304) | (~w20681 & w31304);
assign w23960 = ~pi26 & w23959;
assign w23961 = pi26 & ~w23959;
assign v7559 = ~(w23960 | w23961);
assign w23962 = v7559;
assign v7560 = ~(w23953 | w23962);
assign w23963 = v7560;
assign w23964 = w23953 & w23962;
assign v7561 = ~(w23963 | w23964);
assign w23965 = v7561;
assign w23966 = ~w23908 & w23965;
assign w23967 = w23908 & ~w23965;
assign v7562 = ~(w23966 | w23967);
assign w23968 = v7562;
assign w23969 = w4764 & w20965;
assign w23970 = w4913 & w19989;
assign w23971 = w4763 & ~w19997;
assign w23972 = w4836 & ~w19992;
assign v7563 = ~(w23971 | w23972);
assign w23973 = v7563;
assign w23974 = ~w23970 & w23973;
assign w23975 = ~w23969 & w23974;
assign w23976 = ~pi23 & w23975;
assign w23977 = pi23 & ~w23975;
assign v7564 = ~(w23976 | w23977);
assign w23978 = v7564;
assign w23979 = w23968 & w23978;
assign v7565 = ~(w23968 | w23978);
assign w23980 = v7565;
assign v7566 = ~(w23979 | w23980);
assign w23981 = v7566;
assign w23982 = ~w23907 & w23981;
assign w23983 = w23907 & ~w23981;
assign v7567 = ~(w23982 | w23983);
assign w23984 = v7567;
assign w23985 = w5114 & w20982;
assign w23986 = w5531 & w19983;
assign w23987 = w5610 & w19980;
assign v7568 = ~(w23986 | w23987);
assign w23988 = v7568;
assign w23989 = w5113 & w19986;
assign w23990 = w23988 & ~w23989;
assign w23991 = ~w23985 & w23990;
assign w23992 = pi20 & w23991;
assign v7569 = ~(pi20 | w23991);
assign w23993 = v7569;
assign v7570 = ~(w23992 | w23993);
assign w23994 = v7570;
assign w23995 = w23984 & ~w23994;
assign w23996 = ~w23984 & w23994;
assign v7571 = ~(w23995 | w23996);
assign w23997 = v7571;
assign w23998 = (~w23806 & w23718) | (~w23806 & w30443) | (w23718 & w30443);
assign w23999 = w23997 & ~w23998;
assign w24000 = ~w23997 & w23998;
assign v7572 = ~(w23999 | w24000);
assign w24001 = v7572;
assign w24002 = w5765 & w21385;
assign w24003 = w5983 & ~w19971;
assign w24004 = w6236 & w19966;
assign v7573 = ~(w24003 | w24004);
assign w24005 = v7573;
assign w24006 = w5764 & w19974;
assign w24007 = w24005 & ~w24006;
assign w24008 = ~w24002 & w24007;
assign w24009 = pi17 & w24008;
assign v7574 = ~(pi17 | w24008);
assign w24010 = v7574;
assign v7575 = ~(w24009 | w24010);
assign w24011 = v7575;
assign w24012 = w24001 & ~w24011;
assign w24013 = ~w24001 & w24011;
assign v7576 = ~(w24012 | w24013);
assign w24014 = v7576;
assign w24015 = w23906 & w24014;
assign v7577 = ~(w23906 | w24014);
assign w24016 = v7577;
assign v7578 = ~(w24015 | w24016);
assign w24017 = v7578;
assign w24018 = w23905 & ~w24017;
assign w24019 = ~w23905 & w24017;
assign v7579 = ~(w24018 | w24019);
assign w24020 = v7579;
assign v7580 = ~(w23893 | w24020);
assign w24021 = v7580;
assign w24022 = w23893 & w24020;
assign v7581 = ~(w24021 | w24022);
assign w24023 = v7581;
assign w24024 = w23892 & w24023;
assign v7582 = ~(w23892 | w24023);
assign w24025 = v7582;
assign v7583 = ~(w24024 | w24025);
assign w24026 = v7583;
assign v7584 = ~(w23883 | w24026);
assign w24027 = v7584;
assign w24028 = w23883 & w24026;
assign v7585 = ~(w24027 | w24028);
assign w24029 = v7585;
assign w24030 = w8926 & w19917;
assign w24031 = w8140 & ~w19929;
assign w24032 = w8526 & ~w19923;
assign v7586 = ~(w24031 | w24032);
assign w24033 = v7586;
assign w24034 = ~w24030 & w24033;
assign w24035 = (~w22895 & w28414) | (~w22895 & w28415) | (w28414 & w28415);
assign w24036 = (w22895 & w28416) | (w22895 & w28417) | (w28416 & w28417);
assign v7587 = ~(w24035 | w24036);
assign w24037 = v7587;
assign v7588 = ~(w24029 | w24037);
assign w24038 = v7588;
assign w24039 = w24029 & w24037;
assign v7589 = ~(w24038 | w24039);
assign w24040 = v7589;
assign v7590 = ~(w23882 | w24040);
assign w24041 = v7590;
assign w24042 = w23882 & w24040;
assign v7591 = ~(w24041 | w24042);
assign w24043 = v7591;
assign w24044 = w23881 & w24043;
assign v7592 = ~(w23881 | w24043);
assign w24045 = v7592;
assign v7593 = ~(w24044 | w24045);
assign w24046 = v7593;
assign w24047 = (~w23858 & w23572) | (~w23858 & w31114) | (w23572 & w31114);
assign w24048 = w24046 & w24047;
assign v7594 = ~(w24046 | w24047);
assign w24049 = v7594;
assign v7595 = ~(w24048 | w24049);
assign w24050 = v7595;
assign w24051 = w23607 & w23670;
assign v7596 = ~(w23643 | w23650);
assign w24052 = v7596;
assign w24053 = w23643 & ~w23649;
assign v7597 = ~(w24052 | w24053);
assign w24054 = v7597;
assign v7598 = ~(w23639 | w23641);
assign w24055 = v7598;
assign w24056 = ~pi31 & w32;
assign w24057 = w4061 & w4191;
assign v7599 = ~(w24056 | w24057);
assign w24058 = v7599;
assign w24059 = ~w24055 & w24058;
assign w24060 = w24055 & ~w24058;
assign v7600 = ~(w24059 | w24060);
assign w24061 = v7600;
assign w24062 = w24054 & ~w24061;
assign w24063 = ~w24054 & w24061;
assign v7601 = ~(w24062 | w24063);
assign w24064 = v7601;
assign v7602 = ~(w23655 | w23667);
assign w24065 = v7602;
assign w24066 = ~w23656 & w23667;
assign v7603 = ~(w24065 | w24066);
assign w24067 = v7603;
assign w24068 = w24064 & w24067;
assign v7604 = ~(w24064 | w24067);
assign w24069 = v7604;
assign v7605 = ~(w24068 | w24069);
assign w24070 = v7605;
assign w24071 = (~w23611 & w28582) | (~w23611 & w28583) | (w28582 & w28583);
assign w24072 = (w23611 & w28584) | (w23611 & w28585) | (w28584 & w28585);
assign v7606 = ~(w24071 | w24072);
assign w24073 = v7606;
assign v7607 = ~(w23655 | w23669);
assign w24074 = v7607;
assign w24075 = ~w24064 & w24074;
assign w24076 = w24064 & ~w24074;
assign v7608 = ~(w24075 | w24076);
assign w24077 = v7608;
assign w24078 = w11035 & ~w24077;
assign w24079 = w11023 & w23670;
assign v7609 = ~(w24078 | w24079);
assign w24080 = v7609;
assign w24081 = (w24080 & ~w24073) | (w24080 & w28418) | (~w24073 & w28418);
assign v7610 = ~(pi02 | w24081);
assign w24082 = v7610;
assign w24083 = w10986 & w23607;
assign w24084 = pi02 & ~w24083;
assign w24085 = w24081 & w24084;
assign v7611 = ~(w24082 | w24085);
assign w24086 = v7611;
assign w24087 = w24050 & ~w24086;
assign w24088 = ~w24050 & w24086;
assign v7612 = ~(w24087 | w24088);
assign w24089 = v7612;
assign w24090 = (~w23864 & ~w23866) | (~w23864 & w28089) | (~w23866 & w28089);
assign w24091 = w24089 & ~w24090;
assign w24092 = ~w24089 & w24090;
assign v7613 = ~(w24091 | w24092);
assign w24093 = v7613;
assign w24094 = w23871 & w24093;
assign v7614 = ~(w23871 | w24093);
assign w24095 = v7614;
assign v7615 = ~(w24094 | w24095);
assign w24096 = v7615;
assign w24097 = (~w24087 & w24090) | (~w24087 & w31115) | (w24090 & w31115);
assign w24098 = (~w24045 & ~w24047) | (~w24045 & w28419) | (~w24047 & w28419);
assign w24099 = w9920 & w22936;
assign w24100 = w8926 & w19853;
assign w24101 = w8526 & w19917;
assign w24102 = w8140 & ~w19923;
assign v7616 = ~(w24101 | w24102);
assign w24103 = v7616;
assign w24104 = ~w24100 & w24103;
assign w24105 = pi08 & ~w24104;
assign w24106 = ~pi08 & w24104;
assign w24107 = (w22936 & w28420) | (w22936 & w28421) | (w28420 & w28421);
assign w24108 = ~w24099 & w24107;
assign w24109 = (~w24024 & ~w23883) | (~w24024 & w29950) | (~w23883 & w29950);
assign w24110 = w7178 & ~w22285;
assign w24111 = w7765 & ~w19929;
assign w24112 = w7177 & ~w19939;
assign w24113 = w7466 & w19933;
assign v7617 = ~(w24112 | w24113);
assign w24114 = v7617;
assign w24115 = ~w24111 & w24114;
assign w24116 = ~w24110 & w24115;
assign w24117 = ~pi11 & w24116;
assign w24118 = pi11 & ~w24116;
assign v7618 = ~(w24117 | w24118);
assign w24119 = v7618;
assign w24120 = w7004 & w19954;
assign w24121 = w6871 & w19952;
assign w24122 = w6388 & w19958;
assign v7619 = ~(w24121 | w24122);
assign w24123 = v7619;
assign w24124 = ~w24120 & w24123;
assign w24125 = pi14 & ~w24124;
assign w24126 = w6389 & ~w21866;
assign w24127 = ~pi14 & w24124;
assign w24128 = ~w24126 & w24127;
assign w24129 = w17118 & ~w21866;
assign v7620 = ~(w24128 | w24129);
assign w24130 = v7620;
assign w24131 = ~w24125 & w24130;
assign v7621 = ~(w23995 | w23999);
assign w24132 = v7621;
assign w24133 = (~w23979 & w23907) | (~w23979 & w30729) | (w23907 & w30729);
assign w24134 = (~w23964 & w23908) | (~w23964 & w30909) | (w23908 & w30909);
assign w24135 = (~w23948 & ~w23950) | (~w23948 & w31116) | (~w23950 & w31116);
assign v7622 = ~(w23933 | w23936);
assign w24136 = v7622;
assign w24137 = w2078 & w4975;
assign w24138 = ~w202 & w24137;
assign w24139 = ~w212 & w14315;
assign w24140 = w24138 & w24139;
assign w24141 = w6706 & w24140;
assign w24142 = w2507 & w3051;
assign w24143 = w1542 & w24142;
assign w24144 = w2431 & w24143;
assign w24145 = w2483 & w24144;
assign w24146 = w1359 & w1378;
assign w24147 = w1442 & w24146;
assign w24148 = w2858 & w24147;
assign w24149 = w24145 & w24148;
assign w24150 = w24141 & w24149;
assign w24151 = w4229 & w24150;
assign w24152 = w3406 & ~w20028;
assign w24153 = w3399 & w20031;
assign w24154 = w3402 & ~w20026;
assign v7623 = ~(w24153 | w24154);
assign w24155 = v7623;
assign w24156 = ~w24152 & w24155;
assign w24157 = (w24156 & ~w20431) | (w24156 & w30910) | (~w20431 & w30910);
assign v7624 = ~(w24151 | w24157);
assign w24158 = v7624;
assign w24159 = w24151 & w24157;
assign v7625 = ~(w24158 | w24159);
assign w24160 = v7625;
assign w24161 = ~w24136 & w24160;
assign w24162 = w24136 & ~w24160;
assign v7626 = ~(w24161 | w24162);
assign w24163 = v7626;
assign w24164 = w3529 & w20446;
assign w24165 = w3763 & ~w20011;
assign w24166 = w3760 & ~w20008;
assign v7627 = ~(w24165 | w24166);
assign w24167 = v7627;
assign w24168 = w3767 & w20014;
assign w24169 = w24167 & ~w24168;
assign w24170 = ~w24164 & w24169;
assign w24171 = pi29 & w24170;
assign v7628 = ~(pi29 | w24170);
assign w24172 = v7628;
assign v7629 = ~(w24171 | w24172);
assign w24173 = v7629;
assign w24174 = w24163 & ~w24173;
assign w24175 = ~w24163 & w24173;
assign v7630 = ~(w24174 | w24175);
assign w24176 = v7630;
assign w24177 = ~w24135 & w24176;
assign w24178 = w24135 & ~w24176;
assign v7631 = ~(w24177 | w24178);
assign w24179 = v7631;
assign w24180 = w4153 & w20668;
assign w24181 = w4155 & ~w19997;
assign w24182 = ~w2873 & w20005;
assign w24183 = w4158 & w20000;
assign v7632 = ~(w24182 | w24183);
assign w24184 = v7632;
assign w24185 = ~w24181 & w24184;
assign w24186 = ~w24180 & w24185;
assign w24187 = ~pi26 & w24186;
assign w24188 = pi26 & ~w24186;
assign v7633 = ~(w24187 | w24188);
assign w24189 = v7633;
assign v7634 = ~(w24179 | w24189);
assign w24190 = v7634;
assign w24191 = w24179 & w24189;
assign v7635 = ~(w24190 | w24191);
assign w24192 = v7635;
assign w24193 = ~w24134 & w24192;
assign w24194 = w24134 & ~w24192;
assign v7636 = ~(w24193 | w24194);
assign w24195 = v7636;
assign w24196 = w4764 & w21012;
assign w24197 = w4763 & ~w19992;
assign w24198 = w4913 & w19986;
assign v7637 = ~(w24197 | w24198);
assign w24199 = v7637;
assign w24200 = w4836 & w19989;
assign w24201 = w24199 & ~w24200;
assign w24202 = ~w24196 & w24201;
assign w24203 = pi23 & w24202;
assign v7638 = ~(pi23 | w24202);
assign w24204 = v7638;
assign v7639 = ~(w24203 | w24204);
assign w24205 = v7639;
assign w24206 = w24195 & ~w24205;
assign w24207 = ~w24195 & w24205;
assign v7640 = ~(w24206 | w24207);
assign w24208 = v7640;
assign w24209 = ~w24133 & w24208;
assign w24210 = w24133 & ~w24208;
assign v7641 = ~(w24209 | w24210);
assign w24211 = v7641;
assign w24212 = w5114 & w21362;
assign w24213 = w5531 & w19980;
assign w24214 = w5610 & w19974;
assign v7642 = ~(w24213 | w24214);
assign w24215 = v7642;
assign w24216 = w5113 & w19983;
assign w24217 = w24215 & ~w24216;
assign w24218 = ~w24212 & w24217;
assign w24219 = pi20 & w24218;
assign v7643 = ~(pi20 | w24218);
assign w24220 = v7643;
assign v7644 = ~(w24219 | w24220);
assign w24221 = v7644;
assign w24222 = w24211 & ~w24221;
assign w24223 = ~w24211 & w24221;
assign v7645 = ~(w24222 | w24223);
assign w24224 = v7645;
assign w24225 = w24132 & ~w24224;
assign w24226 = ~w24132 & w24224;
assign v7646 = ~(w24225 | w24226);
assign w24227 = v7646;
assign w24228 = w5765 & w20234;
assign w24229 = w5983 & w19966;
assign w24230 = w6236 & w19961;
assign v7647 = ~(w24229 | w24230);
assign w24231 = v7647;
assign w24232 = w5764 & ~w19971;
assign w24233 = w24231 & ~w24232;
assign w24234 = ~w24228 & w24233;
assign w24235 = pi17 & w24234;
assign v7648 = ~(pi17 | w24234);
assign w24236 = v7648;
assign v7649 = ~(w24235 | w24236);
assign w24237 = v7649;
assign w24238 = w24227 & ~w24237;
assign w24239 = ~w24227 & w24237;
assign v7650 = ~(w24238 | w24239);
assign w24240 = v7650;
assign w24241 = (~w24013 & ~w23906) | (~w24013 & w30444) | (~w23906 & w30444);
assign w24242 = w24240 & w24241;
assign v7651 = ~(w24240 | w24241);
assign w24243 = v7651;
assign v7652 = ~(w24242 | w24243);
assign w24244 = v7652;
assign w24245 = w24131 & w24244;
assign v7653 = ~(w24131 | w24244);
assign w24246 = v7653;
assign v7654 = ~(w24245 | w24246);
assign w24247 = v7654;
assign w24248 = (w23704 & w30091) | (w23704 & w30092) | (w30091 & w30092);
assign w24249 = (~w30092 & w30911) | (~w30092 & w30912) | (w30911 & w30912);
assign w24250 = ~w24247 & w24249;
assign w24251 = w24247 & ~w24249;
assign v7655 = ~(w24250 | w24251);
assign w24252 = v7655;
assign w24253 = w24119 & ~w24252;
assign w24254 = ~w24119 & w24252;
assign v7656 = ~(w24253 | w24254);
assign w24255 = v7656;
assign w24256 = ~w24109 & w24255;
assign w24257 = w24109 & ~w24255;
assign v7657 = ~(w24256 | w24257);
assign w24258 = v7657;
assign v7658 = ~(w24108 | w24258);
assign w24259 = v7658;
assign w24260 = w24108 & w24258;
assign v7659 = ~(w24259 | w24260);
assign w24261 = v7659;
assign w24262 = (~w24038 & ~w23882) | (~w24038 & w28090) | (~w23882 & w28090);
assign w24263 = ~w24261 & w24262;
assign w24264 = w24261 & ~w24262;
assign v7660 = ~(w24263 | w24264);
assign w24265 = v7660;
assign w24266 = w10419 & w23607;
assign w24267 = w9401 & ~w19912;
assign w24268 = w9891 & w20197;
assign v7661 = ~(w24267 | w24268);
assign w24269 = v7661;
assign w24270 = ~w24266 & w24269;
assign w24271 = (~w23614 & w28586) | (~w23614 & w28587) | (w28586 & w28587);
assign w24272 = (w23614 & w28588) | (w23614 & w28589) | (w28588 & w28589);
assign v7662 = ~(w24271 | w24272);
assign w24273 = v7662;
assign w24274 = w24265 & w24273;
assign v7663 = ~(w24265 | w24273);
assign w24275 = v7663;
assign v7664 = ~(w24274 | w24275);
assign w24276 = v7664;
assign w24277 = w24098 & w24276;
assign v7665 = ~(w24098 | w24276);
assign w24278 = v7665;
assign v7666 = ~(w24277 | w24278);
assign w24279 = v7666;
assign w24280 = (~w23611 & w28590) | (~w23611 & w28591) | (w28590 & w28591);
assign w24281 = (w23634 & w28423) | (w23634 & w28424) | (w28423 & w28424);
assign v7667 = ~(w24280 | w24281);
assign w24282 = v7667;
assign w24283 = ~w4 & w24282;
assign w24284 = ~w23670 & w24077;
assign w24285 = w11035 & w24284;
assign w24286 = w11023 & ~w24077;
assign v7668 = ~(w24285 | w24286);
assign w24287 = v7668;
assign w24288 = ~w24283 & w24287;
assign w24289 = pi02 & ~w24288;
assign w24290 = w10986 & w23670;
assign w24291 = pi02 & ~w24290;
assign w24292 = w24288 & ~w24291;
assign v7669 = ~(w24289 | w24292);
assign w24293 = v7669;
assign w24294 = w24279 & ~w24293;
assign w24295 = ~w24279 & w24293;
assign v7670 = ~(w24294 | w24295);
assign w24296 = v7670;
assign w24297 = ~w24097 & w24296;
assign w24298 = w24097 & ~w24296;
assign v7671 = ~(w24297 | w24298);
assign w24299 = v7671;
assign w24300 = w24094 & w24299;
assign v7672 = ~(w24094 | w24299);
assign w24301 = v7672;
assign v7673 = ~(w24300 | w24301);
assign w24302 = v7673;
assign w24303 = w11023 & w24284;
assign w24304 = w24070 & ~w24280;
assign v7674 = ~(w4 | w24304);
assign w24305 = v7674;
assign v7675 = ~(w24303 | w24305);
assign w24306 = v7675;
assign w24307 = pi02 & ~w24306;
assign w24308 = w10986 & ~w24077;
assign w24309 = pi02 & ~w24308;
assign w24310 = w24306 & ~w24309;
assign v7676 = ~(w24307 | w24310);
assign w24311 = v7676;
assign w24312 = w10445 & w23666;
assign w24313 = w10419 & w23670;
assign w24314 = w9891 & w23607;
assign w24315 = w9401 & w20197;
assign v7677 = ~(w24314 | w24315);
assign w24316 = v7677;
assign w24317 = ~w24313 & w24316;
assign w24318 = pi05 & w24317;
assign v7678 = ~(pi05 | w24317);
assign w24319 = v7678;
assign v7679 = ~(w24318 | w24319);
assign w24320 = v7679;
assign w24321 = (w24320 & ~w23666) | (w24320 & w28425) | (~w23666 & w28425);
assign v7680 = ~(w24312 | w24321);
assign w24322 = v7680;
assign w24323 = w9920 & w22917;
assign w24324 = w8926 & ~w19912;
assign w24325 = w8526 & w19853;
assign w24326 = w8140 & w19917;
assign v7681 = ~(w24325 | w24326);
assign w24327 = v7681;
assign w24328 = (pi08 & w24324) | (pi08 & w28426) | (w24324 & w28426);
assign w24329 = ~w24324 & w28427;
assign w24330 = (w22917 & w28236) | (w22917 & w28237) | (w28236 & w28237);
assign w24331 = ~w24323 & w24330;
assign w24332 = w9464 & w22262;
assign w24333 = w7765 & ~w19923;
assign w24334 = w7177 & w19933;
assign w24335 = w7466 & ~w19929;
assign v7682 = ~(w24334 | w24335);
assign w24336 = v7682;
assign w24337 = ~w24333 & w24336;
assign w24338 = pi11 & ~w24337;
assign w24339 = ~pi11 & w24337;
assign w24340 = (w24339 & ~w22262) | (w24339 & w28428) | (~w22262 & w28428);
assign v7683 = ~(w24338 | w24340);
assign w24341 = v7683;
assign w24342 = ~w24332 & w24341;
assign w24343 = (~w24238 & ~w24240) | (~w24238 & w31221) | (~w24240 & w31221);
assign w24344 = (~w24206 & w24133) | (~w24206 & w30913) | (w24133 & w30913);
assign w24345 = (~w24191 & w24134) | (~w24191 & w31117) | (w24134 & w31117);
assign v7684 = ~(w24174 | w24177);
assign w24346 = v7684;
assign w24347 = (~w24158 & w24136) | (~w24158 & w31118) | (w24136 & w31118);
assign w24348 = ~w1108 & w13155;
assign w24349 = w1892 & w1912;
assign w24350 = ~w220 & w2995;
assign w24351 = w24349 & w24350;
assign w24352 = w2363 & w2805;
assign w24353 = w1366 & w24352;
assign w24354 = w24351 & w24353;
assign w24355 = w24348 & w24354;
assign w24356 = w829 & w24355;
assign w24357 = w1028 & w1864;
assign w24358 = w796 & w24357;
assign w24359 = w24356 & w24358;
assign w24360 = w261 & w712;
assign w24361 = w1541 & w24360;
assign w24362 = w2718 & w24361;
assign w24363 = w419 & w2452;
assign w24364 = ~w505 & w1410;
assign w24365 = w24363 & w24364;
assign w24366 = w24362 & w24365;
assign w24367 = ~w338 & w24366;
assign w24368 = w24359 & w24367;
assign w24369 = w1085 & w1981;
assign w24370 = w4650 & w24369;
assign w24371 = w24368 & w24370;
assign w24372 = w928 & w20472;
assign w24373 = w3406 & w20014;
assign w24374 = w3402 & ~w20028;
assign w24375 = w3399 & ~w20026;
assign v7685 = ~(w24374 | w24375);
assign w24376 = v7685;
assign w24377 = ~w24373 & w24376;
assign w24378 = ~w24372 & w24377;
assign v7686 = ~(w24371 | w24378);
assign w24379 = v7686;
assign w24380 = w24371 & w24378;
assign v7687 = ~(w24379 | w24380);
assign w24381 = v7687;
assign w24382 = ~w24347 & w24381;
assign w24383 = w24347 & ~w24381;
assign v7688 = ~(w24382 | w24383);
assign w24384 = v7688;
assign w24385 = w3529 & w20639;
assign w24386 = w3760 & w20005;
assign w24387 = w3763 & ~w20008;
assign w24388 = w3767 & ~w20011;
assign v7689 = ~(w24387 | w24388);
assign w24389 = v7689;
assign w24390 = ~w24386 & w24389;
assign w24391 = ~w24385 & w24390;
assign w24392 = ~pi29 & w24391;
assign w24393 = pi29 & ~w24391;
assign v7690 = ~(w24392 | w24393);
assign w24394 = v7690;
assign w24395 = w24384 & w24394;
assign v7691 = ~(w24384 | w24394);
assign w24396 = v7691;
assign v7692 = ~(w24395 | w24396);
assign w24397 = v7692;
assign w24398 = ~w24346 & w24397;
assign w24399 = w24346 & ~w24397;
assign v7693 = ~(w24398 | w24399);
assign w24400 = v7693;
assign w24401 = w4153 & w20655;
assign w24402 = w4155 & ~w19992;
assign w24403 = w4158 & ~w19997;
assign w24404 = ~w2873 & w20000;
assign v7694 = ~(w24403 | w24404);
assign w24405 = v7694;
assign w24406 = ~w24402 & w24405;
assign w24407 = ~w24401 & w24406;
assign w24408 = ~pi26 & w24407;
assign w24409 = pi26 & ~w24407;
assign v7695 = ~(w24408 | w24409);
assign w24410 = v7695;
assign w24411 = w24400 & w24410;
assign v7696 = ~(w24400 | w24410);
assign w24412 = v7696;
assign v7697 = ~(w24411 | w24412);
assign w24413 = v7697;
assign w24414 = ~w24345 & w24413;
assign w24415 = w24345 & ~w24413;
assign v7698 = ~(w24414 | w24415);
assign w24416 = v7698;
assign w24417 = w4764 & w20997;
assign w24418 = w4913 & w19983;
assign w24419 = w4763 & w19989;
assign w24420 = w4836 & w19986;
assign v7699 = ~(w24419 | w24420);
assign w24421 = v7699;
assign w24422 = ~w24418 & w24421;
assign w24423 = ~w24417 & w24422;
assign w24424 = ~pi23 & w24423;
assign w24425 = pi23 & ~w24423;
assign v7700 = ~(w24424 | w24425);
assign w24426 = v7700;
assign w24427 = w24416 & w24426;
assign v7701 = ~(w24416 | w24426);
assign w24428 = v7701;
assign v7702 = ~(w24427 | w24428);
assign w24429 = v7702;
assign w24430 = ~w24344 & w24429;
assign w24431 = w24344 & ~w24429;
assign v7703 = ~(w24430 | w24431);
assign w24432 = v7703;
assign w24433 = w5114 & w21401;
assign w24434 = w5610 & ~w19971;
assign w24435 = w5113 & w19980;
assign w24436 = w5531 & w19974;
assign v7704 = ~(w24435 | w24436);
assign w24437 = v7704;
assign w24438 = ~w24434 & w24437;
assign w24439 = ~w24433 & w24438;
assign w24440 = ~pi20 & w24439;
assign w24441 = pi20 & ~w24439;
assign v7705 = ~(w24440 | w24441);
assign w24442 = v7705;
assign w24443 = w24432 & w24442;
assign v7706 = ~(w24432 | w24442);
assign w24444 = v7706;
assign v7707 = ~(w24443 | w24444);
assign w24445 = v7707;
assign w24446 = (~w24222 & w24132) | (~w24222 & w30730) | (w24132 & w30730);
assign w24447 = w24445 & ~w24446;
assign w24448 = ~w24445 & w24446;
assign v7708 = ~(w24447 | w24448);
assign w24449 = v7708;
assign w24450 = w5765 & w21716;
assign w24451 = w5983 & w19961;
assign w24452 = w6236 & w19958;
assign v7709 = ~(w24451 | w24452);
assign w24453 = v7709;
assign w24454 = w5764 & w19966;
assign w24455 = w24453 & ~w24454;
assign w24456 = ~w24450 & w24455;
assign w24457 = pi17 & w24456;
assign v7710 = ~(pi17 | w24456);
assign w24458 = v7710;
assign v7711 = ~(w24457 | w24458);
assign w24459 = v7711;
assign w24460 = w24449 & ~w24459;
assign w24461 = ~w24449 & w24459;
assign v7712 = ~(w24460 | w24461);
assign w24462 = v7712;
assign w24463 = w24343 & ~w24462;
assign w24464 = ~w24343 & w24462;
assign v7713 = ~(w24463 | w24464);
assign w24465 = v7713;
assign w24466 = w6389 & w20214;
assign w24467 = w6388 & w19952;
assign w24468 = w7004 & ~w19939;
assign v7714 = ~(w24467 | w24468);
assign w24469 = v7714;
assign w24470 = w6871 & w19954;
assign w24471 = w24469 & ~w24470;
assign w24472 = ~w24466 & w24471;
assign v7715 = ~(pi14 | w24472);
assign w24473 = v7715;
assign w24474 = pi14 & w24472;
assign v7716 = ~(w24473 | w24474);
assign w24475 = v7716;
assign w24476 = ~w24465 & w24475;
assign w24477 = w24465 & ~w24475;
assign v7717 = ~(w24476 | w24477);
assign w24478 = v7717;
assign w24479 = (~w24245 & ~w30445) | (~w24245 & w31222) | (~w30445 & w31222);
assign w24480 = w24478 & ~w24479;
assign w24481 = ~w24478 & w24479;
assign v7718 = ~(w24480 | w24481);
assign w24482 = v7718;
assign v7719 = ~(w24342 | w24482);
assign w24483 = v7719;
assign w24484 = w24342 & w24482;
assign v7720 = ~(w24483 | w24484);
assign w24485 = v7720;
assign w24486 = (~w24254 & ~w24109) | (~w24254 & w30093) | (~w24109 & w30093);
assign w24487 = w24485 & w24486;
assign v7721 = ~(w24485 | w24486);
assign w24488 = v7721;
assign v7722 = ~(w24487 | w24488);
assign w24489 = v7722;
assign v7723 = ~(w24331 | w24489);
assign w24490 = v7723;
assign w24491 = w24331 & w24489;
assign v7724 = ~(w24490 | w24491);
assign w24492 = v7724;
assign w24493 = (~w24260 & ~w24262) | (~w24260 & w29951) | (~w24262 & w29951);
assign w24494 = w24492 & w24493;
assign v7725 = ~(w24492 | w24493);
assign w24495 = v7725;
assign v7726 = ~(w24494 | w24495);
assign w24496 = v7726;
assign w24497 = w24322 & ~w24496;
assign w24498 = ~w24322 & w24496;
assign v7727 = ~(w24497 | w24498);
assign w24499 = v7727;
assign w24500 = w24274 & ~w24499;
assign w24501 = ~w24274 & w24499;
assign v7728 = ~(w24500 | w24501);
assign w24502 = v7728;
assign w24503 = ~w24277 & w24502;
assign w24504 = w24277 & ~w24502;
assign v7729 = ~(w24503 | w24504);
assign w24505 = v7729;
assign w24506 = ~w24311 & w24505;
assign w24507 = w24311 & ~w24505;
assign v7730 = ~(w24506 | w24507);
assign w24508 = v7730;
assign w24509 = (~w24294 & ~w24097) | (~w24294 & w28092) | (~w24097 & w28092);
assign w24510 = w24508 & w24509;
assign v7731 = ~(w24508 | w24509);
assign w24511 = v7731;
assign v7732 = ~(w24510 | w24511);
assign w24512 = v7732;
assign w24513 = w24300 & w24512;
assign v7733 = ~(w24300 | w24512);
assign w24514 = v7733;
assign v7734 = ~(w24513 | w24514);
assign w24515 = v7734;
assign w24516 = (~w24506 & w24509) | (~w24506 & w31223) | (w24509 & w31223);
assign w24517 = w10986 & w24284;
assign w24518 = pi02 & ~w24517;
assign w24519 = (~w24497 & ~w24501) | (~w24497 & w28429) | (~w24501 & w28429);
assign v7735 = ~(w24484 | w24487);
assign w24520 = v7735;
assign w24521 = w7466 & ~w19923;
assign w24522 = w7765 & w19917;
assign v7736 = ~(w24521 | w24522);
assign w24523 = v7736;
assign w24524 = w7177 & ~w19929;
assign w24525 = w24523 & ~w24524;
assign w24526 = (w24525 & w22895) | (w24525 & w28592) | (w22895 & w28592);
assign w24527 = pi11 & w24526;
assign v7737 = ~(pi11 | w24526);
assign w24528 = v7737;
assign v7738 = ~(w24527 | w24528);
assign w24529 = v7738;
assign v7739 = ~(w24477 | w24480);
assign w24530 = v7739;
assign w24531 = (~w24427 & w24344) | (~w24427 & w31119) | (w24344 & w31119);
assign v7740 = ~(w24411 | w24414);
assign w24532 = v7740;
assign v7741 = ~(w24395 | w24398);
assign w24533 = v7741;
assign v7742 = ~(w24379 | w24382);
assign w24534 = v7742;
assign v7743 = ~(w248 | w588);
assign w24535 = v7743;
assign w24536 = w1888 & w24535;
assign w24537 = w4210 & w24536;
assign w24538 = ~w652 & w24537;
assign w24539 = w2412 & w24538;
assign w24540 = w3807 & w24539;
assign w24541 = w14542 & w24540;
assign w24542 = w3200 & w4242;
assign w24543 = w1448 & w3579;
assign w24544 = w24542 & w24543;
assign w24545 = w1142 & w5218;
assign w24546 = w24544 & w24545;
assign w24547 = w5420 & w24546;
assign w24548 = w24541 & w24547;
assign w24549 = w928 & w20459;
assign w24550 = w3406 & ~w20011;
assign w24551 = w3402 & w20014;
assign w24552 = w3399 & ~w20028;
assign v7744 = ~(w24551 | w24552);
assign w24553 = v7744;
assign w24554 = ~w24550 & w24553;
assign w24555 = ~w24549 & w24554;
assign v7745 = ~(w24548 | w24555);
assign w24556 = v7745;
assign w24557 = w24548 & w24555;
assign v7746 = ~(w24556 | w24557);
assign w24558 = v7746;
assign w24559 = ~w24534 & w24558;
assign w24560 = w24534 & ~w24558;
assign v7747 = ~(w24559 | w24560);
assign w24561 = v7747;
assign w24562 = w3529 & w20681;
assign w24563 = w3760 & w20000;
assign w24564 = w3767 & ~w20008;
assign w24565 = w3763 & w20005;
assign v7748 = ~(w24564 | w24565);
assign w24566 = v7748;
assign w24567 = ~w24563 & w24566;
assign w24568 = ~w24562 & w24567;
assign w24569 = ~pi29 & w24568;
assign w24570 = pi29 & ~w24568;
assign v7749 = ~(w24569 | w24570);
assign w24571 = v7749;
assign w24572 = w24561 & w24571;
assign v7750 = ~(w24561 | w24571);
assign w24573 = v7750;
assign v7751 = ~(w24572 | w24573);
assign w24574 = v7751;
assign w24575 = ~w24533 & w24574;
assign w24576 = w24533 & ~w24574;
assign v7752 = ~(w24575 | w24576);
assign w24577 = v7752;
assign w24578 = w4153 & w20965;
assign w24579 = w4158 & ~w19992;
assign w24580 = w4155 & w19989;
assign v7753 = ~(w24579 | w24580);
assign w24581 = v7753;
assign v7754 = ~(w2873 | w19997);
assign w24582 = v7754;
assign w24583 = w24581 & ~w24582;
assign w24584 = ~w24578 & w24583;
assign w24585 = pi26 & w24584;
assign v7755 = ~(pi26 | w24584);
assign w24586 = v7755;
assign v7756 = ~(w24585 | w24586);
assign w24587 = v7756;
assign w24588 = w24577 & ~w24587;
assign w24589 = ~w24577 & w24587;
assign v7757 = ~(w24588 | w24589);
assign w24590 = v7757;
assign w24591 = ~w24532 & w24590;
assign w24592 = w24532 & ~w24590;
assign v7758 = ~(w24591 | w24592);
assign w24593 = v7758;
assign w24594 = w4764 & w20982;
assign w24595 = w4836 & w19983;
assign w24596 = w4913 & w19980;
assign v7759 = ~(w24595 | w24596);
assign w24597 = v7759;
assign w24598 = w4763 & w19986;
assign w24599 = w24597 & ~w24598;
assign w24600 = ~w24594 & w24599;
assign w24601 = pi23 & w24600;
assign v7760 = ~(pi23 | w24600);
assign w24602 = v7760;
assign v7761 = ~(w24601 | w24602);
assign w24603 = v7761;
assign w24604 = w24593 & ~w24603;
assign w24605 = ~w24593 & w24603;
assign v7762 = ~(w24604 | w24605);
assign w24606 = v7762;
assign w24607 = ~w24531 & w24606;
assign w24608 = w24531 & ~w24606;
assign v7763 = ~(w24607 | w24608);
assign w24609 = v7763;
assign w24610 = w5114 & w21385;
assign w24611 = w5531 & ~w19971;
assign w24612 = w5610 & w19966;
assign v7764 = ~(w24611 | w24612);
assign w24613 = v7764;
assign w24614 = w5113 & w19974;
assign w24615 = w24613 & ~w24614;
assign w24616 = ~w24610 & w24615;
assign w24617 = pi20 & w24616;
assign v7765 = ~(pi20 | w24616);
assign w24618 = v7765;
assign v7766 = ~(w24617 | w24618);
assign w24619 = v7766;
assign w24620 = ~w24609 & w24619;
assign w24621 = w24609 & ~w24619;
assign v7767 = ~(w24620 | w24621);
assign w24622 = v7767;
assign w24623 = (~w24443 & w24446) | (~w24443 & w30914) | (w24446 & w30914);
assign w24624 = w24622 & ~w24623;
assign w24625 = ~w24622 & w24623;
assign v7768 = ~(w24624 | w24625);
assign w24626 = v7768;
assign w24627 = w5765 & ~w21882;
assign w24628 = w5983 & w19958;
assign w24629 = w6236 & w19952;
assign v7769 = ~(w24628 | w24629);
assign w24630 = v7769;
assign w24631 = w5764 & w19961;
assign w24632 = w24630 & ~w24631;
assign w24633 = ~w24627 & w24632;
assign w24634 = pi17 & w24633;
assign v7770 = ~(pi17 | w24633);
assign w24635 = v7770;
assign v7771 = ~(w24634 | w24635);
assign w24636 = v7771;
assign w24637 = w24626 & ~w24636;
assign w24638 = ~w24626 & w24636;
assign v7772 = ~(w24637 | w24638);
assign w24639 = v7772;
assign w24640 = (~w24461 & ~w30731) | (~w24461 & w30915) | (~w30731 & w30915);
assign v7773 = ~(w24639 | w24640);
assign w24641 = v7773;
assign w24642 = w24639 & w24640;
assign v7774 = ~(w24641 | w24642);
assign w24643 = v7774;
assign w24644 = w6389 & ~w22304;
assign w24645 = w7004 & w19933;
assign w24646 = w6388 & w19954;
assign w24647 = w6871 & ~w19939;
assign v7775 = ~(w24646 | w24647);
assign w24648 = v7775;
assign w24649 = ~w24645 & w24648;
assign w24650 = ~w24644 & w24649;
assign w24651 = ~pi14 & w24650;
assign w24652 = pi14 & ~w24650;
assign v7776 = ~(w24651 | w24652);
assign w24653 = v7776;
assign w24654 = w24643 & w24653;
assign v7777 = ~(w24643 | w24653);
assign w24655 = v7777;
assign v7778 = ~(w24654 | w24655);
assign w24656 = v7778;
assign v7779 = ~(w24530 | w24656);
assign w24657 = v7779;
assign w24658 = w24530 & w24656;
assign v7780 = ~(w24657 | w24658);
assign w24659 = v7780;
assign v7781 = ~(w24529 | w24659);
assign w24660 = v7781;
assign w24661 = w24529 & w24659;
assign v7782 = ~(w24660 | w24661);
assign w24662 = v7782;
assign w24663 = ~w24520 & w24662;
assign w24664 = w24520 & ~w24662;
assign v7783 = ~(w24663 | w24664);
assign w24665 = v7783;
assign w24666 = w8926 & w20197;
assign w24667 = w8140 & w19853;
assign w24668 = w8526 & ~w19912;
assign v7784 = ~(w24667 | w24668);
assign w24669 = v7784;
assign w24670 = ~w24666 & w24669;
assign w24671 = (~w20203 & w28593) | (~w20203 & w28594) | (w28593 & w28594);
assign w24672 = (w20203 & w28595) | (w20203 & w28596) | (w28595 & w28596);
assign v7785 = ~(w24671 | w24672);
assign w24673 = v7785;
assign w24674 = ~w24665 & w24673;
assign w24675 = w24665 & ~w24673;
assign v7786 = ~(w24674 | w24675);
assign w24676 = v7786;
assign w24677 = (~w24490 & ~w24492) | (~w24490 & w28597) | (~w24492 & w28597);
assign w24678 = w24676 & w24677;
assign v7787 = ~(w24676 | w24677);
assign w24679 = v7787;
assign v7788 = ~(w24678 | w24679);
assign w24680 = v7788;
assign w24681 = w9402 & w24073;
assign w24682 = w9401 & w23607;
assign w24683 = w10419 & ~w24077;
assign v7789 = ~(w24682 | w24683);
assign w24684 = v7789;
assign w24685 = w9891 & w23670;
assign w24686 = w24684 & ~w24685;
assign w24687 = ~w24681 & w24686;
assign v7790 = ~(pi05 | w24687);
assign w24688 = v7790;
assign w24689 = pi05 & w24687;
assign v7791 = ~(w24688 | w24689);
assign w24690 = v7791;
assign w24691 = w24680 & ~w24690;
assign w24692 = ~w24680 & w24690;
assign v7792 = ~(w24691 | w24692);
assign w24693 = v7792;
assign w24694 = w24519 & ~w24693;
assign w24695 = ~w24519 & w24693;
assign v7793 = ~(w24694 | w24695);
assign w24696 = v7793;
assign w24697 = w24518 & w24696;
assign v7794 = ~(w24518 | w24696);
assign w24698 = v7794;
assign v7795 = ~(w24697 | w24698);
assign w24699 = v7795;
assign v7796 = ~(w24516 | w24699);
assign w24700 = v7796;
assign w24701 = w24516 & w24699;
assign v7797 = ~(w24700 | w24701);
assign w24702 = v7797;
assign w24703 = w24513 & w24702;
assign v7798 = ~(w24513 | w24702);
assign w24704 = v7798;
assign v7799 = ~(w24703 | w24704);
assign w24705 = v7799;
assign w24706 = w10445 & w24282;
assign w24707 = w10419 & w24284;
assign w24708 = w9401 & w23670;
assign w24709 = w9891 & ~w24077;
assign v7800 = ~(w24708 | w24709);
assign w24710 = v7800;
assign w24711 = ~w24707 & w24710;
assign w24712 = pi05 & ~w24711;
assign w24713 = w9402 & w24282;
assign w24714 = ~pi05 & w24711;
assign w24715 = ~w24713 & w24714;
assign v7801 = ~(w24712 | w24715);
assign w24716 = v7801;
assign w24717 = ~w24706 & w24716;
assign v7802 = ~(pi02 | w24717);
assign w24718 = v7802;
assign w24719 = pi02 & w24717;
assign v7803 = ~(w24718 | w24719);
assign w24720 = v7803;
assign v7804 = ~(w24675 | w24678);
assign w24721 = v7804;
assign v7805 = ~(w24660 | w24663);
assign w24722 = v7805;
assign w24723 = w7178 & w22936;
assign w24724 = w7466 & w19917;
assign w24725 = w7765 & w19853;
assign v7806 = ~(w24724 | w24725);
assign w24726 = v7806;
assign w24727 = w7177 & ~w19923;
assign w24728 = w24726 & ~w24727;
assign w24729 = ~w24723 & w24728;
assign w24730 = pi11 & w24729;
assign v7807 = ~(pi11 | w24729);
assign w24731 = v7807;
assign v7808 = ~(w24730 | w24731);
assign w24732 = v7808;
assign v7809 = ~(w24637 | w24642);
assign w24733 = v7809;
assign w24734 = w5765 & ~w21866;
assign w24735 = w6236 & w19954;
assign w24736 = w5764 & w19958;
assign w24737 = w5983 & w19952;
assign v7810 = ~(w24736 | w24737);
assign w24738 = v7810;
assign w24739 = ~w24735 & w24738;
assign w24740 = ~w24734 & w24739;
assign w24741 = ~pi17 & w24740;
assign w24742 = pi17 & ~w24740;
assign v7811 = ~(w24741 | w24742);
assign w24743 = v7811;
assign v7812 = ~(w24621 | w24624);
assign w24744 = v7812;
assign v7813 = ~(w24604 | w24607);
assign w24745 = v7813;
assign v7814 = ~(w24588 | w24591);
assign w24746 = v7814;
assign v7815 = ~(w24572 | w24575);
assign w24747 = v7815;
assign v7816 = ~(w24556 | w24559);
assign w24748 = v7816;
assign w24749 = ~w103 & w2180;
assign w24750 = ~w753 & w24749;
assign w24751 = w24147 & w24750;
assign w24752 = ~w405 & w1409;
assign w24753 = ~w272 & w24752;
assign w24754 = w13292 & w24753;
assign w24755 = w24751 & w24754;
assign w24756 = w3019 & w13675;
assign w24757 = ~w202 & w399;
assign w24758 = w2053 & w24757;
assign w24759 = ~w438 & w649;
assign w24760 = w1242 & w24759;
assign w24761 = w24758 & w24760;
assign w24762 = w894 & w1470;
assign w24763 = w1396 & w1574;
assign w24764 = w24762 & w24763;
assign w24765 = w2277 & w24357;
assign w24766 = w24764 & w24765;
assign w24767 = w24761 & w24766;
assign w24768 = w5194 & w24767;
assign w24769 = w24756 & w24768;
assign w24770 = w24755 & w24769;
assign w24771 = w928 & w20446;
assign w24772 = w3406 & ~w20008;
assign w24773 = w3402 & ~w20011;
assign w24774 = w3399 & w20014;
assign v7817 = ~(w24773 | w24774);
assign w24775 = v7817;
assign w24776 = ~w24772 & w24775;
assign w24777 = ~w24771 & w24776;
assign v7818 = ~(w24770 | w24777);
assign w24778 = v7818;
assign w24779 = w24770 & w24777;
assign v7819 = ~(w24778 | w24779);
assign w24780 = v7819;
assign w24781 = ~w24748 & w24780;
assign w24782 = w24748 & ~w24780;
assign v7820 = ~(w24781 | w24782);
assign w24783 = v7820;
assign w24784 = w3529 & w20668;
assign w24785 = w3760 & ~w19997;
assign w24786 = w3767 & w20005;
assign w24787 = w3763 & w20000;
assign v7821 = ~(w24786 | w24787);
assign w24788 = v7821;
assign w24789 = ~w24785 & w24788;
assign w24790 = ~w24784 & w24789;
assign w24791 = ~pi29 & w24790;
assign w24792 = pi29 & ~w24790;
assign v7822 = ~(w24791 | w24792);
assign w24793 = v7822;
assign w24794 = w24783 & w24793;
assign v7823 = ~(w24783 | w24793);
assign w24795 = v7823;
assign v7824 = ~(w24794 | w24795);
assign w24796 = v7824;
assign w24797 = ~w24747 & w24796;
assign w24798 = w24747 & ~w24796;
assign v7825 = ~(w24797 | w24798);
assign w24799 = v7825;
assign w24800 = w4153 & w21012;
assign w24801 = w4155 & w19986;
assign v7826 = ~(w2873 | w19992);
assign w24802 = v7826;
assign w24803 = w4158 & w19989;
assign v7827 = ~(w24802 | w24803);
assign w24804 = v7827;
assign w24805 = ~w24801 & w24804;
assign w24806 = ~w24800 & w24805;
assign w24807 = ~pi26 & w24806;
assign w24808 = pi26 & ~w24806;
assign v7828 = ~(w24807 | w24808);
assign w24809 = v7828;
assign w24810 = w24799 & w24809;
assign v7829 = ~(w24799 | w24809);
assign w24811 = v7829;
assign v7830 = ~(w24810 | w24811);
assign w24812 = v7830;
assign w24813 = ~w24746 & w24812;
assign w24814 = w24746 & ~w24812;
assign v7831 = ~(w24813 | w24814);
assign w24815 = v7831;
assign w24816 = w4764 & w21362;
assign w24817 = w4836 & w19980;
assign w24818 = w4913 & w19974;
assign v7832 = ~(w24817 | w24818);
assign w24819 = v7832;
assign w24820 = w4763 & w19983;
assign w24821 = w24819 & ~w24820;
assign w24822 = ~w24816 & w24821;
assign w24823 = pi23 & w24822;
assign v7833 = ~(pi23 | w24822);
assign w24824 = v7833;
assign v7834 = ~(w24823 | w24824);
assign w24825 = v7834;
assign w24826 = w24815 & ~w24825;
assign w24827 = ~w24815 & w24825;
assign v7835 = ~(w24826 | w24827);
assign w24828 = v7835;
assign w24829 = ~w24745 & w24828;
assign w24830 = w24745 & ~w24828;
assign v7836 = ~(w24829 | w24830);
assign w24831 = v7836;
assign w24832 = w5114 & w20234;
assign w24833 = w5531 & w19966;
assign w24834 = w5610 & w19961;
assign v7837 = ~(w24833 | w24834);
assign w24835 = v7837;
assign w24836 = w5113 & ~w19971;
assign w24837 = w24835 & ~w24836;
assign w24838 = ~w24832 & w24837;
assign w24839 = pi20 & w24838;
assign v7838 = ~(pi20 | w24838);
assign w24840 = v7838;
assign v7839 = ~(w24839 | w24840);
assign w24841 = v7839;
assign w24842 = w24831 & ~w24841;
assign w24843 = ~w24831 & w24841;
assign v7840 = ~(w24842 | w24843);
assign w24844 = v7840;
assign w24845 = w24744 & w24844;
assign v7841 = ~(w24744 | w24844);
assign w24846 = v7841;
assign v7842 = ~(w24845 | w24846);
assign w24847 = v7842;
assign w24848 = w24743 & ~w24847;
assign w24849 = ~w24743 & w24847;
assign v7843 = ~(w24848 | w24849);
assign w24850 = v7843;
assign w24851 = ~w24733 & w24850;
assign w24852 = w24733 & ~w24850;
assign v7844 = ~(w24851 | w24852);
assign w24853 = v7844;
assign w24854 = w6389 & ~w22285;
assign w24855 = w7004 & ~w19929;
assign w24856 = w6388 & ~w19939;
assign w24857 = w6871 & w19933;
assign v7845 = ~(w24856 | w24857);
assign w24858 = v7845;
assign w24859 = ~w24855 & w24858;
assign w24860 = ~w24854 & w24859;
assign w24861 = ~pi14 & w24860;
assign w24862 = pi14 & ~w24860;
assign v7846 = ~(w24861 | w24862);
assign w24863 = v7846;
assign w24864 = w24853 & w24863;
assign v7847 = ~(w24853 | w24863);
assign w24865 = v7847;
assign v7848 = ~(w24864 | w24865);
assign w24866 = v7848;
assign v7849 = ~(w24530 | w24655);
assign w24867 = v7849;
assign v7850 = ~(w24654 | w24867);
assign w24868 = v7850;
assign w24869 = w24866 & w24868;
assign v7851 = ~(w24866 | w24868);
assign w24870 = v7851;
assign v7852 = ~(w24869 | w24870);
assign w24871 = v7852;
assign w24872 = w24732 & w24871;
assign v7853 = ~(w24732 | w24871);
assign w24873 = v7853;
assign v7854 = ~(w24872 | w24873);
assign w24874 = v7854;
assign w24875 = w24722 & w24874;
assign v7855 = ~(w24722 | w24874);
assign w24876 = v7855;
assign v7856 = ~(w24875 | w24876);
assign w24877 = v7856;
assign w24878 = w8141 & w23614;
assign w24879 = w8526 & w20197;
assign w24880 = w8926 & w23607;
assign v7857 = ~(w24879 | w24880);
assign w24881 = v7857;
assign w24882 = w8140 & ~w19912;
assign w24883 = w24881 & ~w24882;
assign w24884 = ~w24878 & w24883;
assign w24885 = pi08 & w24884;
assign v7858 = ~(pi08 | w24884);
assign w24886 = v7858;
assign v7859 = ~(w24885 | w24886);
assign w24887 = v7859;
assign w24888 = w24877 & w24887;
assign v7860 = ~(w24877 | w24887);
assign w24889 = v7860;
assign v7861 = ~(w24888 | w24889);
assign w24890 = v7861;
assign w24891 = ~w24721 & w24890;
assign w24892 = w24721 & ~w24890;
assign v7862 = ~(w24891 | w24892);
assign w24893 = v7862;
assign w24894 = w24720 & w24893;
assign v7863 = ~(w24720 | w24893);
assign w24895 = v7863;
assign v7864 = ~(w24894 | w24895);
assign w24896 = v7864;
assign w24897 = w24519 & ~w24691;
assign v7865 = ~(w24692 | w24897);
assign w24898 = v7865;
assign v7866 = ~(w24896 | w24898);
assign w24899 = v7866;
assign w24900 = w24896 & w24898;
assign v7867 = ~(w24899 | w24900);
assign w24901 = v7867;
assign w24902 = (~w28431 & w31224) | (~w28431 & w31225) | (w31224 & w31225);
assign w24903 = (w28431 & w31226) | (w28431 & w31227) | (w31226 & w31227);
assign v7868 = ~(w24902 | w24903);
assign w24904 = v7868;
assign w24905 = w24703 & ~w24904;
assign w24906 = ~w24703 & w24904;
assign v7869 = ~(w24905 | w24906);
assign w24907 = v7869;
assign v7870 = ~(w24719 | w24894);
assign w24908 = v7870;
assign v7871 = ~(w24889 | w24891);
assign w24909 = v7871;
assign w24910 = w9402 & ~w24304;
assign w24911 = w9891 & w24284;
assign w24912 = w9401 & ~w24077;
assign v7872 = ~(w24911 | w24912);
assign w24913 = v7872;
assign w24914 = ~w24910 & w24913;
assign w24915 = ~pi05 & w24914;
assign w24916 = pi05 & ~w24914;
assign v7873 = ~(w24915 | w24916);
assign w24917 = v7873;
assign w24918 = ~w24909 & w24917;
assign w24919 = w24909 & ~w24917;
assign v7874 = ~(w24918 | w24919);
assign w24920 = v7874;
assign w24921 = w5765 & w20214;
assign w24922 = w5983 & w19954;
assign w24923 = w6236 & ~w19939;
assign v7875 = ~(w24922 | w24923);
assign w24924 = v7875;
assign w24925 = w5764 & w19952;
assign w24926 = w24924 & ~w24925;
assign w24927 = ~w24921 & w24926;
assign w24928 = pi17 & w24927;
assign v7876 = ~(pi17 | w24927);
assign w24929 = v7876;
assign v7877 = ~(w24928 | w24929);
assign w24930 = v7877;
assign w24931 = w24744 & ~w24842;
assign v7878 = ~(w24843 | w24931);
assign w24932 = v7878;
assign w24933 = ~w24930 & w24932;
assign w24934 = w24930 & ~w24932;
assign v7879 = ~(w24933 | w24934);
assign w24935 = v7879;
assign v7880 = ~(w24826 | w24829);
assign w24936 = v7880;
assign v7881 = ~(w24810 | w24813);
assign w24937 = v7881;
assign w24938 = (~w24778 & w24748) | (~w24778 & w31228) | (w24748 & w31228);
assign w24939 = w1113 & w4013;
assign w24940 = w3095 & w24939;
assign w24941 = w6719 & w12565;
assign w24942 = w1201 & w3060;
assign w24943 = w3271 & w24942;
assign w24944 = w2793 & w24943;
assign w24945 = w24941 & w24944;
assign v7882 = ~(w159 | w812);
assign w24946 = v7882;
assign w24947 = ~w427 & w24946;
assign w24948 = ~w267 & w13118;
assign w24949 = w24947 & w24948;
assign w24950 = w13144 & w24949;
assign w24951 = w24945 & w24950;
assign w24952 = w757 & w24951;
assign w24953 = w24940 & w24952;
assign w24954 = w3877 & w24953;
assign w24955 = w3406 & w20005;
assign w24956 = w3399 & ~w20011;
assign w24957 = w3402 & ~w20008;
assign v7883 = ~(w24956 | w24957);
assign w24958 = v7883;
assign w24959 = ~w24955 & w24958;
assign w24960 = (w24959 & ~w31120) | (w24959 & w31229) | (~w31120 & w31229);
assign w24961 = w24954 & w24960;
assign v7884 = ~(w24954 | w24960);
assign w24962 = v7884;
assign v7885 = ~(w24961 | w24962);
assign w24963 = v7885;
assign w24964 = ~pi02 & w24963;
assign w24965 = pi02 & ~w24963;
assign v7886 = ~(w24964 | w24965);
assign w24966 = v7886;
assign v7887 = ~(w24938 | w24966);
assign w24967 = v7887;
assign w24968 = w24938 & w24966;
assign v7888 = ~(w24967 | w24968);
assign w24969 = v7888;
assign w24970 = w3529 & w20655;
assign w24971 = w3760 & ~w19992;
assign w24972 = w3763 & ~w19997;
assign w24973 = w3767 & w20000;
assign v7889 = ~(w24972 | w24973);
assign w24974 = v7889;
assign w24975 = ~w24971 & w24974;
assign w24976 = ~w24970 & w24975;
assign w24977 = ~pi29 & w24976;
assign w24978 = pi29 & ~w24976;
assign v7890 = ~(w24977 | w24978);
assign w24979 = v7890;
assign w24980 = w24969 & w24979;
assign v7891 = ~(w24969 | w24979);
assign w24981 = v7891;
assign v7892 = ~(w24980 | w24981);
assign w24982 = v7892;
assign v7893 = ~(w24794 | w24797);
assign w24983 = v7893;
assign w24984 = w4153 & w20997;
assign w24985 = w4155 & w19983;
assign w24986 = ~w2873 & w19989;
assign w24987 = w4158 & w19986;
assign v7894 = ~(w24986 | w24987);
assign w24988 = v7894;
assign w24989 = ~w24985 & w24988;
assign w24990 = ~w24984 & w24989;
assign w24991 = ~pi26 & w24990;
assign w24992 = pi26 & ~w24990;
assign v7895 = ~(w24991 | w24992);
assign w24993 = v7895;
assign w24994 = w24983 & ~w24993;
assign w24995 = ~w24983 & w24993;
assign v7896 = ~(w24994 | w24995);
assign w24996 = v7896;
assign w24997 = ~w24982 & w24996;
assign w24998 = w24982 & ~w24996;
assign v7897 = ~(w24997 | w24998);
assign w24999 = v7897;
assign v7898 = ~(w24937 | w24999);
assign w25000 = v7898;
assign w25001 = w24937 & w24999;
assign v7899 = ~(w25000 | w25001);
assign w25002 = v7899;
assign w25003 = w4764 & w21401;
assign w25004 = w4836 & w19974;
assign w25005 = w4913 & ~w19971;
assign v7900 = ~(w25004 | w25005);
assign w25006 = v7900;
assign w25007 = w4763 & w19980;
assign w25008 = w25006 & ~w25007;
assign w25009 = ~w25003 & w25008;
assign w25010 = pi23 & w25009;
assign v7901 = ~(pi23 | w25009);
assign w25011 = v7901;
assign v7902 = ~(w25010 | w25011);
assign w25012 = v7902;
assign w25013 = w25002 & ~w25012;
assign w25014 = ~w25002 & w25012;
assign v7903 = ~(w25013 | w25014);
assign w25015 = v7903;
assign w25016 = ~w24936 & w25015;
assign w25017 = w24936 & ~w25015;
assign v7904 = ~(w25016 | w25017);
assign w25018 = v7904;
assign w25019 = w5114 & w21716;
assign w25020 = w5610 & w19958;
assign w25021 = w5531 & w19961;
assign w25022 = w5113 & w19966;
assign v7905 = ~(w25021 | w25022);
assign w25023 = v7905;
assign w25024 = ~w25020 & w25023;
assign w25025 = ~w25019 & w25024;
assign w25026 = ~pi20 & w25025;
assign w25027 = pi20 & ~w25025;
assign v7906 = ~(w25026 | w25027);
assign w25028 = v7906;
assign w25029 = w25018 & w25028;
assign v7907 = ~(w25018 | w25028);
assign w25030 = v7907;
assign v7908 = ~(w25029 | w25030);
assign w25031 = v7908;
assign w25032 = ~w24935 & w25031;
assign w25033 = w24935 & ~w25031;
assign v7909 = ~(w25032 | w25033);
assign w25034 = v7909;
assign v7910 = ~(w24848 | w24851);
assign w25035 = v7910;
assign w25036 = w25034 & w25035;
assign v7911 = ~(w25034 | w25035);
assign w25037 = v7911;
assign v7912 = ~(w25036 | w25037);
assign w25038 = v7912;
assign w25039 = w6389 & w22262;
assign w25040 = w7004 & ~w19923;
assign w25041 = w6388 & w19933;
assign w25042 = w6871 & ~w19929;
assign v7913 = ~(w25041 | w25042);
assign w25043 = v7913;
assign w25044 = ~w25040 & w25043;
assign w25045 = ~w25039 & w25044;
assign w25046 = ~pi14 & w25045;
assign w25047 = pi14 & ~w25045;
assign v7914 = ~(w25046 | w25047);
assign w25048 = v7914;
assign w25049 = ~w25038 & w25048;
assign w25050 = w25038 & ~w25048;
assign v7915 = ~(w25049 | w25050);
assign w25051 = v7915;
assign w25052 = w7466 & w19853;
assign w25053 = w7765 & ~w19912;
assign v7916 = ~(w25052 | w25053);
assign w25054 = v7916;
assign w25055 = w7177 & w19917;
assign w25056 = w25054 & ~w25055;
assign w25057 = (~w22917 & w28844) | (~w22917 & w28845) | (w28844 & w28845);
assign w25058 = (w22917 & w28846) | (w22917 & w28847) | (w28846 & w28847);
assign v7917 = ~(w25057 | w25058);
assign w25059 = v7917;
assign w25060 = ~w24864 & w24868;
assign v7918 = ~(w24865 | w25060);
assign w25061 = v7918;
assign w25062 = ~w25059 & w25061;
assign w25063 = w25059 & ~w25061;
assign v7919 = ~(w25062 | w25063);
assign w25064 = v7919;
assign w25065 = w25051 & ~w25064;
assign w25066 = ~w25051 & w25064;
assign v7920 = ~(w25065 | w25066);
assign w25067 = v7920;
assign w25068 = w8141 & w23666;
assign w25069 = w8140 & w20197;
assign w25070 = w8926 & w23670;
assign v7921 = ~(w25069 | w25070);
assign w25071 = v7921;
assign w25072 = w8526 & w23607;
assign w25073 = w25071 & ~w25072;
assign w25074 = ~w25068 & w25073;
assign v7922 = ~(pi08 | w25074);
assign w25075 = v7922;
assign w25076 = pi08 & w25074;
assign v7923 = ~(w25075 | w25076);
assign w25077 = v7923;
assign w25078 = w25067 & ~w25077;
assign w25079 = ~w25067 & w25077;
assign v7924 = ~(w25078 | w25079);
assign w25080 = v7924;
assign v7925 = ~(w24872 | w24875);
assign w25081 = v7925;
assign w25082 = ~w25080 & w25081;
assign w25083 = w25080 & ~w25081;
assign v7926 = ~(w25082 | w25083);
assign w25084 = v7926;
assign w25085 = w24920 & ~w25084;
assign w25086 = ~w24920 & w25084;
assign v7927 = ~(w25085 | w25086);
assign w25087 = v7927;
assign w25088 = w24908 & ~w25087;
assign w25089 = ~w24908 & w25087;
assign v7928 = ~(w25088 | w25089);
assign w25090 = v7928;
assign w25091 = (~w24701 & w28094) | (~w24701 & w28095) | (w28094 & w28095);
assign w25092 = ~w25090 & w25091;
assign w25093 = w25090 & ~w25091;
assign v7929 = ~(w25092 | w25093);
assign w25094 = v7929;
assign w25095 = w24905 & w25094;
assign v7930 = ~(w24905 | w25094);
assign w25096 = v7930;
assign v7931 = ~(w25095 | w25096);
assign w25097 = v7931;
assign v7932 = ~(w24918 | w25085);
assign w25098 = v7932;
assign w25099 = w9400 & w24284;
assign v7933 = ~(pi05 | w25099);
assign w25100 = v7933;
assign w25101 = w13696 & w24284;
assign v7934 = ~(w25100 | w25101);
assign w25102 = v7934;
assign v7935 = ~(w25062 | w25066);
assign w25103 = v7935;
assign v7936 = ~(w25036 | w25050);
assign w25104 = v7936;
assign w25105 = w7765 & w20197;
assign w25106 = w7177 & w19853;
assign w25107 = w7466 & ~w19912;
assign v7937 = ~(w25106 | w25107);
assign w25108 = v7937;
assign w25109 = ~w25105 & w25108;
assign w25110 = (~w20203 & w28433) | (~w20203 & w28434) | (w28433 & w28434);
assign w25111 = (w20203 & w28435) | (w20203 & w28436) | (w28435 & w28436);
assign v7938 = ~(w25110 | w25111);
assign w25112 = v7938;
assign v7939 = ~(w24967 | w24980);
assign w25113 = v7939;
assign v7940 = ~(pi02 | w24962);
assign w25114 = v7940;
assign w25115 = pi02 & ~w24961;
assign v7941 = ~(w25114 | w25115);
assign w25116 = v7941;
assign v7942 = ~(w56 | w288);
assign w25117 = v7942;
assign w25118 = w2915 & w25117;
assign w25119 = w346 & w25118;
assign w25120 = w2179 & w25119;
assign v7943 = ~(w77 | w176);
assign w25121 = v7943;
assign w25122 = w1154 & w1974;
assign w25123 = w893 & w3947;
assign w25124 = w25122 & w25123;
assign w25125 = w1465 & w21267;
assign w25126 = w25124 & w25125;
assign w25127 = w25121 & w25126;
assign w25128 = w233 & w3051;
assign w25129 = w3223 & w25128;
assign w25130 = w1503 & w25129;
assign w25131 = w2207 & w25130;
assign w25132 = w25127 & w25131;
assign w25133 = w25120 & w25132;
assign w25134 = w2756 & w25133;
assign w25135 = w14605 & w25134;
assign w25136 = w25116 & w25135;
assign v7944 = ~(w25116 | w25135);
assign w25137 = v7944;
assign v7945 = ~(w25136 | w25137);
assign w25138 = v7945;
assign w25139 = w928 & w20681;
assign w25140 = w3406 & w20000;
assign w25141 = w3399 & ~w20008;
assign w25142 = w3402 & w20005;
assign v7946 = ~(w25141 | w25142);
assign w25143 = v7946;
assign w25144 = ~w25140 & w25143;
assign w25145 = ~w25139 & w25144;
assign v7947 = ~(w25138 | w25145);
assign w25146 = v7947;
assign w25147 = w25138 & w25145;
assign v7948 = ~(w25146 | w25147);
assign w25148 = v7948;
assign w25149 = ~w25113 & w25148;
assign w25150 = w25113 & ~w25148;
assign v7949 = ~(w25149 | w25150);
assign w25151 = v7949;
assign w25152 = w4153 & w20982;
assign w25153 = w4155 & w19980;
assign w25154 = ~w2873 & w19986;
assign w25155 = w4158 & w19983;
assign v7950 = ~(w25154 | w25155);
assign w25156 = v7950;
assign w25157 = ~w25153 & w25156;
assign w25158 = ~w25152 & w25157;
assign w25159 = ~pi26 & w25158;
assign w25160 = pi26 & ~w25158;
assign v7951 = ~(w25159 | w25160);
assign w25161 = v7951;
assign w25162 = w3529 & w20965;
assign w25163 = w3760 & w19989;
assign w25164 = w3767 & ~w19997;
assign w25165 = w3763 & ~w19992;
assign v7952 = ~(w25164 | w25165);
assign w25166 = v7952;
assign w25167 = ~w25163 & w25166;
assign w25168 = ~w25162 & w25167;
assign w25169 = ~pi29 & w25168;
assign w25170 = pi29 & ~w25168;
assign v7953 = ~(w25169 | w25170);
assign w25171 = v7953;
assign v7954 = ~(w25161 | w25171);
assign w25172 = v7954;
assign w25173 = w25161 & w25171;
assign v7955 = ~(w25172 | w25173);
assign w25174 = v7955;
assign w25175 = w25151 & ~w25174;
assign w25176 = ~w25151 & w25174;
assign v7956 = ~(w25175 | w25176);
assign w25177 = v7956;
assign v7957 = ~(w24994 | w24997);
assign w25178 = v7957;
assign w25179 = w4764 & w21385;
assign w25180 = w4836 & ~w19971;
assign w25181 = w4913 & w19966;
assign v7958 = ~(w25180 | w25181);
assign w25182 = v7958;
assign w25183 = w4763 & w19974;
assign w25184 = w25182 & ~w25183;
assign w25185 = ~w25179 & w25184;
assign w25186 = pi23 & w25185;
assign v7959 = ~(pi23 | w25185);
assign w25187 = v7959;
assign v7960 = ~(w25186 | w25187);
assign w25188 = v7960;
assign w25189 = w25178 & ~w25188;
assign w25190 = ~w25178 & w25188;
assign v7961 = ~(w25189 | w25190);
assign w25191 = v7961;
assign w25192 = ~w25177 & w25191;
assign w25193 = w25177 & ~w25191;
assign v7962 = ~(w25192 | w25193);
assign w25194 = v7962;
assign v7963 = ~(w25000 | w25013);
assign w25195 = v7963;
assign w25196 = w5114 & ~w21882;
assign w25197 = w5531 & w19958;
assign w25198 = w5610 & w19952;
assign v7964 = ~(w25197 | w25198);
assign w25199 = v7964;
assign w25200 = w5113 & w19961;
assign w25201 = w25199 & ~w25200;
assign w25202 = ~w25196 & w25201;
assign w25203 = pi20 & w25202;
assign v7965 = ~(pi20 | w25202);
assign w25204 = v7965;
assign v7966 = ~(w25203 | w25204);
assign w25205 = v7966;
assign w25206 = w25195 & w25205;
assign v7967 = ~(w25195 | w25205);
assign w25207 = v7967;
assign v7968 = ~(w25206 | w25207);
assign w25208 = v7968;
assign w25209 = ~w25194 & w25208;
assign w25210 = w25194 & ~w25208;
assign v7969 = ~(w25209 | w25210);
assign w25211 = v7969;
assign v7970 = ~(w25016 | w25029);
assign w25212 = v7970;
assign w25213 = w5765 & ~w22304;
assign w25214 = w6236 & w19933;
assign w25215 = w5764 & w19954;
assign w25216 = w5983 & ~w19939;
assign v7971 = ~(w25215 | w25216);
assign w25217 = v7971;
assign w25218 = ~w25214 & w25217;
assign w25219 = ~w25213 & w25218;
assign w25220 = pi17 & w25219;
assign v7972 = ~(pi17 | w25219);
assign w25221 = v7972;
assign v7973 = ~(w25220 | w25221);
assign w25222 = v7973;
assign w25223 = w25212 & w25222;
assign v7974 = ~(w25212 | w25222);
assign w25224 = v7974;
assign v7975 = ~(w25223 | w25224);
assign w25225 = v7975;
assign w25226 = w25211 & w25225;
assign v7976 = ~(w25211 | w25225);
assign w25227 = v7976;
assign v7977 = ~(w25226 | w25227);
assign w25228 = v7977;
assign v7978 = ~(w24934 | w25033);
assign w25229 = v7978;
assign w25230 = ~w25228 & w25229;
assign w25231 = w25228 & ~w25229;
assign v7979 = ~(w25230 | w25231);
assign w25232 = v7979;
assign w25233 = w6389 & ~w22895;
assign w25234 = w7004 & w19917;
assign w25235 = w6388 & ~w19929;
assign w25236 = w6871 & ~w19923;
assign v7980 = ~(w25235 | w25236);
assign w25237 = v7980;
assign w25238 = ~w25234 & w25237;
assign w25239 = ~w25233 & w25238;
assign w25240 = ~pi14 & w25239;
assign w25241 = pi14 & ~w25239;
assign v7981 = ~(w25240 | w25241);
assign w25242 = v7981;
assign w25243 = w25232 & ~w25242;
assign w25244 = ~w25232 & w25242;
assign v7982 = ~(w25243 | w25244);
assign w25245 = v7982;
assign w25246 = ~w25112 & w25245;
assign w25247 = w25112 & ~w25245;
assign v7983 = ~(w25246 | w25247);
assign w25248 = v7983;
assign w25249 = w25104 & ~w25248;
assign w25250 = ~w25104 & w25248;
assign v7984 = ~(w25249 | w25250);
assign w25251 = v7984;
assign v7985 = ~(w25103 | w25251);
assign w25252 = v7985;
assign w25253 = w25103 & w25251;
assign v7986 = ~(w25252 | w25253);
assign w25254 = v7986;
assign w25255 = w8141 & w24073;
assign w25256 = w8526 & w23670;
assign w25257 = w8926 & ~w24077;
assign v7987 = ~(w25256 | w25257);
assign w25258 = v7987;
assign w25259 = w8140 & w23607;
assign w25260 = w25258 & ~w25259;
assign w25261 = ~w25255 & w25260;
assign v7988 = ~(pi08 | w25261);
assign w25262 = v7988;
assign w25263 = pi08 & w25261;
assign v7989 = ~(w25262 | w25263);
assign w25264 = v7989;
assign w25265 = w25254 & w25264;
assign v7990 = ~(w25254 | w25264);
assign w25266 = v7990;
assign v7991 = ~(w25265 | w25266);
assign w25267 = v7991;
assign w25268 = w25102 & ~w25267;
assign w25269 = ~w25102 & w25267;
assign v7992 = ~(w25268 | w25269);
assign w25270 = v7992;
assign v7993 = ~(w25079 | w25083);
assign w25271 = v7993;
assign w25272 = w25270 & w25271;
assign v7994 = ~(w25270 | w25271);
assign w25273 = v7994;
assign v7995 = ~(w25272 | w25273);
assign w25274 = v7995;
assign w25275 = w25098 & ~w25274;
assign w25276 = ~w25098 & w25274;
assign v7996 = ~(w25275 | w25276);
assign w25277 = v7996;
assign w25278 = (~w25089 & w25091) | (~w25089 & w28096) | (w25091 & w28096);
assign w25279 = ~w25277 & w25278;
assign w25280 = w25277 & ~w25278;
assign v7997 = ~(w25279 | w25280);
assign w25281 = v7997;
assign w25282 = w25095 & w25281;
assign v7998 = ~(w25095 | w25281);
assign w25283 = v7998;
assign v7999 = ~(w25282 | w25283);
assign w25284 = v7999;
assign v8000 = ~(w25189 | w25192);
assign w25285 = v8000;
assign w25286 = w5114 & ~w21866;
assign w25287 = w5531 & w19952;
assign w25288 = w5610 & w19954;
assign v8001 = ~(w25287 | w25288);
assign w25289 = v8001;
assign w25290 = w5113 & w19958;
assign w25291 = w25289 & ~w25290;
assign w25292 = ~w25286 & w25291;
assign w25293 = pi20 & w25292;
assign v8002 = ~(pi20 | w25292);
assign w25294 = v8002;
assign v8003 = ~(w25293 | w25294);
assign w25295 = v8003;
assign v8004 = ~(w25285 | w25295);
assign w25296 = v8004;
assign w25297 = w25285 & w25295;
assign v8005 = ~(w25296 | w25297);
assign w25298 = v8005;
assign v8006 = ~(w25146 | w25149);
assign w25299 = v8006;
assign w25300 = ~w454 & w2078;
assign w25301 = w5427 & w25300;
assign w25302 = w290 & ~w414;
assign w25303 = w6657 & w25302;
assign w25304 = w25301 & w25303;
assign w25305 = w1853 & w4989;
assign w25306 = w3786 & w25305;
assign w25307 = w3061 & w25306;
assign w25308 = w25304 & w25307;
assign w25309 = w1751 & w25308;
assign w25310 = w1511 & w5314;
assign w25311 = w2834 & w13961;
assign w25312 = w25310 & w25311;
assign w25313 = w25309 & w25312;
assign w25314 = ~pi02 & w25313;
assign w25315 = pi02 & ~w25313;
assign v8007 = ~(w25314 | w25315);
assign w25316 = v8007;
assign v8008 = ~(w25114 | w25136);
assign w25317 = v8008;
assign w25318 = w25316 & w25317;
assign v8009 = ~(w25316 | w25317);
assign w25319 = v8009;
assign v8010 = ~(w25318 | w25319);
assign w25320 = v8010;
assign w25321 = w928 & w20668;
assign w25322 = w3406 & ~w19997;
assign w25323 = w3399 & w20005;
assign w25324 = w3402 & w20000;
assign v8011 = ~(w25323 | w25324);
assign w25325 = v8011;
assign w25326 = ~w25322 & w25325;
assign w25327 = ~w25321 & w25326;
assign w25328 = ~w25320 & w25327;
assign w25329 = w25320 & ~w25327;
assign v8012 = ~(w25328 | w25329);
assign w25330 = v8012;
assign w25331 = w25299 & w25330;
assign v8013 = ~(w25299 | w25330);
assign w25332 = v8013;
assign v8014 = ~(w25331 | w25332);
assign w25333 = v8014;
assign w25334 = w3529 & w21012;
assign w25335 = w3760 & w19986;
assign w25336 = w3767 & ~w19992;
assign w25337 = w3763 & w19989;
assign v8015 = ~(w25336 | w25337);
assign w25338 = v8015;
assign w25339 = ~w25335 & w25338;
assign w25340 = ~w25334 & w25339;
assign w25341 = ~pi29 & w25340;
assign w25342 = pi29 & ~w25340;
assign v8016 = ~(w25341 | w25342);
assign w25343 = v8016;
assign w25344 = ~w25333 & w25343;
assign w25345 = w25333 & ~w25343;
assign v8017 = ~(w25344 | w25345);
assign w25346 = v8017;
assign w25347 = w4153 & w21362;
assign w25348 = w4155 & w19974;
assign w25349 = ~w2873 & w19983;
assign w25350 = w4158 & w19980;
assign v8018 = ~(w25349 | w25350);
assign w25351 = v8018;
assign w25352 = ~w25348 & w25351;
assign w25353 = ~w25347 & w25352;
assign w25354 = ~pi26 & w25353;
assign w25355 = pi26 & ~w25353;
assign v8019 = ~(w25354 | w25355);
assign w25356 = v8019;
assign w25357 = w25346 & w25356;
assign v8020 = ~(w25346 | w25356);
assign w25358 = v8020;
assign v8021 = ~(w25357 | w25358);
assign w25359 = v8021;
assign v8022 = ~(w25172 | w25176);
assign w25360 = v8022;
assign w25361 = w4764 & w20234;
assign w25362 = w4836 & w19966;
assign w25363 = w4913 & w19961;
assign v8023 = ~(w25362 | w25363);
assign w25364 = v8023;
assign w25365 = w4763 & ~w19971;
assign w25366 = w25364 & ~w25365;
assign w25367 = ~w25361 & w25366;
assign w25368 = pi23 & w25367;
assign v8024 = ~(pi23 | w25367);
assign w25369 = v8024;
assign v8025 = ~(w25368 | w25369);
assign w25370 = v8025;
assign w25371 = w25360 & ~w25370;
assign w25372 = ~w25360 & w25370;
assign v8026 = ~(w25371 | w25372);
assign w25373 = v8026;
assign w25374 = w25359 & w25373;
assign v8027 = ~(w25359 | w25373);
assign w25375 = v8027;
assign v8028 = ~(w25374 | w25375);
assign w25376 = v8028;
assign w25377 = w25298 & ~w25376;
assign w25378 = ~w25298 & w25376;
assign v8029 = ~(w25377 | w25378);
assign w25379 = v8029;
assign v8030 = ~(w25206 | w25209);
assign w25380 = v8030;
assign w25381 = ~w25379 & w25380;
assign w25382 = w25379 & ~w25380;
assign v8031 = ~(w25381 | w25382);
assign w25383 = v8031;
assign w25384 = w5765 & ~w22285;
assign w25385 = w6236 & ~w19929;
assign w25386 = w5764 & ~w19939;
assign w25387 = w5983 & w19933;
assign v8032 = ~(w25386 | w25387);
assign w25388 = v8032;
assign w25389 = ~w25385 & w25388;
assign w25390 = ~w25384 & w25389;
assign w25391 = ~pi17 & w25390;
assign w25392 = pi17 & ~w25390;
assign v8033 = ~(w25391 | w25392);
assign w25393 = v8033;
assign w25394 = ~w25383 & w25393;
assign w25395 = w25383 & ~w25393;
assign v8034 = ~(w25394 | w25395);
assign w25396 = v8034;
assign v8035 = ~(w25223 | w25226);
assign w25397 = v8035;
assign w25398 = w7004 & w19853;
assign w25399 = w6871 & w19917;
assign w25400 = w6388 & ~w19923;
assign v8036 = ~(w25399 | w25400);
assign w25401 = v8036;
assign w25402 = ~w25398 & w25401;
assign w25403 = (~w22936 & w28437) | (~w22936 & w28438) | (w28437 & w28438);
assign w25404 = (w22936 & w28439) | (w22936 & w28440) | (w28439 & w28440);
assign v8037 = ~(w25403 | w25404);
assign w25405 = v8037;
assign w25406 = w25397 & w25405;
assign v8038 = ~(w25397 | w25405);
assign w25407 = v8038;
assign v8039 = ~(w25406 | w25407);
assign w25408 = v8039;
assign w25409 = w25396 & ~w25408;
assign w25410 = ~w25396 & w25408;
assign v8040 = ~(w25409 | w25410);
assign w25411 = v8040;
assign w25412 = ~w25231 & w25242;
assign v8041 = ~(w25230 | w25412);
assign w25413 = v8041;
assign w25414 = w25411 & ~w25413;
assign w25415 = ~w25411 & w25413;
assign v8042 = ~(w25414 | w25415);
assign w25416 = v8042;
assign w25417 = w7765 & w23607;
assign w25418 = w7177 & ~w19912;
assign w25419 = w7466 & w20197;
assign v8043 = ~(w25418 | w25419);
assign w25420 = v8043;
assign w25421 = ~w25417 & w25420;
assign w25422 = (w25421 & ~w23614) | (w25421 & w29124) | (~w23614 & w29124);
assign w25423 = pi11 & w25422;
assign v8044 = ~(pi11 | w25422);
assign w25424 = v8044;
assign v8045 = ~(w25423 | w25424);
assign w25425 = v8045;
assign w25426 = w25416 & ~w25425;
assign w25427 = ~w25416 & w25425;
assign v8046 = ~(w25426 | w25427);
assign w25428 = v8046;
assign w25429 = (~w25246 & ~w25248) | (~w25246 & w28848) | (~w25248 & w28848);
assign w25430 = ~w24281 & w28598;
assign w25431 = w8140 & w23670;
assign w25432 = w8926 & w24284;
assign v8047 = ~(w25431 | w25432);
assign w25433 = v8047;
assign w25434 = w8526 & ~w24077;
assign w25435 = ~w25430 & w28849;
assign w25436 = (~pi08 & w25430) | (~pi08 & w28850) | (w25430 & w28850);
assign v8048 = ~(w25435 | w25436);
assign w25437 = v8048;
assign w25438 = w25429 & ~w25437;
assign w25439 = ~w25429 & w25437;
assign v8049 = ~(w25438 | w25439);
assign w25440 = v8049;
assign w25441 = w25428 & w25440;
assign v8050 = ~(w25428 | w25440);
assign w25442 = v8050;
assign v8051 = ~(w25441 | w25442);
assign w25443 = v8051;
assign w25444 = (~w25253 & ~w25254) | (~w25253 & w28851) | (~w25254 & w28851);
assign v8052 = ~(pi05 | w25444);
assign w25445 = v8052;
assign w25446 = pi05 & w25444;
assign v8053 = ~(w25445 | w25446);
assign w25447 = v8053;
assign v8054 = ~(w25443 | w25447);
assign w25448 = v8054;
assign w25449 = w25443 & w25447;
assign v8055 = ~(w25448 | w25449);
assign w25450 = v8055;
assign w25451 = (~w25268 & ~w25270) | (~w25268 & w28852) | (~w25270 & w28852);
assign w25452 = w25450 & ~w25451;
assign w25453 = ~w25450 & w25451;
assign v8056 = ~(w25452 | w25453);
assign w25454 = v8056;
assign w25455 = (~w25276 & w25278) | (~w25276 & w28097) | (w25278 & w28097);
assign w25456 = (~w25278 & w28599) | (~w25278 & w28600) | (w28599 & w28600);
assign w25457 = (w25278 & w28601) | (w25278 & w28602) | (w28601 & w28602);
assign v8057 = ~(w25456 | w25457);
assign w25458 = v8057;
assign w25459 = w25282 & ~w25458;
assign w25460 = ~w25282 & w25458;
assign v8058 = ~(w25459 | w25460);
assign w25461 = v8058;
assign w25462 = (~w25446 & ~w25447) | (~w25446 & w29125) | (~w25447 & w29125);
assign v8059 = ~(w25414 | w25426);
assign w25463 = v8059;
assign v8060 = ~(w25382 | w25395);
assign w25464 = v8060;
assign v8061 = ~(w25297 | w25377);
assign w25465 = v8061;
assign v8062 = ~(w25371 | w25374);
assign w25466 = v8062;
assign v8063 = ~(w25344 | w25357);
assign w25467 = v8063;
assign w25468 = w1541 & w4485;
assign w25469 = ~w564 & w2465;
assign w25470 = w25468 & w25469;
assign w25471 = w1263 & w2296;
assign w25472 = w25470 & w25471;
assign w25473 = w2636 & w5185;
assign w25474 = ~w108 & w25473;
assign w25475 = w12666 & w25474;
assign w25476 = w25472 & w25475;
assign w25477 = w20890 & w25476;
assign w25478 = w4596 & w25477;
assign w25479 = w1038 & w25478;
assign w25480 = w2522 & w25479;
assign w25481 = pi02 & w25480;
assign v8064 = ~(pi02 | w25480);
assign w25482 = v8064;
assign v8065 = ~(w25481 | w25482);
assign w25483 = v8065;
assign w25484 = pi05 & w25483;
assign v8066 = ~(pi05 | w25483);
assign w25485 = v8066;
assign v8067 = ~(w25484 | w25485);
assign w25486 = v8067;
assign v8068 = ~(w25315 | w25318);
assign w25487 = v8068;
assign v8069 = ~(w25486 | w25487);
assign w25488 = v8069;
assign w25489 = w25486 & w25487;
assign v8070 = ~(w25488 | w25489);
assign w25490 = v8070;
assign w25491 = w928 & w20655;
assign w25492 = w3406 & ~w19992;
assign w25493 = w3402 & ~w19997;
assign w25494 = w3399 & w20000;
assign v8071 = ~(w25493 | w25494);
assign w25495 = v8071;
assign w25496 = ~w25492 & w25495;
assign w25497 = ~w25491 & w25496;
assign w25498 = w25490 & ~w25497;
assign w25499 = ~w25490 & w25497;
assign v8072 = ~(w25498 | w25499);
assign w25500 = v8072;
assign v8073 = ~(w25328 | w25331);
assign w25501 = v8073;
assign v8074 = ~(w25500 | w25501);
assign w25502 = v8074;
assign w25503 = w25500 & w25501;
assign v8075 = ~(w25502 | w25503);
assign w25504 = v8075;
assign w25505 = w3529 & w20997;
assign w25506 = w3760 & w19983;
assign w25507 = w3767 & w19989;
assign w25508 = w3763 & w19986;
assign v8076 = ~(w25507 | w25508);
assign w25509 = v8076;
assign w25510 = ~w25506 & w25509;
assign w25511 = ~w25505 & w25510;
assign w25512 = ~pi29 & w25511;
assign w25513 = pi29 & ~w25511;
assign v8077 = ~(w25512 | w25513);
assign w25514 = v8077;
assign w25515 = w25504 & ~w25514;
assign w25516 = ~w25504 & w25514;
assign v8078 = ~(w25515 | w25516);
assign w25517 = v8078;
assign w25518 = w4153 & w21401;
assign w25519 = w4155 & ~w19971;
assign w25520 = ~w2873 & w19980;
assign w25521 = w4158 & w19974;
assign v8079 = ~(w25520 | w25521);
assign w25522 = v8079;
assign w25523 = ~w25519 & w25522;
assign w25524 = ~w25518 & w25523;
assign w25525 = ~pi26 & w25524;
assign w25526 = pi26 & ~w25524;
assign v8080 = ~(w25525 | w25526);
assign w25527 = v8080;
assign w25528 = ~w25517 & w25527;
assign w25529 = w25517 & ~w25527;
assign v8081 = ~(w25528 | w25529);
assign w25530 = v8081;
assign w25531 = w25467 & w25530;
assign v8082 = ~(w25467 | w25530);
assign w25532 = v8082;
assign v8083 = ~(w25531 | w25532);
assign w25533 = v8083;
assign w25534 = w4764 & w21716;
assign w25535 = w4913 & w19958;
assign w25536 = w4836 & w19961;
assign w25537 = w4763 & w19966;
assign v8084 = ~(w25536 | w25537);
assign w25538 = v8084;
assign w25539 = ~w25535 & w25538;
assign w25540 = ~w25534 & w25539;
assign w25541 = pi23 & ~w25540;
assign w25542 = ~pi23 & w25540;
assign v8085 = ~(w25541 | w25542);
assign w25543 = v8085;
assign w25544 = ~w25533 & w25543;
assign w25545 = w25533 & ~w25543;
assign v8086 = ~(w25544 | w25545);
assign w25546 = v8086;
assign w25547 = ~w25466 & w25546;
assign w25548 = w25466 & ~w25546;
assign v8087 = ~(w25547 | w25548);
assign w25549 = v8087;
assign w25550 = w5114 & w20214;
assign w25551 = w5610 & ~w19939;
assign w25552 = w5113 & w19952;
assign w25553 = w5531 & w19954;
assign v8088 = ~(w25552 | w25553);
assign w25554 = v8088;
assign w25555 = ~w25551 & w25554;
assign w25556 = ~w25550 & w25555;
assign w25557 = ~pi20 & w25556;
assign w25558 = pi20 & ~w25556;
assign v8089 = ~(w25557 | w25558);
assign w25559 = v8089;
assign v8090 = ~(w25549 | w25559);
assign w25560 = v8090;
assign w25561 = w25549 & w25559;
assign v8091 = ~(w25560 | w25561);
assign w25562 = v8091;
assign w25563 = ~w25465 & w25562;
assign w25564 = w25465 & ~w25562;
assign v8092 = ~(w25563 | w25564);
assign w25565 = v8092;
assign w25566 = w5765 & w22262;
assign w25567 = w6236 & ~w19923;
assign w25568 = w5764 & w19933;
assign w25569 = w5983 & ~w19929;
assign v8093 = ~(w25568 | w25569);
assign w25570 = v8093;
assign w25571 = ~w25567 & w25570;
assign w25572 = ~w25566 & w25571;
assign w25573 = ~pi17 & w25572;
assign w25574 = pi17 & ~w25572;
assign v8094 = ~(w25573 | w25574);
assign w25575 = v8094;
assign w25576 = w25565 & ~w25575;
assign w25577 = ~w25565 & w25575;
assign v8095 = ~(w25576 | w25577);
assign w25578 = v8095;
assign v8096 = ~(w25464 | w25578);
assign w25579 = v8096;
assign w25580 = w25464 & w25578;
assign v8097 = ~(w25579 | w25580);
assign w25581 = v8097;
assign w25582 = (~w25406 & ~w25408) | (~w25406 & w28853) | (~w25408 & w28853);
assign w25583 = w6871 & w19853;
assign w25584 = w7004 & ~w19912;
assign v8098 = ~(w25583 | w25584);
assign w25585 = v8098;
assign w25586 = w6388 & w19917;
assign w25587 = w25585 & ~w25586;
assign w25588 = (~w22917 & w29126) | (~w22917 & w29127) | (w29126 & w29127);
assign w25589 = (w22917 & w29128) | (w22917 & w29129) | (w29128 & w29129);
assign v8099 = ~(w25588 | w25589);
assign w25590 = v8099;
assign v8100 = ~(w25582 | w25590);
assign w25591 = v8100;
assign w25592 = w25582 & w25590;
assign v8101 = ~(w25591 | w25592);
assign w25593 = v8101;
assign w25594 = ~w25581 & w25593;
assign w25595 = w25581 & ~w25593;
assign v8102 = ~(w25594 | w25595);
assign w25596 = v8102;
assign w25597 = w7178 & w23666;
assign w25598 = w7765 & w23670;
assign w25599 = w7177 & w20197;
assign w25600 = w7466 & w23607;
assign v8103 = ~(w25599 | w25600);
assign w25601 = v8103;
assign w25602 = ~w25598 & w25601;
assign w25603 = ~w25597 & w25602;
assign w25604 = pi11 & ~w25603;
assign w25605 = ~pi11 & w25603;
assign v8104 = ~(w25604 | w25605);
assign w25606 = v8104;
assign w25607 = ~w25596 & w25606;
assign w25608 = w25596 & ~w25606;
assign v8105 = ~(w25607 | w25608);
assign w25609 = v8105;
assign w25610 = w25463 & ~w25609;
assign w25611 = ~w25463 & w25609;
assign v8106 = ~(w25610 | w25611);
assign w25612 = v8106;
assign w25613 = w8141 & ~w24304;
assign w25614 = w8526 & w24284;
assign w25615 = w8140 & ~w24077;
assign v8107 = ~(w25614 | w25615);
assign w25616 = v8107;
assign w25617 = ~w25613 & w25616;
assign w25618 = ~pi08 & w25617;
assign w25619 = pi08 & ~w25617;
assign v8108 = ~(w25618 | w25619);
assign w25620 = v8108;
assign w25621 = (w25620 & w25441) | (w25620 & w29130) | (w25441 & w29130);
assign w25622 = ~w25441 & w29131;
assign v8109 = ~(w25621 | w25622);
assign w25623 = v8109;
assign v8110 = ~(w25612 | w25623);
assign w25624 = v8110;
assign w25625 = w25612 & w25623;
assign v8111 = ~(w25624 | w25625);
assign w25626 = v8111;
assign w25627 = ~w25462 & w25626;
assign w25628 = w25462 & ~w25626;
assign v8112 = ~(w25627 | w25628);
assign w25629 = v8112;
assign w25630 = (~w25278 & w28855) | (~w25278 & w28856) | (w28855 & w28856);
assign w25631 = (~w25455 & w28603) | (~w25455 & w28604) | (w28603 & w28604);
assign w25632 = (w25455 & w28605) | (w25455 & w28606) | (w28605 & w28606);
assign v8113 = ~(w25631 | w25632);
assign w25633 = v8113;
assign v8114 = ~(w25459 | w25633);
assign w25634 = v8114;
assign w25635 = w25459 & w25633;
assign v8115 = ~(w25634 | w25635);
assign w25636 = v8115;
assign w25637 = (w25455 & w28607) | (w25455 & w28608) | (w28607 & w28608);
assign v8116 = ~(w25621 | w25625);
assign w25638 = v8116;
assign v8117 = ~(w25577 | w25580);
assign w25639 = v8117;
assign w25640 = w7004 & w20197;
assign w25641 = w6388 & w19853;
assign w25642 = w6871 & ~w19912;
assign v8118 = ~(w25641 | w25642);
assign w25643 = v8118;
assign w25644 = ~w25640 & w25643;
assign w25645 = (w25644 & ~w20203) | (w25644 & w29132) | (~w20203 & w29132);
assign w25646 = pi14 & w25645;
assign v8119 = ~(pi14 | w25645);
assign w25647 = v8119;
assign v8120 = ~(w25646 | w25647);
assign w25648 = v8120;
assign v8121 = ~(w25639 | w25648);
assign w25649 = v8121;
assign w25650 = w25639 & w25648;
assign v8122 = ~(w25649 | w25650);
assign w25651 = v8122;
assign v8123 = ~(w25488 | w25498);
assign w25652 = v8123;
assign w25653 = w476 & w14483;
assign w25654 = w1012 & w25653;
assign w25655 = w1635 & w25654;
assign w25656 = w6651 & w25655;
assign w25657 = w1372 & w25656;
assign w25658 = w283 & w2286;
assign w25659 = ~w420 & w1337;
assign w25660 = w3091 & w25659;
assign w25661 = w977 & w1065;
assign w25662 = w25660 & w25661;
assign w25663 = w2325 & w25662;
assign w25664 = w25658 & w25663;
assign w25665 = w25657 & w25664;
assign w25666 = w2051 & w3715;
assign w25667 = w893 & w25666;
assign w25668 = w783 & w1666;
assign w25669 = w2193 & w25668;
assign w25670 = w2182 & w25669;
assign w25671 = w3593 & w25670;
assign w25672 = w6717 & w13223;
assign w25673 = w6069 & w25672;
assign w25674 = w25671 & w25673;
assign w25675 = w25667 & w25674;
assign w25676 = w1607 & w25675;
assign w25677 = w25665 & w25676;
assign w25678 = w928 & w20965;
assign w25679 = w3406 & w19989;
assign w25680 = w3399 & ~w19997;
assign w25681 = w3402 & ~w19992;
assign v8124 = ~(w25680 | w25681);
assign w25682 = v8124;
assign w25683 = ~w25679 & w25682;
assign w25684 = ~w25678 & w25683;
assign w25685 = ~w25677 & w25684;
assign w25686 = w25677 & ~w25684;
assign v8125 = ~(w25685 | w25686);
assign w25687 = v8125;
assign v8126 = ~(w25481 | w25484);
assign w25688 = v8126;
assign w25689 = w25687 & w25688;
assign v8127 = ~(w25687 | w25688);
assign w25690 = v8127;
assign v8128 = ~(w25689 | w25690);
assign w25691 = v8128;
assign w25692 = w3529 & w20982;
assign w25693 = w3760 & w19980;
assign w25694 = w3763 & w19983;
assign w25695 = w3767 & w19986;
assign v8129 = ~(w25694 | w25695);
assign w25696 = v8129;
assign w25697 = ~w25693 & w25696;
assign w25698 = ~w25692 & w25697;
assign w25699 = ~pi29 & w25698;
assign w25700 = pi29 & ~w25698;
assign v8130 = ~(w25699 | w25700);
assign w25701 = v8130;
assign v8131 = ~(w25691 | w25701);
assign w25702 = v8131;
assign w25703 = w25691 & w25701;
assign v8132 = ~(w25702 | w25703);
assign w25704 = v8132;
assign w25705 = w25652 & w25704;
assign v8133 = ~(w25652 | w25704);
assign w25706 = v8133;
assign v8134 = ~(w25705 | w25706);
assign w25707 = v8134;
assign v8135 = ~(w25502 | w25515);
assign w25708 = v8135;
assign w25709 = ~w25707 & w25708;
assign w25710 = w25707 & ~w25708;
assign v8136 = ~(w25709 | w25710);
assign w25711 = v8136;
assign w25712 = w4153 & w21385;
assign w25713 = w4155 & w19966;
assign w25714 = ~w2873 & w19974;
assign w25715 = w4158 & ~w19971;
assign v8137 = ~(w25714 | w25715);
assign w25716 = v8137;
assign w25717 = ~w25713 & w25716;
assign w25718 = ~w25712 & w25717;
assign w25719 = ~pi26 & w25718;
assign w25720 = pi26 & ~w25718;
assign v8138 = ~(w25719 | w25720);
assign w25721 = v8138;
assign w25722 = w25711 & w25721;
assign v8139 = ~(w25711 | w25721);
assign w25723 = v8139;
assign v8140 = ~(w25722 | w25723);
assign w25724 = v8140;
assign v8141 = ~(w25529 | w25531);
assign w25725 = v8141;
assign w25726 = w25724 & w25725;
assign v8142 = ~(w25724 | w25725);
assign w25727 = v8142;
assign v8143 = ~(w25726 | w25727);
assign w25728 = v8143;
assign w25729 = w4764 & ~w21882;
assign w25730 = w4836 & w19958;
assign w25731 = w4913 & w19952;
assign v8144 = ~(w25730 | w25731);
assign w25732 = v8144;
assign w25733 = w4763 & w19961;
assign w25734 = w25732 & ~w25733;
assign w25735 = ~w25729 & w25734;
assign w25736 = pi23 & w25735;
assign v8145 = ~(pi23 | w25735);
assign w25737 = v8145;
assign v8146 = ~(w25736 | w25737);
assign w25738 = v8146;
assign w25739 = w25728 & ~w25738;
assign w25740 = ~w25728 & w25738;
assign v8147 = ~(w25739 | w25740);
assign w25741 = v8147;
assign v8148 = ~(w25544 | w25547);
assign w25742 = v8148;
assign w25743 = w5114 & ~w22304;
assign w25744 = w5610 & w19933;
assign w25745 = w5113 & w19954;
assign w25746 = w5531 & ~w19939;
assign v8149 = ~(w25745 | w25746);
assign w25747 = v8149;
assign w25748 = ~w25744 & w25747;
assign w25749 = ~w25743 & w25748;
assign w25750 = ~pi20 & w25749;
assign w25751 = pi20 & ~w25749;
assign v8150 = ~(w25750 | w25751);
assign w25752 = v8150;
assign w25753 = ~w25742 & w25752;
assign w25754 = w25742 & ~w25752;
assign v8151 = ~(w25753 | w25754);
assign w25755 = v8151;
assign w25756 = w25741 & w25755;
assign v8152 = ~(w25741 | w25755);
assign w25757 = v8152;
assign v8153 = ~(w25756 | w25757);
assign w25758 = v8153;
assign v8154 = ~(w25560 | w25563);
assign w25759 = v8154;
assign w25760 = w5765 & ~w22895;
assign w25761 = w6236 & w19917;
assign w25762 = w5764 & ~w19929;
assign w25763 = w5983 & ~w19923;
assign v8155 = ~(w25762 | w25763);
assign w25764 = v8155;
assign w25765 = ~w25761 & w25764;
assign w25766 = ~w25760 & w25765;
assign w25767 = ~pi17 & w25766;
assign w25768 = pi17 & ~w25766;
assign v8156 = ~(w25767 | w25768);
assign w25769 = v8156;
assign v8157 = ~(w25759 | w25769);
assign w25770 = v8157;
assign w25771 = w25759 & w25769;
assign v8158 = ~(w25770 | w25771);
assign w25772 = v8158;
assign w25773 = w25758 & w25772;
assign v8159 = ~(w25758 | w25772);
assign w25774 = v8159;
assign v8160 = ~(w25773 | w25774);
assign w25775 = v8160;
assign w25776 = w25651 & w25775;
assign v8161 = ~(w25651 | w25775);
assign w25777 = v8161;
assign v8162 = ~(w25776 | w25777);
assign w25778 = v8162;
assign v8163 = ~(w25592 | w25594);
assign w25779 = v8163;
assign w25780 = w7178 & w24073;
assign w25781 = w7765 & ~w24077;
assign w25782 = w7177 & w23607;
assign v8164 = ~(w25781 | w25782);
assign w25783 = v8164;
assign w25784 = w7466 & w23670;
assign w25785 = w25783 & ~w25784;
assign w25786 = ~w25780 & w25785;
assign w25787 = ~pi11 & w25786;
assign w25788 = pi11 & ~w25786;
assign v8165 = ~(w25787 | w25788);
assign w25789 = v8165;
assign w25790 = w25779 & w25789;
assign v8166 = ~(w25779 | w25789);
assign w25791 = v8166;
assign v8167 = ~(w25790 | w25791);
assign w25792 = v8167;
assign w25793 = w25778 & w25792;
assign v8168 = ~(w25778 | w25792);
assign w25794 = v8168;
assign v8169 = ~(w25793 | w25794);
assign w25795 = v8169;
assign w25796 = (~w25607 & ~w25609) | (~w25607 & w29133) | (~w25609 & w29133);
assign w25797 = w8139 & w24284;
assign v8170 = ~(pi08 | w25797);
assign w25798 = v8170;
assign w25799 = w13300 & w24284;
assign v8171 = ~(w25798 | w25799);
assign w25800 = v8171;
assign w25801 = ~w25796 & w25800;
assign w25802 = w25796 & ~w25800;
assign v8172 = ~(w25801 | w25802);
assign w25803 = v8172;
assign w25804 = w25795 & w25803;
assign v8173 = ~(w25795 | w25803);
assign w25805 = v8173;
assign v8174 = ~(w25804 | w25805);
assign w25806 = v8174;
assign w25807 = ~w25638 & w25806;
assign w25808 = w25638 & ~w25806;
assign v8175 = ~(w25807 | w25808);
assign w25809 = v8175;
assign w25810 = (w25455 & w29134) | (w25455 & w29135) | (w29134 & w29135);
assign w25811 = (~w25455 & w29136) | (~w25455 & w29137) | (w29136 & w29137);
assign v8176 = ~(w25810 | w25811);
assign w25812 = v8176;
assign w25813 = w25635 & w25812;
assign v8177 = ~(w25635 | w25812);
assign w25814 = v8177;
assign v8178 = ~(w25813 | w25814);
assign w25815 = v8178;
assign v8179 = ~(w25790 | w25793);
assign w25816 = v8179;
assign w25817 = ~pi08 & w25816;
assign w25818 = pi08 & ~w25816;
assign v8180 = ~(w25817 | w25818);
assign w25819 = v8180;
assign v8181 = ~(w25649 | w25776);
assign w25820 = v8181;
assign v8182 = ~(w25726 | w25739);
assign w25821 = v8182;
assign v8183 = ~(w25709 | w25722);
assign w25822 = v8183;
assign v8184 = ~(w25702 | w25705);
assign w25823 = v8184;
assign w25824 = w928 & w21012;
assign w25825 = w3406 & w19986;
assign w25826 = w3402 & w19989;
assign w25827 = w3399 & ~w19992;
assign v8185 = ~(w25826 | w25827);
assign w25828 = v8185;
assign w25829 = ~w25825 & w25828;
assign w25830 = ~w25824 & w25829;
assign v8186 = ~(w25685 | w25689);
assign w25831 = v8186;
assign w25832 = ~w479 & w936;
assign w25833 = ~w373 & w25832;
assign w25834 = ~w427 & w6542;
assign w25835 = ~w245 & w3317;
assign w25836 = w1928 & w25835;
assign v8187 = ~(w160 | w232);
assign w25837 = v8187;
assign w25838 = ~w414 & w25837;
assign w25839 = ~w326 & w25838;
assign w25840 = w25836 & w25839;
assign w25841 = ~w997 & w3886;
assign w25842 = w769 & w25841;
assign v8188 = ~(w199 | w216);
assign w25843 = v8188;
assign w25844 = w25842 & w25843;
assign w25845 = w25840 & w25844;
assign w25846 = w4273 & w25845;
assign w25847 = w25834 & w25846;
assign w25848 = w25833 & w25847;
assign w25849 = w1840 & w3057;
assign w25850 = w289 & w4367;
assign v8189 = ~(w132 | w202);
assign w25851 = v8189;
assign w25852 = w279 & w25851;
assign w25853 = ~w430 & w25852;
assign w25854 = w25850 & w25853;
assign w25855 = w6561 & w14317;
assign w25856 = w1856 & w25855;
assign w25857 = w665 & w25856;
assign w25858 = w25854 & w25857;
assign w25859 = w25849 & w25858;
assign w25860 = w12646 & w25859;
assign w25861 = w25848 & w25860;
assign w25862 = w25684 & w25861;
assign v8190 = ~(w25684 | w25861);
assign w25863 = v8190;
assign v8191 = ~(w25862 | w25863);
assign w25864 = v8191;
assign w25865 = w25831 & ~w25864;
assign w25866 = ~w25831 & w25864;
assign v8192 = ~(w25865 | w25866);
assign w25867 = v8192;
assign v8193 = ~(w25830 | w25867);
assign w25868 = v8193;
assign w25869 = w25830 & w25867;
assign v8194 = ~(w25868 | w25869);
assign w25870 = v8194;
assign w25871 = w25823 & w25870;
assign v8195 = ~(w25823 | w25870);
assign w25872 = v8195;
assign v8196 = ~(w25871 | w25872);
assign w25873 = v8196;
assign w25874 = w3529 & w21362;
assign w25875 = w3760 & w19974;
assign w25876 = w3763 & w19980;
assign w25877 = w3767 & w19983;
assign v8197 = ~(w25876 | w25877);
assign w25878 = v8197;
assign w25879 = ~w25875 & w25878;
assign w25880 = ~w25874 & w25879;
assign w25881 = pi29 & w25880;
assign v8198 = ~(pi29 | w25880);
assign w25882 = v8198;
assign v8199 = ~(w25881 | w25882);
assign w25883 = v8199;
assign w25884 = w25873 & ~w25883;
assign w25885 = ~w25873 & w25883;
assign v8200 = ~(w25884 | w25885);
assign w25886 = v8200;
assign w25887 = w4153 & w20234;
assign v8201 = ~(w2873 | w19971);
assign w25888 = v8201;
assign w25889 = w4155 & w19961;
assign v8202 = ~(w25888 | w25889);
assign w25890 = v8202;
assign w25891 = w4158 & w19966;
assign w25892 = w25890 & ~w25891;
assign w25893 = ~w25887 & w25892;
assign w25894 = pi26 & w25893;
assign v8203 = ~(pi26 | w25893);
assign w25895 = v8203;
assign v8204 = ~(w25894 | w25895);
assign w25896 = v8204;
assign w25897 = w25886 & ~w25896;
assign w25898 = ~w25886 & w25896;
assign v8205 = ~(w25897 | w25898);
assign w25899 = v8205;
assign w25900 = w4764 & ~w21866;
assign w25901 = w4836 & w19952;
assign w25902 = w4913 & w19954;
assign v8206 = ~(w25901 | w25902);
assign w25903 = v8206;
assign w25904 = w4763 & w19958;
assign w25905 = w25903 & ~w25904;
assign w25906 = ~w25900 & w25905;
assign w25907 = pi23 & w25906;
assign v8207 = ~(pi23 | w25906);
assign w25908 = v8207;
assign v8208 = ~(w25907 | w25908);
assign w25909 = v8208;
assign w25910 = ~w25899 & w25909;
assign w25911 = w25899 & ~w25909;
assign v8209 = ~(w25910 | w25911);
assign w25912 = v8209;
assign w25913 = w25822 & ~w25912;
assign w25914 = ~w25822 & w25912;
assign v8210 = ~(w25913 | w25914);
assign w25915 = v8210;
assign w25916 = ~w25821 & w25915;
assign w25917 = w25821 & ~w25915;
assign v8211 = ~(w25916 | w25917);
assign w25918 = v8211;
assign w25919 = w5114 & ~w22285;
assign w25920 = w5610 & ~w19929;
assign w25921 = w5113 & ~w19939;
assign w25922 = w5531 & w19933;
assign v8212 = ~(w25921 | w25922);
assign w25923 = v8212;
assign w25924 = ~w25920 & w25923;
assign w25925 = ~w25919 & w25924;
assign w25926 = pi20 & ~w25925;
assign w25927 = ~pi20 & w25925;
assign v8213 = ~(w25926 | w25927);
assign w25928 = v8213;
assign w25929 = w25918 & ~w25928;
assign w25930 = ~w25918 & w25928;
assign v8214 = ~(w25929 | w25930);
assign w25931 = v8214;
assign v8215 = ~(w25753 | w25756);
assign w25932 = v8215;
assign w25933 = w6236 & w19853;
assign w25934 = w5983 & w19917;
assign w25935 = w5764 & ~w19923;
assign v8216 = ~(w25934 | w25935);
assign w25936 = v8216;
assign w25937 = ~w25933 & w25936;
assign w25938 = (~w22936 & w28857) | (~w22936 & w28858) | (w28857 & w28858);
assign w25939 = (w22936 & w28240) | (w22936 & w28241) | (w28240 & w28241);
assign w25940 = ~w25938 & w28242;
assign w25941 = (~w25932 & w25938) | (~w25932 & w28243) | (w25938 & w28243);
assign v8217 = ~(w25940 | w25941);
assign w25942 = v8217;
assign w25943 = w25931 & w25942;
assign v8218 = ~(w25931 | w25942);
assign w25944 = v8218;
assign v8219 = ~(w25943 | w25944);
assign w25945 = v8219;
assign v8220 = ~(w25771 | w25773);
assign w25946 = v8220;
assign v8221 = ~(w25945 | w25946);
assign w25947 = v8221;
assign w25948 = w25945 & w25946;
assign v8222 = ~(w25947 | w25948);
assign w25949 = v8222;
assign w25950 = w6389 & w23614;
assign w25951 = w6871 & w20197;
assign w25952 = w7004 & w23607;
assign v8223 = ~(w25951 | w25952);
assign w25953 = v8223;
assign w25954 = w6388 & ~w19912;
assign w25955 = w25953 & ~w25954;
assign w25956 = ~w25950 & w25955;
assign w25957 = pi14 & w25956;
assign v8224 = ~(pi14 | w25956);
assign w25958 = v8224;
assign v8225 = ~(w25957 | w25958);
assign w25959 = v8225;
assign w25960 = w25949 & ~w25959;
assign w25961 = ~w25949 & w25959;
assign v8226 = ~(w25960 | w25961);
assign w25962 = v8226;
assign w25963 = ~w25820 & w25962;
assign w25964 = w25820 & ~w25962;
assign v8227 = ~(w25963 | w25964);
assign w25965 = v8227;
assign w25966 = w7178 & w24282;
assign w25967 = w7177 & w23670;
assign w25968 = w7765 & w24284;
assign w25969 = w7466 & ~w24077;
assign v8228 = ~(w25968 | w25969);
assign w25970 = v8228;
assign w25971 = ~w25967 & w25970;
assign w25972 = ~w25966 & w25971;
assign w25973 = pi11 & ~w25972;
assign w25974 = ~pi11 & w25972;
assign v8229 = ~(w25973 | w25974);
assign w25975 = v8229;
assign w25976 = w25965 & w25975;
assign v8230 = ~(w25965 | w25975);
assign w25977 = v8230;
assign v8231 = ~(w25976 | w25977);
assign w25978 = v8231;
assign v8232 = ~(w25819 | w25978);
assign w25979 = v8232;
assign w25980 = w25819 & w25978;
assign v8233 = ~(w25979 | w25980);
assign w25981 = v8233;
assign v8234 = ~(w25801 | w25804);
assign w25982 = v8234;
assign w25983 = ~w25981 & w25982;
assign w25984 = w25981 & ~w25982;
assign v8235 = ~(w25983 | w25984);
assign w25985 = v8235;
assign w25986 = (w25630 & w28609) | (w25630 & w28610) | (w28609 & w28610);
assign w25987 = (~w25630 & w29138) | (~w25630 & w29139) | (w29138 & w29139);
assign v8236 = ~(w25986 | w25987);
assign w25988 = v8236;
assign w25989 = w25635 & w28859;
assign v8237 = ~(w25813 | w25988);
assign w25990 = v8237;
assign v8238 = ~(w25989 | w25990);
assign w25991 = v8238;
assign w25992 = (~w25818 & ~w25819) | (~w25818 & w28244) | (~w25819 & w28244);
assign v8239 = ~(w25963 | w25976);
assign w25993 = v8239;
assign v8240 = ~(w25947 | w25960);
assign w25994 = v8240;
assign v8241 = ~(w25917 | w25929);
assign w25995 = v8241;
assign v8242 = ~(w25911 | w25914);
assign w25996 = v8242;
assign v8243 = ~(w25884 | w25897);
assign w25997 = v8243;
assign v8244 = ~(w25868 | w25871);
assign w25998 = v8244;
assign w25999 = ~w456 & w2263;
assign w26000 = w2835 & w25999;
assign w26001 = ~w183 & w2699;
assign w26002 = w844 & w2545;
assign w26003 = w114 & w2296;
assign w26004 = w509 & w26003;
assign w26005 = w26002 & w26004;
assign w26006 = w1602 & w12638;
assign w26007 = w26005 & w26006;
assign w26008 = w26001 & w26007;
assign w26009 = w26000 & w26008;
assign w26010 = w1314 & w3228;
assign w26011 = w26009 & w26010;
assign v8245 = ~(w25677 | w26011);
assign w26012 = v8245;
assign w26013 = w25677 & w26011;
assign v8246 = ~(w26012 | w26013);
assign w26014 = v8246;
assign w26015 = ~pi08 & w26014;
assign w26016 = pi08 & ~w26014;
assign v8247 = ~(w26015 | w26016);
assign w26017 = v8247;
assign v8248 = ~(w25677 | w25863);
assign w26018 = v8248;
assign w26019 = w25677 & ~w25862;
assign v8249 = ~(w25688 | w26019);
assign w26020 = v8249;
assign v8250 = ~(w26018 | w26020);
assign w26021 = v8250;
assign v8251 = ~(w26017 | w26021);
assign w26022 = v8251;
assign w26023 = w26017 & w26021;
assign v8252 = ~(w26022 | w26023);
assign w26024 = v8252;
assign w26025 = w928 & w20997;
assign w26026 = w3406 & w19983;
assign w26027 = w3399 & w19989;
assign w26028 = w3402 & w19986;
assign v8253 = ~(w26027 | w26028);
assign w26029 = v8253;
assign w26030 = ~w26026 & w26029;
assign w26031 = ~w26025 & w26030;
assign w26032 = w26024 & ~w26031;
assign w26033 = ~w26024 & w26031;
assign v8254 = ~(w26032 | w26033);
assign w26034 = v8254;
assign w26035 = w3529 & w21401;
assign w26036 = w3760 & ~w19971;
assign w26037 = w3763 & w19974;
assign w26038 = w3767 & w19980;
assign v8255 = ~(w26037 | w26038);
assign w26039 = v8255;
assign w26040 = ~w26036 & w26039;
assign w26041 = ~w26035 & w26040;
assign w26042 = ~pi29 & w26041;
assign w26043 = pi29 & ~w26041;
assign v8256 = ~(w26042 | w26043);
assign w26044 = v8256;
assign w26045 = w26034 & w26044;
assign v8257 = ~(w26034 | w26044);
assign w26046 = v8257;
assign v8258 = ~(w26045 | w26046);
assign w26047 = v8258;
assign w26048 = ~w25998 & w26047;
assign w26049 = w25998 & ~w26047;
assign v8259 = ~(w26048 | w26049);
assign w26050 = v8259;
assign w26051 = w4153 & w21716;
assign w26052 = ~w2873 & w19966;
assign w26053 = w4155 & w19958;
assign v8260 = ~(w26052 | w26053);
assign w26054 = v8260;
assign w26055 = w4158 & w19961;
assign w26056 = w26054 & ~w26055;
assign w26057 = ~w26051 & w26056;
assign w26058 = pi26 & w26057;
assign v8261 = ~(pi26 | w26057);
assign w26059 = v8261;
assign v8262 = ~(w26058 | w26059);
assign w26060 = v8262;
assign w26061 = w26050 & ~w26060;
assign w26062 = ~w26050 & w26060;
assign v8263 = ~(w26061 | w26062);
assign w26063 = v8263;
assign w26064 = ~w25997 & w26063;
assign w26065 = w25997 & ~w26063;
assign v8264 = ~(w26064 | w26065);
assign w26066 = v8264;
assign w26067 = w4764 & w20214;
assign w26068 = w4836 & w19954;
assign w26069 = w4913 & ~w19939;
assign v8265 = ~(w26068 | w26069);
assign w26070 = v8265;
assign w26071 = w4763 & w19952;
assign w26072 = w26070 & ~w26071;
assign w26073 = ~w26067 & w26072;
assign w26074 = pi23 & w26073;
assign v8266 = ~(pi23 | w26073);
assign w26075 = v8266;
assign v8267 = ~(w26074 | w26075);
assign w26076 = v8267;
assign w26077 = w26066 & ~w26076;
assign w26078 = ~w26066 & w26076;
assign v8268 = ~(w26077 | w26078);
assign w26079 = v8268;
assign w26080 = ~w25996 & w26079;
assign w26081 = w25996 & ~w26079;
assign v8269 = ~(w26080 | w26081);
assign w26082 = v8269;
assign w26083 = w5114 & w22262;
assign w26084 = w5610 & ~w19923;
assign w26085 = w5113 & w19933;
assign w26086 = w5531 & ~w19929;
assign v8270 = ~(w26085 | w26086);
assign w26087 = v8270;
assign w26088 = ~w26084 & w26087;
assign w26089 = ~w26083 & w26088;
assign w26090 = ~pi20 & w26089;
assign w26091 = pi20 & ~w26089;
assign v8271 = ~(w26090 | w26091);
assign w26092 = v8271;
assign w26093 = w26082 & w26092;
assign v8272 = ~(w26082 | w26092);
assign w26094 = v8272;
assign v8273 = ~(w26093 | w26094);
assign w26095 = v8273;
assign v8274 = ~(w25995 | w26095);
assign w26096 = v8274;
assign w26097 = w25995 & w26095;
assign v8275 = ~(w26096 | w26097);
assign w26098 = v8275;
assign w26099 = (~w25940 & ~w25942) | (~w25940 & w28860) | (~w25942 & w28860);
assign w26100 = w26098 & w26099;
assign v8276 = ~(w26098 | w26099);
assign w26101 = v8276;
assign v8277 = ~(w26100 | w26101);
assign w26102 = v8277;
assign w26103 = w5765 & w22917;
assign w26104 = w5983 & w19853;
assign w26105 = w6236 & ~w19912;
assign v8278 = ~(w26104 | w26105);
assign w26106 = v8278;
assign w26107 = w5764 & w19917;
assign w26108 = w26106 & ~w26107;
assign w26109 = ~w26103 & w26108;
assign v8279 = ~(pi17 | w26109);
assign w26110 = v8279;
assign w26111 = pi17 & w26109;
assign v8280 = ~(w26110 | w26111);
assign w26112 = v8280;
assign w26113 = ~w26102 & w26112;
assign w26114 = w26102 & ~w26112;
assign v8281 = ~(w26113 | w26114);
assign w26115 = v8281;
assign w26116 = w6389 & w23666;
assign w26117 = w6871 & w23607;
assign w26118 = w7004 & w23670;
assign v8282 = ~(w26117 | w26118);
assign w26119 = v8282;
assign w26120 = w6388 & w20197;
assign w26121 = w26119 & ~w26120;
assign w26122 = ~w26116 & w26121;
assign w26123 = pi14 & w26122;
assign v8283 = ~(pi14 | w26122);
assign w26124 = v8283;
assign v8284 = ~(w26123 | w26124);
assign w26125 = v8284;
assign w26126 = w26115 & ~w26125;
assign w26127 = ~w26115 & w26125;
assign v8285 = ~(w26126 | w26127);
assign w26128 = v8285;
assign w26129 = w25994 & ~w26128;
assign w26130 = ~w25994 & w26128;
assign v8286 = ~(w26129 | w26130);
assign w26131 = v8286;
assign w26132 = w7178 & ~w24304;
assign w26133 = w7466 & w24284;
assign w26134 = w7177 & ~w24077;
assign v8287 = ~(w26133 | w26134);
assign w26135 = v8287;
assign w26136 = ~w26132 & w26135;
assign w26137 = ~pi11 & w26136;
assign w26138 = pi11 & ~w26136;
assign v8288 = ~(w26137 | w26138);
assign w26139 = v8288;
assign w26140 = w26131 & w26139;
assign v8289 = ~(w26131 | w26139);
assign w26141 = v8289;
assign v8290 = ~(w26140 | w26141);
assign w26142 = v8290;
assign w26143 = ~w25993 & w26142;
assign w26144 = w25993 & ~w26142;
assign v8291 = ~(w26143 | w26144);
assign w26145 = v8291;
assign w26146 = ~w25992 & w26145;
assign w26147 = w25992 & ~w26145;
assign v8292 = ~(w26146 | w26147);
assign w26148 = v8292;
assign w26149 = ~w25983 & w26148;
assign w26150 = (~w25455 & w31305) | (~w25455 & w31306) | (w31305 & w31306);
assign v8293 = ~(w25984 | w26148);
assign w26151 = v8293;
assign w26152 = (~w25630 & w29140) | (~w25630 & w29141) | (w29140 & w29141);
assign v8294 = ~(w26150 | w26152);
assign w26153 = v8294;
assign v8295 = ~(w25989 | w26153);
assign w26154 = v8295;
assign w26155 = w25989 & w26153;
assign v8296 = ~(w26154 | w26155);
assign w26156 = v8296;
assign w26157 = (~w26126 & ~w26128) | (~w26126 & w29142) | (~w26128 & w29142);
assign v8297 = ~(w26045 | w26048);
assign w26158 = v8297;
assign v8298 = ~(w26012 | w26015);
assign w26159 = v8298;
assign w26160 = w542 & w1893;
assign w26161 = w14425 & w26160;
assign w26162 = w3235 & w4371;
assign w26163 = w3185 & w4121;
assign w26164 = w26162 & w26163;
assign w26165 = w26161 & w26164;
assign w26166 = w5022 & w26165;
assign w26167 = w3175 & w13147;
assign w26168 = w13935 & w26167;
assign w26169 = w3543 & w26168;
assign w26170 = w26166 & w26169;
assign w26171 = w2461 & w26170;
assign w26172 = ~w26159 & w26171;
assign w26173 = w26159 & ~w26171;
assign v8299 = ~(w26172 | w26173);
assign w26174 = v8299;
assign w26175 = w928 & w20982;
assign w26176 = w3406 & w19980;
assign w26177 = w3402 & w19983;
assign w26178 = w3399 & w19986;
assign v8300 = ~(w26177 | w26178);
assign w26179 = v8300;
assign w26180 = ~w26176 & w26179;
assign w26181 = ~w26175 & w26180;
assign w26182 = ~w26174 & w26181;
assign w26183 = w26174 & ~w26181;
assign v8301 = ~(w26182 | w26183);
assign w26184 = v8301;
assign v8302 = ~(w26023 | w26032);
assign w26185 = v8302;
assign w26186 = ~w26184 & w26185;
assign w26187 = w26184 & ~w26185;
assign v8303 = ~(w26186 | w26187);
assign w26188 = v8303;
assign w26189 = w3529 & w21385;
assign w26190 = w3760 & w19966;
assign w26191 = w3763 & ~w19971;
assign w26192 = w3767 & w19974;
assign v8304 = ~(w26191 | w26192);
assign w26193 = v8304;
assign w26194 = ~w26190 & w26193;
assign w26195 = ~w26189 & w26194;
assign w26196 = pi29 & w26195;
assign v8305 = ~(pi29 | w26195);
assign w26197 = v8305;
assign v8306 = ~(w26196 | w26197);
assign w26198 = v8306;
assign w26199 = w26188 & ~w26198;
assign w26200 = ~w26188 & w26198;
assign v8307 = ~(w26199 | w26200);
assign w26201 = v8307;
assign w26202 = ~w26158 & w26201;
assign w26203 = w26158 & ~w26201;
assign v8308 = ~(w26202 | w26203);
assign w26204 = v8308;
assign w26205 = w4153 & ~w21882;
assign w26206 = w4155 & w19952;
assign w26207 = ~w2873 & w19961;
assign w26208 = w4158 & w19958;
assign v8309 = ~(w26207 | w26208);
assign w26209 = v8309;
assign w26210 = ~w26206 & w26209;
assign w26211 = ~w26205 & w26210;
assign w26212 = ~pi26 & w26211;
assign w26213 = pi26 & ~w26211;
assign v8310 = ~(w26212 | w26213);
assign w26214 = v8310;
assign w26215 = w26204 & w26214;
assign v8311 = ~(w26204 | w26214);
assign w26216 = v8311;
assign v8312 = ~(w26215 | w26216);
assign w26217 = v8312;
assign v8313 = ~(w26061 | w26064);
assign w26218 = v8313;
assign w26219 = ~w26217 & w26218;
assign w26220 = w26217 & ~w26218;
assign v8314 = ~(w26219 | w26220);
assign w26221 = v8314;
assign w26222 = w4764 & ~w22304;
assign w26223 = w4763 & w19954;
assign w26224 = w4913 & w19933;
assign v8315 = ~(w26223 | w26224);
assign w26225 = v8315;
assign w26226 = w4836 & ~w19939;
assign w26227 = w26225 & ~w26226;
assign w26228 = ~w26222 & w26227;
assign w26229 = pi23 & w26228;
assign v8316 = ~(pi23 | w26228);
assign w26230 = v8316;
assign v8317 = ~(w26229 | w26230);
assign w26231 = v8317;
assign w26232 = w26221 & ~w26231;
assign w26233 = ~w26221 & w26231;
assign v8318 = ~(w26232 | w26233);
assign w26234 = v8318;
assign v8319 = ~(w26077 | w26080);
assign w26235 = v8319;
assign w26236 = ~w26234 & w26235;
assign w26237 = w26234 & ~w26235;
assign v8320 = ~(w26236 | w26237);
assign w26238 = v8320;
assign w26239 = w5114 & ~w22895;
assign w26240 = w5610 & w19917;
assign w26241 = w5113 & ~w19929;
assign w26242 = w5531 & ~w19923;
assign v8321 = ~(w26241 | w26242);
assign w26243 = v8321;
assign w26244 = ~w26240 & w26243;
assign w26245 = ~w26239 & w26244;
assign w26246 = ~pi20 & w26245;
assign w26247 = pi20 & ~w26245;
assign v8322 = ~(w26246 | w26247);
assign w26248 = v8322;
assign w26249 = w26238 & w26248;
assign v8323 = ~(w26238 | w26248);
assign w26250 = v8323;
assign v8324 = ~(w26249 | w26250);
assign w26251 = v8324;
assign v8325 = ~(w26093 | w26097);
assign w26252 = v8325;
assign w26253 = ~w26251 & w26252;
assign w26254 = w26251 & ~w26252;
assign v8326 = ~(w26253 | w26254);
assign w26255 = v8326;
assign w26256 = w6236 & w20197;
assign w26257 = w5983 & ~w19912;
assign w26258 = w5764 & w19853;
assign v8327 = ~(w26257 | w26258);
assign w26259 = v8327;
assign w26260 = ~w26256 & w26259;
assign w26261 = (w26260 & ~w20203) | (w26260 & w29143) | (~w20203 & w29143);
assign w26262 = pi17 & w26261;
assign v8328 = ~(pi17 | w26261);
assign w26263 = v8328;
assign v8329 = ~(w26262 | w26263);
assign w26264 = v8329;
assign w26265 = w26255 & ~w26264;
assign w26266 = ~w26255 & w26264;
assign v8330 = ~(w26265 | w26266);
assign w26267 = v8330;
assign w26268 = (~w26100 & ~w26102) | (~w26100 & w29144) | (~w26102 & w29144);
assign w26269 = ~w26267 & w26268;
assign w26270 = w26267 & ~w26268;
assign v8331 = ~(w26269 | w26270);
assign w26271 = v8331;
assign w26272 = w6389 & w24073;
assign w26273 = w6871 & w23670;
assign w26274 = w7004 & ~w24077;
assign v8332 = ~(w26273 | w26274);
assign w26275 = v8332;
assign w26276 = w6388 & w23607;
assign w26277 = w26275 & ~w26276;
assign w26278 = ~w26272 & w26277;
assign v8333 = ~(pi14 | w26278);
assign w26279 = v8333;
assign w26280 = pi14 & w26278;
assign v8334 = ~(w26279 | w26280);
assign w26281 = v8334;
assign w26282 = w26271 & ~w26281;
assign w26283 = ~w26271 & w26281;
assign v8335 = ~(w26282 | w26283);
assign w26284 = v8335;
assign w26285 = ~w26157 & w26284;
assign w26286 = w26157 & ~w26284;
assign v8336 = ~(w26285 | w26286);
assign w26287 = v8336;
assign w26288 = w7176 & w24284;
assign v8337 = ~(pi11 | w26288);
assign w26289 = v8337;
assign w26290 = w13166 & w24284;
assign v8338 = ~(w26289 | w26290);
assign w26291 = v8338;
assign w26292 = w26287 & w26291;
assign v8339 = ~(w26287 | w26291);
assign w26293 = v8339;
assign v8340 = ~(w26292 | w26293);
assign w26294 = v8340;
assign w26295 = (~w26140 & ~w26142) | (~w26140 & w29145) | (~w26142 & w29145);
assign w26296 = w26294 & ~w26295;
assign w26297 = ~w26294 & w26295;
assign v8341 = ~(w26296 | w26297);
assign w26298 = v8341;
assign w26299 = w26146 & ~w26298;
assign w26300 = (~w25637 & w29423) | (~w25637 & w29424) | (w29423 & w29424);
assign w26301 = w25989 & w28245;
assign w26302 = w26150 & ~w26298;
assign v8342 = ~(w26155 | w26302);
assign w26303 = v8342;
assign w26304 = w26300 & w26303;
assign v8343 = ~(w26301 | w26304);
assign w26305 = v8343;
assign v8344 = ~(w26187 | w26199);
assign w26306 = v8344;
assign v8345 = ~(w26172 | w26183);
assign w26307 = v8345;
assign w26308 = ~w21 & w14491;
assign w26309 = w3623 & w26308;
assign w26310 = w12636 & w26309;
assign w26311 = w25675 & w26310;
assign v8346 = ~(w324 | w674);
assign w26312 = v8346;
assign w26313 = w1989 & w26312;
assign w26314 = w2156 & w26313;
assign w26315 = w13912 & w26314;
assign w26316 = w1048 & w1653;
assign w26317 = w3231 & w26316;
assign w26318 = w339 & w3279;
assign w26319 = w26317 & w26318;
assign w26320 = w26315 & w26319;
assign w26321 = w5420 & w26320;
assign w26322 = w26311 & w26321;
assign w26323 = ~w26171 & w26322;
assign w26324 = w26171 & ~w26322;
assign v8347 = ~(w26323 | w26324);
assign w26325 = v8347;
assign w26326 = w26307 & w26325;
assign v8348 = ~(w26307 | w26325);
assign w26327 = v8348;
assign v8349 = ~(w26326 | w26327);
assign w26328 = v8349;
assign w26329 = w928 & w21362;
assign w26330 = w3406 & w19974;
assign w26331 = w3402 & w19980;
assign w26332 = w3399 & w19983;
assign v8350 = ~(w26331 | w26332);
assign w26333 = v8350;
assign w26334 = ~w26330 & w26333;
assign w26335 = ~w26329 & w26334;
assign v8351 = ~(w26328 | w26335);
assign w26336 = v8351;
assign w26337 = w26328 & w26335;
assign v8352 = ~(w26336 | w26337);
assign w26338 = v8352;
assign w26339 = w3529 & w20234;
assign w26340 = w3763 & w19966;
assign w26341 = w3760 & w19961;
assign v8353 = ~(w26340 | w26341);
assign w26342 = v8353;
assign w26343 = w3767 & ~w19971;
assign w26344 = w26342 & ~w26343;
assign w26345 = ~w26339 & w26344;
assign w26346 = pi29 & w26345;
assign v8354 = ~(pi29 | w26345);
assign w26347 = v8354;
assign v8355 = ~(w26346 | w26347);
assign w26348 = v8355;
assign w26349 = w26338 & ~w26348;
assign w26350 = ~w26338 & w26348;
assign v8356 = ~(w26349 | w26350);
assign w26351 = v8356;
assign w26352 = ~w26306 & w26351;
assign w26353 = w26306 & ~w26351;
assign v8357 = ~(w26352 | w26353);
assign w26354 = v8357;
assign w26355 = w4153 & ~w21866;
assign w26356 = w4158 & w19952;
assign w26357 = w4155 & w19954;
assign v8358 = ~(w26356 | w26357);
assign w26358 = v8358;
assign w26359 = ~w2873 & w19958;
assign w26360 = w26358 & ~w26359;
assign w26361 = ~w26355 & w26360;
assign w26362 = pi26 & w26361;
assign v8359 = ~(pi26 | w26361);
assign w26363 = v8359;
assign v8360 = ~(w26362 | w26363);
assign w26364 = v8360;
assign w26365 = w26354 & ~w26364;
assign w26366 = ~w26354 & w26364;
assign v8361 = ~(w26365 | w26366);
assign w26367 = v8361;
assign v8362 = ~(w26202 | w26215);
assign w26368 = v8362;
assign w26369 = ~w26367 & w26368;
assign w26370 = w26367 & ~w26368;
assign v8363 = ~(w26369 | w26370);
assign w26371 = v8363;
assign w26372 = w4913 & ~w19929;
assign w26373 = w4763 & ~w19939;
assign w26374 = w4836 & w19933;
assign v8364 = ~(w26373 | w26374);
assign w26375 = v8364;
assign w26376 = ~w26372 & w26375;
assign w26377 = (w26376 & w22285) | (w26376 & w29146) | (w22285 & w29146);
assign w26378 = ~pi23 & w26377;
assign w26379 = pi23 & ~w26377;
assign v8365 = ~(w26378 | w26379);
assign w26380 = v8365;
assign w26381 = w26371 & w26380;
assign v8366 = ~(w26371 | w26380);
assign w26382 = v8366;
assign v8367 = ~(w26381 | w26382);
assign w26383 = v8367;
assign v8368 = ~(w26220 | w26232);
assign w26384 = v8368;
assign w26385 = ~w26383 & w26384;
assign w26386 = w26383 & ~w26384;
assign v8369 = ~(w26385 | w26386);
assign w26387 = v8369;
assign w26388 = w5610 & w19853;
assign w26389 = w5531 & w19917;
assign w26390 = w5113 & ~w19923;
assign v8370 = ~(w26389 | w26390);
assign w26391 = v8370;
assign w26392 = ~w26388 & w26391;
assign w26393 = (~w22936 & w29147) | (~w22936 & w29148) | (w29147 & w29148);
assign w26394 = (w22936 & w29149) | (w22936 & w29150) | (w29149 & w29150);
assign v8371 = ~(w26393 | w26394);
assign w26395 = v8371;
assign w26396 = w26387 & ~w26395;
assign w26397 = ~w26387 & w26395;
assign v8372 = ~(w26396 | w26397);
assign w26398 = v8372;
assign v8373 = ~(w26237 | w26249);
assign w26399 = v8373;
assign w26400 = ~w26398 & w26399;
assign w26401 = w26398 & ~w26399;
assign v8374 = ~(w26400 | w26401);
assign w26402 = v8374;
assign w26403 = w5983 & w20197;
assign w26404 = w6236 & w23607;
assign v8375 = ~(w26403 | w26404);
assign w26405 = v8375;
assign w26406 = w5764 & ~w19912;
assign w26407 = w26405 & ~w26406;
assign w26408 = (w26407 & ~w23614) | (w26407 & w29151) | (~w23614 & w29151);
assign w26409 = pi17 & w26408;
assign v8376 = ~(pi17 | w26408);
assign w26410 = v8376;
assign v8377 = ~(w26409 | w26410);
assign w26411 = v8377;
assign w26412 = w26402 & ~w26411;
assign w26413 = ~w26402 & w26411;
assign v8378 = ~(w26412 | w26413);
assign w26414 = v8378;
assign v8379 = ~(w26254 | w26265);
assign w26415 = v8379;
assign w26416 = ~w26414 & w26415;
assign w26417 = w26414 & ~w26415;
assign v8380 = ~(w26416 | w26417);
assign w26418 = v8380;
assign w26419 = w6389 & w24282;
assign w26420 = w6388 & w23670;
assign w26421 = w7004 & w24284;
assign w26422 = w6871 & ~w24077;
assign v8381 = ~(w26421 | w26422);
assign w26423 = v8381;
assign w26424 = ~w26420 & w26423;
assign w26425 = ~w26419 & w26424;
assign w26426 = pi14 & ~w26425;
assign w26427 = ~pi14 & w26425;
assign v8382 = ~(w26426 | w26427);
assign w26428 = v8382;
assign w26429 = w26418 & w26428;
assign v8383 = ~(w26418 | w26428);
assign w26430 = v8383;
assign v8384 = ~(w26429 | w26430);
assign w26431 = v8384;
assign v8385 = ~(w26270 | w26282);
assign w26432 = v8385;
assign w26433 = ~pi11 & w26432;
assign w26434 = pi11 & ~w26432;
assign v8386 = ~(w26433 | w26434);
assign w26435 = v8386;
assign v8387 = ~(w26431 | w26435);
assign w26436 = v8387;
assign w26437 = w26431 & w26435;
assign v8388 = ~(w26436 | w26437);
assign w26438 = v8388;
assign v8389 = ~(w26285 | w26292);
assign w26439 = v8389;
assign w26440 = ~w26438 & w26439;
assign w26441 = w26438 & ~w26439;
assign v8390 = ~(w26440 | w26441);
assign w26442 = v8390;
assign w26443 = (~w25637 & w28864) | (~w25637 & w28865) | (w28864 & w28865);
assign w26444 = (w25637 & w31307) | (w25637 & w31308) | (w31307 & w31308);
assign w26445 = (~w25637 & w31309) | (~w25637 & w31310) | (w31309 & w31310);
assign v8391 = ~(w26444 | w26445);
assign w26446 = v8391;
assign w26447 = w25989 & w28611;
assign v8392 = ~(w26301 | w26446);
assign w26448 = v8392;
assign v8393 = ~(w26447 | w26448);
assign w26449 = v8393;
assign w26450 = (~w26434 & ~w26435) | (~w26434 & w28612) | (~w26435 & w28612);
assign v8394 = ~(w26401 | w26412);
assign w26451 = v8394;
assign v8395 = ~(w26370 | w26381);
assign w26452 = v8395;
assign v8396 = ~(w26352 | w26365);
assign w26453 = v8396;
assign v8397 = ~(w26336 | w26349);
assign w26454 = v8397;
assign w26455 = ~w211 & w1667;
assign w26456 = ~w479 & w5197;
assign w26457 = w26455 & w26456;
assign w26458 = w2816 & w26457;
assign w26459 = w803 & w2381;
assign w26460 = ~w73 & w26459;
assign w26461 = w26458 & w26460;
assign w26462 = w1170 & w1736;
assign w26463 = w5167 & w26462;
assign w26464 = w2213 & w26463;
assign w26465 = w210 & w26464;
assign w26466 = w26461 & w26465;
assign w26467 = w2251 & w3631;
assign w26468 = w26466 & w26467;
assign v8398 = ~(w26171 | w26468);
assign w26469 = v8398;
assign w26470 = w26171 & w26468;
assign v8399 = ~(w26469 | w26470);
assign w26471 = v8399;
assign w26472 = ~pi11 & w26471;
assign w26473 = pi11 & ~w26471;
assign v8400 = ~(w26472 | w26473);
assign w26474 = v8400;
assign w26475 = w928 & w21401;
assign w26476 = w3406 & ~w19971;
assign w26477 = w3402 & w19974;
assign w26478 = w3399 & w19980;
assign v8401 = ~(w26477 | w26478);
assign w26479 = v8401;
assign w26480 = ~w26476 & w26479;
assign w26481 = ~w26475 & w26480;
assign w26482 = ~w26474 & w26481;
assign w26483 = w26474 & ~w26481;
assign v8402 = ~(w26482 | w26483);
assign w26484 = v8402;
assign v8403 = ~(w26323 | w26326);
assign w26485 = v8403;
assign w26486 = w26484 & w26485;
assign v8404 = ~(w26484 | w26485);
assign w26487 = v8404;
assign v8405 = ~(w26486 | w26487);
assign w26488 = v8405;
assign w26489 = ~w26454 & w26488;
assign w26490 = w26454 & ~w26488;
assign v8406 = ~(w26489 | w26490);
assign w26491 = v8406;
assign w26492 = w3529 & w21716;
assign w26493 = w3760 & w19958;
assign w26494 = w3763 & w19961;
assign w26495 = w3767 & w19966;
assign v8407 = ~(w26494 | w26495);
assign w26496 = v8407;
assign w26497 = ~w26493 & w26496;
assign w26498 = ~w26492 & w26497;
assign w26499 = pi29 & w26498;
assign v8408 = ~(pi29 | w26498);
assign w26500 = v8408;
assign v8409 = ~(w26499 | w26500);
assign w26501 = v8409;
assign w26502 = w26491 & ~w26501;
assign w26503 = ~w26491 & w26501;
assign v8410 = ~(w26502 | w26503);
assign w26504 = v8410;
assign w26505 = w4153 & w20214;
assign w26506 = w4155 & ~w19939;
assign w26507 = ~w2873 & w19952;
assign w26508 = w4158 & w19954;
assign v8411 = ~(w26507 | w26508);
assign w26509 = v8411;
assign w26510 = ~w26506 & w26509;
assign w26511 = ~w26505 & w26510;
assign w26512 = ~pi26 & w26511;
assign w26513 = pi26 & ~w26511;
assign v8412 = ~(w26512 | w26513);
assign w26514 = v8412;
assign w26515 = w26504 & w26514;
assign v8413 = ~(w26504 | w26514);
assign w26516 = v8413;
assign v8414 = ~(w26515 | w26516);
assign w26517 = v8414;
assign w26518 = w26453 & ~w26517;
assign w26519 = ~w26453 & w26517;
assign v8415 = ~(w26518 | w26519);
assign w26520 = v8415;
assign w26521 = w4913 & ~w19923;
assign w26522 = w4763 & w19933;
assign w26523 = w4836 & ~w19929;
assign v8416 = ~(w26522 | w26523);
assign w26524 = v8416;
assign w26525 = ~w26521 & w26524;
assign w26526 = (w26525 & ~w22262) | (w26525 & w29152) | (~w22262 & w29152);
assign w26527 = ~pi23 & w26526;
assign w26528 = pi23 & ~w26526;
assign v8417 = ~(w26527 | w26528);
assign w26529 = v8417;
assign w26530 = w26520 & w26529;
assign v8418 = ~(w26520 | w26529);
assign w26531 = v8418;
assign v8419 = ~(w26530 | w26531);
assign w26532 = v8419;
assign w26533 = w26452 & ~w26532;
assign w26534 = ~w26452 & w26532;
assign v8420 = ~(w26533 | w26534);
assign w26535 = v8420;
assign w26536 = (~w26386 & w26395) | (~w26386 & w28613) | (w26395 & w28613);
assign w26537 = w5610 & ~w19912;
assign w26538 = w5531 & w19853;
assign w26539 = w5113 & w19917;
assign v8421 = ~(w26538 | w26539);
assign w26540 = v8421;
assign w26541 = ~w26537 & w26540;
assign w26542 = (~w22917 & w28866) | (~w22917 & w28867) | (w28866 & w28867);
assign w26543 = (w22917 & w28868) | (w22917 & w28869) | (w28868 & w28869);
assign v8422 = ~(w26542 | w26543);
assign w26544 = v8422;
assign w26545 = ~w26536 & w26544;
assign w26546 = w26536 & ~w26544;
assign v8423 = ~(w26545 | w26546);
assign w26547 = v8423;
assign v8424 = ~(w26535 | w26547);
assign w26548 = v8424;
assign w26549 = w26535 & w26547;
assign v8425 = ~(w26548 | w26549);
assign w26550 = v8425;
assign w26551 = w5983 & w23607;
assign w26552 = w6236 & w23670;
assign v8426 = ~(w26551 | w26552);
assign w26553 = v8426;
assign w26554 = w5764 & w20197;
assign w26555 = w26553 & ~w26554;
assign w26556 = (w26555 & ~w23666) | (w26555 & w28870) | (~w23666 & w28870);
assign w26557 = pi17 & w26556;
assign v8427 = ~(pi17 | w26556);
assign w26558 = v8427;
assign v8428 = ~(w26557 | w26558);
assign w26559 = v8428;
assign w26560 = w26550 & ~w26559;
assign w26561 = ~w26550 & w26559;
assign v8429 = ~(w26560 | w26561);
assign w26562 = v8429;
assign w26563 = w26451 & ~w26562;
assign w26564 = ~w26451 & w26562;
assign v8430 = ~(w26563 | w26564);
assign w26565 = v8430;
assign w26566 = (~w26417 & ~w26418) | (~w26417 & w28615) | (~w26418 & w28615);
assign w26567 = w6389 & ~w24304;
assign w26568 = w6871 & w24284;
assign w26569 = w6388 & ~w24077;
assign v8431 = ~(w26568 | w26569);
assign w26570 = v8431;
assign w26571 = ~w26567 & w26570;
assign w26572 = ~pi14 & w26571;
assign w26573 = pi14 & ~w26571;
assign v8432 = ~(w26572 | w26573);
assign w26574 = v8432;
assign w26575 = ~w26566 & w26574;
assign w26576 = w26566 & ~w26574;
assign v8433 = ~(w26575 | w26576);
assign w26577 = v8433;
assign v8434 = ~(w26565 | w26577);
assign w26578 = v8434;
assign w26579 = w26565 & w26577;
assign v8435 = ~(w26578 | w26579);
assign w26580 = v8435;
assign w26581 = ~w26450 & w26580;
assign w26582 = w26450 & ~w26580;
assign v8436 = ~(w26581 | w26582);
assign w26583 = v8436;
assign w26584 = (w25637 & w28871) | (w25637 & w28872) | (w28871 & w28872);
assign w26585 = ~w26584 & w28109;
assign w26586 = (~w26583 & ~w26443) | (~w26583 & w28616) | (~w26443 & w28616);
assign w26587 = ~w26441 & w26586;
assign v8437 = ~(w26585 | w26587);
assign w26588 = v8437;
assign w26589 = w26447 & w26588;
assign v8438 = ~(w26447 | w26588);
assign w26590 = v8438;
assign v8439 = ~(w26589 | w26590);
assign w26591 = v8439;
assign w26592 = (~w26560 & ~w26562) | (~w26560 & w29153) | (~w26562 & w29153);
assign v8440 = ~(w26489 | w26502);
assign w26593 = v8440;
assign v8441 = ~(w26483 | w26486);
assign w26594 = v8441;
assign v8442 = ~(w26469 | w26472);
assign w26595 = v8442;
assign w26596 = w3558 & w12424;
assign w26597 = w19863 & w26596;
assign w26598 = w24355 & w26597;
assign w26599 = w3015 & w26598;
assign w26600 = ~w223 & w1130;
assign w26601 = ~w234 & w26600;
assign w26602 = w498 & w3745;
assign w26603 = w567 & w26602;
assign w26604 = w26601 & w26603;
assign v8443 = ~(w53 | w381);
assign w26605 = v8443;
assign w26606 = w24761 & w26605;
assign w26607 = w26604 & w26606;
assign w26608 = w26599 & w26607;
assign w26609 = w806 & w13922;
assign w26610 = w26608 & w26609;
assign w26611 = ~w26595 & w26610;
assign w26612 = w26595 & ~w26610;
assign v8444 = ~(w26611 | w26612);
assign w26613 = v8444;
assign w26614 = w928 & w21385;
assign w26615 = w3406 & w19966;
assign w26616 = w3402 & ~w19971;
assign w26617 = w3399 & w19974;
assign v8445 = ~(w26616 | w26617);
assign w26618 = v8445;
assign w26619 = ~w26615 & w26618;
assign w26620 = ~w26614 & w26619;
assign w26621 = w26613 & w26620;
assign v8446 = ~(w26613 | w26620);
assign w26622 = v8446;
assign v8447 = ~(w26621 | w26622);
assign w26623 = v8447;
assign v8448 = ~(w26594 | w26623);
assign w26624 = v8448;
assign w26625 = w26594 & w26623;
assign v8449 = ~(w26624 | w26625);
assign w26626 = v8449;
assign w26627 = w3529 & ~w21882;
assign w26628 = w3760 & w19952;
assign w26629 = w3763 & w19958;
assign w26630 = w3767 & w19961;
assign v8450 = ~(w26629 | w26630);
assign w26631 = v8450;
assign w26632 = ~w26628 & w26631;
assign w26633 = ~w26627 & w26632;
assign w26634 = ~pi29 & w26633;
assign w26635 = pi29 & ~w26633;
assign v8451 = ~(w26634 | w26635);
assign w26636 = v8451;
assign w26637 = w26626 & w26636;
assign v8452 = ~(w26626 | w26636);
assign w26638 = v8452;
assign v8453 = ~(w26637 | w26638);
assign w26639 = v8453;
assign w26640 = ~w26593 & w26639;
assign w26641 = w26593 & ~w26639;
assign v8454 = ~(w26640 | w26641);
assign w26642 = v8454;
assign w26643 = w4153 & ~w22304;
assign w26644 = ~w2873 & w19954;
assign w26645 = w4155 & w19933;
assign v8455 = ~(w26644 | w26645);
assign w26646 = v8455;
assign w26647 = w4158 & ~w19939;
assign w26648 = w26646 & ~w26647;
assign w26649 = ~w26643 & w26648;
assign w26650 = pi26 & w26649;
assign v8456 = ~(pi26 | w26649);
assign w26651 = v8456;
assign v8457 = ~(w26650 | w26651);
assign w26652 = v8457;
assign w26653 = w26642 & ~w26652;
assign w26654 = ~w26642 & w26652;
assign v8458 = ~(w26653 | w26654);
assign w26655 = v8458;
assign v8459 = ~(w26515 | w26519);
assign w26656 = v8459;
assign w26657 = ~w26655 & w26656;
assign w26658 = w26655 & ~w26656;
assign v8460 = ~(w26657 | w26658);
assign w26659 = v8460;
assign w26660 = w4913 & w19917;
assign w26661 = w4763 & ~w19929;
assign w26662 = w4836 & ~w19923;
assign v8461 = ~(w26661 | w26662);
assign w26663 = v8461;
assign w26664 = ~w26660 & w26663;
assign w26665 = (w26664 & w22895) | (w26664 & w29154) | (w22895 & w29154);
assign w26666 = ~pi23 & w26665;
assign w26667 = pi23 & ~w26665;
assign v8462 = ~(w26666 | w26667);
assign w26668 = v8462;
assign w26669 = w26659 & w26668;
assign v8463 = ~(w26659 | w26668);
assign w26670 = v8463;
assign v8464 = ~(w26669 | w26670);
assign w26671 = v8464;
assign v8465 = ~(w26530 | w26534);
assign w26672 = v8465;
assign w26673 = ~w26671 & w26672;
assign w26674 = w26671 & ~w26672;
assign v8466 = ~(w26673 | w26674);
assign w26675 = v8466;
assign w26676 = w5610 & w20197;
assign w26677 = w5531 & ~w19912;
assign w26678 = w5113 & w19853;
assign v8467 = ~(w26677 | w26678);
assign w26679 = v8467;
assign w26680 = ~w26676 & w26679;
assign w26681 = (~w20203 & w29155) | (~w20203 & w29156) | (w29155 & w29156);
assign w26682 = (w20203 & w29157) | (w20203 & w29158) | (w29157 & w29158);
assign v8468 = ~(w26681 | w26682);
assign w26683 = v8468;
assign w26684 = w26675 & w26683;
assign v8469 = ~(w26675 | w26683);
assign w26685 = v8469;
assign v8470 = ~(w26684 | w26685);
assign w26686 = v8470;
assign w26687 = (~w26545 & ~w26547) | (~w26545 & w29159) | (~w26547 & w29159);
assign w26688 = ~w26686 & w26687;
assign w26689 = w26686 & ~w26687;
assign v8471 = ~(w26688 | w26689);
assign w26690 = v8471;
assign w26691 = w5765 & w24073;
assign w26692 = w5983 & w23670;
assign w26693 = w6236 & ~w24077;
assign v8472 = ~(w26692 | w26693);
assign w26694 = v8472;
assign w26695 = w5764 & w23607;
assign w26696 = w26694 & ~w26695;
assign w26697 = ~w26691 & w26696;
assign v8473 = ~(pi17 | w26697);
assign w26698 = v8473;
assign w26699 = pi17 & w26697;
assign v8474 = ~(w26698 | w26699);
assign w26700 = v8474;
assign w26701 = w26690 & ~w26700;
assign w26702 = ~w26690 & w26700;
assign v8475 = ~(w26701 | w26702);
assign w26703 = v8475;
assign w26704 = ~w26592 & w26703;
assign w26705 = w26592 & ~w26703;
assign v8476 = ~(w26704 | w26705);
assign w26706 = v8476;
assign w26707 = w6387 & w24284;
assign v8477 = ~(pi14 | w26707);
assign w26708 = v8477;
assign w26709 = w12684 & w24284;
assign v8478 = ~(w26708 | w26709);
assign w26710 = v8478;
assign w26711 = w26706 & w26710;
assign v8479 = ~(w26706 | w26710);
assign w26712 = v8479;
assign v8480 = ~(w26711 | w26712);
assign w26713 = v8480;
assign v8481 = ~(w26575 | w26579);
assign w26714 = v8481;
assign w26715 = w26713 & ~w26714;
assign w26716 = ~w26713 & w26714;
assign v8482 = ~(w26715 | w26716);
assign w26717 = v8482;
assign w26718 = (~w26584 & w29160) | (~w26584 & w29161) | (w29160 & w29161);
assign w26719 = (w26584 & w29162) | (w26584 & w29163) | (w29162 & w29163);
assign v8483 = ~(w26718 | w26719);
assign w26720 = v8483;
assign w26721 = w26589 & ~w26720;
assign w26722 = ~w26589 & w26720;
assign v8484 = ~(w26721 | w26722);
assign w26723 = v8484;
assign v8485 = ~(w26640 | w26653);
assign w26724 = v8485;
assign v8486 = ~(w26624 | w26637);
assign w26725 = v8486;
assign v8487 = ~(w26612 | w26621);
assign w26726 = v8487;
assign w26727 = w898 & w3110;
assign v8488 = ~(w699 | w874);
assign w26728 = v8488;
assign w26729 = w26727 & w26728;
assign w26730 = w3965 & w12122;
assign w26731 = ~w132 & w6089;
assign w26732 = w4365 & w26731;
assign w26733 = ~w186 & w5330;
assign w26734 = w26732 & w26733;
assign w26735 = w26730 & w26734;
assign w26736 = ~w128 & w3044;
assign w26737 = ~w428 & w26736;
assign w26738 = w2839 & w26737;
assign w26739 = w3682 & w26738;
assign w26740 = w1126 & w26739;
assign w26741 = w26735 & w26740;
assign w26742 = w26729 & w26741;
assign w26743 = ~w26610 & w26742;
assign w26744 = w26610 & ~w26742;
assign v8489 = ~(w26743 | w26744);
assign w26745 = v8489;
assign w26746 = w928 & w20234;
assign w26747 = w3406 & w19961;
assign w26748 = w3402 & w19966;
assign w26749 = w3399 & ~w19971;
assign v8490 = ~(w26748 | w26749);
assign w26750 = v8490;
assign w26751 = ~w26747 & w26750;
assign w26752 = ~w26746 & w26751;
assign v8491 = ~(w26745 | w26752);
assign w26753 = v8491;
assign w26754 = w26745 & w26752;
assign v8492 = ~(w26753 | w26754);
assign w26755 = v8492;
assign w26756 = ~w26726 & w26755;
assign w26757 = w26726 & ~w26755;
assign v8493 = ~(w26756 | w26757);
assign w26758 = v8493;
assign w26759 = w26725 & ~w26758;
assign w26760 = ~w26725 & w26758;
assign v8494 = ~(w26759 | w26760);
assign w26761 = v8494;
assign w26762 = w3529 & ~w21866;
assign w26763 = w3763 & w19952;
assign w26764 = w3760 & w19954;
assign v8495 = ~(w26763 | w26764);
assign w26765 = v8495;
assign w26766 = w3767 & w19958;
assign w26767 = w26765 & ~w26766;
assign w26768 = ~w26762 & w26767;
assign w26769 = pi29 & w26768;
assign v8496 = ~(pi29 | w26768);
assign w26770 = v8496;
assign v8497 = ~(w26769 | w26770);
assign w26771 = v8497;
assign w26772 = ~w26761 & w26771;
assign w26773 = w26761 & ~w26771;
assign v8498 = ~(w26772 | w26773);
assign w26774 = v8498;
assign w26775 = w4155 & ~w19929;
assign v8499 = ~(w2873 | w19939);
assign w26776 = v8499;
assign w26777 = w4158 & w19933;
assign v8500 = ~(w26776 | w26777);
assign w26778 = v8500;
assign w26779 = ~w26775 & w26778;
assign w26780 = (w26779 & w22285) | (w26779 & w29164) | (w22285 & w29164);
assign w26781 = ~pi26 & w26780;
assign w26782 = pi26 & ~w26780;
assign v8501 = ~(w26781 | w26782);
assign w26783 = v8501;
assign w26784 = w26774 & w26783;
assign v8502 = ~(w26774 | w26783);
assign w26785 = v8502;
assign v8503 = ~(w26784 | w26785);
assign w26786 = v8503;
assign w26787 = ~w26724 & w26786;
assign w26788 = w26724 & ~w26786;
assign v8504 = ~(w26787 | w26788);
assign w26789 = v8504;
assign w26790 = w4913 & w19853;
assign w26791 = w4836 & w19917;
assign w26792 = w4763 & ~w19923;
assign v8505 = ~(w26791 | w26792);
assign w26793 = v8505;
assign w26794 = ~w26790 & w26793;
assign w26795 = (~w22936 & w28874) | (~w22936 & w28875) | (w28874 & w28875);
assign w26796 = (w22936 & w28876) | (w22936 & w28877) | (w28876 & w28877);
assign v8506 = ~(w26795 | w26796);
assign w26797 = v8506;
assign w26798 = w26789 & ~w26797;
assign w26799 = ~w26789 & w26797;
assign v8507 = ~(w26798 | w26799);
assign w26800 = v8507;
assign v8508 = ~(w26658 | w26669);
assign w26801 = v8508;
assign w26802 = ~w26800 & w26801;
assign w26803 = w26800 & ~w26801;
assign v8509 = ~(w26802 | w26803);
assign w26804 = v8509;
assign w26805 = w5531 & w20197;
assign w26806 = w5610 & w23607;
assign v8510 = ~(w26805 | w26806);
assign w26807 = v8510;
assign w26808 = w5113 & ~w19912;
assign w26809 = w26807 & ~w26808;
assign w26810 = (~w23614 & w28878) | (~w23614 & w28879) | (w28878 & w28879);
assign w26811 = (w23614 & w28880) | (w23614 & w28881) | (w28880 & w28881);
assign v8511 = ~(w26810 | w26811);
assign w26812 = v8511;
assign w26813 = w26804 & ~w26812;
assign w26814 = ~w26804 & w26812;
assign v8512 = ~(w26813 | w26814);
assign w26815 = v8512;
assign v8513 = ~(w26674 | w26684);
assign w26816 = v8513;
assign w26817 = ~w26815 & w26816;
assign w26818 = w26815 & ~w26816;
assign v8514 = ~(w26817 | w26818);
assign w26819 = v8514;
assign w26820 = ~w24281 & w28882;
assign w26821 = w5983 & ~w24077;
assign w26822 = w6236 & w24284;
assign w26823 = w5764 & w23670;
assign v8515 = ~(w26822 | w26823);
assign w26824 = v8515;
assign w26825 = ~w26821 & w26824;
assign w26826 = ~w26820 & w26825;
assign w26827 = pi17 & ~w26826;
assign w26828 = ~pi17 & w26826;
assign v8516 = ~(w26827 | w26828);
assign w26829 = v8516;
assign w26830 = w26819 & w26829;
assign v8517 = ~(w26819 | w26829);
assign w26831 = v8517;
assign v8518 = ~(w26830 | w26831);
assign w26832 = v8518;
assign v8519 = ~(w26689 | w26701);
assign w26833 = v8519;
assign w26834 = ~pi14 & w26833;
assign w26835 = pi14 & ~w26833;
assign v8520 = ~(w26834 | w26835);
assign w26836 = v8520;
assign v8521 = ~(w26832 | w26836);
assign w26837 = v8521;
assign w26838 = w26832 & w26836;
assign v8522 = ~(w26837 | w26838);
assign w26839 = v8522;
assign v8523 = ~(w26704 | w26711);
assign w26840 = v8523;
assign w26841 = ~w26839 & w26840;
assign w26842 = w26839 & ~w26840;
assign v8524 = ~(w26841 | w26842);
assign w26843 = v8524;
assign w26844 = (w25637 & w29425) | (w25637 & w29426) | (w29425 & w29426);
assign w26845 = (~w26150 & w29165) | (~w26150 & w29166) | (w29165 & w29166);
assign w26846 = (w26150 & w29167) | (w26150 & w29168) | (w29167 & w29168);
assign v8525 = ~(w26845 | w26846);
assign w26847 = v8525;
assign w26848 = w26589 & w28248;
assign v8526 = ~(w26721 | w26847);
assign w26849 = v8526;
assign v8527 = ~(w26848 | w26849);
assign w26850 = v8527;
assign w26851 = (~w26835 & ~w26836) | (~w26835 & w28249) | (~w26836 & w28249);
assign v8528 = ~(w26803 | w26813);
assign w26852 = v8528;
assign v8529 = ~(w26773 | w26784);
assign w26853 = v8529;
assign v8530 = ~(w26757 | w26760);
assign w26854 = v8530;
assign w26855 = w1019 & w1281;
assign w26856 = ~w481 & w1165;
assign w26857 = w3150 & w26856;
assign w26858 = w26855 & w26857;
assign w26859 = w6697 & w26858;
assign w26860 = w1933 & w26859;
assign w26861 = w1383 & w13209;
assign w26862 = ~w108 & w26861;
assign w26863 = w3450 & w26862;
assign w26864 = w26860 & w26863;
assign w26865 = w12966 & w26864;
assign w26866 = w2155 & w26865;
assign v8531 = ~(w26610 | w26866);
assign w26867 = v8531;
assign w26868 = w26610 & w26866;
assign v8532 = ~(w26867 | w26868);
assign w26869 = v8532;
assign w26870 = ~pi14 & w26869;
assign w26871 = pi14 & ~w26869;
assign v8533 = ~(w26870 | w26871);
assign w26872 = v8533;
assign v8534 = ~(w26743 | w26752);
assign w26873 = v8534;
assign v8535 = ~(w26744 | w26873);
assign w26874 = v8535;
assign w26875 = ~w26872 & w26874;
assign w26876 = w26872 & ~w26874;
assign v8536 = ~(w26875 | w26876);
assign w26877 = v8536;
assign w26878 = w928 & w21716;
assign w26879 = w3406 & w19958;
assign w26880 = w3399 & w19966;
assign w26881 = w3402 & w19961;
assign v8537 = ~(w26880 | w26881);
assign w26882 = v8537;
assign w26883 = ~w26879 & w26882;
assign w26884 = ~w26878 & w26883;
assign w26885 = w26877 & ~w26884;
assign w26886 = ~w26877 & w26884;
assign v8538 = ~(w26885 | w26886);
assign w26887 = v8538;
assign w26888 = w3529 & w20214;
assign w26889 = w3763 & w19954;
assign w26890 = w3760 & ~w19939;
assign v8539 = ~(w26889 | w26890);
assign w26891 = v8539;
assign w26892 = w3767 & w19952;
assign w26893 = w26891 & ~w26892;
assign w26894 = ~w26888 & w26893;
assign w26895 = pi29 & w26894;
assign v8540 = ~(pi29 | w26894);
assign w26896 = v8540;
assign v8541 = ~(w26895 | w26896);
assign w26897 = v8541;
assign w26898 = w26887 & ~w26897;
assign w26899 = ~w26887 & w26897;
assign v8542 = ~(w26898 | w26899);
assign w26900 = v8542;
assign w26901 = w26854 & ~w26900;
assign w26902 = ~w26854 & w26900;
assign v8543 = ~(w26901 | w26902);
assign w26903 = v8543;
assign w26904 = w4155 & ~w19923;
assign w26905 = ~w2873 & w19933;
assign w26906 = w4158 & ~w19929;
assign v8544 = ~(w26905 | w26906);
assign w26907 = v8544;
assign w26908 = ~w26904 & w26907;
assign w26909 = (w26908 & ~w22262) | (w26908 & w29169) | (~w22262 & w29169);
assign w26910 = pi26 & ~w26909;
assign w26911 = ~pi26 & w26909;
assign v8545 = ~(w26910 | w26911);
assign w26912 = v8545;
assign v8546 = ~(w26903 | w26912);
assign w26913 = v8546;
assign w26914 = w26903 & w26912;
assign v8547 = ~(w26913 | w26914);
assign w26915 = v8547;
assign w26916 = w26853 & ~w26915;
assign w26917 = ~w26853 & w26915;
assign v8548 = ~(w26916 | w26917);
assign w26918 = v8548;
assign w26919 = (~w26787 & w26797) | (~w26787 & w29170) | (w26797 & w29170);
assign w26920 = w4913 & ~w19912;
assign w26921 = w4836 & w19853;
assign w26922 = w4763 & w19917;
assign v8549 = ~(w26921 | w26922);
assign w26923 = v8549;
assign w26924 = ~w26920 & w26923;
assign w26925 = (~w22917 & w28883) | (~w22917 & w28884) | (w28883 & w28884);
assign w26926 = (w22917 & w28885) | (w22917 & w28886) | (w28885 & w28886);
assign v8550 = ~(w26925 | w26926);
assign w26927 = v8550;
assign w26928 = ~w26919 & w26927;
assign w26929 = w26919 & ~w26927;
assign v8551 = ~(w26928 | w26929);
assign w26930 = v8551;
assign v8552 = ~(w26918 | w26930);
assign w26931 = v8552;
assign w26932 = w26918 & w26930;
assign v8553 = ~(w26931 | w26932);
assign w26933 = v8553;
assign w26934 = w5531 & w23607;
assign w26935 = w5610 & w23670;
assign v8554 = ~(w26934 | w26935);
assign w26936 = v8554;
assign w26937 = w5113 & w20197;
assign w26938 = w26936 & ~w26937;
assign w26939 = (w26938 & ~w23666) | (w26938 & w28887) | (~w23666 & w28887);
assign w26940 = pi20 & w26939;
assign v8555 = ~(pi20 | w26939);
assign w26941 = v8555;
assign v8556 = ~(w26940 | w26941);
assign w26942 = v8556;
assign w26943 = ~w26933 & w26942;
assign w26944 = w26933 & ~w26942;
assign v8557 = ~(w26943 | w26944);
assign w26945 = v8557;
assign w26946 = w26852 & ~w26945;
assign w26947 = ~w26852 & w26945;
assign v8558 = ~(w26946 | w26947);
assign w26948 = v8558;
assign w26949 = (~w26818 & ~w26819) | (~w26818 & w28250) | (~w26819 & w28250);
assign w26950 = w5765 & ~w24304;
assign w26951 = w5983 & w24284;
assign w26952 = w5764 & ~w24077;
assign v8559 = ~(w26951 | w26952);
assign w26953 = v8559;
assign w26954 = ~w26950 & w26953;
assign w26955 = ~pi17 & w26954;
assign w26956 = pi17 & ~w26954;
assign v8560 = ~(w26955 | w26956);
assign w26957 = v8560;
assign w26958 = ~w26949 & w26957;
assign w26959 = w26949 & ~w26957;
assign v8561 = ~(w26958 | w26959);
assign w26960 = v8561;
assign v8562 = ~(w26948 | w26960);
assign w26961 = v8562;
assign w26962 = w26948 & w26960;
assign v8563 = ~(w26961 | w26962);
assign w26963 = v8563;
assign w26964 = ~w26851 & w26963;
assign w26965 = w26851 & ~w26963;
assign v8564 = ~(w26964 | w26965);
assign w26966 = v8564;
assign w26967 = (w26150 & w28888) | (w26150 & w28889) | (w28888 & w28889);
assign w26968 = ~w26967 & w29171;
assign w26969 = (w26966 & w26967) | (w26966 & w29172) | (w26967 & w29172);
assign v8565 = ~(w26968 | w26969);
assign w26970 = v8565;
assign v8566 = ~(w26848 | w26970);
assign w26971 = v8566;
assign w26972 = w26589 & w28620;
assign v8567 = ~(w26971 | w26972);
assign w26973 = v8567;
assign w26974 = (~w26964 & ~w26842) | (~w26964 & w28251) | (~w26842 & w28251);
assign w26975 = (~w26944 & ~w26945) | (~w26944 & w29173) | (~w26945 & w29173);
assign v8568 = ~(w26898 | w26902);
assign w26976 = v8568;
assign v8569 = ~(w26867 | w26870);
assign w26977 = v8569;
assign w26978 = w2280 & w2955;
assign w26979 = ~w271 & w26978;
assign w26980 = w96 & w2077;
assign w26981 = w3733 & w21734;
assign w26982 = w26980 & w26981;
assign w26983 = w26979 & w26982;
assign w26984 = w5181 & w26983;
assign w26985 = w233 & w3690;
assign w26986 = w14592 & w26985;
assign w26987 = w5854 & w13258;
assign w26988 = w26986 & w26987;
assign w26989 = w3228 & w26988;
assign w26990 = w26984 & w26989;
assign w26991 = ~w26977 & w26990;
assign w26992 = w26977 & ~w26990;
assign v8570 = ~(w26991 | w26992);
assign w26993 = v8570;
assign w26994 = w928 & ~w21882;
assign w26995 = w3406 & w19952;
assign w26996 = w3402 & w19958;
assign w26997 = w3399 & w19961;
assign v8571 = ~(w26996 | w26997);
assign w26998 = v8571;
assign w26999 = ~w26995 & w26998;
assign w27000 = ~w26994 & w26999;
assign w27001 = ~w26993 & w27000;
assign w27002 = w26993 & ~w27000;
assign v8572 = ~(w27001 | w27002);
assign w27003 = v8572;
assign v8573 = ~(w26876 | w26885);
assign w27004 = v8573;
assign w27005 = ~w27003 & w27004;
assign w27006 = w27003 & ~w27004;
assign v8574 = ~(w27005 | w27006);
assign w27007 = v8574;
assign w27008 = w3529 & ~w22304;
assign w27009 = w3760 & w19933;
assign w27010 = w3767 & w19954;
assign w27011 = w3763 & ~w19939;
assign v8575 = ~(w27010 | w27011);
assign w27012 = v8575;
assign w27013 = ~w27009 & w27012;
assign w27014 = ~w27008 & w27013;
assign w27015 = ~pi29 & w27014;
assign w27016 = pi29 & ~w27014;
assign v8576 = ~(w27015 | w27016);
assign w27017 = v8576;
assign w27018 = w27007 & w27017;
assign v8577 = ~(w27007 | w27017);
assign w27019 = v8577;
assign v8578 = ~(w27018 | w27019);
assign w27020 = v8578;
assign w27021 = ~w26976 & w27020;
assign w27022 = w26976 & ~w27020;
assign v8579 = ~(w27021 | w27022);
assign w27023 = v8579;
assign w27024 = w4155 & w19917;
assign v8580 = ~(w2873 | w19929);
assign w27025 = v8580;
assign w27026 = w4158 & ~w19923;
assign v8581 = ~(w27025 | w27026);
assign w27027 = v8581;
assign w27028 = ~w27024 & w27027;
assign w27029 = (w27028 & w22895) | (w27028 & w29174) | (w22895 & w29174);
assign w27030 = ~pi26 & w27029;
assign w27031 = pi26 & ~w27029;
assign v8582 = ~(w27030 | w27031);
assign w27032 = v8582;
assign w27033 = w27023 & w27032;
assign v8583 = ~(w27023 | w27032);
assign w27034 = v8583;
assign v8584 = ~(w27033 | w27034);
assign w27035 = v8584;
assign v8585 = ~(w26914 | w26917);
assign w27036 = v8585;
assign w27037 = ~w27035 & w27036;
assign w27038 = w27035 & ~w27036;
assign v8586 = ~(w27037 | w27038);
assign w27039 = v8586;
assign w27040 = w4913 & w20197;
assign w27041 = w4836 & ~w19912;
assign w27042 = w4763 & w19853;
assign v8587 = ~(w27041 | w27042);
assign w27043 = v8587;
assign w27044 = ~w27040 & w27043;
assign w27045 = (~w20203 & w29175) | (~w20203 & w29176) | (w29175 & w29176);
assign w27046 = (w20203 & w29177) | (w20203 & w29178) | (w29177 & w29178);
assign v8588 = ~(w27045 | w27046);
assign w27047 = v8588;
assign w27048 = w27039 & ~w27047;
assign w27049 = ~w27039 & w27047;
assign v8589 = ~(w27048 | w27049);
assign w27050 = v8589;
assign w27051 = (~w26928 & ~w26930) | (~w26928 & w29179) | (~w26930 & w29179);
assign w27052 = ~w27050 & w27051;
assign w27053 = w27050 & ~w27051;
assign v8590 = ~(w27052 | w27053);
assign w27054 = v8590;
assign w27055 = w5114 & w24073;
assign w27056 = w5531 & w23670;
assign w27057 = w5610 & ~w24077;
assign v8591 = ~(w27056 | w27057);
assign w27058 = v8591;
assign w27059 = w5113 & w23607;
assign w27060 = w27058 & ~w27059;
assign w27061 = ~w27055 & w27060;
assign v8592 = ~(pi20 | w27061);
assign w27062 = v8592;
assign w27063 = pi20 & w27061;
assign v8593 = ~(w27062 | w27063);
assign w27064 = v8593;
assign w27065 = w27054 & ~w27064;
assign w27066 = ~w27054 & w27064;
assign v8594 = ~(w27065 | w27066);
assign w27067 = v8594;
assign w27068 = ~w26975 & w27067;
assign w27069 = w26975 & ~w27067;
assign v8595 = ~(w27068 | w27069);
assign w27070 = v8595;
assign w27071 = w5760 & w24284;
assign v8596 = ~(pi17 | w27071);
assign w27072 = v8596;
assign w27073 = w12581 & w24284;
assign v8597 = ~(w27072 | w27073);
assign w27074 = v8597;
assign w27075 = w27070 & w27074;
assign v8598 = ~(w27070 | w27074);
assign w27076 = v8598;
assign v8599 = ~(w27075 | w27076);
assign w27077 = v8599;
assign v8600 = ~(w26958 | w26962);
assign w27078 = v8600;
assign w27079 = ~w27077 & w27078;
assign w27080 = w27077 & ~w27078;
assign v8601 = ~(w27079 | w27080);
assign w27081 = v8601;
assign w27082 = (~w26150 & w28891) | (~w26150 & w28892) | (w28891 & w28892);
assign w27083 = (w26150 & w28893) | (w26150 & w28894) | (w28893 & w28894);
assign v8602 = ~(w27082 | w27083);
assign w27084 = v8602;
assign w27085 = w26589 & w29180;
assign v8603 = ~(w26972 | w27084);
assign w27086 = v8603;
assign v8604 = ~(w27085 | w27086);
assign w27087 = v8604;
assign v8605 = ~(w27006 | w27018);
assign w27088 = v8605;
assign v8606 = ~(w26991 | w27002);
assign w27089 = v8606;
assign w27090 = ~w248 & w14519;
assign w27091 = w3015 & w3868;
assign w27092 = w27090 & w27091;
assign v8607 = ~(w224 | w488);
assign w27093 = v8607;
assign w27094 = w1026 & w27093;
assign v8608 = ~(w298 | w673);
assign w27095 = v8608;
assign w27096 = ~w120 & w27095;
assign w27097 = w27094 & w27096;
assign w27098 = w1418 & w2671;
assign w27099 = w1372 & w27098;
assign w27100 = w27097 & w27099;
assign w27101 = w5362 & w27100;
assign w27102 = w27092 & w27101;
assign w27103 = w2021 & w3117;
assign w27104 = w11933 & w27103;
assign w27105 = w27102 & w27104;
assign w27106 = ~w584 & w27105;
assign w27107 = ~w26990 & w27106;
assign w27108 = w26990 & ~w27106;
assign v8609 = ~(w27107 | w27108);
assign w27109 = v8609;
assign w27110 = w27089 & w27109;
assign v8610 = ~(w27089 | w27109);
assign w27111 = v8610;
assign v8611 = ~(w27110 | w27111);
assign w27112 = v8611;
assign w27113 = w928 & ~w21866;
assign w27114 = w3406 & w19954;
assign w27115 = w3402 & w19952;
assign w27116 = w3399 & w19958;
assign v8612 = ~(w27115 | w27116);
assign w27117 = v8612;
assign w27118 = ~w27114 & w27117;
assign w27119 = ~w27113 & w27118;
assign v8613 = ~(w27112 | w27119);
assign w27120 = v8613;
assign w27121 = w27112 & w27119;
assign v8614 = ~(w27120 | w27121);
assign w27122 = v8614;
assign w27123 = w3529 & ~w22285;
assign w27124 = w3760 & ~w19929;
assign w27125 = w3767 & ~w19939;
assign w27126 = w3763 & w19933;
assign v8615 = ~(w27125 | w27126);
assign w27127 = v8615;
assign w27128 = ~w27124 & w27127;
assign w27129 = ~w27123 & w27128;
assign w27130 = ~pi29 & w27129;
assign w27131 = pi29 & ~w27129;
assign v8616 = ~(w27130 | w27131);
assign w27132 = v8616;
assign w27133 = w27122 & w27132;
assign v8617 = ~(w27122 | w27132);
assign w27134 = v8617;
assign v8618 = ~(w27133 | w27134);
assign w27135 = v8618;
assign w27136 = ~w27088 & w27135;
assign w27137 = w27088 & ~w27135;
assign v8619 = ~(w27136 | w27137);
assign w27138 = v8619;
assign v8620 = ~(w2873 | w19923);
assign w27139 = v8620;
assign w27140 = w4155 & w19853;
assign v8621 = ~(w27139 | w27140);
assign w27141 = v8621;
assign w27142 = w4158 & w19917;
assign w27143 = w27141 & ~w27142;
assign w27144 = (~w22936 & w29181) | (~w22936 & w29182) | (w29181 & w29182);
assign w27145 = (w22936 & w29183) | (w22936 & w29184) | (w29183 & w29184);
assign v8622 = ~(w27144 | w27145);
assign w27146 = v8622;
assign w27147 = w27138 & ~w27146;
assign w27148 = ~w27138 & w27146;
assign v8623 = ~(w27147 | w27148);
assign w27149 = v8623;
assign v8624 = ~(w27021 | w27033);
assign w27150 = v8624;
assign w27151 = ~w27149 & w27150;
assign w27152 = w27149 & ~w27150;
assign v8625 = ~(w27151 | w27152);
assign w27153 = v8625;
assign w27154 = w4836 & w20197;
assign w27155 = w4913 & w23607;
assign v8626 = ~(w27154 | w27155);
assign w27156 = v8626;
assign w27157 = w4763 & ~w19912;
assign w27158 = w27156 & ~w27157;
assign w27159 = (~w23614 & w29185) | (~w23614 & w29186) | (w29185 & w29186);
assign w27160 = (w23614 & w29187) | (w23614 & w29188) | (w29187 & w29188);
assign v8627 = ~(w27159 | w27160);
assign w27161 = v8627;
assign w27162 = w27153 & ~w27161;
assign w27163 = ~w27153 & w27161;
assign v8628 = ~(w27162 | w27163);
assign w27164 = v8628;
assign v8629 = ~(w27038 | w27048);
assign w27165 = v8629;
assign w27166 = ~w27164 & w27165;
assign w27167 = w27164 & ~w27165;
assign v8630 = ~(w27166 | w27167);
assign w27168 = v8630;
assign w27169 = w5114 & w24282;
assign w27170 = w5113 & w23670;
assign w27171 = w5610 & w24284;
assign w27172 = w5531 & ~w24077;
assign v8631 = ~(w27171 | w27172);
assign w27173 = v8631;
assign w27174 = ~w27170 & w27173;
assign w27175 = ~w27169 & w27174;
assign w27176 = pi20 & ~w27175;
assign w27177 = ~pi20 & w27175;
assign v8632 = ~(w27176 | w27177);
assign w27178 = v8632;
assign w27179 = w27168 & w27178;
assign v8633 = ~(w27168 | w27178);
assign w27180 = v8633;
assign v8634 = ~(w27179 | w27180);
assign w27181 = v8634;
assign v8635 = ~(w27053 | w27065);
assign w27182 = v8635;
assign w27183 = ~pi17 & w27182;
assign w27184 = pi17 & ~w27182;
assign v8636 = ~(w27183 | w27184);
assign w27185 = v8636;
assign v8637 = ~(w27181 | w27185);
assign w27186 = v8637;
assign w27187 = w27181 & w27185;
assign v8638 = ~(w27186 | w27187);
assign w27188 = v8638;
assign v8639 = ~(w27068 | w27075);
assign w27189 = v8639;
assign w27190 = ~w27188 & w27189;
assign w27191 = w27188 & ~w27189;
assign v8640 = ~(w27190 | w27191);
assign w27192 = v8640;
assign w27193 = (~w26150 & w28895) | (~w26150 & w28896) | (w28895 & w28896);
assign w27194 = (w26150 & w28897) | (w26150 & w28898) | (w28897 & w28898);
assign v8641 = ~(w27193 | w27194);
assign w27195 = v8641;
assign w27196 = w26589 & w29189;
assign v8642 = ~(w27085 | w27195);
assign w27197 = v8642;
assign v8643 = ~(w27196 | w27197);
assign w27198 = v8643;
assign v8644 = ~(w27184 | w27187);
assign w27199 = v8644;
assign v8645 = ~(w27152 | w27162);
assign w27200 = v8645;
assign v8646 = ~(w27136 | w27147);
assign w27201 = v8646;
assign w27202 = w4155 & ~w19912;
assign w27203 = ~w2873 & w19917;
assign w27204 = w4158 & w19853;
assign v8647 = ~(w27203 | w27204);
assign w27205 = v8647;
assign w27206 = ~w27202 & w27205;
assign w27207 = (~w22917 & w29190) | (~w22917 & w29191) | (w29190 & w29191);
assign w27208 = (w22917 & w29192) | (w22917 & w29193) | (w29192 & w29193);
assign v8648 = ~(w27207 | w27208);
assign w27209 = v8648;
assign w27210 = ~w27201 & w27209;
assign w27211 = w27201 & ~w27209;
assign v8649 = ~(w27210 | w27211);
assign w27212 = v8649;
assign v8650 = ~(w27120 | w27133);
assign w27213 = v8650;
assign w27214 = w1852 & w3257;
assign w27215 = w1579 & w27214;
assign w27216 = w270 & w1969;
assign w27217 = w27215 & w27216;
assign w27218 = w3443 & w27217;
assign w27219 = ~w42 & w1465;
assign w27220 = w21731 & w27219;
assign w27221 = ~w522 & w27220;
assign w27222 = w941 & w27221;
assign w27223 = w4986 & w27222;
assign w27224 = w27218 & w27223;
assign w27225 = w27105 & w27224;
assign w27226 = ~w584 & w27224;
assign v8651 = ~(w27106 | w27226);
assign w27227 = v8651;
assign v8652 = ~(w27225 | w27227);
assign w27228 = v8652;
assign w27229 = ~pi17 & w27228;
assign w27230 = pi17 & ~w27228;
assign v8653 = ~(w27229 | w27230);
assign w27231 = v8653;
assign w27232 = w928 & w20214;
assign w27233 = w3406 & ~w19939;
assign w27234 = w3402 & w19954;
assign w27235 = w3399 & w19952;
assign v8654 = ~(w27234 | w27235);
assign w27236 = v8654;
assign w27237 = ~w27233 & w27236;
assign w27238 = ~w27232 & w27237;
assign w27239 = ~w27231 & w27238;
assign w27240 = w27231 & ~w27238;
assign v8655 = ~(w27239 | w27240);
assign w27241 = v8655;
assign v8656 = ~(w27108 | w27110);
assign w27242 = v8656;
assign w27243 = w27241 & w27242;
assign v8657 = ~(w27241 | w27242);
assign w27244 = v8657;
assign v8658 = ~(w27243 | w27244);
assign w27245 = v8658;
assign w27246 = ~w27213 & w27245;
assign w27247 = w27213 & ~w27245;
assign v8659 = ~(w27246 | w27247);
assign w27248 = v8659;
assign w27249 = w3529 & w22262;
assign w27250 = w3760 & ~w19923;
assign w27251 = w3767 & w19933;
assign w27252 = w3763 & ~w19929;
assign v8660 = ~(w27251 | w27252);
assign w27253 = v8660;
assign w27254 = ~w27250 & w27253;
assign w27255 = ~w27249 & w27254;
assign w27256 = ~pi29 & w27255;
assign w27257 = pi29 & ~w27255;
assign v8661 = ~(w27256 | w27257);
assign w27258 = v8661;
assign w27259 = w27248 & w27258;
assign v8662 = ~(w27248 | w27258);
assign w27260 = v8662;
assign v8663 = ~(w27259 | w27260);
assign w27261 = v8663;
assign w27262 = w27212 & w27261;
assign v8664 = ~(w27212 | w27261);
assign w27263 = v8664;
assign v8665 = ~(w27262 | w27263);
assign w27264 = v8665;
assign w27265 = w4764 & w23666;
assign w27266 = w4836 & w23607;
assign w27267 = w4913 & w23670;
assign v8666 = ~(w27266 | w27267);
assign w27268 = v8666;
assign w27269 = w4763 & w20197;
assign w27270 = w27268 & ~w27269;
assign w27271 = ~w27265 & w27270;
assign w27272 = pi23 & w27271;
assign v8667 = ~(pi23 | w27271);
assign w27273 = v8667;
assign v8668 = ~(w27272 | w27273);
assign w27274 = v8668;
assign w27275 = ~w27264 & w27274;
assign w27276 = w27264 & ~w27274;
assign v8669 = ~(w27275 | w27276);
assign w27277 = v8669;
assign w27278 = w27200 & ~w27277;
assign w27279 = ~w27200 & w27277;
assign v8670 = ~(w27278 | w27279);
assign w27280 = v8670;
assign v8671 = ~(w27167 | w27179);
assign w27281 = v8671;
assign w27282 = w5114 & ~w24304;
assign w27283 = w5531 & w24284;
assign w27284 = w5113 & ~w24077;
assign v8672 = ~(w27283 | w27284);
assign w27285 = v8672;
assign w27286 = ~w27282 & w27285;
assign w27287 = ~pi20 & w27286;
assign w27288 = pi20 & ~w27286;
assign v8673 = ~(w27287 | w27288);
assign w27289 = v8673;
assign w27290 = ~w27281 & w27289;
assign w27291 = w27281 & ~w27289;
assign v8674 = ~(w27290 | w27291);
assign w27292 = v8674;
assign v8675 = ~(w27280 | w27292);
assign w27293 = v8675;
assign w27294 = w27280 & w27292;
assign v8676 = ~(w27293 | w27294);
assign w27295 = v8676;
assign w27296 = ~w27199 & w27295;
assign w27297 = w27199 & ~w27295;
assign v8677 = ~(w27296 | w27297);
assign w27298 = v8677;
assign w27299 = (w26150 & w29427) | (w26150 & w29428) | (w29427 & w29428);
assign w27300 = (~w26150 & w29429) | (~w26150 & w29430) | (w29429 & w29430);
assign v8678 = ~(w27299 | w27300);
assign w27301 = v8678;
assign v8679 = ~(w27196 | w27301);
assign w27302 = v8679;
assign w27303 = w26589 & w29194;
assign v8680 = ~(w27302 | w27303);
assign w27304 = v8680;
assign v8681 = ~(w27276 | w27279);
assign w27305 = v8681;
assign v8682 = ~(w27246 | w27259);
assign w27306 = v8682;
assign v8683 = ~(w27227 | w27229);
assign w27307 = v8683;
assign w27308 = w1600 & w13928;
assign w27309 = ~w525 & w1603;
assign w27310 = w27308 & w27309;
assign w27311 = w600 & w27310;
assign w27312 = w651 & w27311;
assign w27313 = w3618 & w27312;
assign w27314 = w6484 & w27313;
assign w27315 = ~w108 & w3156;
assign w27316 = ~w192 & w3180;
assign w27317 = ~w338 & w4456;
assign w27318 = w27316 & w27317;
assign w27319 = w27315 & w27318;
assign w27320 = w25859 & w27319;
assign w27321 = w27314 & w27320;
assign w27322 = ~w27307 & w27321;
assign w27323 = w27307 & ~w27321;
assign v8684 = ~(w27322 | w27323);
assign w27324 = v8684;
assign w27325 = w928 & ~w22304;
assign w27326 = w3406 & w19933;
assign w27327 = w3399 & w19954;
assign w27328 = w3402 & ~w19939;
assign v8685 = ~(w27327 | w27328);
assign w27329 = v8685;
assign w27330 = ~w27326 & w27329;
assign w27331 = ~w27325 & w27330;
assign w27332 = ~w27324 & w27331;
assign w27333 = w27324 & ~w27331;
assign v8686 = ~(w27332 | w27333);
assign w27334 = v8686;
assign v8687 = ~(w27240 | w27243);
assign w27335 = v8687;
assign w27336 = ~w27334 & w27335;
assign w27337 = w27334 & ~w27335;
assign v8688 = ~(w27336 | w27337);
assign w27338 = v8688;
assign w27339 = w3760 & w19917;
assign w27340 = w3767 & ~w19929;
assign w27341 = w3763 & ~w19923;
assign v8689 = ~(w27340 | w27341);
assign w27342 = v8689;
assign w27343 = ~w27339 & w27342;
assign w27344 = (w22895 & w29195) | (w22895 & w29196) | (w29195 & w29196);
assign w27345 = (~w22895 & w29197) | (~w22895 & w29198) | (w29197 & w29198);
assign v8690 = ~(w27344 | w27345);
assign w27346 = v8690;
assign w27347 = w27338 & w27346;
assign v8691 = ~(w27338 | w27346);
assign w27348 = v8691;
assign v8692 = ~(w27347 | w27348);
assign w27349 = v8692;
assign w27350 = ~w27306 & w27349;
assign w27351 = w27306 & ~w27349;
assign v8693 = ~(w27350 | w27351);
assign w27352 = v8693;
assign w27353 = w4155 & w20197;
assign w27354 = ~w2873 & w19853;
assign w27355 = w4158 & ~w19912;
assign v8694 = ~(w27354 | w27355);
assign w27356 = v8694;
assign w27357 = ~w27353 & w27356;
assign w27358 = (w27357 & ~w20203) | (w27357 & w29199) | (~w20203 & w29199);
assign w27359 = ~pi26 & w27358;
assign w27360 = pi26 & ~w27358;
assign v8695 = ~(w27359 | w27360);
assign w27361 = v8695;
assign w27362 = w27352 & w27361;
assign v8696 = ~(w27352 | w27361);
assign w27363 = v8696;
assign v8697 = ~(w27362 | w27363);
assign w27364 = v8697;
assign v8698 = ~(w27210 | w27262);
assign w27365 = v8698;
assign w27366 = ~w27364 & w27365;
assign w27367 = w27364 & ~w27365;
assign v8699 = ~(w27366 | w27367);
assign w27368 = v8699;
assign w27369 = w4764 & w24073;
assign w27370 = w4836 & w23670;
assign w27371 = w4913 & ~w24077;
assign v8700 = ~(w27370 | w27371);
assign w27372 = v8700;
assign w27373 = w4763 & w23607;
assign w27374 = w27372 & ~w27373;
assign w27375 = ~w27369 & w27374;
assign w27376 = pi23 & w27375;
assign v8701 = ~(pi23 | w27375);
assign w27377 = v8701;
assign v8702 = ~(w27376 | w27377);
assign w27378 = v8702;
assign w27379 = w27368 & ~w27378;
assign w27380 = ~w27368 & w27378;
assign v8703 = ~(w27379 | w27380);
assign w27381 = v8703;
assign w27382 = ~w27305 & w27381;
assign w27383 = w27305 & ~w27381;
assign v8704 = ~(w27382 | w27383);
assign w27384 = v8704;
assign w27385 = w916 & w24284;
assign v8705 = ~(pi20 | w27385);
assign w27386 = v8705;
assign w27387 = w918 & w24284;
assign v8706 = ~(w27386 | w27387);
assign w27388 = v8706;
assign w27389 = w27384 & w27388;
assign v8707 = ~(w27384 | w27388);
assign w27390 = v8707;
assign v8708 = ~(w27389 | w27390);
assign w27391 = v8708;
assign v8709 = ~(w27290 | w27294);
assign w27392 = v8709;
assign w27393 = w27391 & ~w27392;
assign w27394 = ~w27391 & w27392;
assign v8710 = ~(w27393 | w27394);
assign w27395 = v8710;
assign w27396 = (~w26150 & w29431) | (~w26150 & w29432) | (w29431 & w29432);
assign w27397 = (w26150 & w29433) | (w26150 & w29434) | (w29433 & w29434);
assign v8711 = ~(w27396 | w27397);
assign w27398 = v8711;
assign w27399 = w26972 & w28125;
assign w27400 = ~w27303 & w27398;
assign v8712 = ~(w27399 | w27400);
assign w27401 = v8712;
assign v8713 = ~(w27350 | w27362);
assign w27402 = v8713;
assign v8714 = ~(w27337 | w27347);
assign w27403 = v8714;
assign v8715 = ~(w27322 | w27333);
assign w27404 = v8715;
assign w27405 = w75 & w25119;
assign w27406 = w1607 & w27405;
assign w27407 = w2496 & w27090;
assign w27408 = w3437 & w27407;
assign w27409 = w2951 & w12650;
assign w27410 = w27408 & w27409;
assign w27411 = w6545 & w27410;
assign w27412 = w767 & w4682;
assign w27413 = w751 & w27412;
assign w27414 = w27411 & w27413;
assign w27415 = w27406 & w27414;
assign w27416 = ~w27321 & w27415;
assign w27417 = w27321 & ~w27415;
assign v8716 = ~(w27416 | w27417);
assign w27418 = v8716;
assign w27419 = w928 & ~w22285;
assign w27420 = w3406 & ~w19929;
assign w27421 = w3399 & ~w19939;
assign w27422 = w3402 & w19933;
assign v8717 = ~(w27421 | w27422);
assign w27423 = v8717;
assign w27424 = ~w27420 & w27423;
assign w27425 = ~w27419 & w27424;
assign w27426 = ~w27418 & w27425;
assign w27427 = w27418 & ~w27425;
assign v8718 = ~(w27426 | w27427);
assign w27428 = v8718;
assign w27429 = ~w27404 & w27428;
assign w27430 = w27404 & ~w27428;
assign v8719 = ~(w27429 | w27430);
assign w27431 = v8719;
assign w27432 = w27403 & ~w27431;
assign w27433 = ~w27403 & w27431;
assign v8720 = ~(w27432 | w27433);
assign w27434 = v8720;
assign w27435 = w3529 & w22936;
assign w27436 = w3760 & w19853;
assign w27437 = w3763 & w19917;
assign w27438 = w3767 & ~w19923;
assign v8721 = ~(w27437 | w27438);
assign w27439 = v8721;
assign w27440 = ~w27436 & w27439;
assign w27441 = ~w27435 & w27440;
assign w27442 = pi29 & w27441;
assign v8722 = ~(pi29 | w27441);
assign w27443 = v8722;
assign v8723 = ~(w27442 | w27443);
assign w27444 = v8723;
assign w27445 = ~w27434 & w27444;
assign w27446 = w27434 & ~w27444;
assign v8724 = ~(w27445 | w27446);
assign w27447 = v8724;
assign w27448 = w4155 & w23607;
assign v8725 = ~(w2873 | w19912);
assign w27449 = v8725;
assign w27450 = w4158 & w20197;
assign v8726 = ~(w27449 | w27450);
assign w27451 = v8726;
assign w27452 = ~w27448 & w27451;
assign w27453 = (~w23614 & w29200) | (~w23614 & w29201) | (w29200 & w29201);
assign w27454 = (w23614 & w29202) | (w23614 & w29203) | (w29202 & w29203);
assign v8727 = ~(w27453 | w27454);
assign w27455 = v8727;
assign w27456 = w27447 & w27455;
assign v8728 = ~(w27447 | w27455);
assign w27457 = v8728;
assign v8729 = ~(w27456 | w27457);
assign w27458 = v8729;
assign w27459 = ~w27402 & w27458;
assign w27460 = w27402 & ~w27458;
assign v8730 = ~(w27459 | w27460);
assign w27461 = v8730;
assign w27462 = w4764 & w24282;
assign w27463 = w4763 & w23670;
assign w27464 = w4913 & w24284;
assign v8731 = ~(w27463 | w27464);
assign w27465 = v8731;
assign w27466 = w4836 & ~w24077;
assign w27467 = w27465 & ~w27466;
assign w27468 = ~w27462 & w27467;
assign w27469 = pi23 & w27468;
assign v8732 = ~(pi23 | w27468);
assign w27470 = v8732;
assign v8733 = ~(w27469 | w27470);
assign w27471 = v8733;
assign w27472 = w27461 & ~w27471;
assign w27473 = ~w27461 & w27471;
assign v8734 = ~(w27472 | w27473);
assign w27474 = v8734;
assign v8735 = ~(w27367 | w27379);
assign w27475 = v8735;
assign w27476 = ~pi20 & w27475;
assign w27477 = pi20 & ~w27475;
assign v8736 = ~(w27476 | w27477);
assign w27478 = v8736;
assign v8737 = ~(w27474 | w27478);
assign w27479 = v8737;
assign w27480 = w27474 & w27478;
assign v8738 = ~(w27479 | w27480);
assign w27481 = v8738;
assign v8739 = ~(w27382 | w27389);
assign w27482 = v8739;
assign w27483 = ~w27481 & w27482;
assign w27484 = w27481 & ~w27482;
assign v8740 = ~(w27483 | w27484);
assign w27485 = v8740;
assign w27486 = (w26150 & w28903) | (w26150 & w28904) | (w28903 & w28904);
assign w27487 = (~w26150 & w29435) | (~w26150 & w29436) | (w29435 & w29436);
assign w27488 = (w26150 & w29437) | (w26150 & w29438) | (w29437 & w29438);
assign v8741 = ~(w27487 | w27488);
assign w27489 = v8741;
assign w27490 = w26972 & w28130;
assign w27491 = (~w27489 & ~w26972) | (~w27489 & w29204) | (~w26972 & w29204);
assign v8742 = ~(w27490 | w27491);
assign w27492 = v8742;
assign v8743 = ~(w27477 | w27480);
assign w27493 = v8743;
assign v8744 = ~(w27446 | w27456);
assign w27494 = v8744;
assign w27495 = ~w428 & w3742;
assign w27496 = ~w303 & w1093;
assign w27497 = w900 & w1201;
assign w27498 = w6103 & w27497;
assign w27499 = w27496 & w27498;
assign w27500 = w3291 & w4046;
assign w27501 = w27499 & w27500;
assign w27502 = w27495 & w27501;
assign w27503 = w1547 & w1560;
assign w27504 = w3117 & w27503;
assign w27505 = w13678 & w27504;
assign w27506 = w27502 & w27505;
assign w27507 = w14528 & w27506;
assign w27508 = w157 & w1883;
assign w27509 = w27507 & w27508;
assign v8745 = ~(w27321 | w27509);
assign w27510 = v8745;
assign w27511 = w27321 & w27509;
assign v8746 = ~(w27510 | w27511);
assign w27512 = v8746;
assign w27513 = ~pi20 & w27512;
assign w27514 = pi20 & ~w27512;
assign v8747 = ~(w27513 | w27514);
assign w27515 = v8747;
assign v8748 = ~(w27416 | w27425);
assign w27516 = v8748;
assign v8749 = ~(w27417 | w27516);
assign w27517 = v8749;
assign w27518 = ~w27515 & w27517;
assign w27519 = w27515 & ~w27517;
assign v8750 = ~(w27518 | w27519);
assign w27520 = v8750;
assign w27521 = w928 & w22262;
assign w27522 = w3406 & ~w19923;
assign w27523 = w3399 & w19933;
assign w27524 = w3402 & ~w19929;
assign v8751 = ~(w27523 | w27524);
assign w27525 = v8751;
assign w27526 = ~w27522 & w27525;
assign w27527 = ~w27521 & w27526;
assign w27528 = w27520 & ~w27527;
assign w27529 = ~w27520 & w27527;
assign v8752 = ~(w27528 | w27529);
assign w27530 = v8752;
assign v8753 = ~(w27429 | w27433);
assign w27531 = v8753;
assign w27532 = ~w27530 & w27531;
assign w27533 = w27530 & ~w27531;
assign v8754 = ~(w27532 | w27533);
assign w27534 = v8754;
assign w27535 = w3529 & w22917;
assign w27536 = w3760 & ~w19912;
assign w27537 = w3763 & w19853;
assign w27538 = w3767 & w19917;
assign v8755 = ~(w27537 | w27538);
assign w27539 = v8755;
assign w27540 = ~w27536 & w27539;
assign w27541 = ~w27535 & w27540;
assign w27542 = pi29 & ~w27541;
assign w27543 = ~pi29 & w27541;
assign v8756 = ~(w27542 | w27543);
assign w27544 = v8756;
assign w27545 = w27534 & w27544;
assign v8757 = ~(w27534 | w27544);
assign w27546 = v8757;
assign v8758 = ~(w27545 | w27546);
assign w27547 = v8758;
assign w27548 = w4153 & w23666;
assign w27549 = w4158 & w23607;
assign w27550 = w4155 & w23670;
assign v8759 = ~(w27549 | w27550);
assign w27551 = v8759;
assign w27552 = ~w2873 & w20197;
assign w27553 = w27551 & ~w27552;
assign w27554 = ~w27548 & w27553;
assign v8760 = ~(pi26 | w27554);
assign w27555 = v8760;
assign w27556 = pi26 & w27554;
assign v8761 = ~(w27555 | w27556);
assign w27557 = v8761;
assign w27558 = w27547 & ~w27557;
assign w27559 = ~w27547 & w27557;
assign v8762 = ~(w27558 | w27559);
assign w27560 = v8762;
assign w27561 = w27494 & ~w27560;
assign w27562 = ~w27494 & w27560;
assign v8763 = ~(w27561 | w27562);
assign w27563 = v8763;
assign v8764 = ~(w27459 | w27472);
assign w27564 = v8764;
assign w27565 = w4764 & ~w24304;
assign w27566 = w4836 & w24284;
assign w27567 = w4763 & ~w24077;
assign v8765 = ~(w27566 | w27567);
assign w27568 = v8765;
assign w27569 = ~w27565 & w27568;
assign w27570 = ~pi23 & w27569;
assign w27571 = pi23 & ~w27569;
assign v8766 = ~(w27570 | w27571);
assign w27572 = v8766;
assign w27573 = ~w27564 & w27572;
assign w27574 = w27564 & ~w27572;
assign v8767 = ~(w27573 | w27574);
assign w27575 = v8767;
assign v8768 = ~(w27563 | w27575);
assign w27576 = v8768;
assign w27577 = w27563 & w27575;
assign v8769 = ~(w27576 | w27577);
assign w27578 = v8769;
assign w27579 = ~w27493 & w27578;
assign w27580 = w27493 & ~w27578;
assign v8770 = ~(w27579 | w27580);
assign w27581 = v8770;
assign w27582 = ~w27483 & w27581;
assign w27583 = (w26844 & w28252) | (w26844 & w28253) | (w28252 & w28253);
assign w27584 = w27582 & ~w27583;
assign w27585 = (~w27484 & ~w27486) | (~w27484 & w28254) | (~w27486 & w28254);
assign w27586 = ~w27581 & w27585;
assign v8771 = ~(w27584 | w27586);
assign w27587 = v8771;
assign w27588 = (~w27587 & ~w26972) | (~w27587 & w29205) | (~w26972 & w29205);
assign w27589 = w26972 & w28133;
assign v8772 = ~(w27588 | w27589);
assign w27590 = v8772;
assign v8773 = ~(w27533 | w27545);
assign w27591 = v8773;
assign v8774 = ~(w27510 | w27513);
assign w27592 = v8774;
assign w27593 = w802 & w5364;
assign w27594 = ~w624 & w6072;
assign w27595 = w2732 & w27594;
assign w27596 = w27593 & w27595;
assign w27597 = w1920 & w14597;
assign w27598 = ~w74 & w27597;
assign w27599 = w27596 & w27598;
assign w27600 = w395 & w1017;
assign w27601 = w2345 & w2443;
assign w27602 = w2401 & w27601;
assign w27603 = w826 & w27602;
assign w27604 = w27600 & w27603;
assign w27605 = w3443 & w27604;
assign w27606 = w27599 & w27605;
assign w27607 = ~w27592 & w27606;
assign w27608 = w27592 & ~w27606;
assign v8775 = ~(w27607 | w27608);
assign w27609 = v8775;
assign w27610 = w928 & ~w22895;
assign w27611 = w3406 & w19917;
assign w27612 = w3399 & ~w19929;
assign w27613 = w3402 & ~w19923;
assign v8776 = ~(w27612 | w27613);
assign w27614 = v8776;
assign w27615 = ~w27611 & w27614;
assign w27616 = ~w27610 & w27615;
assign w27617 = ~w27609 & w27616;
assign w27618 = w27609 & ~w27616;
assign v8777 = ~(w27617 | w27618);
assign w27619 = v8777;
assign v8778 = ~(w27519 | w27528);
assign w27620 = v8778;
assign w27621 = ~w27619 & w27620;
assign w27622 = w27619 & ~w27620;
assign v8779 = ~(w27621 | w27622);
assign w27623 = v8779;
assign w27624 = w3763 & ~w19912;
assign w27625 = w3760 & w20197;
assign v8780 = ~(w27624 | w27625);
assign w27626 = v8780;
assign w27627 = w3767 & w19853;
assign w27628 = w27626 & ~w27627;
assign w27629 = (w27628 & ~w20203) | (w27628 & w29206) | (~w20203 & w29206);
assign w27630 = pi29 & w27629;
assign v8781 = ~(pi29 | w27629);
assign w27631 = v8781;
assign v8782 = ~(w27630 | w27631);
assign w27632 = v8782;
assign w27633 = w27623 & ~w27632;
assign w27634 = ~w27623 & w27632;
assign v8783 = ~(w27633 | w27634);
assign w27635 = v8783;
assign w27636 = ~w27591 & w27635;
assign w27637 = w27591 & ~w27635;
assign v8784 = ~(w27636 | w27637);
assign w27638 = v8784;
assign w27639 = w4153 & w24073;
assign w27640 = ~w2873 & w23607;
assign w27641 = w4155 & ~w24077;
assign v8785 = ~(w27640 | w27641);
assign w27642 = v8785;
assign w27643 = w4158 & w23670;
assign w27644 = w27642 & ~w27643;
assign w27645 = ~w27639 & w27644;
assign v8786 = ~(pi26 | w27645);
assign w27646 = v8786;
assign w27647 = pi26 & w27645;
assign v8787 = ~(w27646 | w27647);
assign w27648 = v8787;
assign w27649 = w27638 & ~w27648;
assign w27650 = ~w27638 & w27648;
assign v8788 = ~(w27649 | w27650);
assign w27651 = v8788;
assign v8789 = ~(w27558 | w27562);
assign w27652 = v8789;
assign w27653 = ~w27651 & w27652;
assign w27654 = w27651 & ~w27652;
assign v8790 = ~(w27653 | w27654);
assign w27655 = v8790;
assign w27656 = w11 & w24284;
assign v8791 = ~(pi23 | w27656);
assign w27657 = v8791;
assign w27658 = w13 & w24284;
assign v8792 = ~(w27657 | w27658);
assign w27659 = v8792;
assign w27660 = w27655 & w27659;
assign v8793 = ~(w27655 | w27659);
assign w27661 = v8793;
assign v8794 = ~(w27660 | w27661);
assign w27662 = v8794;
assign v8795 = ~(w27573 | w27577);
assign w27663 = v8795;
assign w27664 = w27662 & ~w27663;
assign w27665 = ~w27662 & w27663;
assign v8796 = ~(w27664 | w27665);
assign w27666 = v8796;
assign w27667 = w27579 & ~w27666;
assign w27668 = ~w27579 & w27666;
assign v8797 = ~(w27667 | w27668);
assign w27669 = v8797;
assign w27670 = (w26972 & w31311) | (w26972 & w31312) | (w31311 & w31312);
assign w27671 = (~w26972 & w31313) | (~w26972 & w31314) | (w31313 & w31314);
assign v8798 = ~(w27670 | w27671);
assign w27672 = v8798;
assign w27673 = w26972 & w28134;
assign v8799 = ~(w27622 | w27633);
assign w27674 = v8799;
assign v8800 = ~(w27607 | w27618);
assign w27675 = v8800;
assign w27676 = w654 & w1476;
assign w27677 = w1048 & w3644;
assign v8801 = ~(w183 | w235);
assign w27678 = v8801;
assign w27679 = w386 & w802;
assign w27680 = w27678 & w27679;
assign w27681 = w27677 & w27680;
assign w27682 = w27676 & w27681;
assign w27683 = w12338 & w27682;
assign w27684 = w4584 & w27683;
assign w27685 = ~w312 & w1722;
assign w27686 = w14437 & w27685;
assign w27687 = ~w605 & w27686;
assign w27688 = w25840 & w27687;
assign w27689 = w20878 & w27688;
assign w27690 = w27684 & w27689;
assign w27691 = ~w27606 & w27690;
assign w27692 = w27606 & ~w27690;
assign v8802 = ~(w27691 | w27692);
assign w27693 = v8802;
assign w27694 = w27675 & ~w27693;
assign w27695 = ~w27675 & w27693;
assign v8803 = ~(w27694 | w27695);
assign w27696 = v8803;
assign w27697 = w928 & w22936;
assign w27698 = w3406 & w19853;
assign w27699 = w3402 & w19917;
assign w27700 = w3399 & ~w19923;
assign v8804 = ~(w27699 | w27700);
assign w27701 = v8804;
assign w27702 = ~w27698 & w27701;
assign w27703 = ~w27697 & w27702;
assign w27704 = ~w27696 & w27703;
assign w27705 = w27696 & ~w27703;
assign v8805 = ~(w27704 | w27705);
assign w27706 = v8805;
assign w27707 = w27674 & ~w27706;
assign w27708 = ~w27674 & w27706;
assign v8806 = ~(w27707 | w27708);
assign w27709 = v8806;
assign w27710 = w3529 & w23614;
assign w27711 = w3763 & w20197;
assign w27712 = w3760 & w23607;
assign v8807 = ~(w27711 | w27712);
assign w27713 = v8807;
assign w27714 = w3767 & ~w19912;
assign w27715 = w27713 & ~w27714;
assign w27716 = ~w27710 & w27715;
assign w27717 = pi29 & w27716;
assign v8808 = ~(pi29 | w27716);
assign w27718 = v8808;
assign v8809 = ~(w27717 | w27718);
assign w27719 = v8809;
assign w27720 = ~w27709 & w27719;
assign w27721 = w27709 & ~w27719;
assign v8810 = ~(w27720 | w27721);
assign w27722 = v8810;
assign w27723 = w4153 & w24282;
assign w27724 = ~w2873 & w23670;
assign w27725 = w4155 & w24284;
assign w27726 = w4158 & ~w24077;
assign v8811 = ~(w27725 | w27726);
assign w27727 = v8811;
assign w27728 = ~w27724 & w27727;
assign w27729 = ~w27723 & w27728;
assign w27730 = pi26 & ~w27729;
assign w27731 = ~pi26 & w27729;
assign v8812 = ~(w27730 | w27731);
assign w27732 = v8812;
assign w27733 = w27722 & w27732;
assign v8813 = ~(w27722 | w27732);
assign w27734 = v8813;
assign v8814 = ~(w27733 | w27734);
assign w27735 = v8814;
assign v8815 = ~(w27636 | w27649);
assign w27736 = v8815;
assign w27737 = ~pi23 & w27736;
assign w27738 = pi23 & ~w27736;
assign v8816 = ~(w27737 | w27738);
assign w27739 = v8816;
assign v8817 = ~(w27735 | w27739);
assign w27740 = v8817;
assign w27741 = w27735 & w27739;
assign v8818 = ~(w27740 | w27741);
assign w27742 = v8818;
assign v8819 = ~(w27654 | w27660);
assign w27743 = v8819;
assign w27744 = ~w27742 & w27743;
assign w27745 = w27742 & ~w27743;
assign v8820 = ~(w27744 | w27745);
assign w27746 = v8820;
assign v8821 = ~(w27579 | w27664);
assign w27747 = v8821;
assign w27748 = (w26844 & w28905) | (w26844 & w28906) | (w28905 & w28906);
assign w27749 = (~w26844 & w28907) | (~w26844 & w28908) | (w28907 & w28908);
assign v8822 = ~(w27748 | w27749);
assign w27750 = v8822;
assign w27751 = w26972 & w31315;
assign w27752 = (~w27750 & ~w26972) | (~w27750 & w31316) | (~w26972 & w31316);
assign v8823 = ~(w27751 | w27752);
assign w27753 = v8823;
assign v8824 = ~(w27738 | w27741);
assign w27754 = v8824;
assign w27755 = w561 & w1358;
assign w27756 = w1946 & w27755;
assign w27757 = ~w425 & w5170;
assign w27758 = w27756 & w27757;
assign w27759 = w3959 & w27758;
assign w27760 = w1228 & w4004;
assign w27761 = w5005 & w27760;
assign w27762 = w4069 & w27761;
assign w27763 = ~w418 & w27762;
assign w27764 = w27759 & w27763;
assign w27765 = w12194 & w27764;
assign v8825 = ~(w27690 | w27765);
assign w27766 = v8825;
assign w27767 = w27690 & w27765;
assign v8826 = ~(w27766 | w27767);
assign w27768 = v8826;
assign w27769 = ~pi23 & w27768;
assign w27770 = pi23 & ~w27768;
assign v8827 = ~(w27769 | w27770);
assign w27771 = v8827;
assign v8828 = ~(w27691 | w27695);
assign w27772 = v8828;
assign w27773 = ~w27771 & w27772;
assign w27774 = w27771 & ~w27772;
assign v8829 = ~(w27773 | w27774);
assign w27775 = v8829;
assign w27776 = w928 & w22917;
assign w27777 = w3406 & ~w19912;
assign w27778 = w3402 & w19853;
assign w27779 = w3399 & w19917;
assign v8830 = ~(w27778 | w27779);
assign w27780 = v8830;
assign w27781 = ~w27777 & w27780;
assign w27782 = ~w27776 & w27781;
assign w27783 = w27775 & ~w27782;
assign w27784 = ~w27775 & w27782;
assign v8831 = ~(w27783 | w27784);
assign w27785 = v8831;
assign v8832 = ~(w27705 | w27708);
assign w27786 = v8832;
assign w27787 = ~w27785 & w27786;
assign w27788 = w27785 & ~w27786;
assign v8833 = ~(w27787 | w27788);
assign w27789 = v8833;
assign w27790 = w3529 & w23666;
assign w27791 = w3767 & w20197;
assign w27792 = w3760 & w23670;
assign v8834 = ~(w27791 | w27792);
assign w27793 = v8834;
assign w27794 = w3763 & w23607;
assign w27795 = w27793 & ~w27794;
assign w27796 = ~w27790 & w27795;
assign w27797 = pi29 & w27796;
assign v8835 = ~(pi29 | w27796);
assign w27798 = v8835;
assign v8836 = ~(w27797 | w27798);
assign w27799 = v8836;
assign w27800 = w27789 & ~w27799;
assign w27801 = ~w27789 & w27799;
assign v8837 = ~(w27800 | w27801);
assign w27802 = v8837;
assign v8838 = ~(w27721 | w27733);
assign w27803 = v8838;
assign w27804 = w4153 & ~w24304;
assign w27805 = w4158 & w24284;
assign v8839 = ~(w2873 | w24077);
assign w27806 = v8839;
assign v8840 = ~(w27805 | w27806);
assign w27807 = v8840;
assign w27808 = ~w27804 & w27807;
assign w27809 = ~pi26 & w27808;
assign w27810 = pi26 & ~w27808;
assign v8841 = ~(w27809 | w27810);
assign w27811 = v8841;
assign w27812 = ~w27803 & w27811;
assign w27813 = w27803 & ~w27811;
assign v8842 = ~(w27812 | w27813);
assign w27814 = v8842;
assign w27815 = w27802 & w27814;
assign v8843 = ~(w27802 | w27814);
assign w27816 = v8843;
assign v8844 = ~(w27815 | w27816);
assign w27817 = v8844;
assign w27818 = ~w27754 & w27817;
assign w27819 = w27754 & ~w27817;
assign v8845 = ~(w27818 | w27819);
assign w27820 = v8845;
assign w27821 = (~w26844 & w28443) | (~w26844 & w28444) | (w28443 & w28444);
assign w27822 = (~w26844 & w28909) | (~w26844 & w28910) | (w28909 & w28910);
assign w27823 = (w26844 & w28911) | (w26844 & w28912) | (w28911 & w28912);
assign v8846 = ~(w27822 | w27823);
assign w27824 = v8846;
assign w27825 = (~w26972 & w31317) | (~w26972 & w31318) | (w31317 & w31318);
assign w27826 = w26972 & w31319;
assign v8847 = ~(w27825 | w27826);
assign w27827 = v8847;
assign v8848 = ~(w27788 | w27800);
assign w27828 = v8848;
assign v8849 = ~(w27766 | w27769);
assign w27829 = v8849;
assign w27830 = w1475 & w2076;
assign w27831 = w13716 & w27830;
assign w27832 = w6581 & w27831;
assign w27833 = w304 & w3723;
assign w27834 = w27832 & w27833;
assign w27835 = w4117 & w27834;
assign v8850 = ~(w300 | w533);
assign w27836 = v8850;
assign w27837 = w6564 & w27836;
assign w27838 = w489 & w2444;
assign w27839 = w990 & w27838;
assign w27840 = w27837 & w27839;
assign w27841 = w3955 & w27840;
assign w27842 = w14453 & w27841;
assign w27843 = w27835 & w27842;
assign w27844 = w20149 & w27843;
assign w27845 = ~w27829 & w27844;
assign w27846 = w27829 & ~w27844;
assign v8851 = ~(w27845 | w27846);
assign w27847 = v8851;
assign w27848 = w928 & w20203;
assign w27849 = w3406 & w20197;
assign w27850 = w3402 & ~w19912;
assign w27851 = w3399 & w19853;
assign v8852 = ~(w27850 | w27851);
assign w27852 = v8852;
assign w27853 = ~w27849 & w27852;
assign w27854 = ~w27848 & w27853;
assign w27855 = ~w27847 & w27854;
assign w27856 = w27847 & ~w27854;
assign v8853 = ~(w27855 | w27856);
assign w27857 = v8853;
assign v8854 = ~(w27774 | w27783);
assign w27858 = v8854;
assign w27859 = ~w27857 & w27858;
assign w27860 = w27857 & ~w27858;
assign v8855 = ~(w27859 | w27860);
assign w27861 = v8855;
assign w27862 = w3529 & w24073;
assign w27863 = w3763 & w23670;
assign w27864 = w3760 & ~w24077;
assign v8856 = ~(w27863 | w27864);
assign w27865 = v8856;
assign w27866 = w3767 & w23607;
assign w27867 = w27865 & ~w27866;
assign w27868 = ~w27862 & w27867;
assign w27869 = pi29 & w27868;
assign v8857 = ~(pi29 | w27868);
assign w27870 = v8857;
assign v8858 = ~(w27869 | w27870);
assign w27871 = v8858;
assign w27872 = w27861 & ~w27871;
assign w27873 = ~w27861 & w27871;
assign v8859 = ~(w27872 | w27873);
assign w27874 = v8859;
assign w27875 = ~w27828 & w27874;
assign w27876 = w27828 & ~w27874;
assign v8860 = ~(w27875 | w27876);
assign w27877 = v8860;
assign w27878 = ~w2873 & w24284;
assign w27879 = pi26 & ~w27878;
assign w27880 = ~pi26 & w27878;
assign v8861 = ~(w27879 | w27880);
assign w27881 = v8861;
assign w27882 = w27877 & ~w27881;
assign w27883 = ~w27877 & w27881;
assign v8862 = ~(w27882 | w27883);
assign w27884 = v8862;
assign v8863 = ~(w27812 | w27815);
assign w27885 = v8863;
assign w27886 = w27884 & ~w27885;
assign w27887 = ~w27884 & w27885;
assign v8864 = ~(w27886 | w27887);
assign w27888 = v8864;
assign w27889 = (w26844 & w29207) | (w26844 & w29208) | (w29207 & w29208);
assign w27890 = (~w26844 & w29209) | (~w26844 & w29210) | (w29209 & w29210);
assign v8865 = ~(w27889 | w27890);
assign w27891 = v8865;
assign w27892 = w26972 & w31320;
assign w27893 = (~w26972 & w31321) | (~w26972 & w31322) | (w31321 & w31322);
assign v8866 = ~(w27892 | w27893);
assign w27894 = v8866;
assign v8867 = ~(w27875 | w27882);
assign w27895 = v8867;
assign v8868 = ~(w27860 | w27872);
assign w27896 = v8868;
assign v8869 = ~(w27845 | w27856);
assign w27897 = v8869;
assign w27898 = w2895 & w3970;
assign w27899 = w4014 & w4058;
assign w27900 = w27898 & w27899;
assign w27901 = w4049 & w12368;
assign w27902 = w27900 & w27901;
assign w27903 = ~w27843 & w27902;
assign w27904 = w27844 & ~w27902;
assign v8870 = ~(w27903 | w27904);
assign w27905 = v8870;
assign w27906 = ~w27897 & w27905;
assign w27907 = w27897 & ~w27905;
assign v8871 = ~(w27906 | w27907);
assign w27908 = v8871;
assign w27909 = w928 & w23614;
assign w27910 = w3406 & w23607;
assign w27911 = w3399 & ~w19912;
assign w27912 = w3402 & w20197;
assign v8872 = ~(w27911 | w27912);
assign w27913 = v8872;
assign w27914 = ~w27910 & w27913;
assign w27915 = ~w27909 & w27914;
assign w27916 = ~w27908 & w27915;
assign w27917 = w27908 & ~w27915;
assign v8873 = ~(w27916 | w27917);
assign w27918 = v8873;
assign w27919 = w27896 & ~w27918;
assign w27920 = ~w27896 & w27918;
assign v8874 = ~(w27919 | w27920);
assign w27921 = v8874;
assign w27922 = w3529 & w24282;
assign w27923 = w3763 & ~w24077;
assign w27924 = w3760 & w24284;
assign w27925 = w3767 & w23670;
assign v8875 = ~(w27924 | w27925);
assign w27926 = v8875;
assign w27927 = ~w27923 & w27926;
assign w27928 = ~w27922 & w27927;
assign w27929 = pi29 & ~w27928;
assign w27930 = ~pi29 & w27928;
assign v8876 = ~(w27929 | w27930);
assign w27931 = v8876;
assign w27932 = pi26 & w27931;
assign v8877 = ~(pi26 | w27931);
assign w27933 = v8877;
assign v8878 = ~(w27932 | w27933);
assign w27934 = v8878;
assign v8879 = ~(w27921 | w27934);
assign w27935 = v8879;
assign w27936 = w27921 & w27934;
assign v8880 = ~(w27935 | w27936);
assign w27937 = v8880;
assign w27938 = ~w27895 & w27937;
assign w27939 = w27895 & ~w27937;
assign v8881 = ~(w27938 | w27939);
assign w27940 = v8881;
assign w27941 = (~w27821 & w28913) | (~w27821 & w28914) | (w28913 & w28914);
assign w27942 = (w27821 & w28915) | (w27821 & w28916) | (w28915 & w28916);
assign v8882 = ~(w27941 | w27942);
assign w27943 = v8882;
assign w27944 = (~w26972 & w31323) | (~w26972 & w31324) | (w31323 & w31324);
assign w27945 = w26972 & w31325;
assign v8883 = ~(w27944 | w27945);
assign w27946 = v8883;
assign v8884 = ~(w27932 | w27936);
assign w27947 = v8884;
assign v8885 = ~(pi26 | pi29);
assign w27948 = v8885;
assign w27949 = pi26 & pi29;
assign v8886 = ~(w27948 | w27949);
assign w27950 = v8886;
assign w27951 = w3529 & ~w24304;
assign w27952 = w3767 & ~w24077;
assign v8887 = ~(w27951 | w27952);
assign w27953 = v8887;
assign w27954 = ~w27950 & w27953;
assign w27955 = w27950 & ~w27953;
assign v8888 = ~(w27954 | w27955);
assign w27956 = v8888;
assign v8889 = ~(w27904 | w27906);
assign w27957 = v8889;
assign w27958 = w4079 & w4187;
assign v8890 = ~(w27957 | w27958);
assign w27959 = v8890;
assign w27960 = w27957 & w27958;
assign v8891 = ~(w27959 | w27960);
assign w27961 = v8891;
assign w27962 = w928 & w23666;
assign w27963 = w3402 & w23607;
assign w27964 = w3406 & w23670;
assign v8892 = ~(w27963 | w27964);
assign w27965 = v8892;
assign w27966 = w3399 & w20197;
assign w27967 = w27965 & ~w27966;
assign w27968 = ~w27962 & w27967;
assign w27969 = w27844 & w27968;
assign v8893 = ~(w27844 | w27968);
assign w27970 = v8893;
assign v8894 = ~(w27969 | w27970);
assign w27971 = v8894;
assign w27972 = ~w27961 & w27971;
assign w27973 = w27961 & ~w27971;
assign v8895 = ~(w27972 | w27973);
assign w27974 = v8895;
assign v8896 = ~(w27956 | w27974);
assign w27975 = v8896;
assign w27976 = w27956 & w27974;
assign v8897 = ~(w27975 | w27976);
assign w27977 = v8897;
assign v8898 = ~(w27917 | w27920);
assign w27978 = v8898;
assign w27979 = ~w27977 & w27978;
assign w27980 = w27977 & ~w27978;
assign v8899 = ~(w27979 | w27980);
assign w27981 = v8899;
assign w27982 = w27947 & w27981;
assign v8900 = ~(w27947 | w27981);
assign w27983 = v8900;
assign v8901 = ~(w27982 | w27983);
assign w27984 = v8901;
assign w27985 = (~w27821 & w28917) | (~w27821 & w28918) | (w28917 & w28918);
assign w27986 = ~w27984 & w27985;
assign w27987 = w27984 & ~w27985;
assign v8902 = ~(w27986 | w27987);
assign w27988 = v8902;
assign w27989 = w27673 & w28261;
assign w27990 = (~w27988 & ~w27673) | (~w27988 & w28262) | (~w27673 & w28262);
assign v8903 = ~(w27989 | w27990);
assign w27991 = v8903;
assign w27992 = w1729 & w2069;
assign w27993 = w1945 & w2084;
assign v8904 = ~(w945 | w978);
assign w27994 = v8904;
assign v8905 = ~(w3337 | w3163);
assign w27995 = v8905;
assign v8906 = ~(w3127 | w3125);
assign w27996 = v8906;
assign v8907 = ~(w9402 | w10843);
assign w27997 = v8907;
assign w27998 = w10852 & pi05;
assign w27999 = w10307 & ~w10879;
assign w28000 = ~w11380 & w10848;
assign w28001 = w7308 & w1;
assign w28002 = ~w11386 & w28449;
assign v8908 = ~(w11392 | w11398);
assign w28003 = v8908;
assign w28004 = w4 & w11403;
assign w28005 = w11364 & ~w11363;
assign w28006 = w11510 & ~w11163;
assign w28007 = w11520 & ~w11085;
assign w28008 = w11523 & ~w11058;
assign w28009 = (~w28182 & w31230) | (~w28182 & w31231) | (w31230 & w31231);
assign w28010 = (~w11805 & ~w11807) | (~w11805 & w30094) | (~w11807 & w30094);
assign w28011 = w11819 & w11790;
assign w28012 = (~w11788 & ~w11774) | (~w11788 & w29439) | (~w11774 & w29439);
assign v8909 = ~(w4437 | w11667);
assign w28013 = v8909;
assign v8910 = ~(w11668 | w11667);
assign w28014 = v8910;
assign v8911 = ~(w11979 | w11667);
assign w28015 = v8911;
assign w28016 = ~w11979 & w28014;
assign v8912 = ~(w12162 | w12159);
assign w28017 = v8912;
assign w28018 = w11715 & ~w11880;
assign v8913 = ~(w11721 | w11876);
assign w28019 = v8913;
assign v8914 = ~(w11727 | w11868);
assign w28020 = v8914;
assign w28021 = w11724 & ~w11872;
assign w28022 = w11738 & ~w11857;
assign w28023 = w11730 & ~w11864;
assign v8915 = ~(w11857 | w11735);
assign w28024 = v8915;
assign v8916 = ~(w11741 | w11853);
assign w28025 = v8916;
assign v8917 = ~(w11843 | w11751);
assign w28026 = v8917;
assign w28027 = w11749 & w14284;
assign v8918 = ~(w11749 | w14284);
assign w28028 = v8918;
assign w28029 = (~w11788 & w11818) | (~w11788 & w28263) | (w11818 & w28263);
assign w28030 = ~w13193 & w9402;
assign w28031 = ~w13513 & w9402;
assign w28032 = w13309 & w9402;
assign w28033 = w13736 & w9402;
assign w28034 = ~w13863 & w9402;
assign w28035 = w13702 & w9402;
assign w28036 = ~w13881 & w9402;
assign w28037 = ~w13947 & w9402;
assign w28038 = ~w11783 & w10419;
assign w28039 = w19082 & w28264;
assign w28040 = (~pi05 & ~w19082) | (~pi05 & w28265) | (~w19082 & w28265);
assign v8919 = ~(w9402 | w19122);
assign w28041 = v8919;
assign w28042 = w19125 & ~w19122;
assign w28043 = w19125 & w28041;
assign w28044 = w19065 & ~w19064;
assign w28045 = w19059 & ~w19058;
assign v8920 = ~(w19144 | w19030);
assign w28046 = v8920;
assign w28047 = w19150 & ~w19008;
assign w28048 = w19174 & ~w18932;
assign w28049 = (w28048 & w29952) | (w28048 & w29953) | (w29952 & w29953);
assign w28050 = (w28049 & w30916) | (w28049 & w30917) | (w30916 & w30917);
assign w28051 = w18847 & ~w18846;
assign v8921 = ~(w19194 | w18831);
assign w28052 = v8921;
assign w28053 = w19197 & ~w18798;
assign w28054 = ~w19259 & w28647;
assign w28055 = w4 & ~w19582;
assign w28056 = w4 & w19613;
assign w28057 = w19616 & w19613;
assign w28058 = w19616 & w28056;
assign w28059 = w19562 & ~w19561;
assign w28060 = (w19256 & ~w20062) | (w19256 & w28450) | (~w20062 & w28450);
assign w28061 = w20062 & w28451;
assign v8922 = ~(w20061 | w20069);
assign w28062 = v8922;
assign w28063 = w20077 & ~w20015;
assign w28064 = (w29043 & w30097) | (w29043 & w30098) | (w30097 & w30098);
assign w28065 = w20118 & ~w19972;
assign v8923 = ~(w20124 | w19962);
assign w28066 = v8923;
assign v8924 = ~(w20126 | w19959);
assign w28067 = v8924;
assign w28068 = w20145 & ~w19913;
assign w28069 = w12535 & ~w19907;
assign w28070 = (~w28062 & w30732) | (~w28062 & w30733) | (w30732 & w30733);
assign w28071 = w22596 & w28145;
assign w28072 = w4 & w22939;
assign w28073 = pi02 & ~w23025;
assign v8925 = ~(w23048 | w23044);
assign w28074 = v8925;
assign v8926 = ~(w11035 | w23058);
assign w28075 = v8926;
assign w28076 = w4 & w23301;
assign w28077 = w23338 & ~w23068;
assign v8927 = ~(w23053 | w23039);
assign w28078 = v8927;
assign w28079 = w23020 & ~w23032;
assign w28080 = w23384 & ~w22946;
assign w28081 = w23407 & ~w23563;
assign v8928 = ~(w20192 | w20191);
assign w28082 = v8928;
assign w28083 = w4 & w23617;
assign v8929 = ~(w23610 | w23608);
assign w28084 = v8929;
assign v8930 = ~(w23623 | w22913);
assign w28085 = v8930;
assign v8931 = ~(w23853 | w23851);
assign w28086 = v8931;
assign w28087 = (~w23680 & ~w23693) | (~w23680 & w28266) | (~w23693 & w28266);
assign w28088 = w23663 & ~w24051;
assign w28089 = w23865 & ~w23864;
assign w28090 = w24039 & ~w24038;
assign w28091 = ~w24324 & w28267;
assign w28092 = w24295 & ~w24294;
assign w28093 = w24697 & ~w24899;
assign w28094 = ~w24900 & w24899;
assign v8932 = ~(w24900 | w28093);
assign w28095 = v8932;
assign w28096 = w25088 & ~w25089;
assign w28097 = w25275 & ~w25276;
assign v8933 = ~(w25454 | w25453);
assign w28098 = v8933;
assign v8934 = ~(w25629 | w25627);
assign w28099 = v8934;
assign w28100 = w25807 & ~w25808;
assign w28101 = ~w25984 & w25808;
assign v8935 = ~(w25984 | w28100);
assign w28102 = v8935;
assign w28103 = w26149 & ~w28101;
assign w28104 = w26149 & ~w28102;
assign w28105 = w26298 & ~w26146;
assign w28106 = (~w26297 & ~w26298) | (~w26297 & w28147) | (~w26298 & w28147);
assign w28107 = ~w26441 & w26297;
assign w28108 = (~w28147 & w28107) | (~w28147 & w29211) | (w28107 & w29211);
assign w28109 = w26583 & ~w26440;
assign w28110 = (~w26581 & ~w26583) | (~w26581 & w28148) | (~w26583 & w28148);
assign w28111 = ~w26716 & w26581;
assign v8936 = ~(w26715 | w28111);
assign w28112 = v8936;
assign w28113 = (w28148 & w28648) | (w28148 & w28649) | (w28648 & w28649);
assign w28114 = ~w26841 & w26966;
assign w28115 = ~w28114 & w26974;
assign w28116 = (~w27080 & w26974) | (~w27080 & w28149) | (w26974 & w28149);
assign w28117 = (~w27080 & w28115) | (~w27080 & w28149) | (w28115 & w28149);
assign w28118 = w27192 & ~w28116;
assign w28119 = (~w28115 & w28269) | (~w28115 & w28270) | (w28269 & w28270);
assign w28120 = w27084 & w27195;
assign w28121 = (~w27191 & w28116) | (~w27191 & w28650) | (w28116 & w28650);
assign w28122 = (w28115 & w29212) | (w28115 & w29213) | (w29212 & w29213);
assign w28123 = w28120 & w27301;
assign v8937 = ~(w27298 | w27296);
assign w28124 = v8937;
assign w28125 = w28123 & ~w27398;
assign v8938 = ~(w27393 | w27296);
assign w28126 = v8938;
assign w28127 = ~w27298 & w28126;
assign v8939 = ~(w27394 | w28126);
assign w28128 = v8939;
assign v8940 = ~(w27394 | w28127);
assign w28129 = v8940;
assign w28130 = w28123 & w28150;
assign w28131 = (~w27484 & w28126) | (~w27484 & w28651) | (w28126 & w28651);
assign w28132 = (~w27484 & w28127) | (~w27484 & w28651) | (w28127 & w28651);
assign w28133 = w28130 & w27587;
assign w28134 = w28130 & w28271;
assign v8941 = ~(w27665 | w27747);
assign w28135 = v8941;
assign w28136 = (~w27665 & w27582) | (~w27665 & w28135) | (w27582 & w28135);
assign w28137 = w27750 & w27824;
assign v8942 = ~(w27820 | w27818);
assign w28138 = v8942;
assign w28139 = w28137 & ~w27891;
assign v8943 = ~(w27888 | w27887);
assign w28140 = v8943;
assign w28141 = w28139 & w27943;
assign v8944 = ~(w27939 | w27887);
assign w28142 = v8944;
assign w28143 = ~w27939 & w28140;
assign w28144 = w19759 & w19341;
assign v8945 = ~(pi05 | w9402);
assign w28145 = v8945;
assign v8946 = ~(pi08 | w8141);
assign w28146 = v8946;
assign w28147 = w26146 & ~w26297;
assign w28148 = w26440 & ~w26581;
assign w28149 = w27079 & ~w27080;
assign w28150 = ~w27398 & w27489;
assign w28151 = ~w822 & w1821;
assign v8947 = ~(w888 | w98);
assign w28152 = v8947;
assign w28153 = w3043 & w3048;
assign w28154 = w1722 & w3078;
assign w28155 = ~w584 & w1263;
assign w28156 = w3122 & w3118;
assign v8948 = ~(w3070 | w3125);
assign w28157 = v8948;
assign w28158 = ~w3127 & w28157;
assign w28159 = (w8926 & ~w3227) | (w8926 & w28452) | (~w3227 & w28452);
assign w28160 = (w8526 & ~w3283) | (w8526 & w28453) | (~w3283 & w28453);
assign w28161 = ~w3284 & w8138;
assign w28162 = ~w10844 & w28454;
assign w28163 = w10846 & w27997;
assign w28164 = (w10419 & ~w3227) | (w10419 & w28455) | (~w3227 & w28455);
assign w28165 = (w9891 & ~w3283) | (w9891 & w28456) | (~w3283 & w28456);
assign w28166 = w27998 & ~w10848;
assign v8949 = ~(w27999 | w10880);
assign w28167 = v8949;
assign w28168 = w10878 & pi05;
assign v8950 = ~(w10878 | pi05);
assign w28169 = v8950;
assign w28170 = w10607 & ~w10606;
assign v8951 = ~(w10964 | w10591);
assign w28171 = v8951;
assign v8952 = ~(w10968 | w10560);
assign w28172 = v8952;
assign w28173 = (~w10529 & w10971) | (~w10529 & w29618) | (w10971 & w29618);
assign v8953 = ~(w10975 | w10494);
assign w28174 = v8953;
assign v8954 = ~(w10978 | w10463);
assign w28175 = v8954;
assign v8955 = ~(w4082 | w10989);
assign w28176 = v8955;
assign w28177 = w4 & ~w11024;
assign w28178 = w4 & w11037;
assign w28179 = w4 & w11357;
assign w28180 = w4 & w11371;
assign w28181 = (w11029 & ~w11032) | (w11029 & w31232) | (~w11032 & w31232);
assign w28182 = w10429 & ~w11535;
assign w28183 = ~w11017 & w11536;
assign w28184 = w9906 & ~w10432;
assign w28185 = w9906 & w28009;
assign w28186 = ~w11778 & w11526;
assign v8956 = ~(w11820 | w11821);
assign w28187 = v8956;
assign w28188 = ~w11824 & w28012;
assign w28189 = ~w18443 & w28457;
assign v8957 = ~(w19571 | w19567);
assign w28190 = v8957;
assign w28191 = w19606 & ~pi02;
assign w28192 = ~w19606 & pi02;
assign v8958 = ~(pi02 | w19613);
assign w28193 = v8958;
assign v8959 = ~(pi02 | w28056);
assign w28194 = v8959;
assign w28195 = ~w19618 & w19623;
assign w28196 = w19523 & ~w19522;
assign w28197 = w19458 & w19471;
assign w28198 = (~w19440 & w19699) | (~w19440 & w30446) | (w19699 & w30446);
assign w28199 = ~w19760 & w29954;
assign w28200 = (~w19335 & w19322) | (~w19335 & w28652) | (w19322 & w28652);
assign v8960 = ~(w19280 | w19267);
assign w28201 = v8960;
assign w28202 = w19786 & ~w19242;
assign v8961 = ~(w20025 | w20024);
assign w28203 = v8961;
assign w28204 = ~w19788 & w29955;
assign w28205 = (~w20034 & ~w19269) | (~w20034 & w20038) | (~w19269 & w20038);
assign w28206 = ~w19269 & w19781;
assign w28207 = w20073 & ~w20029;
assign w28208 = ~w22570 & w28653;
assign w28209 = ~w22581 & w28654;
assign w28210 = ~w22597 & w22591;
assign w28211 = w22597 & ~w22591;
assign v8962 = ~(w22654 | w22576);
assign w28212 = v8962;
assign w28213 = w22656 & ~w22566;
assign w28214 = w22668 & ~w22535;
assign w28215 = w22684 & ~w22491;
assign w28216 = w22704 & ~w22427;
assign w28217 = (~w21379 & ~w21845) | (~w21379 & w30099) | (~w21845 & w30099);
assign w28218 = ~w8141 & w22879;
assign w28219 = w4 & w22920;
assign w28220 = w28082 & ~w20191;
assign w28221 = (~w20191 & w28082) | (~w20191 & ~w19908) | (w28082 & ~w19908);
assign v8963 = ~(w20198 | w23610);
assign w28222 = v8963;
assign w28223 = w20198 & w23610;
assign w28224 = ~w23663 & w23608;
assign w28225 = (~w23663 & w23610) | (~w23663 & w28224) | (w23610 & w28224);
assign w28226 = w23663 & ~w23608;
assign w28227 = ~w23610 & w28226;
assign w28228 = w23846 & w28146;
assign v8964 = ~(w28085 | w23624);
assign w28229 = v8964;
assign w28230 = ~w8141 & w24034;
assign w28231 = w24070 & w24051;
assign w28232 = w24070 & ~w28088;
assign v8965 = ~(w24070 | w24051);
assign w28233 = v8965;
assign w28234 = ~w24070 & w28088;
assign w28235 = w24104 & w28146;
assign v8966 = ~(w24328 | w28091);
assign w28236 = v8966;
assign v8967 = ~(w24328 | w24329);
assign w28237 = v8967;
assign w28238 = ~w25398 & w28655;
assign w28239 = ~w25933 & w28656;
assign v8968 = ~(pi17 | w25937);
assign w28240 = v8968;
assign v8969 = ~(pi17 | w28239);
assign w28241 = v8969;
assign w28242 = ~w25939 & w25932;
assign w28243 = w25939 & ~w25932;
assign v8970 = ~(w25978 | w25818);
assign w28244 = v8970;
assign w28245 = w26153 & ~w26300;
assign w28246 = (w28112 & w28113) | (w28112 & w28107) | (w28113 & w28107);
assign w28247 = (w28112 & w28113) | (w28112 & w28108) | (w28113 & w28108);
assign w28248 = ~w26720 & w26847;
assign v8971 = ~(w26832 | w26835);
assign w28249 = v8971;
assign v8972 = ~(w26829 | w26818);
assign w28250 = v8972;
assign w28251 = w26965 & ~w26964;
assign w28252 = (w28131 & w28132) | (w28131 & w28122) | (w28132 & w28122);
assign w28253 = (w28131 & w28132) | (w28131 & w28121) | (w28132 & w28121);
assign v8973 = ~(w27485 | w27484);
assign w28254 = v8973;
assign w28255 = (~w27584 & ~w28130) | (~w27584 & w28274) | (~w28130 & w28274);
assign w28256 = ~w27744 & w28135;
assign w28257 = ~w27744 & w28136;
assign v8974 = ~(w27750 | w27824);
assign w28258 = v8974;
assign w28259 = ~w28137 & w27891;
assign v8975 = ~(w28139 | w27943);
assign w28260 = v8975;
assign w28261 = w28141 & w27988;
assign v8976 = ~(w28141 | w27988);
assign w28262 = v8976;
assign w28263 = w11814 & ~w11788;
assign w28264 = ~w19083 & pi05;
assign w28265 = w19083 & ~pi05;
assign v8977 = ~(w23857 | w23680);
assign w28266 = v8977;
assign w28267 = w24327 & w28146;
assign w28268 = w26716 & ~w26715;
assign w28269 = w27192 & w27080;
assign w28270 = w27192 & ~w28149;
assign w28271 = ~w27586 & w28458;
assign v8978 = ~(w22572 | w9402);
assign w28272 = v8978;
assign w28273 = ~w22640 & w28657;
assign w28274 = w27586 & ~w27584;
assign v8979 = ~(w3069 | w28157);
assign w28275 = v8979;
assign v8980 = ~(w3069 | w28158);
assign w28276 = v8980;
assign w28277 = w10294 & w28658;
assign w28278 = (~w8141 & w3332) | (~w8141 & w28459) | (w3332 & w28459);
assign w28279 = w10303 & ~w10300;
assign w28280 = w10303 & w28278;
assign w28281 = ~w8141 & w10307;
assign w28282 = w10325 & ~w10299;
assign w28283 = w10329 & ~w10288;
assign w28284 = (~w10395 & w10392) | (~w10395 & w29440) | (w10392 & w29440);
assign w28285 = ~w9402 & w10823;
assign v8981 = ~(w10447 | w10835);
assign w28286 = v8981;
assign w28287 = ~w3284 & w9401;
assign w28288 = ~w3228 & w9891;
assign w28289 = ~w9402 & w10852;
assign w28290 = ~w3228 & w9401;
assign w28291 = ~w10861 & pi05;
assign w28292 = w10861 & ~pi05;
assign w28293 = ~w9402 & w10876;
assign v8982 = ~(w10893 | w10842);
assign w28294 = v8982;
assign w28295 = w4191 & ~pi02;
assign w28296 = w28176 & ~w10989;
assign w28297 = (~w10989 & w28176) | (~w10989 & ~w4083) | (w28176 & ~w4083);
assign w28298 = ~w9402 & w10998;
assign v8983 = ~(pi02 | w11357);
assign w28299 = v8983;
assign v8984 = ~(pi02 | w28179);
assign w28300 = v8984;
assign w28301 = w11360 & w11357;
assign w28302 = w11360 & w28179;
assign w28303 = pi02 & ~w11371;
assign w28304 = pi02 & ~w28180;
assign w28305 = ~w11374 & w11371;
assign w28306 = ~w11374 & w28180;
assign v8985 = ~(pi02 | w10848);
assign w28307 = v8985;
assign v8986 = ~(pi02 | w28000);
assign w28308 = v8986;
assign w28309 = ~w3228 & pi01;
assign w28310 = w11388 & ~pi02;
assign v8987 = ~(w11388 | w10988);
assign w28311 = v8987;
assign w28312 = pi02 & ~w11403;
assign w28313 = pi02 & ~w28004;
assign w28314 = ~w11406 & w11403;
assign w28315 = ~w11406 & w28004;
assign w28316 = w11411 & ~w11377;
assign w28317 = w9904 & w9420;
assign w28318 = (~w10432 & w11018) | (~w10432 & w29956) | (w11018 & w29956);
assign w28319 = ~w11801 & w11798;
assign w28320 = w11020 & w11013;
assign v8988 = ~(w11772 | w11769);
assign w28321 = v8988;
assign v8989 = ~(w11840 | w11763);
assign w28322 = v8989;
assign w28323 = ~w11877 & w30734;
assign w28324 = (~w11892 & w11891) | (~w11892 & w28461) | (w11891 & w28461);
assign w28325 = ~w11581 & w28013;
assign w28326 = ~w17869 & w28659;
assign w28327 = ~w17882 & w28660;
assign w28328 = (pi11 & ~w17895) | (pi11 & w28463) | (~w17895 & w28463);
assign w28329 = w17895 & w28464;
assign w28330 = pi08 & ~w18447;
assign w28331 = pi08 & ~w28189;
assign w28332 = ~pi08 & w18447;
assign w28333 = ~pi08 & w28189;
assign w28334 = (w9402 & ~w12992) | (w9402 & w30278) | (~w12992 & w30278);
assign w28335 = ~w19065 & w19064;
assign v8990 = ~(w19117 | w19087);
assign w28336 = v8990;
assign w28337 = w18816 & ~w18815;
assign w28338 = w18781 & ~w18780;
assign v8991 = ~(w19200 | w18763);
assign w28339 = v8991;
assign w28340 = w18734 & ~w18733;
assign w28341 = w19204 & ~w18714;
assign w28342 = w19212 & ~w18668;
assign v8992 = ~(w12382 | w4);
assign w28343 = v8992;
assign w28344 = ~w12502 & w28661;
assign v8993 = ~(pi02 | w19261);
assign w28345 = v8993;
assign v8994 = ~(pi02 | w28054);
assign w28346 = v8994;
assign w28347 = w19264 & w19261;
assign w28348 = w19264 & w28054;
assign w28349 = ~w19272 & w29958;
assign w28350 = ~w19285 & w29959;
assign w28351 = ~w19296 & w30279;
assign w28352 = w4 & w19313;
assign w28353 = w4 & w19329;
assign v8995 = ~(w11989 | w4);
assign w28354 = v8995;
assign v8996 = ~(w19532 | w19528);
assign w28355 = v8996;
assign w28356 = w4 & w19540;
assign w28357 = w19555 & ~w19557;
assign w28358 = ~w19555 & pi02;
assign w28359 = ~w11767 & w11035;
assign w28360 = w19563 & w19577;
assign w28361 = w19585 & ~w19582;
assign w28362 = w19585 & w28055;
assign v8997 = ~(w19682 | w19471);
assign w28363 = v8997;
assign v8998 = ~(w19682 | w19468);
assign w28364 = v8998;
assign w28365 = w19774 & ~w19323;
assign v8999 = ~(w19225 | w19223);
assign w28366 = v8999;
assign w28367 = w20123 & ~w19967;
assign w28368 = w22111 & w28662;
assign w28369 = w22122 & w28663;
assign w28370 = w22551 & w28664;
assign w28371 = (~pi05 & ~w22551) | (~pi05 & w28665) | (~w22551 & w28665);
assign w28372 = ~w9402 & w22562;
assign v9000 = ~(pi05 | w28208);
assign w28373 = v9000;
assign w28374 = (~pi05 & ~w22571) | (~pi05 & w28666) | (~w22571 & w28666);
assign w28375 = pi05 & w28208;
assign w28376 = w22571 & w28667;
assign w28377 = pi05 & ~w22584;
assign w28378 = pi05 & ~w28209;
assign w28379 = ~pi05 & w22584;
assign w28380 = ~pi05 & w28209;
assign w28381 = (pi05 & w22639) | (pi05 & w28668) | (w22639 & w28668);
assign w28382 = (pi05 & w22639) | (pi05 & w28669) | (w22639 & w28669);
assign w28383 = ~w22639 & w28670;
assign w28384 = ~pi05 & w22643;
assign v9001 = ~(w21854 | w21852);
assign w28385 = v9001;
assign v9002 = ~(w21840 | w21838);
assign w28386 = v9002;
assign w28387 = pi08 & ~w22879;
assign w28388 = pi08 & ~w28218;
assign w28389 = ~pi08 & w22879;
assign w28390 = ~pi08 & w28218;
assign w28391 = ~w9402 & w22903;
assign w28392 = w4 & w23246;
assign w28393 = pi02 & w23265;
assign w28394 = w4 & w23271;
assign w28395 = w22907 & ~w22908;
assign w28396 = ~w8141 & w23412;
assign v9003 = ~(w22874 | w22873);
assign w28397 = v9003;
assign w28398 = (w28221 & w28220) | (w28221 & w19907) | (w28220 & w19907);
assign w28399 = (w28221 & w28220) | (w28221 & ~w28069) | (w28220 & ~w28069);
assign v9004 = ~(pi02 | w23617);
assign w28400 = v9004;
assign v9005 = ~(pi02 | w28083);
assign w28401 = v9005;
assign w28402 = w23620 & w23617;
assign w28403 = w23620 & w28083;
assign w28404 = w4 & w23673;
assign v9006 = ~(w23847 | w28228);
assign w28405 = v9006;
assign v9007 = ~(w23847 | w23848);
assign w28406 = v9007;
assign w28407 = w23682 & ~w23857;
assign w28408 = ~w23682 & w23857;
assign w28409 = pi05 & w23878;
assign w28410 = w23878 & w28465;
assign v9008 = ~(pi05 | w23878);
assign w28411 = v9008;
assign w28412 = (~pi05 & ~w23878) | (~pi05 & w28466) | (~w23878 & w28466);
assign w28413 = ~w7178 & w23888;
assign w28414 = pi08 & ~w24034;
assign w28415 = pi08 & ~w28230;
assign w28416 = ~pi08 & w24034;
assign w28417 = ~pi08 & w28230;
assign w28418 = w4 & w24080;
assign v9009 = ~(w24046 | w24045);
assign w28419 = v9009;
assign v9010 = ~(w24105 | w28235);
assign w28420 = v9010;
assign v9011 = ~(w24105 | w24106);
assign w28421 = v9011;
assign w28422 = ~w9402 & w24270;
assign w28423 = w23670 & ~w28232;
assign w28424 = (w23670 & ~w24070) | (w23670 & w28467) | (~w24070 & w28467);
assign w28425 = ~w10447 & w24320;
assign w28426 = ~w24327 & pi08;
assign w28427 = w24327 & ~pi08;
assign w28428 = ~w7178 & w24339;
assign w28429 = w24098 & w31233;
assign w28430 = ~w8141 & w24670;
assign v9012 = ~(w24699 | w24697);
assign w28431 = v9012;
assign w28432 = w25054 & w28671;
assign w28433 = ~pi11 & w25109;
assign w28434 = w25109 & w17575;
assign w28435 = pi11 & ~w25109;
assign w28436 = (pi11 & ~w25109) | (pi11 & w28672) | (~w25109 & w28672);
assign w28437 = ~pi14 & w25402;
assign w28438 = ~pi14 & w28238;
assign w28439 = pi14 & ~w25402;
assign w28440 = pi14 & ~w28238;
assign w28441 = (~w25808 & w28100) | (~w25808 & w25627) | (w28100 & w25627);
assign w28442 = (~w25808 & w28100) | (~w25808 & ~w28099) | (w28100 & ~w28099);
assign w28443 = (w28256 & w28257) | (w28256 & ~w28253) | (w28257 & ~w28253);
assign w28444 = (w28256 & w28257) | (w28256 & ~w28252) | (w28257 & ~w28252);
assign w28445 = w27745 & w27820;
assign v9013 = ~(w27745 | w27820);
assign w28446 = v9013;
assign w28447 = w28138 & ~w27818;
assign w28448 = (~w27818 & w28138) | (~w27818 & ~w27745) | (w28138 & ~w27745);
assign w28449 = ~w11385 & w3332;
assign w28450 = ~w19785 & w19256;
assign w28451 = w19785 & ~w19256;
assign w28452 = ~w3212 & w8926;
assign w28453 = ~w869 & w8526;
assign v9014 = ~(w10845 | w10843);
assign w28454 = v9014;
assign w28455 = ~w3212 & w10419;
assign w28456 = ~w869 & w9891;
assign w28457 = w18446 & ~w8141;
assign w28458 = (~w27669 & w27583) | (~w27669 & w28919) | (w27583 & w28919);
assign v9015 = ~(w8140 | w8141);
assign w28459 = v9015;
assign w28460 = (~w8141 & w3211) | (~w8141 & w28673) | (w3211 & w28673);
assign w28461 = w11687 & ~w11892;
assign v9016 = ~(w17884 | w7178);
assign w28462 = v9016;
assign w28463 = w17892 & pi11;
assign v9017 = ~(w17892 | pi11);
assign w28464 = v9017;
assign w28465 = ~w9402 & pi05;
assign w28466 = w9402 & ~pi05;
assign w28467 = ~w24051 & w23670;
assign w28468 = ~w103 & w712;
assign w28469 = w713 & w717;
assign v9018 = ~(w731 | w609);
assign w28470 = v9018;
assign v9019 = ~(w68 | w680);
assign w28471 = v9019;
assign w28472 = w3183 & w31121;
assign v9020 = ~(w522 | w168);
assign w28473 = v9020;
assign w28474 = w3202 & w3200;
assign w28475 = w3002 & ~w3001;
assign w28476 = w6548 & ~w3125;
assign w28477 = w6548 & w27996;
assign w28478 = ~w6548 & w3125;
assign v9021 = ~(w6548 | w27996);
assign w28479 = v9021;
assign w28480 = w9772 & w28920;
assign w28481 = w9791 & ~w9787;
assign w28482 = ~w8141 & w10280;
assign w28483 = pi08 & ~w10295;
assign w28484 = pi08 & ~w28277;
assign w28485 = ~pi08 & w10295;
assign w28486 = ~pi08 & w28277;
assign w28487 = ~w3228 & w8526;
assign w28488 = ~w3193 & w8926;
assign w28489 = (~pi08 & ~w10319) | (~pi08 & w28674) | (~w10319 & w28674);
assign w28490 = (~pi08 & ~w10319) | (~pi08 & w28675) | (~w10319 & w28675);
assign w28491 = w10319 & w28676;
assign w28492 = w10319 & w28921;
assign w28493 = w10323 & ~w10314;
assign w28494 = ~w3123 & w9891;
assign v9022 = ~(w10829 | pi05);
assign w28495 = v9022;
assign w28496 = w10829 & pi05;
assign w28497 = ~w3193 & w10419;
assign v9023 = ~(w10897 | w10827);
assign w28498 = v9023;
assign w28499 = w4 & w11345;
assign v9024 = ~(w28002 | w10848);
assign w28500 = v9024;
assign w28501 = w11352 & ~w11340;
assign w28502 = w11328 & ~w11327;
assign v9025 = ~(w11224 | w11487);
assign w28503 = v9025;
assign w28504 = (~w4 & ~w3390) | (~w4 & w29214) | (~w3390 & w29214);
assign v9026 = ~(w9418 | w9420);
assign w28505 = v9026;
assign w28506 = (~w9418 & ~w9420) | (~w9418 & w29441) | (~w9420 & w29441);
assign v9027 = ~(w9904 | w9420);
assign w28507 = v9027;
assign w28508 = (pi11 & w17869) | (pi11 & w28922) | (w17869 & w28922);
assign w28509 = (pi11 & w17869) | (pi11 & w28923) | (w17869 & w28923);
assign w28510 = ~w17869 & w28924;
assign w28511 = ~pi11 & w28326;
assign v9028 = ~(pi11 | w28327);
assign w28512 = v9028;
assign w28513 = (~pi11 & ~w17883) | (~pi11 & w28677) | (~w17883 & w28677);
assign w28514 = pi11 & w28327;
assign w28515 = w17883 & w28678;
assign v9029 = ~(w7178 | w17909);
assign w28516 = v9029;
assign w28517 = (pi11 & ~w17924) | (pi11 & w28679) | (~w17924 & w28679);
assign w28518 = w17924 & w28680;
assign w28519 = w17929 & ~w17899;
assign w28520 = w11770 & w8926;
assign w28521 = w18435 & w28682;
assign w28522 = (~pi08 & ~w18435) | (~pi08 & w28683) | (~w18435 & w28683);
assign w28523 = ~w18476 & pi08;
assign w28524 = w18475 & w28684;
assign w28525 = ~w18490 & w18485;
assign w28526 = w18490 & ~w18485;
assign w28527 = w18505 & w28685;
assign w28528 = w18512 & ~w18451;
assign v9030 = ~(w18530 | w18407);
assign w28529 = v9030;
assign w28530 = w18540 & ~w18371;
assign v9031 = ~(w18557 | w18301);
assign w28531 = v9031;
assign v9032 = ~(w18560 | w18270);
assign w28532 = v9032;
assign v9033 = ~(w18563 | w18239);
assign w28533 = v9033;
assign v9034 = ~(w18570 | w18173);
assign w28534 = v9034;
assign w28535 = ~w12502 & w28686;
assign w28536 = w11770 & w10419;
assign w28537 = ~w19054 & pi05;
assign w28538 = w19054 & ~pi05;
assign w28539 = pi08 & w17900;
assign v9035 = ~(pi02 | w19540);
assign w28540 = v9035;
assign v9036 = ~(pi02 | w28356);
assign w28541 = v9036;
assign w28542 = w19543 & w19540;
assign w28543 = w19543 & w28356;
assign w28544 = w11770 & w11035;
assign v9037 = ~(w19563 | w19577);
assign w28545 = v9037;
assign w28546 = ~w11526 & w11035;
assign w28547 = w19588 & ~w28362;
assign w28548 = w19588 & ~w28361;
assign v9038 = ~(w19590 | w11800);
assign w28549 = v9038;
assign v9039 = ~(w19589 | w19581);
assign w28550 = v9039;
assign v9040 = ~(w19605 | w19603);
assign w28551 = v9040;
assign w28552 = w19549 & ~w19548;
assign w28553 = w19505 & ~w19522;
assign w28554 = w19505 & w19631;
assign w28555 = w4 & w19638;
assign w28556 = w19472 & ~w19457;
assign w28557 = w19385 & ~w19384;
assign w28558 = ~w19743 & w29960;
assign v9041 = ~(pi02 | w19762);
assign w28559 = v9041;
assign v9042 = ~(pi02 | w28199);
assign w28560 = v9042;
assign w28561 = w19765 & w19762;
assign w28562 = w19765 & w28199;
assign v9043 = ~(w19799 | w18628);
assign w28563 = v9043;
assign v9044 = ~(w20012 | w20081);
assign w28564 = v9044;
assign w28565 = ~w21596 & w29961;
assign w28566 = ~w22142 & w30918;
assign v9045 = ~(w22630 | w22602);
assign w28567 = v9045;
assign v9046 = ~(w11035 | w23298);
assign w28568 = v9046;
assign w28569 = pi02 & w23301;
assign w28570 = pi02 & w28076;
assign v9047 = ~(w3 | w23303);
assign w28571 = v9047;
assign w28572 = w23190 & ~w23189;
assign w28573 = w22888 & ~w23407;
assign w28574 = (~w21838 & ~w22855) | (~w21838 & w30100) | (~w22855 & w30100);
assign w28575 = ~w22866 & w28386;
assign w28576 = ~w23562 & w28081;
assign w28577 = w28398 | w28399;
assign w28578 = (w28399 & w28398) | (w28399 & ~w12537) | (w28398 & ~w12537);
assign w28579 = w23557 & ~w23556;
assign w28580 = ~w23562 & w23563;
assign v9048 = ~(w23562 | w28081);
assign w28581 = v9048;
assign w28582 = (w28232 & w28231) | (w28232 & w23608) | (w28231 & w23608);
assign w28583 = (w28232 & w28231) | (w28232 & ~w28084) | (w28231 & ~w28084);
assign w28584 = (w28234 & w28233) | (w28234 & ~w23608) | (w28233 & ~w23608);
assign w28585 = (w28234 & w28233) | (w28234 & w28084) | (w28233 & w28084);
assign w28586 = pi05 & w24270;
assign w28587 = pi05 & w28422;
assign v9049 = ~(pi05 | w24270);
assign w28588 = v9049;
assign v9050 = ~(pi05 | w28422);
assign w28589 = v9050;
assign w28590 = ~w23670 & w28224;
assign w28591 = ~w23670 & w28225;
assign w28592 = ~w7178 & w24525;
assign w28593 = pi08 & w24670;
assign w28594 = pi08 & w28430;
assign v9051 = ~(pi08 | w24670);
assign w28595 = v9051;
assign v9052 = ~(pi08 | w28430);
assign w28596 = v9052;
assign v9053 = ~(w24493 | w24490);
assign w28597 = v9053;
assign w28598 = ~w24280 & w8141;
assign w28599 = ~w25454 & w25276;
assign v9054 = ~(w25454 | w28097);
assign w28600 = v9054;
assign w28601 = w25454 & ~w25276;
assign w28602 = w25454 & w28097;
assign w28603 = w25629 & ~w25453;
assign w28604 = w25629 & w28098;
assign w28605 = ~w25629 & w25453;
assign v9055 = ~(w25629 | w28098);
assign w28606 = v9055;
assign w28607 = (~w25627 & ~w25629) | (~w25627 & w28687) | (~w25629 & w28687);
assign w28608 = (~w25627 & w28099) | (~w25627 & ~w28098) | (w28099 & ~w28098);
assign w28609 = w25985 & w28442;
assign w28610 = w25985 & w28441;
assign w28611 = w28245 & w26446;
assign v9056 = ~(w26431 | w26434);
assign w28612 = v9056;
assign v9057 = ~(w26387 | w26386);
assign w28613 = v9057;
assign w28614 = ~w26537 & w28925;
assign v9058 = ~(w26428 | w26417);
assign w28615 = v9058;
assign v9059 = ~(w26442 | w26583);
assign w28616 = v9059;
assign w28617 = ~w26790 & w28926;
assign w28618 = w26807 & w28927;
assign w28619 = ~w26920 & w28928;
assign w28620 = w28248 & w26970;
assign w28621 = ~w27081 & w26974;
assign w28622 = ~w27081 & w28115;
assign w28623 = w27081 & ~w26974;
assign w28624 = w27081 & ~w28115;
assign w28625 = w27141 & w28929;
assign w28626 = ~w4764 & w27158;
assign w28627 = ~w27192 & w28116;
assign w28628 = ~w27192 & w28117;
assign w28629 = ~w4153 & w27206;
assign w28630 = (~w27296 & w28124) | (~w27296 & w28122) | (w28124 & w28122);
assign w28631 = (~w27296 & w28124) | (~w27296 & w28121) | (w28124 & w28121);
assign w28632 = ~w3529 & w27343;
assign w28633 = ~w4153 & w27452;
assign w28634 = (w28128 & w28129) | (w28128 & ~w28122) | (w28129 & ~w28122);
assign w28635 = (w28128 & w28129) | (w28128 & ~w28121) | (w28129 & ~w28121);
assign w28636 = (~w28122 & w28688) | (~w28122 & w28689) | (w28688 & w28689);
assign w28637 = w27888 & w28448;
assign w28638 = w27888 & w28447;
assign v9060 = ~(w27888 | w28448);
assign w28639 = v9060;
assign v9061 = ~(w27888 | w28447);
assign w28640 = v9061;
assign w28641 = (~w27887 & w28140) | (~w27887 & ~w28448) | (w28140 & ~w28448);
assign w28642 = (~w27887 & w28140) | (~w27887 & ~w28447) | (w28140 & ~w28447);
assign w28643 = (w28142 & w28143) | (w28142 & ~w28448) | (w28143 & ~w28448);
assign w28644 = (w28142 & w28143) | (w28142 & ~w28447) | (w28143 & ~w28447);
assign v9062 = ~(w19019 | w19030);
assign w28645 = v9062;
assign v9063 = ~(w19019 | w19032);
assign w28646 = v9063;
assign w28647 = ~w19260 & w4;
assign w28648 = (~w26715 & w28268) | (~w26715 & ~w26581) | (w28268 & ~w26581);
assign w28649 = (~w26715 & w28268) | (~w26715 & ~w26583) | (w28268 & ~w26583);
assign v9064 = ~(w27192 | w27191);
assign w28650 = v9064;
assign w28651 = w27394 & ~w27484;
assign w28652 = w19318 & ~w19335;
assign w28653 = ~w22569 & w28272;
assign w28654 = w22583 & ~w9402;
assign w28655 = w25401 & ~w6389;
assign w28656 = w25936 & ~w5765;
assign v9065 = ~(w22641 | w9402);
assign w28657 = v9065;
assign v9066 = ~(w10291 | w8141);
assign w28658 = v9066;
assign w28659 = w17872 & ~w7178;
assign w28660 = ~w17881 & w28462;
assign w28661 = ~w12406 & w29962;
assign v9067 = ~(w22112 | w8141);
assign w28662 = v9067;
assign v9068 = ~(w22123 | w8141);
assign w28663 = v9068;
assign w28664 = ~w22552 & pi05;
assign w28665 = w22552 & ~pi05;
assign w28666 = w22572 & ~pi05;
assign w28667 = ~w22572 & pi05;
assign w28668 = ~w28273 & pi05;
assign w28669 = ~w22642 & pi05;
assign w28670 = w28273 & ~pi05;
assign v9069 = ~(w25055 | w7178);
assign w28671 = v9069;
assign w28672 = w7178 & pi11;
assign v9070 = ~(w8526 | w8141);
assign w28673 = v9070;
assign v9071 = ~(w28460 | pi08);
assign w28674 = v9071;
assign w28675 = w10320 & ~pi08;
assign w28676 = w28460 & pi08;
assign w28677 = w17884 & ~pi11;
assign w28678 = ~w17884 & pi11;
assign w28679 = w17921 & pi11;
assign v9072 = ~(w17921 | pi11);
assign w28680 = v9072;
assign w28681 = (~w8141 & w11771) | (~w8141 & w28673) | (w11771 & w28673);
assign w28682 = ~w18436 & pi08;
assign w28683 = w18436 & ~pi08;
assign v9073 = ~(w18472 | pi08);
assign w28684 = v9073;
assign v9074 = ~(w18502 | w8141);
assign w28685 = v9074;
assign w28686 = ~w12406 & w29963;
assign w28687 = ~w25627 & w25453;
assign w28688 = (w28135 & w28136) | (w28135 & ~w28131) | (w28136 & ~w28131);
assign w28689 = (w28135 & w28136) | (w28135 & ~w28132) | (w28136 & ~w28132);
assign w28690 = w2940 & ~w3001;
assign w28691 = w2940 & w28475;
assign w28692 = w9251 & w29215;
assign w28693 = (~w6389 & w3262) | (~w6389 & w29216) | (w3262 & w29216);
assign w28694 = w9267 & ~w9263;
assign w28695 = ~w7178 & w9759;
assign v9075 = ~(pi11 | w9774);
assign w28696 = v9075;
assign v9076 = ~(pi11 | w28480);
assign w28697 = v9076;
assign w28698 = pi11 & w9774;
assign w28699 = pi11 & w28480;
assign w28700 = (w7172 & ~w3283) | (w7172 & w28930) | (~w3283 & w28930);
assign w28701 = (w7466 & ~w3283) | (w7466 & w28931) | (~w3283 & w28931);
assign w28702 = (w7765 & ~w3227) | (w7765 & w28932) | (~w3227 & w28932);
assign w28703 = w9791 & w29217;
assign w28704 = ~w9788 & w29218;
assign w28705 = (~w9262 & w9788) | (~w9262 & w29219) | (w9788 & w29219);
assign w28706 = ~w8141 & w10271;
assign w28707 = pi08 & ~w10280;
assign w28708 = pi08 & ~w28482;
assign w28709 = ~pi08 & w10280;
assign w28710 = ~pi08 & w28482;
assign w28711 = ~w3228 & w8140;
assign v9077 = ~(w10335 | w10275);
assign w28712 = v9077;
assign w28713 = ~w9402 & w10811;
assign v9078 = ~(pi05 | w10823);
assign w28714 = v9078;
assign v9079 = ~(pi05 | w28285);
assign w28715 = v9079;
assign w28716 = pi05 & w10823;
assign w28717 = pi05 & w28285;
assign v9080 = ~(w10905 | w10804);
assign w28718 = v9080;
assign v9081 = ~(w10913 | w10778);
assign w28719 = v9081;
assign w28720 = w10915 & ~w10765;
assign w28721 = w10512 & ~w10511;
assign w28722 = w28295 & ~pi02;
assign w28723 = (~pi02 & w28295) | (~pi02 & w4082) | (w28295 & w4082);
assign w28724 = w28296 | w28297;
assign w28725 = (w28297 & w28296) | (w28297 & ~w4085) | (w28296 & ~w4085);
assign w28726 = pi05 & ~w10998;
assign w28727 = pi05 & ~w28298;
assign w28728 = ~pi05 & w10998;
assign w28729 = ~pi05 & w28298;
assign w28730 = ~pi02 & w11024;
assign v9082 = ~(pi02 | w28177);
assign w28731 = v9082;
assign w28732 = w11027 & ~w11024;
assign w28733 = w11027 & w28177;
assign v9083 = ~(pi02 | w11037);
assign w28734 = v9083;
assign v9084 = ~(pi02 | w28178);
assign w28735 = v9084;
assign w28736 = w11040 & w11037;
assign w28737 = w11040 & w28178;
assign w28738 = w4 & w11052;
assign w28739 = w4 & w11065;
assign w28740 = w4 & w11075;
assign w28741 = w4 & w11090;
assign w28742 = w4 & w11106;
assign w28743 = w4 & w11118;
assign w28744 = w4 & w11128;
assign w28745 = w4 & w11141;
assign w28746 = w4 & w11153;
assign w28747 = ~w11352 & w11340;
assign w28748 = w11435 & ~w11436;
assign w28749 = w8959 & ~w28505;
assign w28750 = w8959 & ~w28506;
assign w28751 = w11761 & ~w11755;
assign v9085 = ~(w11758 | w11843);
assign w28752 = v9085;
assign w28753 = ~w17346 & w29442;
assign w28754 = (pi14 & ~w17359) | (pi14 & w28934) | (~w17359 & w28934);
assign w28755 = w17359 & w28935;
assign w28756 = w11770 & w7765;
assign w28757 = w17861 & w28936;
assign w28758 = (~pi11 & ~w17861) | (~pi11 & w28937) | (~w17861 & w28937);
assign v9086 = ~(w17939 | w17876);
assign w28759 = v9086;
assign w28760 = ~w8141 & w18402;
assign w28761 = w18412 & w29221;
assign w28762 = w18424 & w29222;
assign w28763 = w18424 & w29223;
assign w28764 = (pi08 & ~w18424) | (pi08 & w29224) | (~w18424 & w29224);
assign w28765 = pi08 & ~w18425;
assign v9087 = ~(w8926 | w18488);
assign w28766 = v9087;
assign w28767 = w18501 & ~w28527;
assign w28768 = w18501 & ~w18506;
assign w28769 = ~w18501 & w28527;
assign w28770 = ~w18501 & w18506;
assign v9088 = ~(w18522 | w18429);
assign w28771 = v9088;
assign w28772 = w18222 & ~w18221;
assign w28773 = w18567 & ~w18206;
assign w28774 = w18156 & ~w18155;
assign v9089 = ~(w18576 | w18106);
assign w28775 = v9089;
assign w28776 = w18580 & ~w18076;
assign v9090 = ~(w18582 | w18063);
assign w28777 = v9090;
assign v9091 = ~(w18586 | w18050);
assign w28778 = v9091;
assign w28779 = ~w12382 & w9402;
assign w28780 = w18616 & w28145;
assign w28781 = w18618 & ~w28535;
assign w28782 = ~w9402 & w18635;
assign w28783 = ~w9402 & w18649;
assign w28784 = ~w9402 & w18677;
assign w28785 = ~w9402 & w18710;
assign w28786 = ~w11989 & w10447;
assign w28787 = w18739 & w29964;
assign w28788 = ~w9402 & w19015;
assign w28789 = ~w9402 & w19026;
assign v9092 = ~(w10419 | w19038);
assign w28790 = v9092;
assign w28791 = w19035 & ~w19034;
assign w28792 = ~w19035 & w19034;
assign v9093 = ~(w19139 | w19076);
assign w28793 = v9093;
assign w28794 = w12501 & w28343;
assign w28795 = w19247 & w4;
assign w28796 = w19247 & ~w28344;
assign v9094 = ~(pi02 | w19274);
assign w28797 = v9094;
assign v9095 = ~(pi02 | w28349);
assign w28798 = v9095;
assign w28799 = w19277 & w19274;
assign w28800 = w19277 & w28349;
assign v9096 = ~(pi02 | w19287);
assign w28801 = v9096;
assign v9097 = ~(pi02 | w28350);
assign w28802 = v9097;
assign w28803 = w19290 & w19287;
assign w28804 = w19290 & w28350;
assign v9098 = ~(pi02 | w19298);
assign w28805 = v9098;
assign v9099 = ~(pi02 | w28351);
assign w28806 = v9099;
assign w28807 = w19301 & w19298;
assign w28808 = w19301 & w28351;
assign v9100 = ~(pi02 | w19329);
assign w28809 = v9100;
assign v9101 = ~(pi02 | w28353);
assign w28810 = v9101;
assign w28811 = w19332 & w19329;
assign w28812 = w19332 & w28353;
assign v9102 = ~(w19345 | pi02);
assign w28813 = v9102;
assign w28814 = w19345 & w19348;
assign w28815 = w19770 & ~w19351;
assign v9103 = ~(w18609 | w18607);
assign w28816 = v9103;
assign v9104 = ~(w20009 | w20085);
assign w28817 = v9104;
assign w28818 = ~w8141 & w22103;
assign w28819 = (w29080 & w30919) | (w29080 & w30920) | (w30919 & w30920);
assign w28820 = ~w9402 & w22531;
assign w28821 = ~w9402 & w22541;
assign w28822 = ~pi05 & w22562;
assign w28823 = ~pi05 & w28372;
assign w28824 = pi05 & ~w22562;
assign w28825 = pi05 & ~w28372;
assign w28826 = ~w10419 & w22642;
assign w28827 = w22634 & ~w22651;
assign w28828 = w22660 & ~w22556;
assign w28829 = w22347 & ~w22346;
assign v9105 = ~(w22729 | w22331);
assign w28830 = v9105;
assign v9106 = ~(w22734 | w22275);
assign w28831 = v9106;
assign v9107 = ~(w28217 | w21847);
assign w28832 = v9107;
assign w28833 = w4 & w23183;
assign w28834 = w4 & w23195;
assign w28835 = ~w23206 & pi02;
assign w28836 = w23206 & ~pi02;
assign w28837 = w4 & w23236;
assign v9108 = ~(w11035 | w23270);
assign w28838 = v9108;
assign v9109 = ~(pi02 | w23271);
assign w28839 = v9109;
assign v9110 = ~(pi02 | w28394);
assign w28840 = v9110;
assign w28841 = w23274 & w23271;
assign w28842 = w23274 & w28394;
assign w28843 = w23203 & w23215;
assign w28844 = pi11 & w28432;
assign w28845 = pi11 & w25056;
assign v9111 = ~(pi11 | w28432);
assign w28846 = v9111;
assign v9112 = ~(pi11 | w25056);
assign w28847 = v9112;
assign w28848 = (w25104 & w25112) | (w25104 & w28938) | (w25112 & w28938);
assign w28849 = w25433 & w28939;
assign w28850 = (~pi08 & ~w25433) | (~pi08 & w28940) | (~w25433 & w28940);
assign v9113 = ~(w25264 | w25253);
assign w28851 = v9113;
assign v9114 = ~(w25271 | w25268);
assign w28852 = v9114;
assign w28853 = (w25396 & ~w25405) | (w25396 & w28941) | (~w25405 & w28941);
assign w28854 = w25585 & w28942;
assign w28855 = (~w25453 & w28098) | (~w25453 & w25276) | (w28098 & w25276);
assign w28856 = (~w25453 & w28098) | (~w25453 & ~w28097) | (w28098 & ~w28097);
assign w28857 = pi17 & w28239;
assign w28858 = pi17 & w25937;
assign w28859 = w25812 & w25988;
assign w28860 = (~w25931 & ~w28242) | (~w25931 & w28943) | (~w28242 & w28943);
assign w28861 = (w28105 & ~w26149) | (w28105 & w29225) | (~w26149 & w29225);
assign w28862 = (w28105 & ~w26149) | (w28105 & w29226) | (~w26149 & w29226);
assign w28863 = ~w5114 & w26392;
assign w28864 = (~w26297 & w28106) | (~w26297 & w28104) | (w28106 & w28104);
assign w28865 = (~w26297 & w28106) | (~w26297 & w28103) | (w28106 & w28103);
assign w28866 = ~pi20 & w26541;
assign w28867 = ~pi20 & w28614;
assign w28868 = pi20 & ~w26541;
assign w28869 = pi20 & ~w28614;
assign w28870 = ~w5765 & w26555;
assign w28871 = (w28107 & w28108) | (w28107 & ~w28104) | (w28108 & ~w28104);
assign w28872 = (w28107 & w28108) | (w28107 & ~w28103) | (w28108 & ~w28103);
assign w28873 = ~w5114 & w26680;
assign w28874 = pi23 & w26794;
assign w28875 = pi23 & w28617;
assign v9115 = ~(pi23 | w26794);
assign w28876 = v9115;
assign v9116 = ~(pi23 | w28617);
assign w28877 = v9116;
assign w28878 = pi20 & w26809;
assign w28879 = pi20 & w28618;
assign v9117 = ~(pi20 | w26809);
assign w28880 = v9117;
assign v9118 = ~(pi20 | w28618);
assign w28881 = v9118;
assign w28882 = ~w24280 & w5765;
assign w28883 = ~pi23 & w26924;
assign w28884 = ~pi23 & w28619;
assign w28885 = pi23 & ~w26924;
assign w28886 = pi23 & ~w28619;
assign w28887 = ~w5114 & w26938;
assign v9119 = ~(w26841 | w28247);
assign w28888 = v9119;
assign w28889 = (~w28113 & w28944) | (~w28113 & w28945) | (w28944 & w28945);
assign w28890 = ~w4764 & w27044;
assign w28891 = (w28621 & w28622) | (w28621 & w28247) | (w28622 & w28247);
assign w28892 = (w28113 & w28946) | (w28113 & w28947) | (w28946 & w28947);
assign w28893 = (w28623 & w28624) | (w28623 & ~w28247) | (w28624 & ~w28247);
assign w28894 = (~w28113 & w28948) | (~w28113 & w28949) | (w28948 & w28949);
assign w28895 = (w28627 & w28628) | (w28627 & w28247) | (w28628 & w28247);
assign w28896 = (w28627 & w28628) | (w28627 & w28246) | (w28628 & w28246);
assign w28897 = (w28119 & w28118) | (w28119 & ~w28247) | (w28118 & ~w28247);
assign w28898 = (~w28113 & w28950) | (~w28113 & w28951) | (w28950 & w28951);
assign w28899 = (w28121 & w28122) | (w28121 & w28247) | (w28122 & w28247);
assign w28900 = (w28121 & w28122) | (w28121 & w28246) | (w28122 & w28246);
assign w28901 = (w28631 & w28630) | (w28631 & w28247) | (w28630 & w28247);
assign w28902 = (w28631 & w28630) | (w28631 & w28246) | (w28630 & w28246);
assign w28903 = (w28635 & w28634) | (w28635 & ~w28247) | (w28634 & ~w28247);
assign w28904 = (w28635 & w28634) | (w28635 & ~w28246) | (w28634 & ~w28246);
assign v9120 = ~(w27746 | w28636);
assign w28905 = v9120;
assign w28906 = (w28253 & w28952) | (w28253 & w28953) | (w28952 & w28953);
assign w28907 = w27746 & w28636;
assign w28908 = (~w28253 & w28954) | (~w28253 & w28955) | (w28954 & w28955);
assign w28909 = (w27820 & w28445) | (w27820 & w28444) | (w28445 & w28444);
assign w28910 = (w27820 & w28445) | (w27820 & w28443) | (w28445 & w28443);
assign w28911 = w28446 & ~w28444;
assign w28912 = w28446 & ~w28443;
assign v9121 = ~(w27940 | w28642);
assign w28913 = v9121;
assign v9122 = ~(w27940 | w28641);
assign w28914 = v9122;
assign w28915 = w27940 & w28642;
assign w28916 = w27940 & w28641;
assign v9123 = ~(w27938 | w28644);
assign w28917 = v9123;
assign v9124 = ~(w27938 | w28643);
assign w28918 = v9124;
assign v9125 = ~(w27582 | w27669);
assign w28919 = v9125;
assign v9126 = ~(w9773 | w7178);
assign w28920 = v9126;
assign w28921 = ~w10320 & pi08;
assign w28922 = ~w17872 & pi11;
assign w28923 = ~w28659 & pi11;
assign w28924 = w17872 & ~pi11;
assign w28925 = w26540 & ~w5114;
assign w28926 = w26793 & ~w4764;
assign v9127 = ~(w26808 | w5114);
assign w28927 = v9127;
assign w28928 = w26923 & ~w4764;
assign v9128 = ~(w27142 | w4153);
assign w28929 = v9128;
assign w28930 = ~w869 & w7172;
assign w28931 = ~w869 & w7466;
assign w28932 = ~w3212 & w7765;
assign w28933 = (~w7178 & w3211) | (~w7178 & w29227) | (w3211 & w29227);
assign w28934 = w17356 & pi14;
assign v9129 = ~(w17356 | pi14);
assign w28935 = v9129;
assign w28936 = ~w17862 & pi11;
assign w28937 = w17862 & ~pi11;
assign w28938 = ~w25245 & w25104;
assign w28939 = ~w25434 & pi08;
assign w28940 = w25434 & ~pi08;
assign w28941 = ~w25397 & w25396;
assign v9130 = ~(w25586 | w6389);
assign w28942 = v9130;
assign w28943 = w25938 & ~w25931;
assign v9131 = ~(w26841 | w28107);
assign w28944 = v9131;
assign v9132 = ~(w26841 | w28112);
assign w28945 = v9132;
assign w28946 = (w28621 & w28622) | (w28621 & w28107) | (w28622 & w28107);
assign w28947 = (w28621 & w28622) | (w28621 & w28112) | (w28622 & w28112);
assign w28948 = (w28623 & w28624) | (w28623 & ~w28107) | (w28624 & ~w28107);
assign w28949 = (w28623 & w28624) | (w28623 & ~w28112) | (w28624 & ~w28112);
assign w28950 = (w28119 & w28118) | (w28119 & ~w28107) | (w28118 & ~w28107);
assign w28951 = (w28119 & w28118) | (w28119 & ~w28112) | (w28118 & ~w28112);
assign v9133 = ~(w27746 | w28135);
assign w28952 = v9133;
assign v9134 = ~(w27746 | w28136);
assign w28953 = v9134;
assign w28954 = w27746 & w28135;
assign w28955 = w27746 & w28136;
assign v9135 = ~(w2938 | w28691);
assign w28956 = v9135;
assign w28957 = (~w2938 & ~w2940) | (~w2938 & w29228) | (~w2940 & w29228);
assign w28958 = ~w6389 & w9237;
assign w28959 = pi14 & ~w9252;
assign w28960 = pi14 & ~w28692;
assign w28961 = ~pi14 & w9252;
assign w28962 = ~pi14 & w28692;
assign w28963 = w9260 & ~w9257;
assign w28964 = w9260 & w28693;
assign w28965 = w6383 & pi14;
assign w28966 = (w6871 & ~w3283) | (w6871 & w29229) | (~w3283 & w29229);
assign w28967 = (w7004 & ~w3227) | (w7004 & w29230) | (~w3227 & w29230);
assign w28968 = w9267 & w29443;
assign w28969 = pi11 & ~w9759;
assign w28970 = pi11 & ~w28695;
assign w28971 = ~pi11 & w9759;
assign w28972 = ~pi11 & w28695;
assign w28973 = pi11 & w7172;
assign w28974 = pi11 & w28700;
assign w28975 = w9799 & w29232;
assign w28976 = w9799 & w29233;
assign w28977 = (~pi11 & ~w9799) | (~pi11 & w29234) | (~w9799 & w29234);
assign w28978 = (~pi11 & ~w9799) | (~pi11 & w29444) | (~w9799 & w29444);
assign w28979 = w9803 & ~w9794;
assign w28980 = w9805 & ~w9778;
assign w28981 = ~w8141 & w10259;
assign w28982 = ~pi08 & w10271;
assign w28983 = ~pi08 & w28706;
assign w28984 = pi08 & ~w10271;
assign w28985 = pi08 & ~w28706;
assign v9136 = ~(w10343 | w10252);
assign w28986 = v9136;
assign w28987 = w10109 & ~w10108;
assign w28988 = (w10385 & w29965) | (w10385 & w29966) | (w29965 & w29966);
assign v9137 = ~(w10389 | w10064);
assign w28989 = v9137;
assign w28990 = (w10028 & w10029) | (w10028 & w30280) | (w10029 & w30280);
assign w28991 = w10018 & ~w10017;
assign v9138 = ~(w10397 | w10002);
assign w28992 = v9138;
assign v9139 = ~(w10399 | w9985);
assign w28993 = v9139;
assign v9140 = ~(w10406 | w9935);
assign w28994 = v9140;
assign v9141 = ~(w10408 | w9919);
assign w28995 = v9141;
assign w28996 = ~w9402 & w10423;
assign w28997 = ~w9402 & w10439;
assign w28998 = w11314 & w11448;
assign w28999 = w8957 & ~w8541;
assign v9142 = ~(w11751 | w11749);
assign w29000 = v9142;
assign w29001 = ~w16853 & w29619;
assign w29002 = (pi17 & ~w16866) | (pi17 & w29235) | (~w16866 & w29235);
assign w29003 = w16866 & w29236;
assign w29004 = ~w17332 & w29446;
assign w29005 = (~pi14 & ~w17347) | (~pi14 & w29447) | (~w17347 & w29447);
assign v9143 = ~(pi14 | w28753);
assign w29006 = v9143;
assign w29007 = w17347 & w29448;
assign w29008 = pi14 & w28753;
assign w29009 = (w17392 & ~w17362) | (w17392 & w30281) | (~w17362 & w30281);
assign w29010 = ~w7178 & w17842;
assign w29011 = (~w7765 & ~w11768) | (~w7765 & w29449) | (~w11768 & w29449);
assign w29012 = ~pi11 & w17852;
assign w29013 = w17852 & w17575;
assign w29014 = pi11 & ~w17852;
assign w29015 = (pi11 & ~w17852) | (pi11 & w28672) | (~w17852 & w28672);
assign w29016 = ~w11767 & w7765;
assign v9144 = ~(w17947 | w17856);
assign w29017 = v9144;
assign w29018 = w17799 & ~w17798;
assign v9145 = ~(w17966 | w17783);
assign w29019 = v9145;
assign v9146 = ~(w17969 | w17754);
assign w29020 = v9146;
assign w29021 = (~w17723 & w17972) | (~w17723 & w30921) | (w17972 & w30921);
assign v9147 = ~(w17976 | w17692);
assign w29022 = v9147;
assign v9148 = ~(w17980 | w17661);
assign w29023 = v9148;
assign w29024 = w17615 & ~w17614;
assign w29025 = w17988 & ~w17599;
assign v9149 = ~(w17994 | w17566);
assign w29026 = v9149;
assign w29027 = w17998 & ~w17551;
assign w29028 = w18002 & ~w17536;
assign v9150 = ~(w18006 | w17521);
assign w29029 = v9150;
assign w29030 = w18010 & w29237;
assign v9151 = ~(w19525 | w19530);
assign w29031 = v9151;
assign w29032 = w11770 & w11023;
assign w29033 = w19601 & ~w19600;
assign w29034 = w19579 & ~w19578;
assign w29035 = w19644 & ~w28196;
assign w29036 = w19644 & ~w28553;
assign w29037 = w18609 & w18628;
assign w29038 = (w18609 & w19799) | (w18609 & w29037) | (w19799 & w29037);
assign w29039 = (~w18607 & ~w18609) | (~w18607 & w29238) | (~w18609 & w29238);
assign w29040 = (~w18607 & w28816) | (~w18607 & w28563) | (w28816 & w28563);
assign v9152 = ~(w18609 | w18628);
assign w29041 = v9152;
assign w29042 = ~w19799 & w29041;
assign v9153 = ~(w20006 | w20089);
assign w29043 = v9153;
assign w29044 = w28069 & ~w19907;
assign w29045 = (~w19907 & w28069) | (~w19907 & w12537) | (w28069 & w12537);
assign w29046 = w4 & w20206;
assign v9154 = ~(w20081 | w20015);
assign w29047 = v9154;
assign v9155 = ~(w20081 | w20017);
assign w29048 = v9155;
assign v9156 = ~(w20085 | w20012);
assign w29049 = v9156;
assign w29050 = ~w20085 & w28564;
assign w29051 = ~w20737 & w30101;
assign w29052 = ~w20757 & w30102;
assign w29053 = (w20063 & w30103) | (w20063 & w30104) | (w30103 & w30104);
assign w29054 = ~w20778 & w30105;
assign w29055 = ~w21113 & w29967;
assign w29056 = w21124 & w29968;
assign w29057 = (~pi14 & ~w21124) | (~pi14 & w29969) | (~w21124 & w29969);
assign w29058 = ~w21132 & w30106;
assign w29059 = (w20063 & w30107) | (w20063 & w30108) | (w30107 & w30108);
assign w29060 = ~w21153 & w30109;
assign w29061 = ~w21555 & w29970;
assign w29062 = (w20063 & w29971) | (w20063 & w29972) | (w29971 & w29972);
assign w29063 = ~w20445 & w8141;
assign w29064 = ~w8141 & w22082;
assign w29065 = w22093 & pi08;
assign v9157 = ~(w22093 | pi08);
assign w29066 = v9157;
assign w29067 = pi08 & ~w22103;
assign w29068 = pi08 & ~w28818;
assign w29069 = ~pi08 & w22103;
assign w29070 = ~pi08 & w28818;
assign v9158 = ~(w8926 | w22110);
assign w29071 = v9158;
assign w29072 = pi08 & w28368;
assign w29073 = pi08 & w22113;
assign v9159 = ~(pi08 | w28368);
assign w29074 = v9159;
assign v9160 = ~(pi08 | w22113);
assign w29075 = v9160;
assign w29076 = pi08 & w28369;
assign w29077 = pi08 & w22124;
assign v9161 = ~(pi08 | w28369);
assign w29078 = v9161;
assign v9162 = ~(pi08 | w22124);
assign w29079 = v9162;
assign w29080 = ~w8926 & w22134;
assign w29081 = ~pi08 & w22135;
assign w29082 = ~pi08 & w28819;
assign w29083 = pi08 & ~w22135;
assign w29084 = pi08 & ~w28819;
assign w29085 = pi08 & ~w22145;
assign w29086 = pi08 & ~w28566;
assign w29087 = ~pi08 & w22145;
assign w29088 = ~pi08 & w28566;
assign w29089 = ~w20638 & w9402;
assign w29090 = w28820 | w22531;
assign w29091 = (w22531 & w28820) | (w22531 & w20445) | (w28820 & w20445);
assign v9163 = ~(w22538 | w22540);
assign w29092 = v9163;
assign w29093 = pi05 & w22541;
assign w29094 = pi05 & w28821;
assign v9164 = ~(pi05 | w22541);
assign w29095 = v9164;
assign v9165 = ~(pi05 | w28821);
assign w29096 = v9165;
assign v9166 = ~(w9891 | w22560);
assign w29097 = v9166;
assign v9167 = ~(w10419 | w22569);
assign w29098 = v9167;
assign v9168 = ~(w9891 | w22582);
assign w29099 = v9168;
assign w29100 = ~w9402 & w22625;
assign v9169 = ~(w22502 | w22682);
assign w29101 = v9169;
assign w29102 = w4 & w23171;
assign w29103 = w28833 | w23183;
assign w29104 = (w23183 & w28833) | (w23183 & w20638) | (w28833 & w20638);
assign w29105 = w28834 | w23195;
assign w29106 = (w23195 & w28834) | (w23195 & w20445) | (w28834 & w20445);
assign v9170 = ~(w11035 | w23218);
assign w29107 = v9170;
assign v9171 = ~(w23224 | w23220);
assign w29108 = v9171;
assign w29109 = pi02 & ~w23236;
assign w29110 = pi02 & ~w28837;
assign w29111 = ~w23239 & w23236;
assign w29112 = ~w23239 & w28837;
assign v9172 = ~(w11035 | w23245);
assign w29113 = v9172;
assign v9173 = ~(pi02 | w23246);
assign w29114 = v9173;
assign v9174 = ~(pi02 | w28392);
assign w29115 = v9174;
assign w29116 = w23249 & w23246;
assign w29117 = w23249 & w28392;
assign v9175 = ~(w1 | w23262);
assign w29118 = v9175;
assign w29119 = w23261 & ~w23265;
assign w29120 = w23261 & ~w28393;
assign v9176 = ~(w23267 | w23258);
assign w29121 = v9176;
assign w29122 = w23325 & ~w23202;
assign v9177 = ~(w20200 | w20198);
assign w29123 = v9177;
assign w29124 = ~w7178 & w25421;
assign v9178 = ~(w25443 | w25446);
assign w29125 = v9178;
assign w29126 = pi14 & w28854;
assign w29127 = pi14 & w25587;
assign v9179 = ~(pi14 | w28854);
assign w29128 = v9179;
assign v9180 = ~(pi14 | w25587);
assign w29129 = v9180;
assign w29130 = w25438 & w25620;
assign v9181 = ~(w25438 | w25620);
assign w29131 = v9181;
assign w29132 = ~w6389 & w25644;
assign w29133 = w25463 & ~w25607;
assign w29134 = ~w25809 & w28607;
assign w29135 = ~w25809 & w28608;
assign w29136 = w25809 & ~w28607;
assign w29137 = w25809 & ~w28608;
assign v9182 = ~(w25985 | w28442);
assign w29138 = v9182;
assign v9183 = ~(w25985 | w28441);
assign w29139 = v9183;
assign w29140 = w26151 & ~w28610;
assign w29141 = w26151 & ~w28609;
assign w29142 = w25994 & ~w26126;
assign w29143 = ~w5765 & w26260;
assign w29144 = w26112 & ~w26100;
assign w29145 = w25993 & ~w26140;
assign w29146 = ~w4764 & w26376;
assign w29147 = pi20 & w26392;
assign w29148 = pi20 & w28863;
assign v9184 = ~(pi20 | w26392);
assign w29149 = v9184;
assign v9185 = ~(pi20 | w28863);
assign w29150 = v9185;
assign w29151 = ~w5765 & w26407;
assign w29152 = ~w4764 & w26525;
assign w29153 = w26451 & ~w26560;
assign w29154 = ~w4764 & w26664;
assign w29155 = ~pi20 & w26680;
assign w29156 = ~pi20 & w28873;
assign w29157 = pi20 & ~w26680;
assign w29158 = pi20 & ~w28873;
assign v9186 = ~(w26535 | w26545);
assign w29159 = v9186;
assign w29160 = ~w26717 & w26581;
assign v9187 = ~(w26717 | w28110);
assign w29161 = v9187;
assign w29162 = w26717 & ~w26581;
assign w29163 = w26717 & w28110;
assign w29164 = ~w4153 & w26779;
assign w29165 = ~w26843 & w28246;
assign w29166 = ~w26843 & w28247;
assign w29167 = w26843 & ~w28246;
assign w29168 = w26843 & ~w28247;
assign w29169 = ~w4153 & w26908;
assign v9188 = ~(w26789 | w26787);
assign w29170 = v9188;
assign v9189 = ~(w26842 | w26966);
assign w29171 = v9189;
assign w29172 = w26842 & w26966;
assign w29173 = w26852 & ~w26944;
assign w29174 = ~w4153 & w27028;
assign w29175 = pi23 & w27044;
assign w29176 = pi23 & w28890;
assign v9190 = ~(pi23 | w27044);
assign w29177 = v9190;
assign v9191 = ~(pi23 | w28890);
assign w29178 = v9191;
assign v9192 = ~(w26918 | w26928);
assign w29179 = v9192;
assign w29180 = w28620 & w27084;
assign w29181 = pi26 & w28625;
assign w29182 = pi26 & w27143;
assign v9193 = ~(pi26 | w28625);
assign w29183 = v9193;
assign v9194 = ~(pi26 | w27143);
assign w29184 = v9194;
assign w29185 = pi23 & w27158;
assign w29186 = pi23 & w28626;
assign v9195 = ~(pi23 | w27158);
assign w29187 = v9195;
assign v9196 = ~(pi23 | w28626);
assign w29188 = v9196;
assign w29189 = w28620 & w28120;
assign w29190 = ~pi26 & w27206;
assign w29191 = ~pi26 & w28629;
assign w29192 = pi26 & ~w27206;
assign w29193 = pi26 & ~w28629;
assign w29194 = w28620 & w28123;
assign w29195 = ~pi29 & w27343;
assign w29196 = ~pi29 & w28632;
assign w29197 = pi29 & ~w27343;
assign w29198 = pi29 & ~w28632;
assign w29199 = ~w4153 & w27357;
assign w29200 = ~pi26 & w27452;
assign w29201 = ~pi26 & w28633;
assign w29202 = pi26 & ~w27452;
assign w29203 = pi26 & ~w28633;
assign v9197 = ~(w28125 | w27489);
assign w29204 = v9197;
assign v9198 = ~(w28130 | w27587);
assign w29205 = v9198;
assign w29206 = ~w3529 & w27628;
assign w29207 = (w28638 & w28637) | (w28638 & ~w28443) | (w28637 & ~w28443);
assign w29208 = (w28638 & w28637) | (w28638 & ~w28444) | (w28637 & ~w28444);
assign w29209 = (w28640 & w28639) | (w28640 & w28443) | (w28639 & w28443);
assign w29210 = (w28640 & w28639) | (w28640 & w28444) | (w28639 & w28444);
assign w29211 = ~w26441 & w26298;
assign v9199 = ~(w27191 | w28270);
assign w29212 = v9199;
assign v9200 = ~(w27191 | w28269);
assign w29213 = v9200;
assign w29214 = w3492 & ~w4;
assign v9201 = ~(w9248 | w6389);
assign w29215 = v9201;
assign v9202 = ~(w6871 | w6389);
assign w29216 = v9202;
assign w29217 = ~w9787 & pi11;
assign w29218 = w28703 & w9262;
assign v9203 = ~(w28703 | w9262);
assign w29219 = v9203;
assign v9204 = ~(w17348 | w6389);
assign w29220 = v9204;
assign v9205 = ~(w18413 | w8141);
assign w29221 = v9205;
assign w29222 = w28681 & ~pi08;
assign v9206 = ~(w18421 | pi08);
assign w29223 = v9206;
assign w29224 = ~w28681 & pi08;
assign w29225 = w28102 & w28105;
assign w29226 = w28101 & w28105;
assign v9207 = ~(w7466 | w7178);
assign w29227 = v9207;
assign w29228 = w3001 & ~w2938;
assign w29229 = ~w869 & w6871;
assign w29230 = ~w3212 & w7004;
assign w29231 = (~w6389 & w3211) | (~w6389 & w29216) | (w3211 & w29216);
assign w29232 = w28933 & pi11;
assign w29233 = ~w9800 & pi11;
assign v9208 = ~(w28933 | pi11);
assign w29234 = v9208;
assign w29235 = w16863 & pi17;
assign v9209 = ~(w16863 | pi17);
assign w29236 = v9209;
assign v9210 = ~(w18011 | w8141);
assign w29237 = v9210;
assign v9211 = ~(w18607 | w18628);
assign w29238 = v9211;
assign w29239 = w2218 & w2215;
assign w29240 = w2851 & w2859;
assign w29241 = w2860 & w2849;
assign w29242 = ~w640 & w1945;
assign w29243 = w2888 & ~w488;
assign v9212 = ~(w451 | w566);
assign w29244 = v9212;
assign w29245 = w8803 & w29620;
assign w29246 = w8822 & ~w8818;
assign v9213 = ~(pi14 | w9237);
assign w29247 = v9213;
assign v9214 = ~(pi14 | w28958);
assign w29248 = v9214;
assign w29249 = pi14 & w9237;
assign w29250 = pi14 & w28958;
assign w29251 = ~w3193 & w7004;
assign w29252 = ~w3284 & w6388;
assign w29253 = ~w3284 & w28965;
assign w29254 = w9277 & w29451;
assign w29255 = w9277 & w29452;
assign w29256 = (~pi14 & ~w9277) | (~pi14 & w29453) | (~w9277 & w29453);
assign w29257 = (~pi14 & ~w9277) | (~pi14 & w29621) | (~w9277 & w29621);
assign w29258 = w9281 & ~w9272;
assign w29259 = w9283 & ~w9256;
assign w29260 = ~w7178 & w9750;
assign w29261 = ~w3228 & w7177;
assign v9215 = ~(w9815 | w9754);
assign w29262 = v9215;
assign v9216 = ~(w9823 | w9731);
assign w29263 = v9216;
assign w29264 = (~w9875 & w9872) | (~w9875 & w30571) | (w9872 & w30571);
assign w29265 = ~w9402 & w9893;
assign w29266 = ~w3342 & w9402;
assign v9217 = ~(w10921 | w10752);
assign w29267 = v9217;
assign v9218 = ~(pi02 | w11052);
assign w29268 = v9218;
assign v9219 = ~(pi02 | w28738);
assign w29269 = v9219;
assign w29270 = w11055 & w11052;
assign w29271 = w11055 & w28738;
assign w29272 = w11312 & ~w11311;
assign w29273 = (w11533 & w31234) | (w11533 & w31235) | (w31234 & w31235);
assign v9220 = ~(w8957 | w28749);
assign w29274 = v9220;
assign w29275 = (~w11533 & w31236) | (~w11533 & w31237) | (w31236 & w31237);
assign w29276 = (~w8541 & w28999) | (~w8541 & w28749) | (w28999 & w28749);
assign w29277 = ~w9906 & w10432;
assign v9221 = ~(w9906 | w28009);
assign w29278 = v9221;
assign w29279 = (w11758 & w11840) | (w11758 & w29973) | (w11840 & w29973);
assign w29280 = w28752 & ~w11843;
assign w29281 = (~w11843 & w28752) | (~w11843 & w28322) | (w28752 & w28322);
assign w29282 = w11838 & ~w11758;
assign w29283 = ~w16842 & w30922;
assign w29284 = (w16842 & w30923) | (w16842 & w30924) | (w30923 & w30924);
assign w29285 = ~w11533 & w29456;
assign w29286 = (w17324 & w29622) | (w17324 & w29623) | (w29622 & w29623);
assign w29287 = ~w17324 & w29624;
assign w29288 = ~w11767 & w7004;
assign w29289 = ~pi14 & w17336;
assign w29290 = ~pi14 & w29004;
assign w29291 = pi14 & ~w17336;
assign w29292 = pi14 & ~w29004;
assign w29293 = (pi14 & ~w17387) | (pi14 & w29459) | (~w17387 & w29459);
assign w29294 = w17387 & w29460;
assign w29295 = w28760 & w18402;
assign w29296 = (w18402 & w28760) | (w18402 & ~w14330) | (w28760 & ~w14330);
assign v9222 = ~(pi08 | w28761);
assign w29297 = v9222;
assign v9223 = ~(pi08 | w18414);
assign w29298 = v9223;
assign w29299 = pi08 & w28761;
assign w29300 = pi08 & w18414;
assign w29301 = w18516 & ~w18440;
assign v9224 = ~(w18526 | w18418);
assign w29302 = v9224;
assign v9225 = ~(w18383 | w18538);
assign w29303 = v9225;
assign w29304 = w18317 & ~w18316;
assign w29305 = w12501 & w28779;
assign w29306 = w18602 & ~w18591;
assign w29307 = pi05 & w19015;
assign w29308 = pi05 & w28788;
assign v9226 = ~(pi05 | w19015);
assign w29309 = v9226;
assign v9227 = ~(pi05 | w28788);
assign w29310 = v9227;
assign v9228 = ~(pi05 | w19026);
assign w29311 = v9228;
assign v9229 = ~(pi05 | w28789);
assign w29312 = v9229;
assign w29313 = pi05 & w19026;
assign w29314 = pi05 & w28789;
assign v9230 = ~(w19053 | w19051);
assign w29315 = v9230;
assign w29316 = ~w11767 & w10419;
assign v9231 = ~(w18996 | w19156);
assign w29317 = v9231;
assign w29318 = w14330 & w1;
assign w29319 = w19633 & ~w19657;
assign w29320 = w19658 & w19674;
assign w29321 = ~w17504 & w19809;
assign v9232 = ~(w19998 | w20095);
assign w29322 = v9232;
assign w29323 = ~w20445 & w5765;
assign w29324 = w20730 & pi17;
assign v9233 = ~(w20730 | pi17);
assign w29325 = v9233;
assign w29326 = pi17 & ~w20740;
assign w29327 = pi17 & ~w29051;
assign w29328 = ~pi17 & w20740;
assign w29329 = ~pi17 & w29051;
assign w29330 = ~w20748 & w30110;
assign w29331 = pi17 & w20750;
assign w29332 = w20750 & w30111;
assign v9234 = ~(pi17 | w20750);
assign w29333 = v9234;
assign w29334 = (~pi17 & ~w20750) | (~pi17 & w30112) | (~w20750 & w30112);
assign w29335 = pi17 & ~w20760;
assign w29336 = pi17 & ~w29052;
assign w29337 = ~pi17 & w20760;
assign w29338 = ~pi17 & w29052;
assign w29339 = (w29556 & w30735) | (w29556 & w30736) | (w30735 & w30736);
assign w29340 = pi17 & ~w20771;
assign w29341 = pi17 & ~w29053;
assign w29342 = ~pi17 & w20771;
assign w29343 = ~pi17 & w29053;
assign w29344 = ~pi17 & w20781;
assign w29345 = ~pi17 & w29054;
assign w29346 = pi17 & ~w20781;
assign w29347 = pi17 & ~w29054;
assign w29348 = ~w20445 & w6389;
assign w29349 = w21106 & pi14;
assign v9235 = ~(w21106 | pi14);
assign w29350 = v9235;
assign w29351 = pi14 & ~w21116;
assign w29352 = pi14 & ~w29055;
assign w29353 = ~pi14 & w21116;
assign w29354 = ~pi14 & w29055;
assign v9236 = ~(w7004 | w21123);
assign w29355 = v9236;
assign w29356 = pi14 & ~w21135;
assign w29357 = pi14 & ~w29058;
assign w29358 = ~pi14 & w21135;
assign w29359 = ~pi14 & w29058;
assign w29360 = (w29574 & w30737) | (w29574 & w30738) | (w30737 & w30738);
assign w29361 = pi14 & ~w21146;
assign w29362 = pi14 & ~w29059;
assign w29363 = ~pi14 & w21146;
assign w29364 = ~pi14 & w29059;
assign w29365 = pi14 & ~w21156;
assign w29366 = pi14 & ~w29060;
assign w29367 = ~pi14 & w21156;
assign w29368 = ~pi14 & w29060;
assign w29369 = w21201 & ~w21129;
assign w29370 = ~w20445 & w7178;
assign w29371 = w21548 & pi11;
assign v9237 = ~(w21548 | pi11);
assign w29372 = v9237;
assign w29373 = pi11 & w21558;
assign w29374 = pi11 & w29061;
assign v9238 = ~(pi11 | w21558);
assign w29375 = v9238;
assign v9239 = ~(pi11 | w29061);
assign w29376 = v9239;
assign w29377 = ~w21566 & w29974;
assign w29378 = ~pi11 & w21568;
assign w29379 = w21568 & w17575;
assign w29380 = pi11 & ~w21568;
assign w29381 = (pi11 & ~w21568) | (pi11 & w28672) | (~w21568 & w28672);
assign v9240 = ~(w21575 | w21577);
assign w29382 = v9240;
assign w29383 = pi11 & w21578;
assign w29384 = w21578 & w29975;
assign v9241 = ~(pi11 | w21578);
assign w29385 = v9241;
assign w29386 = (~pi11 & ~w21578) | (~pi11 & w29976) | (~w21578 & w29976);
assign w29387 = (w29589 & w30925) | (w29589 & w30926) | (w30925 & w30926);
assign w29388 = ~pi11 & w21589;
assign w29389 = ~pi11 & w29062;
assign w29390 = pi11 & ~w21589;
assign w29391 = pi11 & ~w29062;
assign w29392 = ~pi11 & w21599;
assign w29393 = ~pi11 & w28565;
assign w29394 = pi11 & ~w21599;
assign w29395 = pi11 & ~w28565;
assign w29396 = ~w20638 & w8141;
assign w29397 = w22072 & pi08;
assign v9242 = ~(w22072 | pi08);
assign w29398 = v9242;
assign w29399 = ~pi08 & w22082;
assign w29400 = ~pi08 & w29064;
assign w29401 = pi08 & ~w22082;
assign w29402 = pi08 & ~w29064;
assign v9243 = ~(w8926 | w22090);
assign w29403 = v9243;
assign v9244 = ~(w8526 | w22101);
assign w29404 = v9244;
assign v9245 = ~(w22112 | w22110);
assign w29405 = v9245;
assign w29406 = ~w22112 & w29071;
assign v9246 = ~(w22120 | w22123);
assign w29407 = v9246;
assign v9247 = ~(w8526 | w22133);
assign w29408 = v9247;
assign w29409 = ~w8141 & w22171;
assign w29410 = w22176 & ~w22149;
assign w29411 = w22180 & ~w22139;
assign w29412 = w22184 & ~w22128;
assign w29413 = w22188 & ~w22117;
assign w29414 = w22196 & ~w22097;
assign w29415 = ~w9402 & w22498;
assign v9248 = ~(w22478 | w22690);
assign w29416 = v9248;
assign w29417 = pi02 & w23160;
assign v9249 = ~(pi02 | w23171);
assign w29418 = v9249;
assign v9250 = ~(pi02 | w29102);
assign w29419 = v9250;
assign w29420 = w23174 & w23171;
assign w29421 = w23174 & w29102;
assign w29422 = w23178 & ~w23177;
assign v9251 = ~(w26299 | w28862);
assign w29423 = v9251;
assign v9252 = ~(w26299 | w28861);
assign w29424 = v9252;
assign w29425 = (w28247 & w28246) | (w28247 & ~w28104) | (w28246 & ~w28104);
assign w29426 = (w28247 & w28246) | (w28247 & ~w28103) | (w28246 & ~w28103);
assign w29427 = w27298 & ~w28900;
assign w29428 = w27298 & ~w28899;
assign w29429 = ~w27298 & w28900;
assign w29430 = ~w27298 & w28899;
assign w29431 = w27395 & w28902;
assign w29432 = w27395 & w28901;
assign v9253 = ~(w27395 | w28902);
assign w29433 = v9253;
assign v9254 = ~(w27395 | w28901);
assign w29434 = v9254;
assign v9255 = ~(w27485 | w28904);
assign w29435 = v9255;
assign v9256 = ~(w27485 | w28903);
assign w29436 = v9256;
assign w29437 = w27485 & w28904;
assign w29438 = w27485 & w28903;
assign v9257 = ~(w11776 | w11788);
assign w29439 = v9257;
assign w29440 = (w10048 & ~w28990) | (w10048 & w30572) | (~w28990 & w30572);
assign v9258 = ~(w9904 | w9418);
assign w29441 = v9258;
assign w29442 = ~w17345 & w29220;
assign w29443 = ~w9263 & pi14;
assign w29444 = w9800 & ~pi11;
assign v9259 = ~(w16855 | w5765);
assign w29445 = v9259;
assign w29446 = w17335 & ~w6389;
assign w29447 = w17348 & ~pi14;
assign w29448 = ~w17348 & pi14;
assign v9260 = ~(w7177 | w7765);
assign w29449 = v9260;
assign v9261 = ~(w2938 | w2848);
assign w29450 = v9261;
assign w29451 = w29231 & pi14;
assign w29452 = ~w9278 & pi14;
assign v9262 = ~(w29231 | pi14);
assign w29453 = v9262;
assign w29454 = ~w16843 & pi17;
assign w29455 = w16843 & ~pi17;
assign w29456 = ~w11764 & w7004;
assign w29457 = w17325 & ~pi14;
assign w29458 = ~w17325 & pi14;
assign w29459 = w17384 & pi14;
assign v9263 = ~(w17384 | pi14);
assign w29460 = v9263;
assign w29461 = (~w2847 & w28691) | (~w2847 & w29625) | (w28691 & w29625);
assign w29462 = (~w2847 & ~w28957) | (~w2847 & w29827) | (~w28957 & w29827);
assign w29463 = ~w2940 & w3001;
assign v9264 = ~(w2940 | w28475);
assign w29464 = v9264;
assign w29465 = ~w5765 & w8790;
assign w29466 = pi17 & w8805;
assign w29467 = pi17 & w29245;
assign v9265 = ~(pi17 | w8805);
assign w29468 = v9265;
assign v9266 = ~(pi17 | w29245);
assign w29469 = v9266;
assign w29470 = (w5756 & ~w3283) | (w5756 & w29626) | (~w3283 & w29626);
assign w29471 = (w6236 & ~w3227) | (w6236 & w29627) | (~w3227 & w29627);
assign w29472 = (w5983 & ~w3283) | (w5983 & w29628) | (~w3283 & w29628);
assign w29473 = w8822 & w29977;
assign w29474 = ~w8819 & w29978;
assign w29475 = (~w8374 & w8819) | (~w8374 & w29979) | (w8819 & w29979);
assign w29476 = w8831 & w29629;
assign w29477 = ~w6389 & w9228;
assign w29478 = ~w3228 & w6388;
assign v9267 = ~(w9293 | w9232);
assign w29479 = v9267;
assign w29480 = ~w7178 & w9738;
assign w29481 = pi11 & w9750;
assign w29482 = pi11 & w29260;
assign v9268 = ~(pi11 | w9750);
assign w29483 = v9268;
assign v9269 = ~(pi11 | w29260);
assign w29484 = v9269;
assign v9270 = ~(w9831 | w9705);
assign w29485 = v9270;
assign v9271 = ~(w10351 | w10226);
assign w29486 = v9271;
assign v9272 = ~(w10929 | w10726);
assign w29487 = v9272;
assign w29488 = w11284 & ~w11283;
assign w29489 = w11254 & ~w11253;
assign w29490 = w4 & w11476;
assign w29491 = ~w28504 & w11502;
assign w29492 = w8540 & w8157;
assign v9273 = ~(w11833 | w28012);
assign w29493 = v9273;
assign v9274 = ~(w11833 | w28188);
assign w29494 = v9274;
assign w29495 = w11850 & ~w11746;
assign w29496 = w11833 & w28012;
assign w29497 = w11833 & w28188;
assign w29498 = w16821 & w29630;
assign w29499 = ~w11533 & w29631;
assign v9275 = ~(pi17 | w29001);
assign w29500 = v9275;
assign w29501 = (~pi17 & ~w16854) | (~pi17 & w29632) | (~w16854 & w29632);
assign w29502 = pi17 & w29001;
assign w29503 = w16854 & w29633;
assign w29504 = ~w16895 & pi17;
assign w29505 = w16894 & w29634;
assign w29506 = (w16900 & ~w16869) | (w16900 & w29980) | (~w16869 & w29980);
assign w29507 = ~w6389 & w17305;
assign w29508 = ~pi14 & w17316;
assign w29509 = w17316 & w29635;
assign w29510 = pi14 & ~w17316;
assign w29511 = (pi14 & ~w17316) | (pi14 & w29636) | (~w17316 & w29636);
assign v9276 = ~(w6389 | w17372);
assign w29512 = v9276;
assign v9277 = ~(w17382 | w17380);
assign w29513 = v9277;
assign v9278 = ~(w17406 | w17329);
assign w29514 = v9278;
assign w29515 = w14330 & w7178;
assign w29516 = pi11 & ~w17842;
assign w29517 = pi11 & ~w29010;
assign w29518 = ~pi11 & w17842;
assign w29519 = ~pi11 & w29010;
assign v9279 = ~(w17943 | w17866);
assign w29520 = v9279;
assign v9280 = ~(w17951 | w17846);
assign w29521 = v9280;
assign v9281 = ~(w17963 | w17811);
assign w29522 = v9281;
assign w29523 = pi08 & w29030;
assign w29524 = pi08 & w18012;
assign v9282 = ~(pi08 | w29030);
assign w29525 = v9282;
assign v9283 = ~(pi08 | w18012);
assign w29526 = v9283;
assign v9284 = ~(w18018 | w18016);
assign w29527 = v9284;
assign w29528 = ~w11989 & w8141;
assign w29529 = ~w8141 & w18116;
assign w29530 = ~w8141 & w18131;
assign w29531 = ~w8141 & w18149;
assign w29532 = ~w8141 & w18378;
assign v9285 = ~(w18358 | w18546);
assign w29533 = v9285;
assign w29534 = ~w9402 & w18991;
assign w29535 = (~w19019 & ~w19148) | (~w19019 & w28646) | (~w19148 & w28646);
assign w29536 = (~w19019 & ~w19148) | (~w19019 & w28645) | (~w19148 & w28645);
assign v9286 = ~(w18971 | w19164);
assign w29537 = v9286;
assign w29538 = w19680 & ~w19503;
assign w29539 = w17007 & w17015;
assign w29540 = w17016 & w19812;
assign v9287 = ~(w17016 | w19812);
assign w29541 = v9287;
assign v9288 = ~(w19993 | w19995);
assign w29542 = v9288;
assign w29543 = ~w20525 & w30114;
assign v9289 = ~(w20095 | w20001);
assign w29544 = v9289;
assign v9290 = ~(w20095 | w20003);
assign w29545 = v9290;
assign w29546 = ~w20638 & w5765;
assign w29547 = w20708 & ~pi17;
assign w29548 = ~w20708 & pi17;
assign w29549 = ~pi17 & w20719;
assign w29550 = w20719 & w30115;
assign w29551 = pi17 & ~w20719;
assign w29552 = (pi17 & ~w20719) | (pi17 & w30116) | (~w20719 & w30116);
assign v9291 = ~(w6236 | w20727);
assign w29553 = v9291;
assign v9292 = ~(w5983 | w20738);
assign w29554 = v9292;
assign v9293 = ~(w5983 | w20758);
assign w29555 = v9293;
assign v9294 = ~(w5983 | w20769);
assign w29556 = v9294;
assign w29557 = ~w5765 & w20809;
assign w29558 = w20814 & ~w20785;
assign w29559 = w20818 & ~w20775;
assign w29560 = w20822 & ~w20764;
assign w29561 = w20826 & ~w20754;
assign w29562 = w20834 & ~w20734;
assign w29563 = ~w20638 & w6389;
assign w29564 = w21084 & w30117;
assign w29565 = (~pi14 & ~w21084) | (~pi14 & w30118) | (~w21084 & w30118);
assign v9295 = ~(w21092 | w21094);
assign w29566 = v9295;
assign w29567 = pi14 & w21095;
assign w29568 = w21095 & w30119;
assign v9296 = ~(pi14 | w21095);
assign w29569 = v9296;
assign w29570 = (~pi14 & ~w21095) | (~pi14 & w30120) | (~w21095 & w30120);
assign v9297 = ~(w7004 | w21103);
assign w29571 = v9297;
assign v9298 = ~(w6871 | w21114);
assign w29572 = v9298;
assign v9299 = ~(w6871 | w21133);
assign w29573 = v9299;
assign v9300 = ~(w6871 | w21144);
assign w29574 = v9300;
assign w29575 = ~w6389 & w21184;
assign w29576 = w21189 & ~w21160;
assign w29577 = w21193 & ~w21150;
assign w29578 = w21197 & ~w21139;
assign v9301 = ~(w21215 | w21099);
assign w29579 = v9301;
assign w29580 = ~w20638 & w7178;
assign w29581 = w21525 & w29981;
assign w29582 = (~pi11 & ~w21525) | (~pi11 & w29982) | (~w21525 & w29982);
assign w29583 = ~pi11 & w21537;
assign w29584 = w21537 & w17575;
assign w29585 = pi11 & ~w21537;
assign w29586 = (pi11 & ~w21537) | (pi11 & w28672) | (~w21537 & w28672);
assign v9302 = ~(w7765 | w21545);
assign w29587 = v9302;
assign v9303 = ~(w7466 | w21556);
assign w29588 = v9303;
assign v9304 = ~(w7466 | w21587);
assign w29589 = v9304;
assign w29590 = ~w7178 & w21627;
assign w29591 = w21632 & ~w21603;
assign w29592 = w21636 & ~w21593;
assign w29593 = w21640 & ~w21582;
assign w29594 = w21644 & ~w21572;
assign w29595 = w21652 & ~w21552;
assign w29596 = ~w8141 & w22050;
assign w29597 = w22061 & ~pi08;
assign w29598 = ~w22061 & pi08;
assign v9305 = ~(w8526 | w22080);
assign w29599 = v9305;
assign v9306 = ~(w8141 | w22158);
assign w29600 = v9306;
assign v9307 = ~(w8926 | w22170);
assign w29601 = v9307;
assign w29602 = ~pi08 & w22171;
assign w29603 = ~pi08 & w29409;
assign w29604 = pi08 & ~w22171;
assign w29605 = pi08 & ~w29409;
assign v9308 = ~(w22210 | w22065);
assign w29606 = v9308;
assign w29607 = ~w9402 & w22473;
assign w29608 = ~w9402 & w22509;
assign w29609 = ~w22521 & pi05;
assign w29610 = w22521 & ~pi05;
assign v9309 = ~(w22525 | w22674);
assign w29611 = v9309;
assign w29612 = pi02 & w23131;
assign w29613 = ~w20654 & w1;
assign v9310 = ~(w1 | w23157);
assign w29614 = v9310;
assign w29615 = w23156 & ~w23160;
assign w29616 = w23156 & ~w29417;
assign w29617 = w23137 & ~w23136;
assign w29618 = (w10544 & w10528) | (w10544 & w30282) | (w10528 & w30282);
assign w29619 = ~w16852 & w29445;
assign v9311 = ~(w8804 | w5765);
assign w29620 = v9311;
assign w29621 = w9278 & ~pi14;
assign w29622 = w29457 | ~pi14;
assign w29623 = (~pi14 & w29457) | (~pi14 & w17323) | (w29457 & w17323);
assign w29624 = ~w17323 & w29458;
assign v9312 = ~(w29450 | w2847);
assign w29625 = v9312;
assign w29626 = ~w869 & w5756;
assign w29627 = ~w3212 & w6236;
assign w29628 = ~w869 & w5983;
assign w29629 = (~w5765 & w3162) | (~w5765 & w29983) | (w3162 & w29983);
assign v9313 = ~(w16822 | w5765);
assign w29630 = v9313;
assign w29631 = ~w11764 & w6236;
assign w29632 = w16855 & ~pi17;
assign w29633 = ~w16855 & pi17;
assign v9314 = ~(w16891 | pi17);
assign w29634 = v9314;
assign v9315 = ~(w6389 | pi14);
assign w29635 = v9315;
assign w29636 = w6389 & pi14;
assign v9316 = ~(w215 | w167);
assign w29637 = v9316;
assign w29638 = w1340 & ~w291;
assign w29639 = w121 & ~w822;
assign v9317 = ~(w88 | w110);
assign w29640 = v9317;
assign w29641 = ~w438 & w884;
assign v9318 = ~(w2814 | w2812);
assign w29642 = v9318;
assign w29643 = w8362 & w29984;
assign w29644 = (~w5114 & w3262) | (~w5114 & w29985) | (w3262 & w29985);
assign w29645 = w8379 & ~w8375;
assign v9319 = ~(pi17 | w8790);
assign w29646 = v9319;
assign v9320 = ~(pi17 | w29465);
assign w29647 = v9320;
assign w29648 = pi17 & w8790;
assign w29649 = pi17 & w29465;
assign w29650 = pi17 & w5756;
assign w29651 = pi17 & w29470;
assign w29652 = pi17 & ~w29476;
assign w29653 = pi17 & ~w8832;
assign w29654 = ~pi17 & w29476;
assign w29655 = ~pi17 & w8832;
assign v9321 = ~(w8835 | w8825);
assign w29656 = v9321;
assign w29657 = w8837 & ~w8809;
assign w29658 = ~w6389 & w9216;
assign w29659 = pi14 & w9228;
assign w29660 = pi14 & w29477;
assign v9322 = ~(pi14 | w9228);
assign w29661 = v9322;
assign v9323 = ~(pi14 | w29477);
assign w29662 = v9323;
assign v9324 = ~(w9301 | w9209);
assign w29663 = v9324;
assign v9325 = ~(w9839 | w9679);
assign w29664 = v9325;
assign v9326 = ~(w10359 | w10200);
assign w29665 = v9326;
assign v9327 = ~(w10937 | w10700);
assign w29666 = v9327;
assign w29667 = w28723 | w28722;
assign w29668 = (w28722 & w28723) | (w28722 & w4083) | (w28723 & w4083);
assign w29669 = w28724 | w28725;
assign w29670 = (w28725 & w28724) | (w28725 & w4135) | (w28724 & w4135);
assign v9328 = ~(pi02 | w11065);
assign w29671 = v9328;
assign v9329 = ~(pi02 | w28739);
assign w29672 = v9329;
assign w29673 = w11068 & w11065;
assign w29674 = w11068 & w28739;
assign v9330 = ~(pi02 | w11075);
assign w29675 = v9330;
assign v9331 = ~(pi02 | w28740);
assign w29676 = v9331;
assign w29677 = w11078 & w11075;
assign w29678 = w11078 & w28740;
assign v9332 = ~(pi02 | w11090);
assign w29679 = v9332;
assign v9333 = ~(pi02 | w28741);
assign w29680 = v9333;
assign w29681 = w11093 & w11090;
assign w29682 = w11093 & w28741;
assign v9334 = ~(pi02 | w11106);
assign w29683 = v9334;
assign v9335 = ~(pi02 | w28742);
assign w29684 = v9335;
assign w29685 = w11109 & w11106;
assign w29686 = w11109 & w28742;
assign v9336 = ~(pi02 | w11118);
assign w29687 = v9336;
assign v9337 = ~(pi02 | w28743);
assign w29688 = v9337;
assign w29689 = w11121 & w11118;
assign w29690 = w11121 & w28743;
assign v9338 = ~(pi02 | w11128);
assign w29691 = v9338;
assign v9339 = ~(pi02 | w28744);
assign w29692 = v9339;
assign w29693 = w11131 & w11128;
assign w29694 = w11131 & w28744;
assign v9340 = ~(pi02 | w11141);
assign w29695 = v9340;
assign v9341 = ~(pi02 | w28745);
assign w29696 = v9341;
assign w29697 = w11144 & w11141;
assign w29698 = w11144 & w28745;
assign v9342 = ~(pi02 | w11153);
assign w29699 = v9342;
assign v9343 = ~(pi02 | w28746);
assign w29700 = v9343;
assign w29701 = w11156 & w11153;
assign w29702 = w11156 & w28746;
assign w29703 = w4 & w11168;
assign w29704 = w4 & w11181;
assign w29705 = w4 & w11191;
assign w29706 = w4 & w11204;
assign w29707 = w4 & w11218;
assign w29708 = ~w11240 & w11227;
assign w29709 = w11240 & ~w11227;
assign w29710 = w11213 & ~w11491;
assign w29711 = ~w11511 & w11158;
assign w29712 = w11150 & ~w11149;
assign w29713 = w11113 & ~w11112;
assign v9344 = ~(w8155 | w8157);
assign w29714 = v9344;
assign v9345 = ~(w8155 | w29492);
assign w29715 = v9345;
assign v9346 = ~(w11058 | w11524);
assign w29716 = v9346;
assign w29717 = (~w11741 & ~w11850) | (~w11741 & w29986) | (~w11850 & w29986);
assign w29718 = ~w16388 & w30927;
assign w29719 = ~w16402 & pi20;
assign w29720 = w16402 & ~pi20;
assign w29721 = ~w5765 & w16812;
assign w29722 = pi17 & w29498;
assign w29723 = pi17 & w16823;
assign v9347 = ~(pi17 | w29498);
assign w29724 = v9347;
assign v9348 = ~(pi17 | w16823);
assign w29725 = v9348;
assign v9349 = ~(w16831 | w16833);
assign w29726 = v9349;
assign v9350 = ~(w16834 | pi17);
assign w29727 = v9350;
assign w29728 = w16834 & pi17;
assign v9351 = ~(w5765 | w16879);
assign w29729 = v9351;
assign w29730 = ~w5765 & w29505;
assign v9352 = ~(w16889 | w16887);
assign w29731 = v9352;
assign v9353 = ~(w16914 | w16838);
assign w29732 = v9353;
assign w29733 = w14330 & w6389;
assign w29734 = pi14 & w17305;
assign w29735 = pi14 & w29507;
assign v9354 = ~(pi14 | w17305);
assign w29736 = v9354;
assign v9355 = ~(pi14 | w29507);
assign w29737 = v9355;
assign v9356 = ~(w17418 | w17298);
assign w29738 = v9356;
assign v9357 = ~(w17426 | w17273);
assign w29739 = v9357;
assign v9358 = ~(w17442 | w17157);
assign w29740 = v9358;
assign w29741 = ~w7178 & w17620;
assign w29742 = ~w11851 & w7178;
assign w29743 = ~w7178 & w17806;
assign w29744 = ~w7178 & w17818;
assign w29745 = w17831 & pi11;
assign v9359 = ~(w17831 | pi11);
assign w29746 = v9359;
assign v9360 = ~(w17959 | w17823);
assign w29747 = v9360;
assign w29748 = w17770 & ~w17769;
assign w29749 = ~w8141 & w18390;
assign v9361 = ~(w18395 | w18534);
assign w29750 = v9361;
assign v9362 = ~(w18345 | w18550);
assign w29751 = v9362;
assign w29752 = w9402 & ~w11851;
assign w29753 = w11845 & w19003;
assign v9363 = ~(w18984 | w19160);
assign w29754 = v9363;
assign v9364 = ~(w18958 | w19168);
assign w29755 = v9364;
assign v9365 = ~(w19488 | w19503);
assign w29756 = v9365;
assign w29757 = ~w19488 & w29538;
assign w29758 = w19681 & ~w19472;
assign w29759 = w19695 & w19457;
assign w29760 = w19695 & ~w28556;
assign v9366 = ~(w16562 | w19812);
assign w29761 = v9366;
assign w29762 = (~w16562 & ~w17016) | (~w16562 & w29761) | (~w17016 & w29761);
assign v9367 = ~(w19990 | w20101);
assign w29763 = v9367;
assign w29764 = ~w20494 & w30739;
assign w29765 = ~w20494 & w30928;
assign w29766 = (pi20 & w20494) | (pi20 & w30740) | (w20494 & w30740);
assign w29767 = (pi20 & w20494) | (pi20 & w30929) | (w20494 & w30929);
assign w29768 = ~pi20 & w20508;
assign w29769 = w20508 & w30121;
assign w29770 = pi20 & ~w20508;
assign w29771 = (pi20 & ~w20508) | (pi20 & w30122) | (~w20508 & w30122);
assign w29772 = ~w5610 & w20517;
assign w29773 = pi20 & ~w20518;
assign w29774 = (pi20 & ~w20518) | (pi20 & w30122) | (~w20518 & w30122);
assign w29775 = ~pi20 & w20518;
assign w29776 = w20518 & w30121;
assign w29777 = pi20 & ~w20528;
assign w29778 = pi20 & ~w29543;
assign w29779 = ~pi20 & w20528;
assign w29780 = ~pi20 & w29543;
assign v9368 = ~(w5765 | w20794);
assign w29781 = v9368;
assign w29782 = pi17 & ~w20809;
assign w29783 = pi17 & ~w29557;
assign w29784 = ~pi17 & w20809;
assign w29785 = ~pi17 & w29557;
assign v9369 = ~(w20840 | w20723);
assign w29786 = v9369;
assign v9370 = ~(w19995 | w19998);
assign w29787 = v9370;
assign w29788 = ~w19995 & w29322;
assign w29789 = w20086 & w21075;
assign w29790 = ~w6389 & w29056;
assign w29791 = w29057 & ~pi14;
assign w29792 = (~pi14 & w29057) | (~pi14 & w6389) | (w29057 & w6389);
assign w29793 = w20086 & w21516;
assign v9371 = ~(w7178 | w21612);
assign w29794 = v9371;
assign w29795 = pi11 & w21627;
assign w29796 = pi11 & w29590;
assign v9372 = ~(pi11 | w21627);
assign w29797 = v9372;
assign v9373 = ~(pi11 | w29590);
assign w29798 = v9373;
assign v9374 = ~(w21658 | w21541);
assign w29799 = v9374;
assign w29800 = ~w20654 & w8141;
assign w29801 = w22037 & w29989;
assign w29802 = w20086 & w29597;
assign w29803 = w29598 & pi08;
assign w29804 = (pi08 & w29598) | (pi08 & ~w20086) | (w29598 & ~w20086);
assign v9375 = ~(w22202 | w22086);
assign w29805 = v9375;
assign w29806 = w29607 | w22473;
assign w29807 = (w22473 & w29607) | (w22473 & w20964) | (w29607 & w20964);
assign w29808 = ~w20654 & w9402;
assign w29809 = ~pi05 & w22498;
assign w29810 = ~pi05 & w29415;
assign w29811 = pi05 & ~w22498;
assign w29812 = pi05 & ~w29415;
assign w29813 = w29609 & pi05;
assign w29814 = (pi05 & w29609) | (pi05 & ~w20086) | (w29609 & ~w20086);
assign w29815 = w20086 & w29610;
assign v9376 = ~(w22545 | w22666);
assign w29816 = v9376;
assign w29817 = w4 & w23115;
assign v9377 = ~(w23128 | w23131);
assign w29818 = v9377;
assign v9378 = ~(w23128 | w29612);
assign w29819 = v9378;
assign v9379 = ~(pi02 | w20086);
assign w29820 = v9379;
assign v9380 = ~(pi02 | w29103);
assign w29821 = v9380;
assign w29822 = w23186 & w20086;
assign w29823 = w23186 & w29103;
assign v9381 = ~(w23321 | w23215);
assign w29824 = v9381;
assign v9382 = ~(w23321 | w23212);
assign w29825 = v9382;
assign w29826 = w23166 & ~w23165;
assign w29827 = w2848 & ~w2847;
assign w29828 = (~w2812 & w29642) | (~w2812 & w29462) | (w29642 & w29462);
assign w29829 = (~w2812 & w29642) | (~w2812 & w29461) | (w29642 & w29461);
assign v9383 = ~(w2727 | w2725);
assign w29830 = v9383;
assign w29831 = ~w5114 & w8347;
assign w29832 = pi20 & w8364;
assign w29833 = pi20 & w29643;
assign v9384 = ~(pi20 | w8364);
assign w29834 = v9384;
assign v9385 = ~(pi20 | w29643);
assign w29835 = v9385;
assign w29836 = w8372 & ~w8369;
assign w29837 = w8372 & w29644;
assign w29838 = w912 & pi20;
assign w29839 = (w5531 & ~w3283) | (w5531 & w29990) | (~w3283 & w29990);
assign w29840 = (w5610 & ~w3227) | (w5610 & w29991) | (~w3227 & w29991);
assign w29841 = w8379 & w30124;
assign w29842 = ~w5765 & w8781;
assign w29843 = ~w3228 & w5764;
assign w29844 = ~w3193 & w5983;
assign v9386 = ~(w8847 | w8785);
assign w29845 = v9386;
assign v9387 = ~(w9309 | w9183);
assign w29846 = v9387;
assign v9388 = ~(w9847 | w9653);
assign w29847 = v9388;
assign w29848 = w9588 & ~w9587;
assign v9389 = ~(w9866 | w9572);
assign w29849 = v9389;
assign w29850 = w9869 & ~w9543;
assign w29851 = ~w9509 & w9507;
assign w29852 = w9497 & ~w9496;
assign v9390 = ~(w9877 | w9479);
assign w29853 = v9390;
assign w29854 = ~pi05 & w9893;
assign w29855 = ~pi05 & w29265;
assign w29856 = pi05 & ~w9893;
assign w29857 = pi05 & ~w29265;
assign v9391 = ~(w10367 | w10174);
assign w29858 = v9391;
assign w29859 = w9953 & ~w9952;
assign v9392 = ~(w10945 | w10674);
assign w29860 = v9392;
assign w29861 = w10479 & ~w10478;
assign w29862 = w7798 & ~w29714;
assign w29863 = w7798 & ~w29715;
assign w29864 = (~pi20 & ~w16389) | (~pi20 & w30930) | (~w16389 & w30930);
assign v9393 = ~(pi20 | w29718);
assign w29865 = v9393;
assign w29866 = w16389 & w30931;
assign w29867 = pi20 & w29718;
assign w29868 = w5610 & w28186;
assign w29869 = w5610 & ~w11783;
assign w29870 = w16436 & ~w16406;
assign v9394 = ~(w16918 | w16827);
assign w29871 = v9394;
assign w29872 = w29286 & ~pi14;
assign w29873 = (~pi14 & w29286) | (~pi14 & w6389) | (w29286 & w6389);
assign w29874 = ~w6389 & w29287;
assign v9395 = ~(w17402 | w17340);
assign w29875 = v9395;
assign v9396 = ~(w17410 | w17320);
assign w29876 = v9396;
assign v9397 = ~(w17422 | w17285);
assign w29877 = v9397;
assign v9398 = ~(w17955 | w17835);
assign w29878 = v9398;
assign v9399 = ~(w18332 | w18554);
assign w29879 = v9399;
assign v9400 = ~(w18945 | w19172);
assign w29880 = v9400;
assign w29881 = w19457 & ~w19472;
assign w29882 = w19457 & ~w19683;
assign w29883 = w19698 & ~w19455;
assign w29884 = w19399 & ~w19398;
assign w29885 = w19371 & ~w19384;
assign w29886 = w19371 & w19703;
assign w29887 = w4 & w19729;
assign w29888 = w28558 | w19745;
assign w29889 = (w19745 & w28558) | (w19745 & w11895) | (w28558 & w11895);
assign w29890 = (~w19771 & ~w19350) | (~w19771 & ~w19767) | (~w19350 & ~w19767);
assign w29891 = (~w19771 & ~w19350) | (~w19771 & w19341) | (~w19350 & w19341);
assign v9401 = ~(w19776 | w19308);
assign w29892 = v9401;
assign w29893 = (~w19254 & ~w19785) | (~w19254 & w31122) | (~w19785 & w31122);
assign w29894 = ~w19230 & w19225;
assign w29895 = w19799 & ~w19223;
assign w29896 = w19799 & w28366;
assign w29897 = w16136 & w29761;
assign w29898 = w16136 & w29762;
assign w29899 = ~w19799 & w19223;
assign v9402 = ~(w19799 | w28366);
assign w29900 = v9402;
assign w29901 = w19230 & ~w19225;
assign w29902 = w20023 & ~w20076;
assign v9403 = ~(w19987 | w20104);
assign w29903 = v9403;
assign w29904 = ~w20474 & w30283;
assign w29905 = pi20 & ~w20487;
assign w29906 = (pi20 & ~w20487) | (pi20 & w30122) | (~w20487 & w30122);
assign w29907 = ~pi20 & w20487;
assign w29908 = w20487 & w30121;
assign w29909 = w19790 & w5610;
assign w29910 = w20082 & w29547;
assign w29911 = w29548 & pi17;
assign w29912 = (pi17 & w29548) | (pi17 & ~w20082) | (w29548 & ~w20082);
assign w29913 = w20082 & w29564;
assign w29914 = w29565 & ~pi14;
assign w29915 = (~pi14 & w29565) | (~pi14 & ~w20082) | (w29565 & ~w20082);
assign w29916 = w29355 & ~w21123;
assign w29917 = (~w21123 & w29355) | (~w21123 & ~w19790) | (w29355 & ~w19790);
assign v9404 = ~(w6389 | w21169);
assign w29918 = v9404;
assign w29919 = w21209 & ~w21110;
assign w29920 = w20082 & w29581;
assign w29921 = w29582 & ~pi11;
assign w29922 = (~pi11 & w29582) | (~pi11 & ~w20082) | (w29582 & ~w20082);
assign w29923 = w20082 & w29397;
assign w29924 = w29398 & ~pi08;
assign w29925 = (~pi08 & w29398) | (~pi08 & ~w20082) | (w29398 & ~w20082);
assign v9405 = ~(w22214 | w22054);
assign w29926 = v9405;
assign v9406 = ~(w22528 | w22530);
assign w29927 = v9406;
assign v9407 = ~(pi05 | w20082);
assign w29928 = v9407;
assign v9408 = ~(pi05 | w29090);
assign w29929 = v9408;
assign w29930 = pi05 & w20082;
assign w29931 = pi05 & w29090;
assign v9409 = ~(w22514 | w22678);
assign w29932 = v9409;
assign v9410 = ~(w22453 | w22698);
assign w29933 = v9410;
assign w29934 = w23123 & ~w23122;
assign w29935 = w23336 & ~w23096;
assign w29936 = w23065 & ~w23339;
assign w29937 = w23054 & ~w23053;
assign v9411 = ~(w23344 | w23037);
assign w29938 = v9411;
assign w29939 = (w30719 & w31238) | (w30719 & w31239) | (w31238 & w31239);
assign v9412 = ~(w22820 | w22818);
assign w29940 = v9412;
assign v9413 = ~(w23564 | w23407);
assign w29941 = v9413;
assign w29942 = ~w23564 & w28573;
assign v9414 = ~(w23505 | w23503);
assign w29943 = v9414;
assign w29944 = w23853 & ~w28580;
assign w29945 = w23853 & ~w28581;
assign w29946 = ~w23853 & w28580;
assign w29947 = ~w23853 & w28581;
assign w29948 = w23828 & ~w23829;
assign v9415 = ~(w23824 | w23822);
assign w29949 = v9415;
assign v9416 = ~(w24026 | w24024);
assign w29950 = v9416;
assign w29951 = w24259 & ~w24260;
assign w29952 = (~w18932 & ~w18908) | (~w18932 & w30932) | (~w18908 & w30932);
assign v9417 = ~(w18919 | w19176);
assign w29953 = v9417;
assign w29954 = ~w19761 & w4;
assign w29955 = (w19254 & w19785) | (w19254 & w31123) | (w19785 & w31123);
assign v9418 = ~(w11531 | w10432);
assign w29956 = v9418;
assign w29957 = (~w11712 & ~w11700) | (~w11712 & w30284) | (~w11700 & w30284);
assign w29958 = ~w19273 & w4;
assign w29959 = ~w19286 & w4;
assign w29960 = ~w19744 & w4;
assign w29961 = w21598 & ~w7178;
assign w29962 = w12381 & ~w4;
assign w29963 = w12381 & w9402;
assign v9419 = ~(w18740 | w9402);
assign w29964 = v9419;
assign w29965 = (w10108 & ~w10082) | (w10108 & w30126) | (~w10082 & w30126);
assign v9420 = ~(w10093 | w28987);
assign w29966 = v9420;
assign w29967 = w21115 & ~w6389;
assign w29968 = ~w21125 & pi14;
assign w29969 = w21125 & ~pi14;
assign w29970 = w21557 & ~w7178;
assign w29971 = ~w7178 & w21588;
assign w29972 = ~w7178 & w29387;
assign w29973 = w11763 & w11758;
assign v9421 = ~(w21565 | w7765);
assign w29974 = v9421;
assign w29975 = ~w7178 & pi11;
assign w29976 = w7178 & ~pi11;
assign w29977 = ~w8818 & pi17;
assign w29978 = w29473 & w8374;
assign v9422 = ~(w29473 | w8374);
assign w29979 = v9422;
assign w29980 = (~w16898 & w30933) | (~w16898 & w30934) | (w30933 & w30934);
assign w29981 = ~w21526 & pi11;
assign w29982 = w21526 & ~pi11;
assign v9423 = ~(w6236 | w5765);
assign w29983 = v9423;
assign v9424 = ~(w8363 | w5114);
assign w29984 = v9424;
assign v9425 = ~(w5531 | w5114);
assign w29985 = v9425;
assign w29986 = w11746 & ~w11741;
assign w29987 = w16377 & ~w5114;
assign v9426 = ~(w16390 | w5114);
assign w29988 = v9426;
assign v9427 = ~(w22038 | w8141);
assign w29989 = v9427;
assign w29990 = ~w869 & w5531;
assign w29991 = ~w3212 & w5610;
assign w29992 = (~w5114 & w3162) | (~w5114 & w30127) | (w3162 & w30127);
assign w29993 = ~w475 & w1448;
assign v9428 = ~(w31 | w128);
assign w29994 = v9428;
assign w29995 = w3350 & w2725;
assign w29996 = w3350 & ~w29830;
assign w29997 = w7979 & w30285;
assign w29998 = w7990 & pi23;
assign w29999 = (~w4764 & w3211) | (~w4764 & w30286) | (w3211 & w30286);
assign w30000 = pi20 & w8347;
assign w30001 = pi20 & w29831;
assign v9429 = ~(pi20 | w8347);
assign w30002 = v9429;
assign v9430 = ~(pi20 | w29831);
assign w30003 = v9430;
assign w30004 = ~w3193 & w5610;
assign w30005 = ~w3284 & w5113;
assign w30006 = ~w3284 & w29838;
assign w30007 = (pi20 & ~w8390) | (pi20 & w30128) | (~w8390 & w30128);
assign w30008 = (pi20 & ~w8390) | (pi20 & w30129) | (~w8390 & w30129);
assign w30009 = w8390 & w30130;
assign w30010 = ~pi20 & w8391;
assign v9431 = ~(w8394 | w8384);
assign w30011 = v9431;
assign w30012 = w8396 & ~w8368;
assign w30013 = ~w5765 & w8769;
assign w30014 = pi17 & w8781;
assign w30015 = pi17 & w29842;
assign v9432 = ~(pi17 | w8781);
assign w30016 = v9432;
assign v9433 = ~(pi17 | w29842);
assign w30017 = v9433;
assign v9434 = ~(w8855 | w8762);
assign w30018 = v9434;
assign v9435 = ~(w9317 | w9157);
assign w30019 = v9435;
assign w30020 = w9064 & ~w9063;
assign v9436 = ~(w9342 | w9048);
assign w30021 = v9436;
assign w30022 = w9347 & ~w9006;
assign w30023 = ~w4082 & w9402;
assign w30024 = ~w8141 & w9429;
assign v9437 = ~(w10375 | w10148);
assign w30025 = v9437;
assign v9438 = ~(w10648 | w10953);
assign w30026 = v9438;
assign v9439 = ~(w7796 | w29862);
assign w30027 = v9439;
assign w30028 = (~w7796 & w29715) | (~w7796 & w30131) | (w29715 & w30131);
assign v9440 = ~(w8540 | w8157);
assign w30029 = v9440;
assign w30030 = w11853 & w11741;
assign w30031 = w11853 & ~w29717;
assign v9441 = ~(w11769 | w28011);
assign w30032 = v9441;
assign v9442 = ~(w11769 | w29493);
assign w30033 = v9442;
assign w30034 = ~w15954 & w30935;
assign w30035 = (pi23 & ~w15967) | (pi23 & w30132) | (~w15967 & w30132);
assign w30036 = w15967 & w30133;
assign w30037 = w16367 & pi20;
assign w30038 = (~pi20 & ~w16365) | (~pi20 & w30134) | (~w16365 & w30134);
assign w30039 = ~w16374 & w30135;
assign w30040 = ~w16374 & w30136;
assign w30041 = (pi20 & w16374) | (pi20 & w30137) | (w16374 & w30137);
assign w30042 = pi20 & ~w16378;
assign w30043 = w16429 & w30936;
assign v9443 = ~(w16446 | w16382);
assign w30044 = v9443;
assign w30045 = w14330 & w5765;
assign w30046 = pi17 & w16812;
assign w30047 = pi17 & w29721;
assign v9444 = ~(pi17 | w16812);
assign w30048 = v9444;
assign v9445 = ~(pi17 | w29721);
assign w30049 = v9445;
assign v9446 = ~(w16926 | w16805);
assign w30050 = v9446;
assign w30051 = ~w6389 & w17268;
assign w30052 = ~w6389 & w17280;
assign w30053 = w17261 & ~w17260;
assign w30054 = (~w17754 & ~w17727) | (~w17754 & w30937) | (~w17727 & w30937);
assign v9447 = ~(w17739 | w17756);
assign w30055 = v9447;
assign w30056 = w18286 & ~w18285;
assign w30057 = w19441 & ~w19427;
assign w30058 = (w30217 & w30938) | (w30217 & w30939) | (w30938 & w30939);
assign w30059 = (~w30217 & w30940) | (~w30217 & w30941) | (w30940 & w30941);
assign w30060 = w18862 & w19736;
assign v9448 = ~(w18862 | w19736);
assign w30061 = v9448;
assign v9449 = ~(pi02 | w12593);
assign w30062 = v9449;
assign v9450 = ~(pi02 | w29888);
assign w30063 = v9450;
assign w30064 = w19748 & w12593;
assign w30065 = w19748 & w29888;
assign w30066 = (w19750 & ~w19739) | (w19750 & w30741) | (~w19739 & w30741);
assign w30067 = (~w16134 & ~w29761) | (~w16134 & w30138) | (~w29761 & w30138);
assign w30068 = (~w16134 & ~w29762) | (~w16134 & w30138) | (~w29762 & w30138);
assign w30069 = w17504 & ~w19809;
assign v9451 = ~(w19790 | w20031);
assign w30070 = v9451;
assign v9452 = ~(w20038 | w20059);
assign w30071 = v9452;
assign v9453 = ~(w20001 | w20003);
assign w30072 = v9453;
assign w30073 = ~w7178 & w21494;
assign w30074 = ~w7178 & w21505;
assign w30075 = w21616 & pi11;
assign v9454 = ~(w21670 | w21509);
assign w30076 = v9454;
assign w30077 = ~w20093 & w30139;
assign w30078 = pi08 & w29801;
assign w30079 = pi08 & w22039;
assign v9455 = ~(pi08 | w29801);
assign w30080 = v9455;
assign v9456 = ~(pi08 | w22039);
assign w30081 = v9456;
assign w30082 = pi08 & ~w22050;
assign w30083 = pi08 & ~w29596;
assign w30084 = ~pi08 & w22050;
assign w30085 = ~pi08 & w29596;
assign v9457 = ~(w22218 | w22043);
assign w30086 = v9457;
assign v9458 = ~(w22466 | w22694);
assign w30087 = v9458;
assign v9459 = ~(w21793 | w21791);
assign w30088 = v9459;
assign v9460 = ~(w22836 | w22834);
assign w30089 = v9460;
assign v9461 = ~(w23521 | w23519);
assign w30090 = v9461;
assign w30091 = (w23829 & w24017) | (w23829 & w30742) | (w24017 & w30742);
assign v9462 = ~(w24018 | w29948);
assign w30092 = v9462;
assign w30093 = w24253 & ~w24254;
assign w30094 = (~w11803 & ~w28319) | (~w11803 & w30288) | (~w28319 & w30288);
assign v9463 = ~(w18893 | w18906);
assign w30095 = v9463;
assign v9464 = ~(w18893 | w19184);
assign w30096 = v9464;
assign v9465 = ~(w20001 | w20006);
assign w30097 = v9465;
assign w30098 = ~w20001 & w20087;
assign w30099 = (~w21722 & ~w21378) | (~w21722 & w31124) | (~w21378 & w31124);
assign w30100 = (~w22865 & ~w21827) | (~w22865 & w30942) | (~w21827 & w30942);
assign w30101 = w20739 & ~w5765;
assign w30102 = w20759 & ~w5765;
assign w30103 = ~w5765 & w20770;
assign w30104 = ~w5765 & w29339;
assign w30105 = w20780 & ~w5765;
assign w30106 = w21134 & ~w6389;
assign w30107 = ~w6389 & w21145;
assign w30108 = ~w6389 & w29360;
assign w30109 = w21155 & ~w6389;
assign v9466 = ~(w20747 | w6236);
assign w30110 = v9466;
assign w30111 = ~w5765 & pi17;
assign w30112 = w5765 & ~pi17;
assign w30113 = ~w20496 & w30743;
assign w30114 = w20527 & ~w5114;
assign v9467 = ~(w5765 | pi17);
assign w30115 = v9467;
assign w30116 = w5765 & pi17;
assign w30117 = ~w21085 & pi14;
assign w30118 = w21085 & ~pi14;
assign w30119 = ~w6389 & pi14;
assign w30120 = w6389 & ~pi14;
assign v9468 = ~(w5114 | pi20);
assign w30121 = v9468;
assign w30122 = w5114 & pi20;
assign w30123 = w20085 & w20697;
assign w30124 = ~w8375 & pi20;
assign v9469 = ~(w20476 | w5114);
assign w30125 = v9469;
assign w30126 = ~w10097 & w30289;
assign v9470 = ~(w5610 | w5114);
assign w30127 = v9470;
assign w30128 = ~w29992 & pi20;
assign w30129 = w8387 & pi20;
assign w30130 = w29992 & ~pi20;
assign v9471 = ~(w7798 | w7796);
assign w30131 = v9471;
assign w30132 = w15964 & pi23;
assign v9472 = ~(w15964 | pi23);
assign w30133 = v9472;
assign w30134 = w16366 & ~pi20;
assign w30135 = w29987 & ~pi20;
assign w30136 = w16377 & ~pi20;
assign w30137 = ~w29987 & pi20;
assign v9473 = ~(w16136 | w16134);
assign w30138 = v9473;
assign w30139 = w20095 & w22028;
assign w30140 = (~w2670 & ~w3350) | (~w2670 & w30447) | (~w3350 & w30447);
assign w30141 = (~w2670 & w29830) | (~w2670 & w30290) | (w29830 & w30290);
assign w30142 = ~w4764 & w7964;
assign v9474 = ~(pi23 | w7981);
assign w30143 = v9474;
assign v9475 = ~(pi23 | w29997);
assign w30144 = v9475;
assign w30145 = pi23 & w7981;
assign w30146 = pi23 & w29997;
assign w30147 = (w4913 & ~w3227) | (w4913 & w30291) | (~w3227 & w30291);
assign w30148 = (w4836 & ~w3283) | (w4836 & w30292) | (~w3283 & w30292);
assign w30149 = w29998 & ~w7986;
assign w30150 = w7996 & ~w7993;
assign w30151 = w7996 & w29999;
assign w30152 = ~w5114 & w8338;
assign w30153 = ~w3228 & w5113;
assign w30154 = ~w3193 & w5531;
assign v9476 = ~(w8406 | w8342);
assign w30155 = v9476;
assign v9477 = ~(w8863 | w8736);
assign w30156 = v9477;
assign v9478 = ~(w9855 | w9627);
assign w30157 = v9478;
assign v9479 = ~(w10383 | w10122);
assign w30158 = v9479;
assign v9480 = ~(w10961 | w10622);
assign w30159 = v9480;
assign w30160 = w11201 & ~w11200;
assign w30161 = w11176 & ~w11175;
assign v9481 = ~(w7481 | w30028);
assign w30162 = v9481;
assign w30163 = (~w7481 & w29862) | (~w7481 & w30294) | (w29862 & w30294);
assign w30164 = ~w7798 & w29714;
assign w30165 = ~w7798 & w29715;
assign w30166 = w11017 & ~w11764;
assign w30167 = (~w11738 & w29717) | (~w11738 & w30448) | (w29717 & w30448);
assign w30168 = (~w11738 & ~w11853) | (~w11738 & w30295) | (~w11853 & w30295);
assign v9482 = ~(w11850 | w14284);
assign w30169 = v9482;
assign v9483 = ~(w11850 | w28027);
assign w30170 = v9483;
assign w30171 = (~pi23 & ~w15955) | (~pi23 & w30943) | (~w15955 & w30943);
assign v9484 = ~(pi23 | w30034);
assign w30172 = v9484;
assign w30173 = w15955 & w30944;
assign w30174 = pi23 & w30034;
assign w30175 = w16001 & ~w15971;
assign w30176 = ~w5114 & w16344;
assign w30177 = w16354 & w30297;
assign w30178 = w11770 & w5610;
assign w30179 = w30038 & ~pi20;
assign w30180 = (~pi20 & w30038) | (~pi20 & w5114) | (w30038 & w5114);
assign w30181 = ~w11767 & w5610;
assign v9485 = ~(w16454 | w16359);
assign w30182 = v9485;
assign w30183 = ~w5765 & w16788;
assign w30184 = w16801 & ~pi17;
assign w30185 = ~w16801 & pi17;
assign v9486 = ~(w16934 | w16781);
assign w30186 = v9486;
assign w30187 = w17232 & ~w17231;
assign v9487 = ~(w17708 | w17723);
assign w30188 = v9487;
assign v9488 = ~(w17708 | w17725);
assign w30189 = v9488;
assign w30190 = w18255 & ~w18254;
assign w30191 = ~w18222 & w18239;
assign w30192 = ~w18222 & w18241;
assign w30193 = w18191 & ~w18190;
assign w30194 = w12503 & w10445;
assign w30195 = w12404 & w10419;
assign v9489 = ~(w9891 | w18614);
assign w30196 = v9489;
assign w30197 = ~w18612 & w13657;
assign w30198 = w18612 & ~w13657;
assign w30199 = ~w9402 & w18664;
assign w30200 = pi05 & w18710;
assign w30201 = pi05 & w28785;
assign v9490 = ~(pi05 | w18710);
assign w30202 = v9490;
assign v9491 = ~(pi05 | w28785);
assign w30203 = v9491;
assign v9492 = ~(pi05 | w28787);
assign w30204 = v9492;
assign v9493 = ~(pi05 | w18741);
assign w30205 = v9493;
assign w30206 = pi05 & w28787;
assign w30207 = pi05 & w18741;
assign w30208 = w18878 & ~w18877;
assign v9494 = ~(w19218 | w18640);
assign w30209 = v9494;
assign v9495 = ~(pi02 | w19313);
assign w30210 = v9495;
assign v9496 = ~(pi02 | w28352);
assign w30211 = v9496;
assign w30212 = w19316 & w19313;
assign w30213 = w19316 & w28352;
assign w30214 = w4 & w19354;
assign w30215 = w19412 & ~w19701;
assign w30216 = ~w19371 & w19384;
assign v9497 = ~(w19371 | w19703);
assign w30217 = v9497;
assign w30218 = (w29762 & w30298) | (w29762 & w30299) | (w30298 & w30299);
assign w30219 = w19816 & ~w30067;
assign v9498 = ~(w16136 | w29761);
assign w30220 = v9498;
assign v9499 = ~(w16136 | w29762);
assign w30221 = v9499;
assign w30222 = w20101 & w19993;
assign w30223 = w20101 & ~w29542;
assign w30224 = w20104 & w19990;
assign w30225 = w20104 & ~w29763;
assign v9500 = ~(w19984 | w20108);
assign w30226 = v9500;
assign w30227 = ~w20314 & w30945;
assign w30228 = (w20314 & w30946) | (w20314 & w30947) | (w30946 & w30947);
assign w30229 = ~w20350 & w30449;
assign w30230 = w20449 & w30450;
assign w30231 = pi20 & w29904;
assign w30232 = w20475 & w30304;
assign v9501 = ~(pi20 | w29904);
assign w30233 = v9501;
assign w30234 = (~pi20 & ~w20475) | (~pi20 & w30305) | (~w20475 & w30305);
assign w30235 = ~w5114 & w20556;
assign w30236 = w20561 & ~w20532;
assign w30237 = w20565 & ~w20522;
assign w30238 = w20569 & ~w20512;
assign w30239 = w20573 & ~w20501;
assign w30240 = ~w5765 & w20673;
assign w30241 = ~w5765 & w20686;
assign w30242 = ~pi17 & w20697;
assign w30243 = w30123 & w31125;
assign w30244 = pi17 & ~w20697;
assign w30245 = (pi17 & ~w30123) | (pi17 & w31126) | (~w30123 & w31126);
assign v9502 = ~(w20848 | w20701);
assign w30246 = v9502;
assign v9503 = ~(w20104 | w19990);
assign w30247 = v9503;
assign w30248 = ~w20104 & w29763;
assign v9504 = ~(w20101 | w19993);
assign w30249 = v9504;
assign w30250 = ~w20101 & w29542;
assign w30251 = w21051 & w30451;
assign w30252 = ~w6389 & w21064;
assign w30253 = ~pi14 & w21184;
assign w30254 = ~pi14 & w29575;
assign w30255 = pi14 & ~w21184;
assign w30256 = pi14 & ~w29575;
assign v9505 = ~(w21227 | w21068);
assign w30257 = v9505;
assign w30258 = ~w7178 & w21483;
assign w30259 = pi11 & w21494;
assign w30260 = pi11 & w30073;
assign v9506 = ~(pi11 | w21494);
assign w30261 = v9506;
assign v9507 = ~(pi11 | w30073);
assign w30262 = v9507;
assign w30263 = ~pi11 & w21505;
assign w30264 = ~pi11 & w30074;
assign w30265 = pi11 & ~w21505;
assign w30266 = pi11 & ~w30074;
assign v9508 = ~(w21674 | w21498);
assign w30267 = v9508;
assign w30268 = ~w8141 & w22016;
assign w30269 = pi08 & w22028;
assign w30270 = pi08 & w30077;
assign v9509 = ~(pi08 | w22028);
assign w30271 = v9509;
assign v9510 = ~(pi08 | w30077);
assign w30272 = v9510;
assign v9511 = ~(w22230 | w22009);
assign w30273 = v9511;
assign v9512 = ~(w22414 | w22710);
assign w30274 = v9512;
assign v9513 = ~(w21779 | w21777);
assign w30275 = v9513;
assign w30276 = w23344 & w23037;
assign w30277 = (w30276 & w30948) | (w30276 & w30949) | (w30948 & w30949);
assign w30278 = w11882 & w9402;
assign w30279 = ~w19297 & w4;
assign w30280 = (~w29849 & w30744) | (~w29849 & w30745) | (w30744 & w30745);
assign w30281 = ~w17354 & w17392;
assign w30282 = ~w10533 & w30950;
assign w30283 = ~w20473 & w30125;
assign v9514 = ~(w11708 | w11712);
assign w30284 = v9514;
assign v9515 = ~(w7980 | w4764);
assign w30285 = v9515;
assign v9516 = ~(w4913 | w4764);
assign w30286 = v9516;
assign v9517 = ~(w15956 | w4764);
assign w30287 = v9517;
assign v9518 = ~(w11803 | w11798);
assign w30288 = v9518;
assign w30289 = ~w10107 & w10092;
assign v9519 = ~(w3350 | w2670);
assign w30290 = v9519;
assign w30291 = ~w3212 & w4913;
assign w30292 = ~w869 & w4836;
assign w30293 = (~w4764 & w3162) | (~w4764 & w30286) | (w3162 & w30286);
assign w30294 = w7796 & ~w7481;
assign v9520 = ~(w11741 | w11738);
assign w30295 = v9520;
assign w30296 = w15943 & ~w4764;
assign v9521 = ~(w16351 | w5114);
assign w30297 = v9521;
assign w30298 = w19816 & w16134;
assign w30299 = w19816 & ~w30138;
assign w30300 = ~w20315 & pi23;
assign w30301 = w20315 & ~pi23;
assign w30302 = ~w20342 & w30746;
assign v9522 = ~(w20434 | w4764);
assign w30303 = v9522;
assign w30304 = ~w20476 & pi20;
assign w30305 = w20476 & ~pi20;
assign w30306 = w3354 & ~w30141;
assign w30307 = w3354 & ~w30140;
assign w30308 = w7624 & w30573;
assign w30309 = w7634 & pi26;
assign w30310 = (~w4153 & w3262) | (~w4153 & w30574) | (w3262 & w30574);
assign v9523 = ~(pi23 | w7964);
assign w30311 = v9523;
assign v9524 = ~(pi23 | w30142);
assign w30312 = v9524;
assign w30313 = pi23 & w7964;
assign w30314 = pi23 & w30142;
assign w30315 = ~w3228 & w4836;
assign w30316 = ~w3284 & w4763;
assign w30317 = w8004 & w30452;
assign w30318 = w8004 & w30453;
assign w30319 = (~pi23 & ~w8004) | (~pi23 & w30454) | (~w8004 & w30454);
assign v9525 = ~(pi23 | w8006);
assign w30320 = v9525;
assign w30321 = w8009 & ~w7999;
assign w30322 = w8011 & ~w7985;
assign w30323 = ~w5114 & w8326;
assign w30324 = ~pi20 & w8338;
assign w30325 = ~pi20 & w30152;
assign w30326 = pi20 & ~w8338;
assign w30327 = pi20 & ~w30152;
assign v9526 = ~(w8414 | w8319);
assign w30328 = v9526;
assign v9527 = ~(w8871 | w8710);
assign w30329 = v9527;
assign v9528 = ~(w9325 | w9131);
assign w30330 = v9528;
assign v9529 = ~(w9863 | w9601);
assign w30331 = v9529;
assign w30332 = w10080 & ~w10079;
assign v9530 = ~(w10576 | w10591);
assign w30333 = v9530;
assign v9531 = ~(w10576 | w10593);
assign w30334 = v9531;
assign w30335 = w10545 & ~w10544;
assign w30336 = w11125 & ~w11124;
assign w30337 = w7480 & w7196;
assign v9532 = ~(w11731 | w30028);
assign w30338 = v9532;
assign v9533 = ~(w11731 | w30027);
assign w30339 = v9533;
assign w30340 = w11731 & w30028;
assign w30341 = w11731 & w30027;
assign w30342 = ~w11857 & w11860;
assign w30343 = ~w15561 & w30951;
assign w30344 = (pi26 & ~w15574) | (pi26 & w30455) | (~w15574 & w30455);
assign w30345 = w15574 & w30456;
assign w30346 = w15933 & pi23;
assign w30347 = (~pi23 & ~w15931) | (~pi23 & w30457) | (~w15931 & w30457);
assign w30348 = ~w15940 & w30458;
assign w30349 = ~w15940 & w30459;
assign w30350 = (pi23 & w15940) | (pi23 & w30460) | (w15940 & w30460);
assign w30351 = pi23 & ~w15944;
assign w30352 = w15994 & w30952;
assign v9534 = ~(w16011 | w15948);
assign w30353 = v9534;
assign w30354 = w14330 & w5114;
assign w30355 = pi20 & ~w16344;
assign w30356 = pi20 & ~w30176;
assign w30357 = ~pi20 & w16344;
assign w30358 = ~pi20 & w30176;
assign w30359 = ~pi20 & w30177;
assign w30360 = ~pi20 & w16355;
assign w30361 = pi20 & ~w30177;
assign w30362 = pi20 & ~w16355;
assign v9535 = ~(w16462 | w16337);
assign w30363 = v9535;
assign w30364 = ~w5765 & w16776;
assign w30365 = w16769 & ~w16768;
assign w30366 = (~w17216 & ~w17190) | (~w17216 & w30953) | (~w17190 & w30953);
assign w30367 = ~w7178 & w28757;
assign w30368 = w28758 & ~pi11;
assign w30369 = (~pi11 & w28758) | (~pi11 & w7178) | (w28758 & w7178);
assign v9536 = ~(w17677 | w17692);
assign w30370 = v9536;
assign v9537 = ~(w17677 | w17694);
assign w30371 = v9537;
assign w30372 = w18746 & ~w18745;
assign w30373 = (~w15752 & w30067) | (~w15752 & w30461) | (w30067 & w30461);
assign v9538 = ~(w15752 | w30218);
assign w30374 = v9538;
assign w30375 = (~w19987 & ~w20104) | (~w19987 & w30462) | (~w20104 & w30462);
assign w30376 = (~w19987 & w29903) | (~w19987 & w29763) | (w29903 & w29763);
assign w30377 = ~pi23 & w20328;
assign w30378 = w20328 & w30463;
assign w30379 = pi23 & ~w20328;
assign w30380 = (pi23 & ~w20328) | (pi23 & w30464) | (~w20328 & w30464);
assign w30381 = ~w20340 & w30747;
assign w30382 = ~w20340 & w30465;
assign w30383 = (pi23 & w20340) | (pi23 & w30466) | (w20340 & w30466);
assign w30384 = (pi23 & w20340) | (pi23 & w30467) | (w20340 & w30467);
assign w30385 = ~pi23 & w20353;
assign w30386 = ~pi23 & w30229;
assign w30387 = pi23 & ~w20353;
assign w30388 = pi23 & ~w30229;
assign w30389 = w20398 & ~w20319;
assign w30390 = w20433 & w30468;
assign w30391 = w20433 & w30469;
assign w30392 = (~pi23 & ~w20433) | (~pi23 & w30470) | (~w20433 & w30470);
assign v9539 = ~(pi23 | w20435);
assign w30393 = v9539;
assign w30394 = pi20 & w20451;
assign w30395 = pi20 & w30230;
assign v9540 = ~(pi20 | w20451);
assign w30396 = v9540;
assign v9541 = ~(pi20 | w30230);
assign w30397 = v9541;
assign w30398 = ~pi20 & w20464;
assign w30399 = w20464 & w30121;
assign w30400 = pi20 & ~w20464;
assign w30401 = (pi20 & ~w20464) | (pi20 & w30122) | (~w20464 & w30122);
assign v9542 = ~(w5114 | w20541);
assign w30402 = v9542;
assign w30403 = ~pi20 & w20556;
assign w30404 = ~pi20 & w30235;
assign w30405 = pi20 & ~w20556;
assign w30406 = pi20 & ~w30235;
assign v9543 = ~(w20591 | w20455);
assign w30407 = v9543;
assign w30408 = ~w20626 & w30748;
assign w30409 = ~w5114 & w20644;
assign w30410 = ~w5765 & w20660;
assign w30411 = ~pi17 & w20673;
assign w30412 = ~pi17 & w30240;
assign w30413 = pi17 & ~w20673;
assign w30414 = pi17 & ~w30240;
assign w30415 = ~pi17 & w20686;
assign w30416 = ~pi17 & w30241;
assign w30417 = pi17 & ~w20686;
assign w30418 = pi17 & ~w30241;
assign v9544 = ~(w20860 | w20664);
assign w30419 = v9544;
assign w30420 = ~w6389 & w21042;
assign w30421 = pi14 & w21053;
assign w30422 = pi14 & w30251;
assign v9545 = ~(pi14 | w21053);
assign w30423 = v9545;
assign v9546 = ~(pi14 | w30251);
assign w30424 = v9546;
assign w30425 = ~pi14 & w21064;
assign w30426 = ~pi14 & w30252;
assign w30427 = pi14 & ~w21064;
assign w30428 = pi14 & ~w30252;
assign v9547 = ~(w21231 | w21057);
assign w30429 = v9547;
assign w30430 = ~w7178 & w21471;
assign w30431 = pi11 & w21483;
assign w30432 = pi11 & w30258;
assign v9548 = ~(pi11 | w21483);
assign w30433 = v9548;
assign v9549 = ~(pi11 | w30258);
assign w30434 = v9549;
assign v9550 = ~(w21686 | w21464);
assign w30435 = v9550;
assign v9551 = ~(w22234 | w21996);
assign w30436 = v9551;
assign v9552 = ~(w22401 | w22714);
assign w30437 = v9552;
assign w30438 = (~w30276 & w30954) | (~w30276 & w30955) | (w30954 & w30955);
assign w30439 = (w23033 & w23017) | (w23033 & w31240) | (w23017 & w31240);
assign w30440 = ~w23019 & w23379;
assign v9553 = ~(w22806 | w22805);
assign w30441 = v9553;
assign v9554 = ~(w23489 | w23487);
assign w30442 = v9554;
assign v9555 = ~(w23808 | w23806);
assign w30443 = v9555;
assign w30444 = w24012 & ~w24013;
assign w30445 = (~w24019 & w24244) | (~w24019 & w31241) | (w24244 & w31241);
assign w30446 = w19442 & ~w19440;
assign v9556 = ~(w2725 | w2670);
assign w30447 = v9556;
assign v9557 = ~(w11853 | w11738);
assign w30448 = v9557;
assign w30449 = w20352 & ~w4764;
assign v9558 = ~(w20450 | w5114);
assign w30450 = v9558;
assign v9559 = ~(w21052 | w6389);
assign w30451 = v9559;
assign w30452 = w30293 & pi23;
assign w30453 = ~w8005 & pi23;
assign v9560 = ~(w30293 | pi23);
assign w30454 = v9560;
assign w30455 = w15571 & pi26;
assign v9561 = ~(w15571 | pi26);
assign w30456 = v9561;
assign w30457 = w15932 & ~pi23;
assign w30458 = w30296 & ~pi23;
assign w30459 = w15943 & ~pi23;
assign w30460 = ~w30296 & pi23;
assign v9562 = ~(w19816 | w15752);
assign w30461 = v9562;
assign v9563 = ~(w19987 | w19990);
assign w30462 = v9563;
assign v9564 = ~(w4764 | pi23);
assign w30463 = v9564;
assign w30464 = w4764 & pi23;
assign w30465 = w20343 & ~pi23;
assign w30466 = ~w30302 & pi23;
assign w30467 = ~w20343 & pi23;
assign w30468 = w30303 & pi23;
assign w30469 = ~w20434 & pi23;
assign v9565 = ~(w30303 | pi23);
assign w30470 = v9565;
assign v9566 = ~(w20628 | w4764);
assign w30471 = v9566;
assign v9567 = ~(w1032 | w56);
assign w30472 = v9567;
assign w30473 = w2639 & w30576;
assign v9568 = ~(w2597 | w30307);
assign w30474 = v9568;
assign w30475 = (~w2597 & w30141) | (~w2597 & w30577) | (w30141 & w30577);
assign w30476 = ~w4153 & w7608;
assign v9569 = ~(pi26 | w7625);
assign w30477 = v9569;
assign v9570 = ~(pi26 | w30308);
assign w30478 = v9570;
assign w30479 = pi26 & w7625;
assign w30480 = pi26 & w30308;
assign w30481 = (w4158 & ~w3283) | (w4158 & w30578) | (~w3283 & w30578);
assign w30482 = (w4155 & ~w3227) | (w4155 & w30579) | (~w3227 & w30579);
assign w30483 = w30309 & ~w7630;
assign w30484 = w7640 & ~w7637;
assign w30485 = w7640 & w30310;
assign w30486 = ~w4764 & w7955;
assign w30487 = ~w3193 & w4836;
assign w30488 = ~w3228 & w4763;
assign v9571 = ~(w8021 | w7959);
assign w30489 = v9571;
assign v9572 = ~(w8422 | w8293);
assign w30490 = v9572;
assign v9573 = ~(w8877 | w8682);
assign w30491 = v9573;
assign v9574 = ~(w9333 | w9105);
assign w30492 = v9574;
assign v9575 = ~(w10049 | w10064);
assign w30493 = v9575;
assign v9576 = ~(w10049 | w10066);
assign w30494 = v9576;
assign w30495 = w11099 & ~w11098;
assign v9577 = ~(w7194 | w7196);
assign w30496 = v9577;
assign v9578 = ~(w7194 | w30337);
assign w30497 = v9578;
assign w30498 = ~w11735 & w11860;
assign w30499 = ~w11735 & w30342;
assign w30500 = (~pi26 & ~w15562) | (~pi26 & w30956) | (~w15562 & w30956);
assign v9579 = ~(pi26 | w30343);
assign w30501 = v9579;
assign w30502 = w15562 & w30957;
assign w30503 = pi26 & w30343;
assign w30504 = w15608 & ~w15578;
assign w30505 = ~w4764 & w15910;
assign w30506 = w15920 & w30582;
assign w30507 = w11770 & w4913;
assign w30508 = w30347 & ~pi23;
assign w30509 = (~pi23 & w30347) | (~pi23 & w4764) | (w30347 & w4764);
assign w30510 = ~w11767 & w4913;
assign v9580 = ~(w4764 | w15980);
assign w30511 = v9580;
assign w30512 = ~w11526 & w4913;
assign v9581 = ~(w16019 | w15925);
assign w30513 = v9581;
assign w30514 = ~w5114 & w16320;
assign w30515 = w16333 & ~pi20;
assign w30516 = ~w16333 & pi20;
assign v9582 = ~(w5114 | w16415);
assign w30517 = v9582;
assign w30518 = ~w11526 & w5610;
assign v9583 = ~(w16470 | w16313);
assign w30519 = v9583;
assign w30520 = w16883 & pi17;
assign w30521 = w16740 & ~w16739;
assign w30522 = w17376 & pi14;
assign v9584 = ~(w17188 | w17173);
assign w30523 = v9584;
assign w30524 = w17644 & ~w17643;
assign w30525 = w18123 & ~w18122;
assign v9585 = ~(w19295 | w19293);
assign w30526 = v9585;
assign w30527 = w20380 & w30749;
assign w30528 = w20281 & ~w20303;
assign v9586 = ~(w4913 | w20432);
assign w30529 = v9586;
assign v9587 = ~(w5531 | w20526);
assign w30530 = v9587;
assign w30531 = w20545 & pi20;
assign v9588 = ~(w20551 | w20549);
assign w30532 = v9588;
assign w30533 = pi23 & w30408;
assign w30534 = w20627 & w30751;
assign v9589 = ~(pi23 | w30408);
assign w30535 = v9589;
assign w30536 = (~pi23 & ~w20627) | (~pi23 & w30752) | (~w20627 & w30752);
assign w30537 = ~pi20 & w20644;
assign w30538 = ~pi20 & w30409;
assign w30539 = pi20 & ~w20644;
assign w30540 = pi20 & ~w30409;
assign w30541 = pi17 & w20660;
assign w30542 = pi17 & w30410;
assign v9590 = ~(pi17 | w20660);
assign w30543 = v9590;
assign v9591 = ~(pi17 | w30410);
assign w30544 = v9591;
assign v9592 = ~(w5983 | w20779);
assign w30545 = v9592;
assign w30546 = w20798 & pi17;
assign v9593 = ~(w20804 | w20802);
assign w30547 = v9593;
assign v9594 = ~(w20634 | w20633);
assign w30548 = v9594;
assign w30549 = ~w20925 & w30958;
assign w30550 = (w20925 & w30959) | (w20925 & w30960) | (w30959 & w30960);
assign w30551 = ~w5114 & w20954;
assign w30552 = ~w5765 & w20970;
assign w30553 = ~w6389 & w21030;
assign w30554 = ~pi14 & w21042;
assign w30555 = ~pi14 & w30420;
assign w30556 = pi14 & ~w21042;
assign w30557 = pi14 & ~w30420;
assign v9595 = ~(w6871 | w21154);
assign w30558 = v9595;
assign w30559 = w21173 & pi14;
assign v9596 = ~(w21179 | w21177);
assign w30560 = v9596;
assign v9597 = ~(w21239 | w21035);
assign w30561 = v9597;
assign v9598 = ~(w20960 | w20958);
assign w30562 = v9598;
assign w30563 = w21319 & w30961;
assign w30564 = ~w5114 & w21335;
assign v9599 = ~(w7466 | w21597);
assign w30565 = v9599;
assign v9600 = ~(w21622 | w21620);
assign w30566 = v9600;
assign v9601 = ~(w21690 | w21451);
assign w30567 = v9601;
assign v9602 = ~(w21357 | w21355);
assign w30568 = v9602;
assign v9603 = ~(w21957 | w21955);
assign w30569 = v9603;
assign v9604 = ~(w22362 | w22726);
assign w30570 = v9604;
assign w30571 = (w9527 & ~w29851) | (w9527 & w30962) | (~w29851 & w30962);
assign w30572 = w10031 & w10048;
assign v9605 = ~(w7621 | w4153);
assign w30573 = v9605;
assign v9606 = ~(w4158 | w4153);
assign w30574 = v9606;
assign v9607 = ~(w15563 | w4153);
assign w30575 = v9607;
assign w30576 = w2633 & w1536;
assign v9608 = ~(w3354 | w2597);
assign w30577 = v9608;
assign w30578 = ~w869 & w4158;
assign w30579 = ~w3212 & w4155;
assign w30580 = (~w4153 & w3262) | (~w4153 & w30756) | (w3262 & w30756);
assign w30581 = w15552 & ~w4153;
assign v9609 = ~(w15917 | w4764);
assign w30582 = v9609;
assign w30583 = (~w30141 & w30757) | (~w30141 & w30963) | (w30757 & w30963);
assign w30584 = (w3358 & w30307) | (w3358 & w30757) | (w30307 & w30757);
assign w30585 = (w3331 & w31127) | (w3331 & w31128) | (w31127 & w31128);
assign w30586 = w7317 & w30965;
assign w30587 = w7329 & pi29;
assign w30588 = (~w3529 & w3262) | (~w3529 & w30966) | (w3262 & w30966);
assign v9610 = ~(pi26 | w7608);
assign w30589 = v9610;
assign v9611 = ~(pi26 | w30476);
assign w30590 = v9611;
assign w30591 = pi26 & w7608;
assign w30592 = pi26 & w30476;
assign v9612 = ~(w3284 | w2873);
assign w30593 = v9612;
assign w30594 = ~w3193 & w4155;
assign w30595 = w7648 & w30758;
assign w30596 = w7648 & w30759;
assign w30597 = (~pi26 & ~w7648) | (~pi26 & w30760) | (~w7648 & w30760);
assign w30598 = (~pi26 & ~w7648) | (~pi26 & w30967) | (~w7648 & w30967);
assign w30599 = w7652 & ~w7643;
assign w30600 = w7654 & ~w7629;
assign w30601 = ~w4764 & w7943;
assign w30602 = pi23 & w7955;
assign w30603 = pi23 & w30486;
assign v9613 = ~(pi23 | w7955);
assign w30604 = v9613;
assign v9614 = ~(pi23 | w30486);
assign w30605 = v9614;
assign v9615 = ~(w8029 | w7936);
assign w30606 = v9615;
assign v9616 = ~(w8430 | w8267);
assign w30607 = v9616;
assign v9617 = ~(w8885 | w8656);
assign w30608 = v9617;
assign v9618 = ~(w9079 | w9077);
assign w30609 = v9618;
assign w30610 = w9559 & ~w9558;
assign v9619 = ~(w10545 | w10560);
assign w30611 = v9619;
assign v9620 = ~(w10545 | w10562);
assign w30612 = v9620;
assign w30613 = w11072 & ~w11071;
assign w30614 = w11550 & ~w30496;
assign w30615 = w11550 & ~w30497;
assign w30616 = w15201 & w30968;
assign w30617 = (pi29 & ~w15214) | (pi29 & w30761) | (~w15214 & w30761);
assign w30618 = w15214 & w30762;
assign w30619 = (pi26 & ~w15542) | (pi26 & w30969) | (~w15542 & w30969);
assign w30620 = w15542 & w30763;
assign w30621 = ~w15549 & w30764;
assign w30622 = ~w15549 & w30765;
assign w30623 = (pi26 & w15549) | (pi26 & w30766) | (w15549 & w30766);
assign w30624 = pi26 & ~w15553;
assign w30625 = w15601 & w30970;
assign v9621 = ~(w15618 | w15557);
assign w30626 = v9621;
assign w30627 = w14330 & w4764;
assign w30628 = pi23 & w15910;
assign w30629 = pi23 & w30505;
assign v9622 = ~(pi23 | w15910);
assign w30630 = v9622;
assign v9623 = ~(pi23 | w30505);
assign w30631 = v9623;
assign w30632 = ~pi23 & w30506;
assign w30633 = ~pi23 & w15921;
assign w30634 = pi23 & ~w30506;
assign w30635 = pi23 & ~w15921;
assign v9624 = ~(w16027 | w15903);
assign w30636 = v9624;
assign w30637 = ~w5114 & w16308;
assign w30638 = w16301 & ~w16300;
assign w30639 = (w16724 & w16697) | (w16724 & w30971) | (w16697 & w30971);
assign v9625 = ~(w17446 | w17142);
assign w30640 = v9625;
assign w30641 = w17630 & ~w17986;
assign v9626 = ~(w18139 | w18141);
assign w30642 = v9626;
assign v9627 = ~(w18701 | w18703);
assign w30643 = v9627;
assign w30644 = w19819 & ~w15392;
assign v9628 = ~(w19976 | w19819);
assign w30645 = v9628;
assign w30646 = ~w19816 & w30067;
assign w30647 = ~w19816 & w30068;
assign v9629 = ~(w20033 | w20069);
assign w30648 = v9629;
assign v9630 = ~(w20033 | w20067);
assign w30649 = v9630;
assign v9631 = ~(w19981 | w20112);
assign w30650 = v9631;
assign w30651 = ~w20274 & w30972;
assign w30652 = w20071 & w30768;
assign w30653 = w20041 & ~w20059;
assign v9632 = ~(w4836 | w20351);
assign w30654 = v9632;
assign w30655 = ~w20362 & w30769;
assign v9633 = ~(w4764 | w20367);
assign w30656 = v9633;
assign v9634 = ~(w4913 | w20379);
assign w30657 = v9634;
assign w30658 = ~pi23 & w20381;
assign w30659 = ~pi23 & w30527;
assign w30660 = pi23 & ~w20381;
assign w30661 = pi23 & ~w30527;
assign w30662 = w20386 & ~w20357;
assign w30663 = w29764 & w29765;
assign w30664 = (w29765 & w29764) | (w29765 & ~w20310) | (w29764 & ~w20310);
assign w30665 = w29766 | w29767;
assign w30666 = (w29767 & w29766) | (w29767 & w20310) | (w29766 & w20310);
assign v9635 = ~(w20583 | w20480);
assign w30667 = v9635;
assign w30668 = w29331 & w29332;
assign w30669 = (w29332 & w29331) | (w29332 & ~w20310) | (w29331 & ~w20310);
assign w30670 = w29333 | w29334;
assign w30671 = (w29334 & w29333) | (w29334 & w20310) | (w29333 & w20310);
assign w30672 = w20840 & w20734;
assign w30673 = w20840 & w20836;
assign v9636 = ~(w20844 | w20712);
assign w30674 = v9636;
assign v9637 = ~(w20852 | w20690);
assign w30675 = v9637;
assign w30676 = w20071 & w30770;
assign v9638 = ~(w20840 | w20734);
assign w30677 = v9638;
assign v9639 = ~(w20840 | w20836);
assign w30678 = v9639;
assign w30679 = w29790 & w29056;
assign w30680 = (w29056 & w29790) | (w29056 & ~w20310) | (w29790 & ~w20310);
assign w30681 = w29791 | w29792;
assign w30682 = (w29792 & w29791) | (w29792 & w20310) | (w29791 & w20310);
assign w30683 = w21215 & w21110;
assign w30684 = w21215 & w21211;
assign v9640 = ~(w21219 | w21089);
assign w30685 = v9640;
assign v9641 = ~(w21235 | w21046);
assign w30686 = v9641;
assign v9642 = ~(w21243 | w21023);
assign w30687 = v9642;
assign v9643 = ~(w21215 | w21110);
assign w30688 = v9643;
assign v9644 = ~(w21215 | w21211);
assign w30689 = v9644;
assign w30690 = w29378 & w29379;
assign w30691 = (w29379 & w29378) | (w29379 & ~w20310) | (w29378 & ~w20310);
assign w30692 = w29380 | w29381;
assign w30693 = (w29381 & w29380) | (w29381 & w20310) | (w29380 & w20310);
assign w30694 = w21658 & w21552;
assign w30695 = w21658 & w21654;
assign v9645 = ~(w21662 | w21530);
assign w30696 = v9645;
assign v9646 = ~(w21678 | w21487);
assign w30697 = v9646;
assign v9647 = ~(w21694 | w21438);
assign w30698 = v9647;
assign w30699 = ~w928 & w21749;
assign v9648 = ~(w21658 | w21552);
assign w30700 = v9648;
assign v9649 = ~(w21658 | w21654);
assign w30701 = v9649;
assign v9650 = ~(w8526 | w22143);
assign w30702 = v9650;
assign w30703 = w22162 & pi08;
assign v9651 = ~(w22169 | w22170);
assign w30704 = v9651;
assign w30705 = ~w22169 & w29601;
assign v9652 = ~(w22168 | w22166);
assign w30706 = v9652;
assign w30707 = w22202 & w22097;
assign w30708 = w22202 & w22198;
assign v9653 = ~(w22222 | w22032);
assign w30709 = v9653;
assign v9654 = ~(w22238 | w21983);
assign w30710 = v9654;
assign v9655 = ~(w22202 | w22097);
assign w30711 = v9655;
assign v9656 = ~(w22202 | w22198);
assign w30712 = v9656;
assign v9657 = ~(w22440 | w22702);
assign w30713 = v9657;
assign v9658 = ~(w22388 | w22718);
assign w30714 = v9658;
assign w30715 = w20071 & w30771;
assign w30716 = ~w28078 & w23354;
assign w30717 = w23355 & w23365;
assign v9659 = ~(w23035 | w23376);
assign w30718 = v9659;
assign v9660 = ~(w23035 | w23366);
assign w30719 = v9660;
assign w30720 = ~w23018 & w29939;
assign v9661 = ~(w23018 | w30439);
assign w30721 = v9661;
assign w30722 = w23005 & ~w23004;
assign w30723 = ~w4153 & w23467;
assign w30724 = ~w4764 & w23482;
assign v9662 = ~(w23459 | w23457);
assign w30725 = v9662;
assign v9663 = ~(w23445 | w23443);
assign w30726 = v9663;
assign v9664 = ~(w23777 | w23776);
assign w30727 = v9664;
assign w30728 = w20310 & w928;
assign v9665 = ~(w23981 | w23979);
assign w30729 = v9665;
assign v9666 = ~(w24224 | w24222);
assign w30730 = v9666;
assign v9667 = ~(w24238 | w24460);
assign w30731 = v9667;
assign w30732 = w20033 & w20069;
assign w30733 = w20033 & w20067;
assign w30734 = ~w11715 & w29957;
assign v9668 = ~(w6236 | w20769);
assign w30735 = v9668;
assign w30736 = ~w6236 & w20038;
assign v9669 = ~(w7004 | w21144);
assign w30737 = v9669;
assign w30738 = ~w7004 & w20038;
assign w30739 = w20497 & ~pi20;
assign w30740 = ~w20497 & pi20;
assign w30741 = w19735 & w19750;
assign w30742 = ~w23827 & w31242;
assign v9670 = ~(w20495 | w5114);
assign w30743 = v9670;
assign w30744 = w10028 & w9572;
assign w30745 = w10028 & w9574;
assign v9671 = ~(w20341 | w4764);
assign w30746 = v9671;
assign w30747 = w30302 & ~pi23;
assign w30748 = ~w20625 & w30471;
assign v9672 = ~(w20378 | w4764);
assign w30749 = v9672;
assign w30750 = ~w20415 & w30973;
assign w30751 = ~w20628 & pi23;
assign w30752 = w20628 & ~pi23;
assign w30753 = ~w20926 & pi26;
assign w30754 = w20926 & ~pi26;
assign v9673 = ~(w21307 | w4153);
assign w30755 = v9673;
assign w30756 = w2873 & ~w4153;
assign w30757 = w2597 & w3358;
assign w30758 = w30580 & pi26;
assign w30759 = ~w7649 & pi26;
assign v9674 = ~(w30580 | pi26);
assign w30760 = v9674;
assign w30761 = w15211 & pi29;
assign v9675 = ~(w15211 | pi29);
assign w30762 = v9675;
assign v9676 = ~(w15539 | pi26);
assign w30763 = v9676;
assign w30764 = w30581 & ~pi26;
assign w30765 = w15552 & ~pi26;
assign w30766 = ~w30581 & pi26;
assign v9677 = ~(w20273 | w4153);
assign w30767 = v9677;
assign w30768 = ~w20032 & w4764;
assign v9678 = ~(w20361 | w20359);
assign w30769 = v9678;
assign w30770 = ~w20032 & w4153;
assign w30771 = ~w20032 & w3529;
assign v9679 = ~(w201 | w90);
assign w30772 = v9679;
assign w30773 = w1446 & w1443;
assign w30774 = w1904 & w1391;
assign w30775 = w1912 & w1916;
assign w30776 = w2185 & w2188;
assign w30777 = w2369 & w1287;
assign w30778 = w1535 & w2518;
assign w30779 = w2540 & ~w533;
assign v9680 = ~(w263 | w753);
assign w30780 = v9680;
assign w30781 = w2191 & w2594;
assign w30782 = w1441 & w2598;
assign w30783 = w2602 & ~w74;
assign w30784 = w2699 & w2722;
assign w30785 = w2569 & w3362;
assign v9681 = ~(w928 | w6642);
assign w30786 = v9681;
assign w30787 = w6680 & ~w6677;
assign w30788 = w6680 & w30585;
assign w30789 = ~w3529 & w7303;
assign v9682 = ~(pi29 | w7319);
assign w30790 = v9682;
assign v9683 = ~(pi29 | w30586);
assign w30791 = v9683;
assign w30792 = pi29 & w7319;
assign w30793 = pi29 & w30586;
assign w30794 = (w3760 & ~w3227) | (w3760 & w30974) | (~w3227 & w30974);
assign w30795 = (w3763 & ~w3283) | (w3763 & w30975) | (~w3283 & w30975);
assign w30796 = w30587 & ~w7325;
assign w30797 = w7335 & ~w7332;
assign w30798 = w7335 & w30588;
assign w30799 = ~w4153 & w7599;
assign w30800 = ~w3193 & w4158;
assign v9684 = ~(w7664 | w7603);
assign w30801 = v9684;
assign v9685 = ~(w8037 | w7910);
assign w30802 = v9685;
assign v9686 = ~(w8438 | w8241);
assign w30803 = v9686;
assign v9687 = ~(w8893 | w8630);
assign w30804 = v9687;
assign w30805 = w9345 & ~w9035;
assign v9688 = ~(w9528 | w9543);
assign w30806 = v9688;
assign v9689 = ~(w9528 | w9545);
assign w30807 = v9689;
assign v9690 = ~(w28320 | w11014);
assign w30808 = v9690;
assign w30809 = ~w15190 & w31243;
assign v9691 = ~(w15622 | w15546);
assign w30810 = v9691;
assign v9692 = ~(w16015 | w15937);
assign w30811 = v9692;
assign v9693 = ~(w16031 | w15890);
assign w30812 = v9693;
assign v9694 = ~(w16450 | w16371);
assign w30813 = v9694;
assign v9695 = ~(w16466 | w16325);
assign w30814 = v9695;
assign v9696 = ~(w16473 | w16285);
assign w30815 = v9696;
assign w30816 = ~w5765 & w29283;
assign w30817 = w29284 & ~pi17;
assign w30818 = (~pi17 & w29284) | (~pi17 & w5765) | (w29284 & w5765);
assign v9697 = ~(w16930 | w16793);
assign w30819 = v9697;
assign v9698 = ~(w16937 | w16753);
assign w30820 = v9698;
assign w30821 = ~w16708 & w16709;
assign v9699 = ~(w16708 | w16941);
assign w30822 = v9699;
assign v9700 = ~(w17429 | w17245);
assign w30823 = v9700;
assign w30824 = w17433 & ~w17201;
assign v9701 = ~(w17723 | w17725);
assign w30825 = v9701;
assign v9702 = ~(w17707 | w30189);
assign w30826 = v9702;
assign v9703 = ~(w17707 | w30188);
assign w30827 = v9703;
assign v9704 = ~(w18906 | w19184);
assign w30828 = v9704;
assign w30829 = (~w18893 & ~w19188) | (~w18893 & w30096) | (~w19188 & w30096);
assign w30830 = (~w18893 & ~w19188) | (~w18893 & w30095) | (~w19188 & w30095);
assign w30831 = w19713 & ~w28557;
assign w30832 = w19713 & ~w29885;
assign v9705 = ~(w19724 | w19367);
assign w30833 = v9705;
assign v9706 = ~(w19724 | w19714);
assign w30834 = v9706;
assign w30835 = w19725 & w19753;
assign w30836 = w15065 & ~w15392;
assign w30837 = w15065 & w30644;
assign v9707 = ~(w19975 | w20116);
assign w30838 = v9707;
assign w30839 = ~w20248 & w30978;
assign v9708 = ~(w4153 | w20258);
assign w30840 = v9708;
assign w30841 = ~pi26 & w30651;
assign w30842 = w20276 & w30979;
assign w30843 = pi26 & ~w30651;
assign w30844 = (pi26 & ~w20276) | (pi26 & w30980) | (~w20276 & w30980);
assign w30845 = ~pi26 & w20299;
assign w30846 = w20299 & w30981;
assign w30847 = pi26 & ~w20299;
assign w30848 = (pi26 & ~w20299) | (pi26 & w30982) | (~w20299 & w30982);
assign w30849 = ~w30655 & pi23;
assign w30850 = ~w20366 & pi23;
assign v9709 = ~(w20377 | w20375);
assign w30851 = v9709;
assign w30852 = ~w20414 & w30983;
assign w30853 = ~w20414 & w30984;
assign w30854 = (pi26 & w20414) | (pi26 & w30985) | (w20414 & w30985);
assign w30855 = pi26 & ~w20418;
assign v9710 = ~(w20587 | w20468);
assign w30856 = v9710;
assign w30857 = ~w20602 & w31129;
assign w30858 = ~pi26 & w20615;
assign w30859 = w20615 & w30981;
assign w30860 = pi26 & ~w20615;
assign w30861 = (pi26 & ~w20615) | (pi26 & w30982) | (~w20615 & w30982);
assign v9711 = ~(w20856 | w20677);
assign w30862 = v9711;
assign w30863 = pi29 & w20913;
assign w30864 = w20913 & w30987;
assign v9712 = ~(pi29 | w20913);
assign w30865 = v9712;
assign w30866 = (~pi29 & ~w20913) | (~pi29 & w30988) | (~w20913 & w30988);
assign w30867 = ~pi23 & w20940;
assign w30868 = w20940 & w30463;
assign w30869 = pi23 & ~w20940;
assign w30870 = (pi23 & ~w20940) | (pi23 & w30464) | (~w20940 & w30464);
assign w30871 = ~pi20 & w20954;
assign w30872 = ~pi20 & w30551;
assign w30873 = pi20 & ~w20954;
assign w30874 = pi20 & ~w30551;
assign v9713 = ~(w21247 | w21008);
assign w30875 = v9713;
assign v9714 = ~(w20946 | w20945);
assign w30876 = v9714;
assign w30877 = (~pi29 & ~w21293) | (~pi29 & w30989) | (~w21293 & w30989);
assign w30878 = w21293 & w30990;
assign w30879 = (~pi26 & ~w21306) | (~pi26 & w31130) | (~w21306 & w31130);
assign w30880 = (~pi26 & ~w21306) | (~pi26 & w30991) | (~w21306 & w30991);
assign w30881 = w21306 & w30992;
assign w30882 = w21306 & w30993;
assign w30883 = pi23 & w21321;
assign w30884 = pi23 & w30563;
assign v9715 = ~(pi23 | w21321);
assign w30885 = v9715;
assign v9716 = ~(pi23 | w30563);
assign w30886 = v9716;
assign w30887 = pi20 & w21335;
assign w30888 = pi20 & w30564;
assign v9717 = ~(pi20 | w21335);
assign w30889 = v9717;
assign v9718 = ~(pi20 | w30564);
assign w30890 = v9718;
assign v9719 = ~(w21702 | w21412);
assign w30891 = v9719;
assign v9720 = ~(w21341 | w21340);
assign w30892 = v9720;
assign w30893 = ~w21783 & w31131;
assign w30894 = ~w5114 & w21801;
assign w30895 = w21942 & ~w21941;
assign w30896 = w22316 & ~w22315;
assign v9721 = ~(w21824 | w21822);
assign w30897 = v9721;
assign w30898 = ~w22798 & w31132;
assign w30899 = ~w22867 & w21842;
assign v9722 = ~(w22867 | w28574);
assign w30900 = v9722;
assign w30901 = ~w928 & w23744;
assign w30902 = w23754 & w31244;
assign w30903 = ~w4153 & w23770;
assign w30904 = ~w4764 & w23785;
assign v9723 = ~(w23762 | w23761);
assign w30905 = v9723;
assign v9724 = ~(w23748 | w23746);
assign w30906 = v9724;
assign w30907 = w23931 & ~w928;
assign w30908 = w23931 & ~w20309;
assign v9725 = ~(w23965 | w23964);
assign w30909 = v9725;
assign w30910 = ~w928 & w24156;
assign v9726 = ~(w24019 | w23704);
assign w30911 = v9726;
assign v9727 = ~(w24019 | w30091);
assign w30912 = v9727;
assign v9728 = ~(w24208 | w24206);
assign w30913 = v9728;
assign v9729 = ~(w24445 | w24443);
assign w30914 = v9729;
assign w30915 = w24242 & ~w24461;
assign v9730 = ~(w18906 | w18919);
assign w30916 = v9730;
assign v9731 = ~(w18906 | w19180);
assign w30917 = v9731;
assign w30918 = w22144 & ~w8141;
assign w30919 = ~w8141 & w22134;
assign w30920 = ~w8141 & w20063;
assign w30921 = w17738 & ~w17723;
assign w30922 = ~w16841 & w29454;
assign w30923 = w29455 | ~pi17;
assign w30924 = (~pi17 & w29455) | (~pi17 & w16841) | (w29455 & w16841);
assign v9732 = ~(w7765 | w21587);
assign w30925 = v9732;
assign w30926 = ~w7765 & w20038;
assign w30927 = ~w16387 & w29988;
assign w30928 = w30113 & ~pi20;
assign w30929 = ~w30113 & pi20;
assign w30930 = w16390 & ~pi20;
assign w30931 = ~w16390 & pi20;
assign w30932 = w18918 & ~w18932;
assign v9733 = ~(w16861 | w16887);
assign w30933 = v9733;
assign w30934 = ~w16861 & w29731;
assign w30935 = ~w15953 & w30287;
assign v9734 = ~(w16426 | w5114);
assign w30936 = v9734;
assign v9735 = ~(w17737 | w17754);
assign w30937 = v9735;
assign w30938 = w19367 & ~w28557;
assign w30939 = w19367 & w30216;
assign w30940 = ~w19367 & w28557;
assign v9736 = ~(w19367 | w30216);
assign w30941 = v9736;
assign w30942 = w21837 & ~w22865;
assign w30943 = w15956 & ~pi23;
assign w30944 = ~w15956 & pi23;
assign w30945 = ~w20313 & w30300;
assign w30946 = w30301 | ~pi23;
assign w30947 = (~pi23 & w30301) | (~pi23 & w20313) | (w30301 & w20313);
assign w30948 = w23376 & w23037;
assign w30949 = w23376 & w23355;
assign v9737 = ~(w10543 | w10524);
assign w30950 = v9737;
assign w30951 = ~w15560 & w30575;
assign v9738 = ~(w15991 | w4764);
assign w30952 = v9738;
assign v9739 = ~(w17200 | w17216);
assign w30953 = v9739;
assign v9740 = ~(w23376 | w23037);
assign w30954 = v9740;
assign v9741 = ~(w23376 | w23355);
assign w30955 = v9741;
assign w30956 = w15563 & ~pi26;
assign w30957 = ~w15563 & pi26;
assign w30958 = ~w20924 & w30753;
assign w30959 = w30754 | ~pi26;
assign w30960 = (~pi26 & w30754) | (~pi26 & w20924) | (w30754 & w20924);
assign v9742 = ~(w21320 | w4764);
assign w30961 = v9742;
assign w30962 = w9510 & w9527;
assign w30963 = w3358 & ~w30577;
assign v9743 = ~(w3399 | w928);
assign w30964 = v9743;
assign v9744 = ~(w7318 | w3529);
assign w30965 = v9744;
assign v9745 = ~(w3763 | w3529);
assign w30966 = v9745;
assign w30967 = w7649 & ~pi26;
assign v9746 = ~(w15202 | w3529);
assign w30968 = v9746;
assign w30969 = w15539 & pi26;
assign v9747 = ~(w15598 | w4153);
assign w30970 = v9747;
assign w30971 = ~w16707 & w16724;
assign w30972 = ~w20275 & w30767;
assign v9748 = ~(w20416 | w4153);
assign w30973 = v9748;
assign w30974 = ~w3212 & w3760;
assign w30975 = ~w869 & w3763;
assign w30976 = (~w3529 & w3162) | (~w3529 & w31133) | (w3162 & w31133);
assign v9749 = ~(w15192 | w3529);
assign w30977 = v9749;
assign v9750 = ~(w20249 | w20243);
assign w30978 = v9750;
assign v9751 = ~(w20273 | pi26);
assign w30979 = v9751;
assign w30980 = w20273 & pi26;
assign v9752 = ~(w4153 | pi26);
assign w30981 = v9752;
assign w30982 = w4153 & pi26;
assign w30983 = w30750 & ~pi26;
assign w30984 = w20417 & ~pi26;
assign w30985 = ~w30750 & pi26;
assign v9753 = ~(w20601 | w3529);
assign w30986 = v9753;
assign w30987 = ~w3529 & pi29;
assign w30988 = w3529 & ~pi29;
assign w30989 = w21294 & ~pi29;
assign w30990 = ~w21294 & pi29;
assign w30991 = w21307 & ~pi26;
assign w30992 = w30755 & pi26;
assign w30993 = ~w21307 & pi26;
assign v9754 = ~(w21772 | w4153);
assign w30994 = v9754;
assign v9755 = ~(w22800 | w4153);
assign w30995 = v9755;
assign w30996 = (w30307 & w31245) | (w30307 & w31246) | (w31245 & w31246);
assign w30997 = (w3362 & w30785) | (w3362 & w30583) | (w30785 & w30583);
assign w30998 = w6645 & ~w6642;
assign w30999 = w6645 & w30786;
assign w31000 = (w3406 & ~w3179) | (w3406 & w31247) | (~w3179 & w31247);
assign w31001 = (w3402 & ~w3227) | (w3402 & w31134) | (~w3227 & w31134);
assign w31002 = (~w6672 & ~w6680) | (~w6672 & w31135) | (~w6680 & w31135);
assign w31003 = (~w6672 & ~w6680) | (~w6672 & w31248) | (~w6680 & w31248);
assign v9756 = ~(w928 | w6736);
assign w31004 = v9756;
assign v9757 = ~(pi29 | w7303);
assign w31005 = v9757;
assign v9758 = ~(pi29 | w30789);
assign w31006 = v9758;
assign w31007 = pi29 & w7303;
assign w31008 = pi29 & w30789;
assign w31009 = ~w3284 & w3767;
assign w31010 = ~w3193 & w3760;
assign w31011 = (pi29 & ~w7344) | (pi29 & w31136) | (~w7344 & w31136);
assign w31012 = (pi29 & ~w7344) | (pi29 & w31137) | (~w7344 & w31137);
assign w31013 = w7344 & w31138;
assign w31014 = ~pi29 & w7345;
assign v9759 = ~(w7348 | w7338);
assign w31015 = v9759;
assign w31016 = w7350 & ~w7323;
assign w31017 = ~w4153 & w7587;
assign w31018 = pi26 & w7599;
assign w31019 = pi26 & w30799;
assign v9760 = ~(pi26 | w7599);
assign w31020 = v9760;
assign v9761 = ~(pi26 | w30799);
assign w31021 = v9761;
assign v9762 = ~(w7672 | w7580);
assign w31022 = v9762;
assign v9763 = ~(w8045 | w7884);
assign w31023 = v9763;
assign v9764 = ~(w8446 | w8215);
assign w31024 = v9764;
assign v9765 = ~(w8617 | w8604);
assign w31025 = v9765;
assign w31026 = w9022 & ~w9021;
assign v9766 = ~(w9970 | w9972);
assign w31027 = v9766;
assign v9767 = ~(w10444 | w10982);
assign w31028 = v9767;
assign v9768 = ~(w11528 | w11030);
assign w31029 = v9768;
assign v9769 = ~(w28183 | w11765);
assign w31030 = v9769;
assign w31031 = ~w11787 & w28186;
assign v9770 = ~(w11787 | w11783);
assign w31032 = v9770;
assign w31033 = w28187 | ~w11821;
assign w31034 = (~w11821 & w28187) | (~w11821 & w11526) | (w28187 & w11526);
assign v9771 = ~(w11830 | w11764);
assign w31035 = v9771;
assign w31036 = w11830 & w11764;
assign v9772 = ~(pi29 | w30616);
assign w31037 = v9772;
assign v9773 = ~(pi29 | w15203);
assign w31038 = v9773;
assign w31039 = pi29 & w30616;
assign w31040 = pi29 & w15203;
assign w31041 = w15250 & ~w15218;
assign w31042 = ~w4153 & w15531;
assign v9774 = ~(w4153 | w15587);
assign w31043 = v9774;
assign v9775 = ~(w15626 | w15535);
assign w31044 = v9775;
assign v9776 = ~(w16035 | w15877);
assign w31045 = v9776;
assign w31046 = w16272 & ~w16271;
assign v9777 = ~(w16847 | w16910);
assign w31047 = v9777;
assign w31048 = w16695 & ~w16694;
assign v9778 = ~(w17449 | w17127);
assign w31049 = v9778;
assign w31050 = ~w17446 & w17624;
assign w31051 = ~w18015 & w17521;
assign w31052 = ~w18015 & w17523;
assign w31053 = w18015 & ~w17521;
assign w31054 = w18015 & ~w17523;
assign v9779 = ~(w18684 | w19210);
assign w31055 = v9779;
assign v9780 = ~(w19754 | w19753);
assign w31056 = v9780;
assign w31057 = ~w19754 & w19741;
assign v9781 = ~(w18035 | w19804);
assign w31058 = v9781;
assign w31059 = ~w30839 & pi26;
assign w31060 = ~w20253 & pi26;
assign v9782 = ~(w20268 | w20266);
assign w31061 = v9782;
assign w31062 = ~w20284 & w31139;
assign v9783 = ~(w3529 | w20405);
assign w31063 = v9783;
assign w31064 = w4155 & ~w28206;
assign w31065 = w4155 & w19782;
assign v9784 = ~(w20491 | w20579);
assign w31066 = v9784;
assign v9785 = ~(w20441 | w20439);
assign w31067 = v9785;
assign w31068 = pi29 & w30857;
assign w31069 = w20604 & w31140;
assign v9786 = ~(pi29 | w30857);
assign w31070 = v9786;
assign w31071 = (~pi29 & ~w20604) | (~pi29 & w31141) | (~w20604 & w31141);
assign v9787 = ~(w20744 | w20832);
assign w31072 = v9787;
assign v9788 = ~(w20650 | w20649);
assign w31073 = v9788;
assign w31074 = pi14 & w21075;
assign w31075 = pi14 & w29789;
assign v9789 = ~(pi14 | w21075);
assign w31076 = v9789;
assign v9790 = ~(pi14 | w29789);
assign w31077 = v9790;
assign v9791 = ~(w21120 | w21207);
assign w31078 = v9791;
assign v9792 = ~(w21223 | w21079);
assign w31079 = v9792;
assign v9793 = ~(w20977 | w20975);
assign w31080 = v9793;
assign w31081 = w20866 & ~w20917;
assign w31082 = pi11 & w21516;
assign w31083 = pi11 & w29793;
assign v9794 = ~(pi11 | w21516);
assign w31084 = v9794;
assign v9795 = ~(pi11 | w29793);
assign w31085 = v9795;
assign v9796 = ~(w21562 | w21650);
assign w31086 = v9796;
assign v9797 = ~(w21666 | w21520);
assign w31087 = v9797;
assign v9798 = ~(w21682 | w21476);
assign w31088 = v9798;
assign v9799 = ~(w21698 | w21425);
assign w31089 = v9799;
assign v9800 = ~(w21313 | w21311);
assign w31090 = v9800;
assign w31091 = w21258 & ~w21298;
assign w31092 = ~pi29 & w21760;
assign w31093 = w21760 & w31142;
assign w31094 = pi29 & ~w21760;
assign w31095 = (pi29 & ~w21760) | (pi29 & w31143) | (~w21760 & w31143);
assign w31096 = w30893 | w21787;
assign w31097 = (w21787 & w30893) | (w21787 & w20086) | (w30893 & w20086);
assign v9801 = ~(w20993 | w21373);
assign w31098 = v9801;
assign v9802 = ~(w22107 | w22194);
assign w31099 = v9802;
assign v9803 = ~(w22226 | w22021);
assign w31100 = v9803;
assign v9804 = ~(w22242 | w21970);
assign w31101 = v9804;
assign v9805 = ~(w21926 | w21911);
assign w31102 = v9805;
assign v9806 = ~(w22375 | w22722);
assign w31103 = v9806;
assign w31104 = w22786 & w31144;
assign w31105 = (~pi29 & ~w22786) | (~pi29 & w31145) | (~w22786 & w31145);
assign v9807 = ~(pi26 | w30898);
assign w31106 = v9807;
assign w31107 = (~pi26 & ~w22799) | (~pi26 & w31146) | (~w22799 & w31146);
assign w31108 = pi26 & w30898;
assign w31109 = w22799 & w31147;
assign w31110 = ~w4764 & w22814;
assign w31111 = w22991 & ~w22990;
assign w31112 = ~w23680 & w23570;
assign v9808 = ~(w23540 | w23537);
assign w31113 = v9808;
assign v9809 = ~(w23858 | w28087);
assign w31114 = v9809;
assign v9810 = ~(w24089 | w24087);
assign w31115 = v9810;
assign w31116 = w23909 & ~w23948;
assign v9811 = ~(w24192 | w24191);
assign w31117 = v9811;
assign v9812 = ~(w24160 | w24158);
assign w31118 = v9812;
assign v9813 = ~(w24429 | w24427);
assign w31119 = v9813;
assign w31120 = ~w20086 & w928;
assign v9814 = ~(w428 | w239);
assign w31121 = v9814;
assign v9815 = ~(w19256 | w19254);
assign w31122 = v9815;
assign w31123 = w19256 & w19254;
assign v9816 = ~(w20240 | w21722);
assign w31124 = v9816;
assign v9817 = ~(w20083 | pi17);
assign w31125 = v9817;
assign w31126 = w20083 & pi17;
assign w31127 = w30964 & ~w928;
assign w31128 = (~w928 & w30964) | (~w928 & w3284) | (w30964 & w3284);
assign w31129 = ~w20603 & w30986;
assign v9818 = ~(w30755 | pi26);
assign w31130 = v9818;
assign w31131 = w21786 & ~w4764;
assign w31132 = ~w22797 & w30995;
assign v9819 = ~(w3760 | w3529);
assign w31133 = v9819;
assign w31134 = ~w3212 & w3402;
assign v9820 = ~(w30585 | w6672);
assign w31135 = v9820;
assign w31136 = ~w30976 & pi29;
assign w31137 = w7341 & pi29;
assign w31138 = w30976 & ~pi29;
assign v9821 = ~(w20285 | w20282);
assign w31139 = v9821;
assign w31140 = ~w20601 & pi29;
assign w31141 = w20601 & ~pi29;
assign v9822 = ~(w3529 | pi29);
assign w31142 = v9822;
assign w31143 = w3529 & pi29;
assign w31144 = ~w22787 & pi29;
assign w31145 = w22787 & ~pi29;
assign w31146 = w22800 & ~pi26;
assign w31147 = ~w22800 & pi26;
assign v9823 = ~(w428 | w812);
assign w31148 = v9823;
assign w31149 = w855 & w2460;
assign w31150 = w2502 & w846;
assign w31151 = w2494 & ~w291;
assign w31152 = w1469 & w1103;
assign w31153 = w2560 & w1344;
assign v9824 = ~(w652 | w303);
assign w31154 = v9824;
assign w31155 = w3180 & ~w630;
assign w31156 = w28472 & w3190;
assign w31157 = w2493 & w3366;
assign w31158 = ~w928 & w6608;
assign v9825 = ~(w6639 | w30999);
assign w31159 = v9825;
assign v9826 = ~(w6639 | w30998);
assign w31160 = v9826;
assign w31161 = ~w3284 & w3399;
assign w31162 = w6739 & ~w6736;
assign w31163 = w6739 & w31004;
assign w31164 = w6740 & ~w6729;
assign w31165 = w6639 & w30999;
assign w31166 = w6639 & w30998;
assign w31167 = ~w3529 & w7291;
assign w31168 = ~w3228 & w3767;
assign w31169 = ~w3193 & w3763;
assign v9827 = ~(w7360 | w7296);
assign w31170 = v9827;
assign v9828 = ~(w7680 | w7554);
assign w31171 = v9828;
assign v9829 = ~(w8053 | w7858);
assign w31172 = v9829;
assign v9830 = ~(w8454 | w8189);
assign w31173 = v9830;
assign w31174 = w8590 & ~w8589;
assign w31175 = (w30615 & w30614) | (w30615 & w30163) | (w30614 & w30163);
assign w31176 = (w30615 & w30614) | (w30615 & w30162) | (w30614 & w30162);
assign w31177 = pi29 & w30809;
assign w31178 = w15191 & w31249;
assign v9831 = ~(pi29 | w30809);
assign w31179 = v9831;
assign w31180 = (~pi29 & ~w15191) | (~pi29 & w31250) | (~w15191 & w31250);
assign w31181 = w15225 & ~w15221;
assign v9832 = ~(w3529 | w15229);
assign w31182 = v9832;
assign w31183 = ~w15245 & pi29;
assign w31184 = w15245 & ~pi29;
assign v9833 = ~(w15260 | w15196);
assign w31185 = v9833;
assign w31186 = ~w4153 & w15519;
assign w31187 = ~pi26 & w15531;
assign w31188 = ~pi26 & w31042;
assign w31189 = pi26 & ~w15531;
assign w31190 = pi26 & ~w31042;
assign v9834 = ~(w15634 | w15512);
assign w31191 = v9834;
assign w31192 = w15864 & ~w15863;
assign v9835 = ~(w16256 | w16241);
assign w31193 = v9835;
assign w31194 = w16679 & ~w16678;
assign w31195 = w17109 & ~w17108;
assign v9836 = ~(w17582 | w17992);
assign w31196 = v9836;
assign v9837 = ~(w18091 | w18093);
assign w31197 = v9837;
assign v9838 = ~(w18654 | w19216);
assign w31198 = v9838;
assign v9839 = ~(w19793 | w19230);
assign w31199 = v9839;
assign w31200 = w20081 & w20015;
assign w31201 = w20081 & w20017;
assign w31202 = ~w31062 & pi29;
assign w31203 = ~w20404 & pi29;
assign v9840 = ~(w20600 | w20598);
assign w31204 = v9840;
assign w31205 = w21397 & ~w21396;
assign w31206 = w21705 & ~w21379;
assign w31207 = w21771 & w31251;
assign w31208 = w21771 & w31252;
assign w31209 = (~pi26 & ~w21771) | (~pi26 & w31253) | (~w21771 & w31253);
assign v9841 = ~(pi26 | w21773);
assign w31210 = v9841;
assign w31211 = ~pi23 & w31096;
assign w31212 = ~pi23 & w20638;
assign w31213 = pi23 & ~w31096;
assign w31214 = pi23 & ~w20638;
assign v9842 = ~(w21895 | w21893);
assign w31215 = v9842;
assign v9843 = ~(w22296 | w22298);
assign w31216 = v9843;
assign w31217 = pi29 & ~w23453;
assign w31218 = (pi29 & ~w23453) | (pi29 & w31143) | (~w23453 & w31143);
assign w31219 = ~pi29 & w23453;
assign w31220 = w23453 & w31142;
assign v9844 = ~(w24241 | w24238);
assign w31221 = v9844;
assign w31222 = w24248 & ~w24245;
assign w31223 = w24507 & ~w24506;
assign w31224 = ~w24901 & w24697;
assign w31225 = ~w24901 & w24516;
assign w31226 = w24901 & ~w24697;
assign w31227 = w24901 & ~w24516;
assign v9845 = ~(w24780 | w24778);
assign w31228 = v9845;
assign w31229 = w20638 & w24959;
assign w31230 = ~w10432 & w10431;
assign w31231 = ~w10432 & w11535;
assign w31232 = w11042 & w11029;
assign w31233 = w24276 & ~w24497;
assign v9846 = ~(w8957 | w28184);
assign w31234 = v9846;
assign v9847 = ~(w8957 | w28185);
assign w31235 = v9847;
assign w31236 = (~w8541 & w28999) | (~w8541 & w28184) | (w28999 & w28184);
assign w31237 = (~w8541 & w28999) | (~w8541 & w28185) | (w28999 & w28185);
assign w31238 = ~w23033 & w30718;
assign v9848 = ~(w23033 | w30277);
assign w31239 = v9848;
assign w31240 = ~w23015 & w23033;
assign w31241 = w24131 & ~w24019;
assign v9849 = ~(w23716 | w23905);
assign w31242 = v9849;
assign w31243 = ~w15189 & w30977;
assign v9850 = ~(w23755 | w3529);
assign w31244 = v9850;
assign w31245 = (w3362 & w30785) | (w3362 & w3358) | (w30785 & w3358);
assign w31246 = (w3362 & w30785) | (w3362 & w30757) | (w30785 & w30757);
assign w31247 = ~w3192 & w3406;
assign w31248 = w6677 & ~w6672;
assign w31249 = ~w15192 & pi29;
assign w31250 = w15192 & ~pi29;
assign w31251 = w30994 & pi26;
assign w31252 = ~w21772 & pi26;
assign v9851 = ~(w30994 | pi26);
assign w31253 = v9851;
assign v9852 = ~(w2425 | w3366);
assign w31254 = v9852;
assign v9853 = ~(w2425 | w31157);
assign w31255 = v9853;
assign v9854 = ~(w6599 | w6608);
assign w31256 = v9854;
assign v9855 = ~(w6599 | w31158);
assign w31257 = v9855;
assign w31258 = ~w6728 & w31003;
assign w31259 = ~w6728 & w31002;
assign w31260 = w6728 & ~w31003;
assign w31261 = w6728 & ~w31002;
assign w31262 = w6599 & w6608;
assign w31263 = w6599 & w31158;
assign v9856 = ~(w6748 | w6609);
assign w31264 = v9856;
assign w31265 = (w9420 & w28317) | (w9420 & w28184) | (w28317 & w28184);
assign w31266 = (w9420 & w28317) | (w9420 & w28185) | (w28317 & w28185);
assign w31267 = w28507 & ~w28184;
assign w31268 = w28507 & ~w28185;
assign w31269 = ~w28321 & w11838;
assign v9857 = ~(w928 | w14505);
assign w31270 = v9857;
assign v9858 = ~(w928 | w14548);
assign w31271 = v9858;
assign v9859 = ~(w928 | w14570);
assign w31272 = v9859;
assign w31273 = ~w3529 & w15169;
assign w31274 = w15182 & pi29;
assign v9860 = ~(w15182 | pi29);
assign w31275 = v9860;
assign v9861 = ~(w15264 | w15186);
assign w31276 = v9861;
assign v9862 = ~(w15638 | w15499);
assign w31277 = v9862;
assign v9863 = ~(w15848 | w15835);
assign w31278 = v9863;
assign w31279 = w16649 & ~w16648;
assign w31280 = w19804 & ~w19797;
assign w31281 = w19804 & w29039;
assign w31282 = (w30837 & w30836) | (w30837 & ~w30373) | (w30836 & ~w30373);
assign w31283 = (w30837 & w30836) | (w30837 & ~w30374) | (w30836 & ~w30374);
assign w31284 = ~w19804 & w19797;
assign v9864 = ~(w19804 | w29039);
assign w31285 = v9864;
assign w31286 = w20085 & w20012;
assign w31287 = w20085 & ~w28564;
assign v9865 = ~(w21744 | w21749);
assign w31288 = v9865;
assign v9866 = ~(w21744 | w30699);
assign w31289 = v9866;
assign w31290 = w21744 & w21749;
assign w31291 = w21744 & w30699;
assign v9867 = ~(w4155 | w21770);
assign w31292 = v9867;
assign w31293 = ~w928 & w22775;
assign w31294 = ~pi23 & w22814;
assign w31295 = ~pi23 & w31110;
assign w31296 = pi23 & ~w22814;
assign w31297 = pi23 & ~w31110;
assign w31298 = w22975 & ~w22974;
assign w31299 = pi29 & w30902;
assign w31300 = pi29 & w23756;
assign v9868 = ~(pi29 | w30902);
assign w31301 = v9868;
assign v9869 = ~(pi29 | w23756);
assign w31302 = v9869;
assign w31303 = ~w3529 & w23943;
assign w31304 = ~w4153 & w23958;
assign w31305 = (w28104 & w28103) | (w28104 & ~w28607) | (w28103 & ~w28607);
assign w31306 = (w28104 & w28103) | (w28104 & ~w28608) | (w28103 & ~w28608);
assign v9870 = ~(w26442 | w28865);
assign w31307 = v9870;
assign v9871 = ~(w26442 | w28864);
assign w31308 = v9871;
assign w31309 = w26442 & w28865;
assign w31310 = w26442 & w28864;
assign w31311 = ~w27669 & w27584;
assign v9872 = ~(w27669 | w28255);
assign w31312 = v9872;
assign w31313 = w27669 & ~w27584;
assign w31314 = w27669 & w28255;
assign w31315 = w28134 & w27750;
assign v9873 = ~(w28134 | w27750);
assign w31316 = v9873;
assign w31317 = w28258 | ~w27824;
assign w31318 = (~w27824 & w28258) | (~w27824 & ~w28134) | (w28258 & ~w28134);
assign w31319 = w28134 & w28137;
assign w31320 = w28134 & w28139;
assign w31321 = w28259 | w27891;
assign w31322 = (w27891 & w28259) | (w27891 & ~w28134) | (w28259 & ~w28134);
assign w31323 = w28260 | ~w27943;
assign w31324 = (~w27943 & w28260) | (~w27943 & ~w28134) | (w28260 & ~w28134);
assign w31325 = w28134 & w28141;
assign one = 1;
assign po00 = w23631;// level 183
assign po01 = w23873;// level 185
assign po02 = w24096;// level 186
assign po03 = w24302;// level 188
assign po04 = w24515;// level 189
assign po05 = w24705;// level 190
assign po06 = w24907;// level 191
assign po07 = w25097;// level 192
assign po08 = w25284;// level 193
assign po09 = w25461;// level 194
assign po10 = w25636;// level 195
assign po11 = w25815;// level 196
assign po12 = w25991;// level 197
assign po13 = w26156;// level 197
assign po14 = w26305;// level 199
assign po15 = w26449;// level 198
assign po16 = w26591;// level 198
assign po17 = w26723;// level 199
assign po18 = w26850;// level 200
assign po19 = w26973;// level 200
assign po20 = w27087;// level 200
assign po21 = w27198;// level 200
assign po22 = w27304;// level 200
assign po23 = w27401;// level 200
assign po24 = w27492;// level 200
assign po25 = w27590;// level 200
assign po26 = w27672;// level 200
assign po27 = w27753;// level 200
assign po28 = w27827;// level 200
assign po29 = w27894;// level 200
assign po30 = w27946;// level 200
assign po31 = ~w27991;// level 201
endmodule
