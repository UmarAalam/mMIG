// Benchmark "sqrt32" written by ABC on Wed Apr 29 17:20:33 2015

module sqrt32 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15;
  wire n50, n51, n52, n53, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
    n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
    n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
    n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n783, n784, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
    n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
    n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160;
  assign po15 = pi30 | pi31;
  assign n50 = ~pi28 & ~pi29;
  assign n51 = pi30 & ~n50;
  assign n52 = ~n50 & ~n51;
  assign n53 = pi30 & pi31;
  assign po14 = n52 | n53;
  assign n55 = ~pi26 & ~pi27;
  assign n56 = po14 & n55;
  assign n57 = pi28 & ~po14;
  assign n58 = ~pi28 & po14;
  assign n59 = ~n57 & ~n58;
  assign n60 = ~po14 & ~n55;
  assign n61 = ~n56 & ~n60;
  assign n62 = n59 & n61;
  assign n63 = ~n56 & ~n62;
  assign n64 = po15 & ~n63;
  assign n65 = ~po15 & n63;
  assign n66 = ~n64 & ~n65;
  assign n67 = pi29 & ~n58;
  assign n68 = n50 & po14;
  assign n69 = ~n67 & ~n68;
  assign n70 = n66 & n69;
  assign n71 = ~po15 & ~n70;
  assign n72 = ~pi30 & n50;
  assign n73 = po15 & n72;
  assign n74 = ~n71 & ~n73;
  assign n75 = n63 & ~n70;
  assign n76 = n51 & po14;
  assign n77 = ~n75 & ~n76;
  assign po13 = ~n74 | ~n77;
  assign n79 = n70 & po13;
  assign n80 = ~pi24 & ~pi25;
  assign n81 = po13 & n80;
  assign n82 = pi26 & ~po13;
  assign n83 = ~pi26 & po13;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~po13 & ~n80;
  assign n86 = ~n81 & ~n85;
  assign n87 = n84 & n86;
  assign n88 = ~n81 & ~n87;
  assign n89 = po14 & ~n88;
  assign n90 = ~po14 & n88;
  assign n91 = ~n89 & ~n90;
  assign n92 = pi27 & ~n83;
  assign n93 = n55 & po13;
  assign n94 = ~n92 & ~n93;
  assign n95 = n91 & n94;
  assign n96 = ~n89 & ~n95;
  assign n97 = po15 & ~n96;
  assign n98 = ~po15 & n96;
  assign n99 = ~n97 & ~n98;
  assign n100 = n61 & po13;
  assign n101 = ~n59 & ~n100;
  assign n102 = n62 & po13;
  assign n103 = ~n101 & ~n102;
  assign n104 = n99 & n103;
  assign n105 = ~n97 & ~n104;
  assign n106 = n64 & ~n69;
  assign n107 = ~n105 & ~n106;
  assign po12 = n79 | ~n107;
  assign n109 = n104 & po12;
  assign n110 = ~pi22 & ~pi23;
  assign n111 = po12 & n110;
  assign n112 = pi24 & ~po12;
  assign n113 = ~pi24 & po12;
  assign n114 = ~n112 & ~n113;
  assign n115 = ~po12 & ~n110;
  assign n116 = ~n111 & ~n115;
  assign n117 = n114 & n116;
  assign n118 = ~n111 & ~n117;
  assign n119 = po13 & ~n118;
  assign n120 = ~po13 & n118;
  assign n121 = ~n119 & ~n120;
  assign n122 = pi25 & ~n113;
  assign n123 = n80 & po12;
  assign n124 = ~n122 & ~n123;
  assign n125 = n121 & n124;
  assign n126 = ~n119 & ~n125;
  assign n127 = po14 & ~n126;
  assign n128 = ~po14 & n126;
  assign n129 = ~n127 & ~n128;
  assign n130 = n86 & po12;
  assign n131 = ~n84 & ~n130;
  assign n132 = n87 & po12;
  assign n133 = ~n131 & ~n132;
  assign n134 = n129 & n133;
  assign n135 = ~n127 & ~n134;
  assign n136 = po15 & ~n135;
  assign n137 = ~po15 & n135;
  assign n138 = ~n136 & ~n137;
  assign n139 = n91 & po12;
  assign n140 = ~n94 & ~n139;
  assign n141 = n95 & po12;
  assign n142 = ~n140 & ~n141;
  assign n143 = n138 & n142;
  assign n144 = ~n136 & ~n143;
  assign n145 = po15 & ~n103;
  assign n146 = ~n96 & n145;
  assign n147 = ~n144 & ~n146;
  assign po11 = n109 | ~n147;
  assign n149 = n143 & po11;
  assign n150 = ~pi20 & ~pi21;
  assign n151 = po11 & n150;
  assign n152 = pi22 & ~po11;
  assign n153 = ~pi22 & po11;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~po11 & ~n150;
  assign n156 = ~n151 & ~n155;
  assign n157 = n154 & n156;
  assign n158 = ~n151 & ~n157;
  assign n159 = po12 & ~n158;
  assign n160 = ~po12 & n158;
  assign n161 = ~n159 & ~n160;
  assign n162 = pi23 & ~n153;
  assign n163 = n110 & po11;
  assign n164 = ~n162 & ~n163;
  assign n165 = n161 & n164;
  assign n166 = ~n159 & ~n165;
  assign n167 = po13 & ~n166;
  assign n168 = ~po13 & n166;
  assign n169 = ~n167 & ~n168;
  assign n170 = n116 & po11;
  assign n171 = ~n114 & ~n170;
  assign n172 = n117 & po11;
  assign n173 = ~n171 & ~n172;
  assign n174 = n169 & n173;
  assign n175 = ~n167 & ~n174;
  assign n176 = po14 & ~n175;
  assign n177 = ~po14 & n175;
  assign n178 = ~n176 & ~n177;
  assign n179 = n121 & po11;
  assign n180 = ~n124 & ~n179;
  assign n181 = n125 & po11;
  assign n182 = ~n180 & ~n181;
  assign n183 = n178 & n182;
  assign n184 = ~n176 & ~n183;
  assign n185 = po15 & ~n184;
  assign n186 = ~po15 & n184;
  assign n187 = ~n185 & ~n186;
  assign n188 = n129 & po11;
  assign n189 = ~n133 & ~n188;
  assign n190 = n134 & po11;
  assign n191 = ~n189 & ~n190;
  assign n192 = n187 & n191;
  assign n193 = ~n185 & ~n192;
  assign n194 = po15 & ~n142;
  assign n195 = ~n135 & n194;
  assign n196 = ~n193 & ~n195;
  assign po10 = n149 | ~n196;
  assign n198 = ~pi18 & ~pi19;
  assign n199 = po10 & n198;
  assign n200 = pi20 & ~po10;
  assign n201 = ~pi20 & po10;
  assign n202 = ~n200 & ~n201;
  assign n203 = ~po10 & ~n198;
  assign n204 = ~n199 & ~n203;
  assign n205 = n202 & n204;
  assign n206 = ~n199 & ~n205;
  assign n207 = po11 & ~n206;
  assign n208 = ~po11 & n206;
  assign n209 = ~n207 & ~n208;
  assign n210 = pi21 & ~n201;
  assign n211 = n150 & po10;
  assign n212 = ~n210 & ~n211;
  assign n213 = n209 & n212;
  assign n214 = ~n207 & ~n213;
  assign n215 = po12 & ~n214;
  assign n216 = ~po12 & n214;
  assign n217 = ~n215 & ~n216;
  assign n218 = n156 & po10;
  assign n219 = ~n154 & ~n218;
  assign n220 = n157 & po10;
  assign n221 = ~n219 & ~n220;
  assign n222 = n217 & n221;
  assign n223 = ~n215 & ~n222;
  assign n224 = po13 & ~n223;
  assign n225 = ~po13 & n223;
  assign n226 = ~n224 & ~n225;
  assign n227 = n161 & po10;
  assign n228 = ~n164 & ~n227;
  assign n229 = n165 & po10;
  assign n230 = ~n228 & ~n229;
  assign n231 = n226 & n230;
  assign n232 = ~n224 & ~n231;
  assign n233 = po14 & ~n232;
  assign n234 = ~po14 & n232;
  assign n235 = ~n233 & ~n234;
  assign n236 = n169 & po10;
  assign n237 = ~n173 & ~n236;
  assign n238 = n174 & po10;
  assign n239 = ~n237 & ~n238;
  assign n240 = n235 & n239;
  assign n241 = ~n233 & ~n240;
  assign n242 = po15 & ~n241;
  assign n243 = ~po15 & n241;
  assign n244 = ~n242 & ~n243;
  assign n245 = n178 & po10;
  assign n246 = ~n182 & ~n245;
  assign n247 = n183 & po10;
  assign n248 = ~n246 & ~n247;
  assign n249 = n244 & n248;
  assign n250 = n192 & po10;
  assign n251 = ~n242 & ~n249;
  assign n252 = ~n187 & ~n191;
  assign n253 = ~n251 & ~n252;
  assign po09 = n250 | ~n253;
  assign n255 = n249 & po09;
  assign n256 = ~pi16 & ~pi17;
  assign n257 = po09 & n256;
  assign n258 = pi18 & ~po09;
  assign n259 = ~pi18 & po09;
  assign n260 = ~n258 & ~n259;
  assign n261 = ~po09 & ~n256;
  assign n262 = ~n257 & ~n261;
  assign n263 = n260 & n262;
  assign n264 = ~n257 & ~n263;
  assign n265 = po10 & ~n264;
  assign n266 = ~po10 & n264;
  assign n267 = ~n265 & ~n266;
  assign n268 = pi19 & ~n259;
  assign n269 = n198 & po09;
  assign n270 = ~n268 & ~n269;
  assign n271 = n267 & n270;
  assign n272 = ~n265 & ~n271;
  assign n273 = po11 & ~n272;
  assign n274 = ~po11 & n272;
  assign n275 = ~n273 & ~n274;
  assign n276 = n204 & po09;
  assign n277 = ~n202 & ~n276;
  assign n278 = n205 & po09;
  assign n279 = ~n277 & ~n278;
  assign n280 = n275 & n279;
  assign n281 = ~n273 & ~n280;
  assign n282 = po12 & ~n281;
  assign n283 = ~po12 & n281;
  assign n284 = ~n282 & ~n283;
  assign n285 = n209 & po09;
  assign n286 = ~n212 & ~n285;
  assign n287 = n213 & po09;
  assign n288 = ~n286 & ~n287;
  assign n289 = n284 & n288;
  assign n290 = ~n282 & ~n289;
  assign n291 = po13 & ~n290;
  assign n292 = ~po13 & n290;
  assign n293 = ~n291 & ~n292;
  assign n294 = n217 & po09;
  assign n295 = ~n221 & ~n294;
  assign n296 = n222 & po09;
  assign n297 = ~n295 & ~n296;
  assign n298 = n293 & n297;
  assign n299 = ~n291 & ~n298;
  assign n300 = po14 & ~n299;
  assign n301 = ~po14 & n299;
  assign n302 = ~n300 & ~n301;
  assign n303 = n226 & po09;
  assign n304 = ~n230 & ~n303;
  assign n305 = n231 & po09;
  assign n306 = ~n304 & ~n305;
  assign n307 = n302 & n306;
  assign n308 = ~n300 & ~n307;
  assign n309 = po15 & ~n308;
  assign n310 = ~po15 & n308;
  assign n311 = ~n309 & ~n310;
  assign n312 = n235 & po09;
  assign n313 = ~n239 & ~n312;
  assign n314 = n240 & po09;
  assign n315 = ~n313 & ~n314;
  assign n316 = n311 & n315;
  assign n317 = ~n309 & ~n316;
  assign n318 = ~n244 & ~n248;
  assign n319 = ~n317 & ~n318;
  assign po08 = n255 | ~n319;
  assign n321 = pi16 & ~po08;
  assign n322 = ~pi16 & po08;
  assign n323 = ~n321 & ~n322;
  assign n324 = ~pi14 & ~pi15;
  assign n325 = po08 & n324;
  assign n326 = ~po08 & ~n324;
  assign n327 = ~n325 & ~n326;
  assign n328 = n316 & po08;
  assign n329 = n323 & n327;
  assign n330 = ~n325 & ~n329;
  assign n331 = po09 & ~n330;
  assign n332 = ~po09 & n330;
  assign n333 = ~n331 & ~n332;
  assign n334 = pi17 & ~n322;
  assign n335 = n256 & po08;
  assign n336 = ~n334 & ~n335;
  assign n337 = n333 & n336;
  assign n338 = ~n331 & ~n337;
  assign n339 = po10 & ~n338;
  assign n340 = ~po10 & n338;
  assign n341 = ~n339 & ~n340;
  assign n342 = n262 & po08;
  assign n343 = ~n260 & ~n342;
  assign n344 = n263 & po08;
  assign n345 = ~n343 & ~n344;
  assign n346 = n341 & n345;
  assign n347 = ~n339 & ~n346;
  assign n348 = po11 & ~n347;
  assign n349 = ~po11 & n347;
  assign n350 = ~n348 & ~n349;
  assign n351 = n267 & po08;
  assign n352 = ~n270 & ~n351;
  assign n353 = n271 & po08;
  assign n354 = ~n352 & ~n353;
  assign n355 = n350 & n354;
  assign n356 = ~n348 & ~n355;
  assign n357 = po12 & ~n356;
  assign n358 = ~po12 & n356;
  assign n359 = ~n357 & ~n358;
  assign n360 = n275 & po08;
  assign n361 = ~n279 & ~n360;
  assign n362 = n280 & po08;
  assign n363 = ~n361 & ~n362;
  assign n364 = n359 & n363;
  assign n365 = ~n357 & ~n364;
  assign n366 = po13 & ~n365;
  assign n367 = ~po13 & n365;
  assign n368 = ~n366 & ~n367;
  assign n369 = n284 & po08;
  assign n370 = ~n288 & ~n369;
  assign n371 = n289 & po08;
  assign n372 = ~n370 & ~n371;
  assign n373 = n368 & n372;
  assign n374 = ~n366 & ~n373;
  assign n375 = po14 & ~n374;
  assign n376 = ~po14 & n374;
  assign n377 = ~n375 & ~n376;
  assign n378 = n293 & po08;
  assign n379 = ~n297 & ~n378;
  assign n380 = n298 & po08;
  assign n381 = ~n379 & ~n380;
  assign n382 = n377 & n381;
  assign n383 = ~n375 & ~n382;
  assign n384 = po15 & ~n383;
  assign n385 = ~po15 & n383;
  assign n386 = ~n384 & ~n385;
  assign n387 = n302 & po08;
  assign n388 = ~n306 & ~n387;
  assign n389 = n307 & po08;
  assign n390 = ~n388 & ~n389;
  assign n391 = n386 & n390;
  assign n392 = ~n384 & ~n391;
  assign n393 = ~n311 & ~n315;
  assign n394 = ~n392 & ~n393;
  assign po07 = n328 | ~n394;
  assign n396 = n327 & po07;
  assign n397 = ~n323 & ~n396;
  assign n398 = n329 & po07;
  assign n399 = ~n397 & ~n398;
  assign n400 = ~pi12 & ~pi13;
  assign n401 = po07 & n400;
  assign n402 = pi14 & ~po07;
  assign n403 = ~pi14 & po07;
  assign n404 = ~n402 & ~n403;
  assign n405 = ~po07 & ~n400;
  assign n406 = ~n401 & ~n405;
  assign n407 = n404 & n406;
  assign n408 = ~n401 & ~n407;
  assign n409 = po08 & ~n408;
  assign n410 = ~po08 & n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = pi15 & ~n403;
  assign n413 = n324 & po07;
  assign n414 = ~n412 & ~n413;
  assign n415 = n411 & n414;
  assign n416 = ~n409 & ~n415;
  assign n417 = po09 & ~n416;
  assign n418 = ~po09 & n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = n391 & po07;
  assign n421 = n399 & n419;
  assign n422 = ~n417 & ~n421;
  assign n423 = po10 & ~n422;
  assign n424 = ~po10 & n422;
  assign n425 = ~n423 & ~n424;
  assign n426 = n333 & po07;
  assign n427 = ~n336 & ~n426;
  assign n428 = n337 & po07;
  assign n429 = ~n427 & ~n428;
  assign n430 = n425 & n429;
  assign n431 = ~n423 & ~n430;
  assign n432 = po11 & ~n431;
  assign n433 = ~po11 & n431;
  assign n434 = ~n432 & ~n433;
  assign n435 = n341 & po07;
  assign n436 = ~n345 & ~n435;
  assign n437 = n346 & po07;
  assign n438 = ~n436 & ~n437;
  assign n439 = n434 & n438;
  assign n440 = ~n432 & ~n439;
  assign n441 = po12 & ~n440;
  assign n442 = ~po12 & n440;
  assign n443 = ~n441 & ~n442;
  assign n444 = n350 & po07;
  assign n445 = ~n354 & ~n444;
  assign n446 = n355 & po07;
  assign n447 = ~n445 & ~n446;
  assign n448 = n443 & n447;
  assign n449 = ~n441 & ~n448;
  assign n450 = po13 & ~n449;
  assign n451 = ~po13 & n449;
  assign n452 = ~n450 & ~n451;
  assign n453 = n359 & po07;
  assign n454 = ~n363 & ~n453;
  assign n455 = n364 & po07;
  assign n456 = ~n454 & ~n455;
  assign n457 = n452 & n456;
  assign n458 = ~n450 & ~n457;
  assign n459 = po14 & ~n458;
  assign n460 = ~po14 & n458;
  assign n461 = ~n459 & ~n460;
  assign n462 = n368 & po07;
  assign n463 = ~n372 & ~n462;
  assign n464 = n373 & po07;
  assign n465 = ~n463 & ~n464;
  assign n466 = n461 & n465;
  assign n467 = ~n459 & ~n466;
  assign n468 = po15 & ~n467;
  assign n469 = ~po15 & n467;
  assign n470 = ~n468 & ~n469;
  assign n471 = n377 & po07;
  assign n472 = ~n381 & ~n471;
  assign n473 = n382 & po07;
  assign n474 = ~n472 & ~n473;
  assign n475 = n470 & n474;
  assign n476 = ~n468 & ~n475;
  assign n477 = ~n386 & ~n390;
  assign n478 = ~n476 & ~n477;
  assign po06 = n420 | ~n478;
  assign n480 = n419 & po06;
  assign n481 = ~n399 & ~n480;
  assign n482 = n421 & po06;
  assign n483 = ~n481 & ~n482;
  assign n484 = ~pi10 & ~pi11;
  assign n485 = ~n476 & n484;
  assign n486 = pi12 & ~po06;
  assign n487 = ~pi12 & po06;
  assign n488 = ~n486 & ~n487;
  assign n489 = n476 & ~n484;
  assign n490 = ~n485 & ~n489;
  assign n491 = n488 & n490;
  assign n492 = ~n485 & ~n491;
  assign n493 = ~n392 & ~n492;
  assign n494 = n392 & n492;
  assign n495 = ~n493 & ~n494;
  assign n496 = pi13 & ~n487;
  assign n497 = n400 & po06;
  assign n498 = ~n496 & ~n497;
  assign n499 = n495 & n498;
  assign n500 = ~n493 & ~n499;
  assign n501 = po08 & ~n500;
  assign n502 = ~po08 & n500;
  assign n503 = ~n501 & ~n502;
  assign n504 = n406 & po06;
  assign n505 = ~n404 & ~n504;
  assign n506 = n407 & po06;
  assign n507 = ~n505 & ~n506;
  assign n508 = n503 & n507;
  assign n509 = ~n501 & ~n508;
  assign n510 = po09 & ~n509;
  assign n511 = ~po09 & n509;
  assign n512 = ~n510 & ~n511;
  assign n513 = n411 & po06;
  assign n514 = ~n414 & ~n513;
  assign n515 = n415 & po06;
  assign n516 = ~n514 & ~n515;
  assign n517 = n512 & n516;
  assign n518 = ~n510 & ~n517;
  assign n519 = po10 & ~n518;
  assign n520 = ~po10 & n518;
  assign n521 = ~n519 & ~n520;
  assign n522 = n475 & po06;
  assign n523 = n483 & n521;
  assign n524 = ~n519 & ~n523;
  assign n525 = po11 & ~n524;
  assign n526 = ~po11 & n524;
  assign n527 = ~n525 & ~n526;
  assign n528 = n425 & po06;
  assign n529 = ~n429 & ~n528;
  assign n530 = n430 & po06;
  assign n531 = ~n529 & ~n530;
  assign n532 = n527 & n531;
  assign n533 = ~n525 & ~n532;
  assign n534 = po12 & ~n533;
  assign n535 = ~po12 & n533;
  assign n536 = ~n534 & ~n535;
  assign n537 = n434 & po06;
  assign n538 = ~n438 & ~n537;
  assign n539 = n439 & po06;
  assign n540 = ~n538 & ~n539;
  assign n541 = n536 & n540;
  assign n542 = ~n534 & ~n541;
  assign n543 = po13 & ~n542;
  assign n544 = ~po13 & n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = n443 & po06;
  assign n547 = ~n447 & ~n546;
  assign n548 = n448 & po06;
  assign n549 = ~n547 & ~n548;
  assign n550 = n545 & n549;
  assign n551 = ~n543 & ~n550;
  assign n552 = po14 & ~n551;
  assign n553 = ~po14 & n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = n452 & po06;
  assign n556 = ~n456 & ~n555;
  assign n557 = n457 & po06;
  assign n558 = ~n556 & ~n557;
  assign n559 = n554 & n558;
  assign n560 = ~n552 & ~n559;
  assign n561 = po15 & ~n560;
  assign n562 = ~po15 & n560;
  assign n563 = ~n561 & ~n562;
  assign n564 = n461 & po06;
  assign n565 = ~n465 & ~n564;
  assign n566 = n466 & po06;
  assign n567 = ~n565 & ~n566;
  assign n568 = n563 & n567;
  assign n569 = ~n561 & ~n568;
  assign n570 = ~n470 & ~n474;
  assign n571 = ~n569 & ~n570;
  assign po05 = n522 | ~n571;
  assign n573 = n521 & po05;
  assign n574 = ~n483 & ~n573;
  assign n575 = n523 & po05;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~pi08 & ~pi09;
  assign n578 = po05 & n577;
  assign n579 = pi10 & ~po05;
  assign n580 = ~pi10 & po05;
  assign n581 = ~n579 & ~n580;
  assign n582 = ~po05 & ~n577;
  assign n583 = ~n578 & ~n582;
  assign n584 = n581 & n583;
  assign n585 = ~n578 & ~n584;
  assign n586 = po06 & ~n585;
  assign n587 = ~po06 & n585;
  assign n588 = ~n586 & ~n587;
  assign n589 = pi11 & ~n580;
  assign n590 = n484 & po05;
  assign n591 = ~n589 & ~n590;
  assign n592 = n588 & n591;
  assign n593 = ~n586 & ~n592;
  assign n594 = po07 & ~n593;
  assign n595 = ~po07 & n593;
  assign n596 = ~n594 & ~n595;
  assign n597 = n490 & po05;
  assign n598 = ~n488 & ~n597;
  assign n599 = n491 & po05;
  assign n600 = ~n598 & ~n599;
  assign n601 = n596 & n600;
  assign n602 = ~n594 & ~n601;
  assign n603 = po08 & ~n602;
  assign n604 = ~po08 & n602;
  assign n605 = ~n603 & ~n604;
  assign n606 = n495 & po05;
  assign n607 = ~n498 & ~n606;
  assign n608 = n499 & po05;
  assign n609 = ~n607 & ~n608;
  assign n610 = n605 & n609;
  assign n611 = ~n603 & ~n610;
  assign n612 = po09 & ~n611;
  assign n613 = ~po09 & n611;
  assign n614 = ~n612 & ~n613;
  assign n615 = n503 & po05;
  assign n616 = ~n507 & ~n615;
  assign n617 = n508 & po05;
  assign n618 = ~n616 & ~n617;
  assign n619 = n614 & n618;
  assign n620 = ~n612 & ~n619;
  assign n621 = po10 & ~n620;
  assign n622 = ~po10 & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = n512 & po05;
  assign n625 = ~n516 & ~n624;
  assign n626 = n517 & po05;
  assign n627 = ~n625 & ~n626;
  assign n628 = n623 & n627;
  assign n629 = ~n621 & ~n628;
  assign n630 = po11 & ~n629;
  assign n631 = ~po11 & n629;
  assign n632 = ~n630 & ~n631;
  assign n633 = n568 & po05;
  assign n634 = n576 & n632;
  assign n635 = ~n630 & ~n634;
  assign n636 = po12 & ~n635;
  assign n637 = ~po12 & n635;
  assign n638 = ~n636 & ~n637;
  assign n639 = n527 & po05;
  assign n640 = ~n531 & ~n639;
  assign n641 = n532 & po05;
  assign n642 = ~n640 & ~n641;
  assign n643 = n638 & n642;
  assign n644 = ~n636 & ~n643;
  assign n645 = po13 & ~n644;
  assign n646 = ~po13 & n644;
  assign n647 = ~n645 & ~n646;
  assign n648 = n536 & po05;
  assign n649 = ~n540 & ~n648;
  assign n650 = n541 & po05;
  assign n651 = ~n649 & ~n650;
  assign n652 = n647 & n651;
  assign n653 = ~n645 & ~n652;
  assign n654 = po14 & ~n653;
  assign n655 = ~po14 & n653;
  assign n656 = ~n654 & ~n655;
  assign n657 = n545 & po05;
  assign n658 = ~n549 & ~n657;
  assign n659 = n550 & po05;
  assign n660 = ~n658 & ~n659;
  assign n661 = n656 & n660;
  assign n662 = ~n654 & ~n661;
  assign n663 = po15 & ~n662;
  assign n664 = ~po15 & n662;
  assign n665 = ~n663 & ~n664;
  assign n666 = n554 & po05;
  assign n667 = ~n558 & ~n666;
  assign n668 = n559 & po05;
  assign n669 = ~n667 & ~n668;
  assign n670 = n665 & n669;
  assign n671 = ~n663 & ~n670;
  assign n672 = ~n563 & ~n567;
  assign n673 = ~n671 & ~n672;
  assign po04 = n633 | ~n673;
  assign n675 = n632 & po04;
  assign n676 = ~n576 & ~n675;
  assign n677 = n634 & po04;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~pi06 & ~pi07;
  assign n680 = po04 & n679;
  assign n681 = pi08 & ~po04;
  assign n682 = ~pi08 & po04;
  assign n683 = ~n681 & ~n682;
  assign n684 = ~po04 & ~n679;
  assign n685 = ~n680 & ~n684;
  assign n686 = n683 & n685;
  assign n687 = ~n680 & ~n686;
  assign n688 = po05 & ~n687;
  assign n689 = ~po05 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = pi09 & ~n682;
  assign n692 = n577 & po04;
  assign n693 = ~n691 & ~n692;
  assign n694 = n690 & n693;
  assign n695 = ~n688 & ~n694;
  assign n696 = po06 & ~n695;
  assign n697 = ~po06 & n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = n583 & po04;
  assign n700 = ~n581 & ~n699;
  assign n701 = n584 & po04;
  assign n702 = ~n700 & ~n701;
  assign n703 = n698 & n702;
  assign n704 = ~n696 & ~n703;
  assign n705 = po07 & ~n704;
  assign n706 = ~po07 & n704;
  assign n707 = ~n705 & ~n706;
  assign n708 = n588 & po04;
  assign n709 = ~n591 & ~n708;
  assign n710 = n592 & po04;
  assign n711 = ~n709 & ~n710;
  assign n712 = n707 & n711;
  assign n713 = ~n705 & ~n712;
  assign n714 = po08 & ~n713;
  assign n715 = ~po08 & n713;
  assign n716 = ~n714 & ~n715;
  assign n717 = n596 & po04;
  assign n718 = ~n600 & ~n717;
  assign n719 = n601 & po04;
  assign n720 = ~n718 & ~n719;
  assign n721 = n716 & n720;
  assign n722 = ~n714 & ~n721;
  assign n723 = po09 & ~n722;
  assign n724 = ~po09 & n722;
  assign n725 = ~n723 & ~n724;
  assign n726 = n605 & po04;
  assign n727 = ~n609 & ~n726;
  assign n728 = n610 & po04;
  assign n729 = ~n727 & ~n728;
  assign n730 = n725 & n729;
  assign n731 = ~n723 & ~n730;
  assign n732 = po10 & ~n731;
  assign n733 = ~po10 & n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = n614 & po04;
  assign n736 = ~n618 & ~n735;
  assign n737 = n619 & po04;
  assign n738 = ~n736 & ~n737;
  assign n739 = n734 & n738;
  assign n740 = ~n732 & ~n739;
  assign n741 = po11 & ~n740;
  assign n742 = ~po11 & n740;
  assign n743 = ~n741 & ~n742;
  assign n744 = n623 & po04;
  assign n745 = ~n627 & ~n744;
  assign n746 = n628 & po04;
  assign n747 = ~n745 & ~n746;
  assign n748 = n743 & n747;
  assign n749 = ~n741 & ~n748;
  assign n750 = po12 & ~n749;
  assign n751 = ~po12 & n749;
  assign n752 = ~n750 & ~n751;
  assign n753 = n670 & po04;
  assign n754 = n678 & n752;
  assign n755 = ~n750 & ~n754;
  assign n756 = po13 & ~n755;
  assign n757 = ~po13 & n755;
  assign n758 = ~n756 & ~n757;
  assign n759 = n638 & po04;
  assign n760 = ~n642 & ~n759;
  assign n761 = n643 & po04;
  assign n762 = ~n760 & ~n761;
  assign n763 = n758 & n762;
  assign n764 = ~n756 & ~n763;
  assign n765 = po14 & ~n764;
  assign n766 = ~po14 & n764;
  assign n767 = ~n765 & ~n766;
  assign n768 = n647 & po04;
  assign n769 = ~n651 & ~n768;
  assign n770 = n652 & po04;
  assign n771 = ~n769 & ~n770;
  assign n772 = n767 & n771;
  assign n773 = ~n765 & ~n772;
  assign n774 = po15 & ~n773;
  assign n775 = ~po15 & n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = n656 & po04;
  assign n778 = ~n660 & ~n777;
  assign n779 = n661 & po04;
  assign n780 = ~n778 & ~n779;
  assign n781 = n776 & n780;
  assign n782 = ~n774 & ~n781;
  assign n783 = ~n665 & ~n669;
  assign n784 = ~n782 & ~n783;
  assign po03 = n753 | ~n784;
  assign n786 = n752 & po03;
  assign n787 = ~n678 & ~n786;
  assign n788 = n754 & po03;
  assign n789 = ~n787 & ~n788;
  assign n790 = ~pi04 & ~pi05;
  assign n791 = po03 & n790;
  assign n792 = pi06 & ~po03;
  assign n793 = ~pi06 & po03;
  assign n794 = ~n792 & ~n793;
  assign n795 = ~po03 & ~n790;
  assign n796 = ~n791 & ~n795;
  assign n797 = n794 & n796;
  assign n798 = ~n791 & ~n797;
  assign n799 = po04 & ~n798;
  assign n800 = ~po04 & n798;
  assign n801 = ~n799 & ~n800;
  assign n802 = pi07 & ~n793;
  assign n803 = n679 & po03;
  assign n804 = ~n802 & ~n803;
  assign n805 = n801 & n804;
  assign n806 = ~n799 & ~n805;
  assign n807 = po05 & ~n806;
  assign n808 = ~po05 & n806;
  assign n809 = ~n807 & ~n808;
  assign n810 = n685 & po03;
  assign n811 = ~n683 & ~n810;
  assign n812 = n686 & po03;
  assign n813 = ~n811 & ~n812;
  assign n814 = n809 & n813;
  assign n815 = ~n807 & ~n814;
  assign n816 = po06 & ~n815;
  assign n817 = ~po06 & n815;
  assign n818 = ~n816 & ~n817;
  assign n819 = n690 & po03;
  assign n820 = ~n693 & ~n819;
  assign n821 = n694 & po03;
  assign n822 = ~n820 & ~n821;
  assign n823 = n818 & n822;
  assign n824 = ~n816 & ~n823;
  assign n825 = po07 & ~n824;
  assign n826 = ~po07 & n824;
  assign n827 = ~n825 & ~n826;
  assign n828 = n698 & po03;
  assign n829 = ~n702 & ~n828;
  assign n830 = n703 & po03;
  assign n831 = ~n829 & ~n830;
  assign n832 = n827 & n831;
  assign n833 = ~n825 & ~n832;
  assign n834 = po08 & ~n833;
  assign n835 = ~po08 & n833;
  assign n836 = ~n834 & ~n835;
  assign n837 = n707 & po03;
  assign n838 = ~n711 & ~n837;
  assign n839 = n712 & po03;
  assign n840 = ~n838 & ~n839;
  assign n841 = n836 & n840;
  assign n842 = ~n834 & ~n841;
  assign n843 = po09 & ~n842;
  assign n844 = ~po09 & n842;
  assign n845 = ~n843 & ~n844;
  assign n846 = n716 & po03;
  assign n847 = ~n720 & ~n846;
  assign n848 = n721 & po03;
  assign n849 = ~n847 & ~n848;
  assign n850 = n845 & n849;
  assign n851 = ~n843 & ~n850;
  assign n852 = po10 & ~n851;
  assign n853 = ~po10 & n851;
  assign n854 = ~n852 & ~n853;
  assign n855 = n725 & po03;
  assign n856 = ~n729 & ~n855;
  assign n857 = n730 & po03;
  assign n858 = ~n856 & ~n857;
  assign n859 = n854 & n858;
  assign n860 = ~n852 & ~n859;
  assign n861 = po11 & ~n860;
  assign n862 = ~po11 & n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = n734 & po03;
  assign n865 = ~n738 & ~n864;
  assign n866 = n739 & po03;
  assign n867 = ~n865 & ~n866;
  assign n868 = n863 & n867;
  assign n869 = ~n861 & ~n868;
  assign n870 = po12 & ~n869;
  assign n871 = ~po12 & n869;
  assign n872 = ~n870 & ~n871;
  assign n873 = n743 & po03;
  assign n874 = ~n747 & ~n873;
  assign n875 = n748 & po03;
  assign n876 = ~n874 & ~n875;
  assign n877 = n872 & n876;
  assign n878 = ~n870 & ~n877;
  assign n879 = po13 & ~n878;
  assign n880 = ~po13 & n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = n781 & po03;
  assign n883 = n789 & n881;
  assign n884 = ~n879 & ~n883;
  assign n885 = po14 & ~n884;
  assign n886 = ~po14 & n884;
  assign n887 = ~n885 & ~n886;
  assign n888 = n758 & po03;
  assign n889 = ~n762 & ~n888;
  assign n890 = n763 & po03;
  assign n891 = ~n889 & ~n890;
  assign n892 = n887 & n891;
  assign n893 = ~n885 & ~n892;
  assign n894 = po15 & ~n893;
  assign n895 = ~po15 & n893;
  assign n896 = ~n894 & ~n895;
  assign n897 = n767 & po03;
  assign n898 = ~n771 & ~n897;
  assign n899 = n772 & po03;
  assign n900 = ~n898 & ~n899;
  assign n901 = n896 & n900;
  assign n902 = ~n894 & ~n901;
  assign n903 = ~n776 & ~n780;
  assign n904 = ~n902 & ~n903;
  assign po02 = n882 | ~n904;
  assign n906 = n881 & po02;
  assign n907 = ~n789 & ~n906;
  assign n908 = n883 & po02;
  assign n909 = ~n907 & ~n908;
  assign n910 = ~pi02 & ~pi03;
  assign n911 = po02 & n910;
  assign n912 = pi04 & ~po02;
  assign n913 = ~pi04 & po02;
  assign n914 = ~n912 & ~n913;
  assign n915 = ~po02 & ~n910;
  assign n916 = ~n911 & ~n915;
  assign n917 = n914 & n916;
  assign n918 = ~n911 & ~n917;
  assign n919 = po03 & ~n918;
  assign n920 = ~po03 & n918;
  assign n921 = ~n919 & ~n920;
  assign n922 = pi05 & ~n913;
  assign n923 = n790 & po02;
  assign n924 = ~n922 & ~n923;
  assign n925 = n921 & n924;
  assign n926 = ~n919 & ~n925;
  assign n927 = po04 & ~n926;
  assign n928 = ~po04 & n926;
  assign n929 = ~n927 & ~n928;
  assign n930 = n796 & po02;
  assign n931 = ~n794 & ~n930;
  assign n932 = n797 & po02;
  assign n933 = ~n931 & ~n932;
  assign n934 = n929 & n933;
  assign n935 = ~n927 & ~n934;
  assign n936 = po05 & ~n935;
  assign n937 = ~po05 & n935;
  assign n938 = ~n936 & ~n937;
  assign n939 = n801 & po02;
  assign n940 = ~n804 & ~n939;
  assign n941 = n805 & po02;
  assign n942 = ~n940 & ~n941;
  assign n943 = n938 & n942;
  assign n944 = ~n936 & ~n943;
  assign n945 = po06 & ~n944;
  assign n946 = ~po06 & n944;
  assign n947 = ~n945 & ~n946;
  assign n948 = n809 & po02;
  assign n949 = ~n813 & ~n948;
  assign n950 = n814 & po02;
  assign n951 = ~n949 & ~n950;
  assign n952 = n947 & n951;
  assign n953 = ~n945 & ~n952;
  assign n954 = po07 & ~n953;
  assign n955 = ~po07 & n953;
  assign n956 = ~n954 & ~n955;
  assign n957 = n818 & po02;
  assign n958 = ~n822 & ~n957;
  assign n959 = n823 & po02;
  assign n960 = ~n958 & ~n959;
  assign n961 = n956 & n960;
  assign n962 = ~n954 & ~n961;
  assign n963 = po08 & ~n962;
  assign n964 = ~po08 & n962;
  assign n965 = ~n963 & ~n964;
  assign n966 = n827 & po02;
  assign n967 = ~n831 & ~n966;
  assign n968 = n832 & po02;
  assign n969 = ~n967 & ~n968;
  assign n970 = n965 & n969;
  assign n971 = ~n963 & ~n970;
  assign n972 = po09 & ~n971;
  assign n973 = ~po09 & n971;
  assign n974 = ~n972 & ~n973;
  assign n975 = n836 & po02;
  assign n976 = ~n840 & ~n975;
  assign n977 = n841 & po02;
  assign n978 = ~n976 & ~n977;
  assign n979 = n974 & n978;
  assign n980 = ~n972 & ~n979;
  assign n981 = po10 & ~n980;
  assign n982 = ~po10 & n980;
  assign n983 = ~n981 & ~n982;
  assign n984 = n845 & po02;
  assign n985 = ~n849 & ~n984;
  assign n986 = n850 & po02;
  assign n987 = ~n985 & ~n986;
  assign n988 = n983 & n987;
  assign n989 = ~n981 & ~n988;
  assign n990 = po11 & ~n989;
  assign n991 = ~po11 & n989;
  assign n992 = ~n990 & ~n991;
  assign n993 = n854 & po02;
  assign n994 = ~n858 & ~n993;
  assign n995 = n859 & po02;
  assign n996 = ~n994 & ~n995;
  assign n997 = n992 & n996;
  assign n998 = ~n990 & ~n997;
  assign n999 = po12 & ~n998;
  assign n1000 = ~po12 & n998;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = n863 & po02;
  assign n1003 = ~n867 & ~n1002;
  assign n1004 = n868 & po02;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = n1001 & n1005;
  assign n1007 = ~n999 & ~n1006;
  assign n1008 = po13 & ~n1007;
  assign n1009 = ~po13 & n1007;
  assign n1010 = ~n1008 & ~n1009;
  assign n1011 = n872 & po02;
  assign n1012 = ~n876 & ~n1011;
  assign n1013 = n877 & po02;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = n1010 & n1014;
  assign n1016 = ~n1008 & ~n1015;
  assign n1017 = po14 & ~n1016;
  assign n1018 = ~po14 & n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n901 & po02;
  assign n1021 = n909 & n1019;
  assign n1022 = ~n1017 & ~n1021;
  assign n1023 = po15 & ~n1022;
  assign n1024 = ~po15 & n1022;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n887 & po02;
  assign n1027 = ~n891 & ~n1026;
  assign n1028 = n892 & po02;
  assign n1029 = ~n1027 & ~n1028;
  assign n1030 = n1025 & n1029;
  assign n1031 = ~n1023 & ~n1030;
  assign n1032 = ~n896 & ~n900;
  assign n1033 = ~n1031 & ~n1032;
  assign po01 = n1020 | ~n1033;
  assign n1035 = n1019 & po01;
  assign n1036 = ~n909 & ~n1035;
  assign n1037 = n1021 & po01;
  assign n1038 = ~n1036 & ~n1037;
  assign n1039 = n1010 & po01;
  assign n1040 = ~n1014 & ~n1039;
  assign n1041 = n1015 & po01;
  assign n1042 = ~n1040 & ~n1041;
  assign n1043 = n1001 & po01;
  assign n1044 = ~n1005 & ~n1043;
  assign n1045 = n1006 & po01;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = n992 & po01;
  assign n1048 = ~n996 & ~n1047;
  assign n1049 = n997 & po01;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = n983 & po01;
  assign n1052 = ~n987 & ~n1051;
  assign n1053 = n988 & po01;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n974 & po01;
  assign n1056 = ~n978 & ~n1055;
  assign n1057 = n979 & po01;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = n965 & po01;
  assign n1060 = ~n969 & ~n1059;
  assign n1061 = n970 & po01;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n956 & po01;
  assign n1064 = ~n960 & ~n1063;
  assign n1065 = n961 & po01;
  assign n1066 = ~n1064 & ~n1065;
  assign n1067 = n947 & po01;
  assign n1068 = ~n951 & ~n1067;
  assign n1069 = n952 & po01;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = n938 & po01;
  assign n1072 = ~n942 & ~n1071;
  assign n1073 = n943 & po01;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = n929 & po01;
  assign n1076 = ~n933 & ~n1075;
  assign n1077 = n934 & po01;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n921 & po01;
  assign n1080 = ~n924 & ~n1079;
  assign n1081 = n925 & po01;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = n916 & po01;
  assign n1084 = ~n914 & ~n1083;
  assign n1085 = n917 & po01;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~pi02 & po01;
  assign n1088 = pi03 & ~n1087;
  assign n1089 = n910 & po01;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = pi02 & po01;
  assign n1092 = ~pi02 & ~po01;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = ~po01 & n1093;
  assign n1095 = ~pi00 & ~pi01;
  assign n1096 = ~n1094 & n1095;
  assign n1097 = po01 & ~n1093;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = ~n1090 & n1098;
  assign n1100 = po02 & ~n1099;
  assign n1101 = n1090 & ~n1098;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = ~n1086 & n1102;
  assign n1104 = po03 & ~n1103;
  assign n1105 = n1086 & ~n1102;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n1082 & n1106;
  assign n1108 = po04 & ~n1107;
  assign n1109 = n1082 & ~n1106;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1078 & n1110;
  assign n1112 = po05 & ~n1111;
  assign n1113 = n1078 & ~n1110;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = ~n1074 & n1114;
  assign n1116 = po06 & ~n1115;
  assign n1117 = n1074 & ~n1114;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = ~n1070 & n1118;
  assign n1120 = po07 & ~n1119;
  assign n1121 = n1070 & ~n1118;
  assign n1122 = ~n1120 & ~n1121;
  assign n1123 = ~n1066 & n1122;
  assign n1124 = po08 & ~n1123;
  assign n1125 = n1066 & ~n1122;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = ~n1062 & n1126;
  assign n1128 = po09 & ~n1127;
  assign n1129 = n1062 & ~n1126;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1058 & n1130;
  assign n1132 = po10 & ~n1131;
  assign n1133 = n1058 & ~n1130;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = ~n1054 & n1134;
  assign n1136 = po11 & ~n1135;
  assign n1137 = n1054 & ~n1134;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = ~n1050 & n1138;
  assign n1140 = po12 & ~n1139;
  assign n1141 = n1050 & ~n1138;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = ~n1046 & n1142;
  assign n1144 = po13 & ~n1143;
  assign n1145 = n1046 & ~n1142;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = ~n1042 & n1146;
  assign n1148 = po14 & ~n1147;
  assign n1149 = n1042 & ~n1146;
  assign n1150 = ~n1148 & ~n1149;
  assign n1151 = n1022 & ~n1029;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n1038 & n1152;
  assign n1154 = ~po15 & ~n1153;
  assign n1155 = ~n1022 & ~n1029;
  assign n1156 = po15 & n1155;
  assign n1157 = ~n1154 & ~n1156;
  assign n1158 = ~n1038 & n1150;
  assign n1159 = n1030 & po01;
  assign n1160 = ~n1158 & ~n1159;
  assign po00 = ~n1157 | ~n1160;
endmodule


