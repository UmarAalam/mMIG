//Written by the Majority Logic Package Wed Apr 29 22:50:58 2015
module top (
            pi00000, pi00001, pi00002, pi00003, pi00004, pi00005, pi00006, pi00007, pi00008, pi00009, pi00010, pi00011, pi00012, pi00013, pi00014, pi00015, pi00016, pi00017, pi00018, pi00019, pi00020, pi00021, pi00022, pi00023, pi00024, pi00025, pi00026, pi00027, pi00028, pi00029, pi00030, pi00031, pi00032, pi00033, pi00034, pi00035, pi00036, pi00037, pi00038, pi00039, pi00040, pi00041, pi00042, pi00043, pi00044, pi00045, pi00046, pi00047, pi00048, pi00049, pi00050, pi00051, pi00052, pi00053, pi00054, pi00055, pi00056, pi00057, pi00058, pi00059, pi00060, pi00061, pi00062, pi00063, pi00064, pi00065, pi00066, pi00067, pi00068, pi00069, pi00070, pi00071, pi00072, pi00073, pi00074, pi00075, pi00076, pi00077, pi00078, pi00079, pi00080, pi00081, pi00082, pi00083, pi00084, pi00085, pi00086, pi00087, pi00088, pi00089, pi00090, pi00091, pi00092, pi00093, pi00094, pi00095, pi00096, pi00097, pi00098, pi00099, pi00100, pi00101, pi00102, pi00103, pi00104, pi00105, pi00106, pi00107, pi00108, pi00109, pi00110, pi00111, pi00112, pi00113, pi00114, pi00115, pi00116, pi00117, pi00118, pi00119, pi00120, pi00121, pi00122, pi00123, pi00124, pi00125, pi00126, pi00127, pi00128, pi00129, pi00130, pi00131, pi00132, pi00133, pi00134, pi00135, pi00136, pi00137, pi00138, pi00139, pi00140, pi00141, pi00142, pi00143, pi00144, pi00145, pi00146, pi00147, pi00148, pi00149, pi00150, pi00151, pi00152, pi00153, pi00154, pi00155, pi00156, pi00157, pi00158, pi00159, pi00160, pi00161, pi00162, pi00163, pi00164, pi00165, pi00166, pi00167, pi00168, pi00169, pi00170, pi00171, pi00172, pi00173, pi00174, pi00175, pi00176, pi00177, pi00178, pi00179, pi00180, pi00181, pi00182, pi00183, pi00184, pi00185, pi00186, pi00187, pi00188, pi00189, pi00190, pi00191, pi00192, pi00193, pi00194, pi00195, pi00196, pi00197, pi00198, pi00199, pi00200, pi00201, pi00202, pi00203, pi00204, pi00205, pi00206, pi00207, pi00208, pi00209, pi00210, pi00211, pi00212, pi00213, pi00214, pi00215, pi00216, pi00217, pi00218, pi00219, pi00220, pi00221, pi00222, pi00223, pi00224, pi00225, pi00226, pi00227, pi00228, pi00229, pi00230, pi00231, pi00232, pi00233, pi00234, pi00235, pi00236, pi00237, pi00238, pi00239, pi00240, pi00241, pi00242, pi00243, pi00244, pi00245, pi00246, pi00247, pi00248, pi00249, pi00250, pi00251, pi00252, pi00253, pi00254, pi00255, pi00256, pi00257, pi00258, pi00259, pi00260, pi00261, pi00262, pi00263, pi00264, pi00265, pi00266, pi00267, pi00268, pi00269, pi00270, pi00271, pi00272, pi00273, pi00274, pi00275, pi00276, pi00277, pi00278, pi00279, pi00280, pi00281, pi00282, pi00283, pi00284, pi00285, pi00286, pi00287, pi00288, pi00289, pi00290, pi00291, pi00292, pi00293, pi00294, pi00295, pi00296, pi00297, pi00298, pi00299, pi00300, pi00301, pi00302, pi00303, pi00304, pi00305, pi00306, pi00307, pi00308, pi00309, pi00310, pi00311, pi00312, pi00313, pi00314, pi00315, pi00316, pi00317, pi00318, pi00319, pi00320, pi00321, pi00322, pi00323, pi00324, pi00325, pi00326, pi00327, pi00328, pi00329, pi00330, pi00331, pi00332, pi00333, pi00334, pi00335, pi00336, pi00337, pi00338, pi00339, pi00340, pi00341, pi00342, pi00343, pi00344, pi00345, pi00346, pi00347, pi00348, pi00349, pi00350, pi00351, pi00352, pi00353, pi00354, pi00355, pi00356, pi00357, pi00358, pi00359, pi00360, pi00361, pi00362, pi00363, pi00364, pi00365, pi00366, pi00367, pi00368, pi00369, pi00370, pi00371, pi00372, pi00373, pi00374, pi00375, pi00376, pi00377, pi00378, pi00379, pi00380, pi00381, pi00382, pi00383, pi00384, pi00385, pi00386, pi00387, pi00388, pi00389, pi00390, pi00391, pi00392, pi00393, pi00394, pi00395, pi00396, pi00397, pi00398, pi00399, pi00400, pi00401, pi00402, pi00403, pi00404, pi00405, pi00406, pi00407, pi00408, pi00409, pi00410, pi00411, pi00412, pi00413, pi00414, pi00415, pi00416, pi00417, pi00418, pi00419, pi00420, pi00421, pi00422, pi00423, pi00424, pi00425, pi00426, pi00427, pi00428, pi00429, pi00430, pi00431, pi00432, pi00433, pi00434, pi00435, pi00436, pi00437, pi00438, pi00439, pi00440, pi00441, pi00442, pi00443, pi00444, pi00445, pi00446, pi00447, pi00448, pi00449, pi00450, pi00451, pi00452, pi00453, pi00454, pi00455, pi00456, pi00457, pi00458, pi00459, pi00460, pi00461, pi00462, pi00463, pi00464, pi00465, pi00466, pi00467, pi00468, pi00469, pi00470, pi00471, pi00472, pi00473, pi00474, pi00475, pi00476, pi00477, pi00478, pi00479, pi00480, pi00481, pi00482, pi00483, pi00484, pi00485, pi00486, pi00487, pi00488, pi00489, pi00490, pi00491, pi00492, pi00493, pi00494, pi00495, pi00496, pi00497, pi00498, pi00499, pi00500, pi00501, pi00502, pi00503, pi00504, pi00505, pi00506, pi00507, pi00508, pi00509, pi00510, pi00511, pi00512, pi00513, pi00514, pi00515, pi00516, pi00517, pi00518, pi00519, pi00520, pi00521, pi00522, pi00523, pi00524, pi00525, pi00526, pi00527, pi00528, pi00529, pi00530, pi00531, pi00532, pi00533, pi00534, pi00535, pi00536, pi00537, pi00538, pi00539, pi00540, pi00541, pi00542, pi00543, pi00544, pi00545, pi00546, pi00547, pi00548, pi00549, pi00550, pi00551, pi00552, pi00553, pi00554, pi00555, pi00556, pi00557, pi00558, pi00559, pi00560, pi00561, pi00562, pi00563, pi00564, pi00565, pi00566, pi00567, pi00568, pi00569, pi00570, pi00571, pi00572, pi00573, pi00574, pi00575, pi00576, pi00577, pi00578, pi00579, pi00580, pi00581, pi00582, pi00583, pi00584, pi00585, pi00586, pi00587, pi00588, pi00589, pi00590, pi00591, pi00592, pi00593, pi00594, pi00595, pi00596, pi00597, pi00598, pi00599, pi00600, pi00601, pi00602, pi00603, pi00604, pi00605, pi00606, pi00607, pi00608, pi00609, pi00610, pi00611, pi00612, pi00613, pi00614, pi00615, pi00616, pi00617, pi00618, pi00619, pi00620, pi00621, pi00622, pi00623, pi00624, pi00625, pi00626, pi00627, pi00628, pi00629, pi00630, pi00631, pi00632, pi00633, pi00634, pi00635, pi00636, pi00637, pi00638, pi00639, pi00640, pi00641, pi00642, pi00643, pi00644, pi00645, pi00646, pi00647, pi00648, pi00649, pi00650, pi00651, pi00652, pi00653, pi00654, pi00655, pi00656, pi00657, pi00658, pi00659, pi00660, pi00661, pi00662, pi00663, pi00664, pi00665, pi00666, pi00667, pi00668, pi00669, pi00670, pi00671, pi00672, pi00673, pi00674, pi00675, pi00676, pi00677, pi00678, pi00679, pi00680, pi00681, pi00682, pi00683, pi00684, pi00685, pi00686, pi00687, pi00688, pi00689, pi00690, pi00691, pi00692, pi00693, pi00694, pi00695, pi00696, pi00697, pi00698, pi00699, pi00700, pi00701, pi00702, pi00703, pi00704, pi00705, pi00706, pi00707, pi00708, pi00709, pi00710, pi00711, pi00712, pi00713, pi00714, pi00715, pi00716, pi00717, pi00718, pi00719, pi00720, pi00721, pi00722, pi00723, pi00724, pi00725, pi00726, pi00727, pi00728, pi00729, pi00730, pi00731, pi00732, pi00733, pi00734, pi00735, pi00736, pi00737, pi00738, pi00739, pi00740, pi00741, pi00742, pi00743, pi00744, pi00745, pi00746, pi00747, pi00748, pi00749, pi00750, pi00751, pi00752, pi00753, pi00754, pi00755, pi00756, pi00757, pi00758, pi00759, pi00760, pi00761, pi00762, pi00763, pi00764, pi00765, pi00766, pi00767, pi00768, pi00769, pi00770, pi00771, pi00772, pi00773, pi00774, pi00775, pi00776, pi00777, pi00778, pi00779, pi00780, pi00781, pi00782, pi00783, pi00784, pi00785, pi00786, pi00787, pi00788, pi00789, pi00790, pi00791, pi00792, pi00793, pi00794, pi00795, pi00796, pi00797, pi00798, pi00799, pi00800, pi00801, pi00802, pi00803, pi00804, pi00805, pi00806, pi00807, pi00808, pi00809, pi00810, pi00811, pi00812, pi00813, pi00814, pi00815, pi00816, pi00817, pi00818, pi00819, pi00820, pi00821, pi00822, pi00823, pi00824, pi00825, pi00826, pi00827, pi00828, pi00829, pi00830, pi00831, pi00832, pi00833, pi00834, pi00835, pi00836, pi00837, pi00838, pi00839, pi00840, pi00841, pi00842, pi00843, pi00844, pi00845, pi00846, pi00847, pi00848, pi00849, pi00850, pi00851, pi00852, pi00853, pi00854, pi00855, pi00856, pi00857, pi00858, pi00859, pi00860, pi00861, pi00862, pi00863, pi00864, pi00865, pi00866, pi00867, pi00868, pi00869, pi00870, pi00871, pi00872, pi00873, pi00874, pi00875, pi00876, pi00877, pi00878, pi00879, pi00880, pi00881, pi00882, pi00883, pi00884, pi00885, pi00886, pi00887, pi00888, pi00889, pi00890, pi00891, pi00892, pi00893, pi00894, pi00895, pi00896, pi00897, pi00898, pi00899, pi00900, pi00901, pi00902, pi00903, pi00904, pi00905, pi00906, pi00907, pi00908, pi00909, pi00910, pi00911, pi00912, pi00913, pi00914, pi00915, pi00916, pi00917, pi00918, pi00919, pi00920, pi00921, pi00922, pi00923, pi00924, pi00925, pi00926, pi00927, pi00928, pi00929, pi00930, pi00931, pi00932, pi00933, pi00934, pi00935, pi00936, pi00937, pi00938, pi00939, pi00940, pi00941, pi00942, pi00943, pi00944, pi00945, pi00946, pi00947, pi00948, pi00949, pi00950, pi00951, pi00952, pi00953, pi00954, pi00955, pi00956, pi00957, pi00958, pi00959, pi00960, pi00961, pi00962, pi00963, pi00964, pi00965, pi00966, pi00967, pi00968, pi00969, pi00970, pi00971, pi00972, pi00973, pi00974, pi00975, pi00976, pi00977, pi00978, pi00979, pi00980, pi00981, pi00982, pi00983, pi00984, pi00985, pi00986, pi00987, pi00988, pi00989, pi00990, pi00991, pi00992, pi00993, pi00994, pi00995, pi00996, pi00997, pi00998, pi00999, pi01000, pi01001, pi01002, pi01003, pi01004, pi01005, pi01006, pi01007, pi01008, pi01009, pi01010, pi01011, pi01012, pi01013, pi01014, pi01015, pi01016, pi01017, pi01018, pi01019, pi01020, pi01021, pi01022, pi01023, pi01024, pi01025, pi01026, pi01027, pi01028, pi01029, pi01030, pi01031, pi01032, pi01033, pi01034, pi01035, pi01036, pi01037, pi01038, pi01039, pi01040, pi01041, pi01042, pi01043, pi01044, pi01045, pi01046, pi01047, pi01048, pi01049, pi01050, pi01051, pi01052, pi01053, pi01054, pi01055, pi01056, pi01057, pi01058, pi01059, pi01060, pi01061, pi01062, pi01063, pi01064, pi01065, pi01066, pi01067, pi01068, pi01069, pi01070, pi01071, pi01072, pi01073, pi01074, pi01075, pi01076, pi01077, pi01078, pi01079, pi01080, pi01081, pi01082, pi01083, pi01084, pi01085, pi01086, pi01087, pi01088, pi01089, pi01090, pi01091, pi01092, pi01093, pi01094, pi01095, pi01096, pi01097, pi01098, pi01099, pi01100, pi01101, pi01102, pi01103, pi01104, pi01105, pi01106, pi01107, pi01108, pi01109, pi01110, pi01111, pi01112, pi01113, pi01114, pi01115, pi01116, pi01117, pi01118, pi01119, pi01120, pi01121, pi01122, pi01123, pi01124, pi01125, pi01126, pi01127, pi01128, pi01129, pi01130, pi01131, pi01132, pi01133, pi01134, pi01135, pi01136, pi01137, pi01138, pi01139, pi01140, pi01141, pi01142, pi01143, pi01144, pi01145, pi01146, pi01147, pi01148, pi01149, pi01150, pi01151, pi01152, pi01153, pi01154, pi01155, pi01156, pi01157, pi01158, pi01159, pi01160, pi01161, pi01162, pi01163, pi01164, pi01165, pi01166, pi01167, pi01168, pi01169, pi01170, pi01171, pi01172, pi01173, pi01174, pi01175, pi01176, pi01177, pi01178, pi01179, pi01180, pi01181, pi01182, pi01183, pi01184, pi01185, pi01186, pi01187, pi01188, pi01189, pi01190, pi01191, pi01192, pi01193, pi01194, pi01195, pi01196, pi01197, pi01198, pi01199, pi01200, pi01201, pi01202, pi01203, pi01204, pi01205, pi01206, pi01207, pi01208, pi01209, pi01210, pi01211, pi01212, pi01213, pi01214, pi01215, pi01216, pi01217, pi01218, pi01219, pi01220, pi01221, pi01222, pi01223, pi01224, pi01225, pi01226, pi01227, pi01228, pi01229, pi01230, pi01231, pi01232, pi01233, pi01234, pi01235, pi01236, pi01237, pi01238, pi01239, pi01240, pi01241, pi01242, pi01243, pi01244, pi01245, pi01246, pi01247, pi01248, pi01249, pi01250, pi01251, pi01252, pi01253, pi01254, pi01255, pi01256, pi01257, pi01258, pi01259, pi01260, pi01261, pi01262, pi01263, pi01264, pi01265, pi01266, pi01267, pi01268, pi01269, pi01270, pi01271, pi01272, pi01273, pi01274, pi01275, pi01276, pi01277, pi01278, pi01279, pi01280, pi01281, pi01282, pi01283, pi01284, pi01285, pi01286, pi01287, pi01288, pi01289, pi01290, pi01291, pi01292, pi01293, pi01294, pi01295, pi01296, pi01297, pi01298, pi01299, pi01300, pi01301, pi01302, pi01303, pi01304, pi01305, pi01306, pi01307, pi01308, pi01309, pi01310, pi01311, pi01312, pi01313, pi01314, pi01315, pi01316, pi01317, pi01318, pi01319, pi01320, pi01321, pi01322, pi01323, pi01324, pi01325, pi01326, pi01327, pi01328, pi01329, pi01330, pi01331, pi01332, pi01333, pi01334, pi01335, pi01336, pi01337, pi01338, pi01339, pi01340, pi01341, pi01342, pi01343, pi01344, pi01345, pi01346, pi01347, pi01348, pi01349, pi01350, pi01351, pi01352, pi01353, pi01354, pi01355, pi01356, pi01357, pi01358, pi01359, pi01360, pi01361, pi01362, pi01363, pi01364, pi01365, pi01366, pi01367, pi01368, pi01369, pi01370, pi01371, pi01372, pi01373, pi01374, pi01375, pi01376, pi01377, pi01378, pi01379, pi01380, pi01381, pi01382, pi01383, pi01384, pi01385, pi01386, pi01387, pi01388, pi01389, pi01390, pi01391, pi01392, pi01393, pi01394, pi01395, pi01396, pi01397, pi01398, pi01399, pi01400, pi01401, pi01402, pi01403, pi01404, pi01405, pi01406, pi01407, pi01408, pi01409, pi01410, pi01411, pi01412, pi01413, pi01414, pi01415, pi01416, pi01417, pi01418, pi01419, pi01420, pi01421, pi01422, pi01423, pi01424, pi01425, pi01426, pi01427, pi01428, pi01429, pi01430, pi01431, pi01432, pi01433, pi01434, pi01435, pi01436, pi01437, pi01438, pi01439, pi01440, pi01441, pi01442, pi01443, pi01444, pi01445, pi01446, pi01447, pi01448, pi01449, pi01450, pi01451, pi01452, pi01453, pi01454, pi01455, pi01456, pi01457, pi01458, pi01459, pi01460, pi01461, pi01462, pi01463, pi01464, pi01465, pi01466, pi01467, pi01468, pi01469, pi01470, pi01471, pi01472, pi01473, pi01474, pi01475, pi01476, pi01477, pi01478, pi01479, pi01480, pi01481, pi01482, pi01483, pi01484, pi01485, pi01486, pi01487, pi01488, pi01489, pi01490, pi01491, pi01492, pi01493, pi01494, pi01495, pi01496, pi01497, pi01498, pi01499, pi01500, pi01501, pi01502, pi01503, pi01504, pi01505, pi01506, pi01507, pi01508, pi01509, pi01510, pi01511, pi01512, pi01513, pi01514, pi01515, pi01516, pi01517, pi01518, pi01519, pi01520, pi01521, pi01522, pi01523, pi01524, pi01525, pi01526, pi01527, pi01528, pi01529, pi01530, pi01531, pi01532, pi01533, pi01534, pi01535, pi01536, pi01537, pi01538, pi01539, pi01540, pi01541, pi01542, pi01543, pi01544, pi01545, pi01546, pi01547, pi01548, pi01549, pi01550, pi01551, pi01552, pi01553, pi01554, pi01555, pi01556, pi01557, pi01558, pi01559, pi01560, pi01561, pi01562, pi01563, pi01564, pi01565, pi01566, pi01567, pi01568, pi01569, pi01570, pi01571, pi01572, pi01573, pi01574, pi01575, pi01576, pi01577, pi01578, pi01579, pi01580, pi01581, pi01582, pi01583, pi01584, pi01585, pi01586, pi01587, pi01588, pi01589, pi01590, pi01591, pi01592, pi01593, pi01594, pi01595, pi01596, pi01597, pi01598, pi01599, pi01600, pi01601, pi01602, pi01603, pi01604, pi01605, pi01606, pi01607, pi01608, pi01609, pi01610, pi01611, pi01612, pi01613, pi01614, pi01615, pi01616, pi01617, pi01618, pi01619, pi01620, pi01621, pi01622, pi01623, pi01624, pi01625, pi01626, pi01627, pi01628, pi01629, pi01630, pi01631, pi01632, pi01633, pi01634, pi01635, pi01636, pi01637, pi01638, pi01639, pi01640, pi01641, pi01642, pi01643, pi01644, pi01645, pi01646, pi01647, pi01648, pi01649, pi01650, pi01651, pi01652, pi01653, pi01654, pi01655, pi01656, pi01657, pi01658, pi01659, pi01660, pi01661, pi01662, pi01663, pi01664, pi01665, pi01666, pi01667, pi01668, pi01669, pi01670, pi01671, pi01672, pi01673, pi01674, pi01675, pi01676, pi01677, pi01678, pi01679, pi01680, pi01681, pi01682, pi01683, pi01684, pi01685, pi01686, pi01687, pi01688, pi01689, pi01690, pi01691, pi01692, pi01693, pi01694, pi01695, pi01696, pi01697, pi01698, pi01699, pi01700, pi01701, pi01702, pi01703, pi01704, pi01705, pi01706, pi01707, pi01708, pi01709, pi01710, pi01711, pi01712, pi01713, pi01714, pi01715, pi01716, pi01717, pi01718, pi01719, pi01720, pi01721, pi01722, pi01723, pi01724, pi01725, pi01726, pi01727, pi01728, pi01729, pi01730, pi01731, pi01732, pi01733, pi01734, pi01735, pi01736, pi01737, pi01738, pi01739, pi01740, pi01741, pi01742, pi01743, pi01744, pi01745, pi01746, pi01747, pi01748, pi01749, pi01750, pi01751, pi01752, pi01753, pi01754, pi01755, pi01756, pi01757, pi01758, pi01759, pi01760, pi01761, pi01762, pi01763, pi01764, pi01765, pi01766, pi01767, pi01768, pi01769, pi01770, pi01771, pi01772, pi01773, pi01774, pi01775, pi01776, pi01777, pi01778, pi01779, pi01780, pi01781, pi01782, pi01783, pi01784, pi01785, pi01786, pi01787, pi01788, pi01789, pi01790, pi01791, pi01792, pi01793, pi01794, pi01795, pi01796, pi01797, pi01798, pi01799, pi01800, pi01801, pi01802, pi01803, pi01804, pi01805, pi01806, pi01807, pi01808, pi01809, pi01810, pi01811, pi01812, pi01813, pi01814, pi01815, pi01816, pi01817, pi01818, pi01819, pi01820, pi01821, pi01822, pi01823, pi01824, pi01825, pi01826, pi01827, pi01828, pi01829, pi01830, pi01831, pi01832, pi01833, pi01834, pi01835, pi01836, pi01837, pi01838, pi01839, pi01840, pi01841, pi01842, pi01843, pi01844, pi01845, pi01846, pi01847, pi01848, pi01849, pi01850, pi01851, pi01852, pi01853, pi01854, pi01855, pi01856, pi01857, pi01858, pi01859, pi01860, pi01861, pi01862, pi01863, pi01864, pi01865, pi01866, pi01867, pi01868, pi01869, pi01870, pi01871, pi01872, pi01873, pi01874, pi01875, pi01876, pi01877, pi01878, pi01879, pi01880, pi01881, pi01882, pi01883, pi01884, pi01885, pi01886, pi01887, pi01888, pi01889, pi01890, pi01891, pi01892, pi01893, pi01894, pi01895, pi01896, pi01897, pi01898, pi01899, pi01900, pi01901, pi01902, pi01903, pi01904, pi01905, pi01906, pi01907, pi01908, pi01909, pi01910, pi01911, pi01912, pi01913, pi01914, pi01915, pi01916, pi01917, pi01918, pi01919, pi01920, pi01921, pi01922, pi01923, pi01924, pi01925, pi01926, pi01927, pi01928, pi01929, pi01930, pi01931, pi01932, pi01933, pi01934, pi01935, pi01936, pi01937, pi01938, pi01939, pi01940, pi01941, pi01942, pi01943, pi01944, pi01945, pi01946, pi01947, pi01948, pi01949, pi01950, pi01951, pi01952, pi01953, pi01954, pi01955, pi01956, pi01957, pi01958, pi01959, pi01960, pi01961, pi01962, pi01963, pi01964, pi01965, pi01966, pi01967, pi01968, pi01969, pi01970, pi01971, pi01972, pi01973, pi01974, pi01975, pi01976, pi01977, pi01978, pi01979, pi01980, pi01981, pi01982, pi01983, pi01984, pi01985, pi01986, pi01987, pi01988, pi01989, pi01990, pi01991, pi01992, pi01993, pi01994, pi01995, pi01996, pi01997, pi01998, pi01999, pi02000, pi02001, pi02002, pi02003, pi02004, pi02005, pi02006, pi02007, pi02008, pi02009, pi02010, pi02011, pi02012, pi02013, pi02014, pi02015, pi02016, pi02017, pi02018, pi02019, pi02020, pi02021, pi02022, pi02023, pi02024, pi02025, pi02026, pi02027, pi02028, pi02029, pi02030, pi02031, pi02032, pi02033, pi02034, pi02035, pi02036, pi02037, pi02038, pi02039, pi02040, pi02041, pi02042, pi02043, pi02044, pi02045, pi02046, pi02047, pi02048, pi02049, pi02050, pi02051, pi02052, pi02053, pi02054, pi02055, pi02056, pi02057, pi02058, pi02059, pi02060, pi02061, pi02062, pi02063, pi02064, pi02065, pi02066, pi02067, pi02068, pi02069, pi02070, pi02071, pi02072, pi02073, pi02074, pi02075, pi02076, pi02077, pi02078, pi02079, pi02080, pi02081, pi02082, pi02083, pi02084, pi02085, pi02086, pi02087, pi02088, pi02089, pi02090, pi02091, pi02092, pi02093, pi02094, pi02095, pi02096, pi02097, pi02098, pi02099, pi02100, pi02101, pi02102, pi02103, pi02104, pi02105, pi02106, pi02107, pi02108, pi02109, pi02110, pi02111, pi02112, pi02113, pi02114, pi02115, pi02116, pi02117, pi02118, pi02119, pi02120, pi02121, pi02122, pi02123, pi02124, pi02125, pi02126, pi02127, pi02128, pi02129, pi02130, pi02131, pi02132, pi02133, pi02134, pi02135, pi02136, pi02137, pi02138, pi02139, pi02140, pi02141, pi02142, pi02143, pi02144, pi02145, pi02146, pi02147, pi02148, pi02149, pi02150, pi02151, pi02152, pi02153, pi02154, pi02155, pi02156, pi02157, pi02158, pi02159, pi02160, pi02161, pi02162, pi02163, pi02164, pi02165, pi02166, pi02167, pi02168, pi02169, pi02170, pi02171, pi02172, pi02173, pi02174, pi02175, pi02176, pi02177, pi02178, pi02179, pi02180, pi02181, pi02182, pi02183, pi02184, pi02185, pi02186, pi02187, pi02188, pi02189, pi02190, pi02191, pi02192, pi02193, pi02194, pi02195, pi02196, pi02197, pi02198, pi02199, pi02200, pi02201, pi02202, pi02203, pi02204, pi02205, pi02206, pi02207, pi02208, pi02209, pi02210, pi02211, pi02212, pi02213, pi02214, pi02215, pi02216, pi02217, pi02218, pi02219, pi02220, pi02221, pi02222, pi02223, pi02224, pi02225, pi02226, pi02227, pi02228, pi02229, pi02230, pi02231, pi02232, pi02233, pi02234, pi02235, pi02236, pi02237, pi02238, pi02239, pi02240, pi02241, pi02242, pi02243, pi02244, pi02245, pi02246, pi02247, pi02248, pi02249, pi02250, pi02251, pi02252, pi02253, pi02254, pi02255, pi02256, pi02257, pi02258, pi02259, pi02260, pi02261, pi02262, pi02263, pi02264, pi02265, pi02266, pi02267, pi02268, pi02269, pi02270, pi02271, pi02272, pi02273, pi02274, pi02275, pi02276, pi02277, pi02278, pi02279, pi02280, pi02281, pi02282, pi02283, pi02284, pi02285, pi02286, pi02287, pi02288, pi02289, pi02290, pi02291, pi02292, pi02293, pi02294, pi02295, pi02296, pi02297, pi02298, pi02299, pi02300, pi02301, pi02302, pi02303, pi02304, pi02305, pi02306, pi02307, pi02308, pi02309, pi02310, pi02311, pi02312, pi02313, pi02314, pi02315, pi02316, pi02317, pi02318, pi02319, pi02320, pi02321, pi02322, pi02323, pi02324, pi02325, pi02326, pi02327, pi02328, pi02329, pi02330, pi02331, pi02332, pi02333, pi02334, pi02335, pi02336, pi02337, pi02338, pi02339, pi02340, pi02341, pi02342, pi02343, pi02344, pi02345, pi02346, pi02347, pi02348, pi02349, pi02350, pi02351, pi02352, pi02353, pi02354, pi02355, pi02356, pi02357, pi02358, pi02359, pi02360, pi02361, pi02362, pi02363, pi02364, pi02365, pi02366, pi02367, pi02368, pi02369, pi02370, pi02371, pi02372, pi02373, pi02374, pi02375, pi02376, pi02377, pi02378, pi02379, pi02380, pi02381, pi02382, pi02383, pi02384, pi02385, pi02386, pi02387, pi02388, pi02389, pi02390, pi02391, pi02392, pi02393, pi02394, pi02395, pi02396, pi02397, pi02398, pi02399, pi02400, pi02401, pi02402, pi02403, pi02404, pi02405, pi02406, pi02407, pi02408, pi02409, pi02410, pi02411, pi02412, pi02413, pi02414, pi02415, pi02416, pi02417, pi02418, pi02419, pi02420, pi02421, pi02422, pi02423, pi02424, pi02425, pi02426, pi02427, pi02428, pi02429, pi02430, pi02431, pi02432, pi02433, pi02434, pi02435, pi02436, pi02437, pi02438, pi02439, pi02440, pi02441, pi02442, pi02443, pi02444, pi02445, pi02446, pi02447, pi02448, pi02449, pi02450, pi02451, pi02452, pi02453, pi02454, pi02455, pi02456, pi02457, pi02458, pi02459, pi02460, pi02461, pi02462, pi02463, pi02464, pi02465, pi02466, pi02467, pi02468, pi02469, pi02470, pi02471, pi02472, pi02473, pi02474, pi02475, pi02476, pi02477, pi02478, pi02479, pi02480, pi02481, pi02482, pi02483, pi02484, pi02485, pi02486, pi02487, pi02488, pi02489, pi02490, pi02491, pi02492, pi02493, pi02494, pi02495, pi02496, pi02497, pi02498, pi02499, pi02500, pi02501, pi02502, pi02503, pi02504, pi02505, pi02506, pi02507, pi02508, pi02509, pi02510, pi02511, pi02512, pi02513, pi02514, pi02515, pi02516, pi02517, pi02518, pi02519, pi02520, pi02521, pi02522, pi02523, pi02524, pi02525, pi02526, pi02527, pi02528, pi02529, pi02530, pi02531, pi02532, pi02533, pi02534, pi02535, pi02536, pi02537, pi02538, pi02539, pi02540, pi02541, pi02542, pi02543, pi02544, pi02545, pi02546, pi02547, pi02548, pi02549, pi02550, pi02551, pi02552, pi02553, pi02554, pi02555, pi02556, pi02557, pi02558, pi02559, pi02560, pi02561, pi02562, pi02563, pi02564, pi02565, pi02566, pi02567, pi02568, pi02569, pi02570, pi02571, pi02572, pi02573, pi02574, pi02575, pi02576, pi02577, pi02578, pi02579, pi02580, pi02581, pi02582, pi02583, pi02584, pi02585, pi02586, pi02587, pi02588, pi02589, pi02590, pi02591, pi02592, pi02593, pi02594, pi02595, pi02596, pi02597, pi02598, pi02599, pi02600, pi02601, pi02602, pi02603, pi02604, pi02605, pi02606, pi02607, pi02608, pi02609, pi02610, pi02611, pi02612, pi02613, pi02614, pi02615, pi02616, pi02617, pi02618, pi02619, pi02620, pi02621, pi02622, pi02623, pi02624, pi02625, pi02626, pi02627, pi02628, pi02629, pi02630, pi02631, pi02632, pi02633, pi02634, pi02635, pi02636, pi02637, pi02638, pi02639, pi02640, pi02641, pi02642, pi02643, pi02644, pi02645, pi02646, pi02647, pi02648, pi02649, pi02650, pi02651, pi02652, pi02653, pi02654, pi02655, pi02656, pi02657, pi02658, pi02659, pi02660, pi02661, pi02662, pi02663, pi02664, pi02665, pi02666, pi02667, pi02668, pi02669, pi02670, pi02671, pi02672, pi02673, pi02674, pi02675, pi02676, pi02677, pi02678, pi02679, pi02680, pi02681, pi02682, pi02683, pi02684, pi02685, pi02686, pi02687, pi02688, pi02689, pi02690, pi02691, pi02692, pi02693, pi02694, pi02695, pi02696, pi02697, pi02698, pi02699, pi02700, pi02701, pi02702, pi02703, pi02704, pi02705, pi02706, pi02707, pi02708, pi02709, pi02710, pi02711, pi02712, pi02713, pi02714, pi02715, pi02716, pi02717, pi02718, pi02719, pi02720, pi02721, pi02722, pi02723, pi02724, pi02725, pi02726, pi02727, pi02728, pi02729, pi02730, pi02731, pi02732, pi02733, pi02734, pi02735, pi02736, pi02737, pi02738, pi02739, pi02740, pi02741, pi02742, pi02743, pi02744, pi02745, pi02746, pi02747, pi02748, pi02749, pi02750, pi02751, pi02752, pi02753, pi02754, pi02755, pi02756, pi02757, pi02758, pi02759, pi02760, pi02761, pi02762, pi02763, pi02764, pi02765, pi02766, pi02767, pi02768, pi02769, pi02770, pi02771, pi02772, pi02773, pi02774, pi02775, pi02776, pi02777, pi02778, pi02779, pi02780, pi02781, pi02782, pi02783, pi02784, pi02785, pi02786, pi02787, pi02788, pi02789, pi02790, pi02791, pi02792, pi02793, pi02794, pi02795, pi02796, pi02797, pi02798, pi02799, pi02800, pi02801, pi02802, pi02803, pi02804, pi02805, pi02806, pi02807, pi02808, pi02809, pi02810, pi02811, pi02812, pi02813, pi02814, pi02815, pi02816, pi02817, pi02818, pi02819, pi02820, pi02821, pi02822, pi02823, pi02824, pi02825, pi02826, pi02827, pi02828, pi02829, pi02830, pi02831, pi02832, pi02833, pi02834, pi02835, pi02836, pi02837, pi02838, pi02839, pi02840, pi02841, pi02842, pi02843, pi02844, pi02845, pi02846, pi02847, pi02848, pi02849, pi02850, pi02851, pi02852, pi02853, pi02854, pi02855, pi02856, pi02857, pi02858, pi02859, pi02860, pi02861, pi02862, pi02863, pi02864, pi02865, pi02866, pi02867, pi02868, pi02869, pi02870, pi02871, pi02872, pi02873, pi02874, pi02875, pi02876, pi02877, pi02878, pi02879, pi02880, pi02881, pi02882, pi02883, pi02884, pi02885, pi02886, pi02887, pi02888, pi02889, pi02890, pi02891, pi02892, pi02893, pi02894, pi02895, pi02896, pi02897, pi02898, pi02899, pi02900, pi02901, pi02902, pi02903, pi02904, pi02905, pi02906, pi02907, pi02908, pi02909, pi02910, pi02911, pi02912, pi02913, pi02914, pi02915, pi02916, pi02917, pi02918, pi02919, pi02920, pi02921, pi02922, pi02923, pi02924, pi02925, pi02926, pi02927, pi02928, pi02929, pi02930, pi02931, pi02932, pi02933, pi02934, pi02935, pi02936, pi02937, pi02938, pi02939, pi02940, pi02941, pi02942, pi02943, pi02944, pi02945, pi02946, pi02947, pi02948, pi02949, pi02950, pi02951, pi02952, pi02953, pi02954, pi02955, pi02956, pi02957, pi02958, pi02959, pi02960, pi02961, pi02962, pi02963, pi02964, pi02965, pi02966, pi02967, pi02968, pi02969, pi02970, pi02971, pi02972, pi02973, pi02974, pi02975, pi02976, pi02977, pi02978, pi02979, pi02980, pi02981, pi02982, pi02983, pi02984, pi02985, pi02986, pi02987, pi02988, pi02989, pi02990, pi02991, pi02992, pi02993, pi02994, pi02995, pi02996, pi02997, pi02998, pi02999, pi03000, pi03001, pi03002, pi03003, pi03004, pi03005, pi03006, pi03007, pi03008, pi03009, pi03010, pi03011, pi03012, pi03013, pi03014, pi03015, pi03016, pi03017, pi03018, pi03019, pi03020, pi03021, pi03022, pi03023, pi03024, pi03025, pi03026, pi03027, pi03028, pi03029, pi03030, pi03031, pi03032, pi03033, pi03034, pi03035, pi03036, pi03037, pi03038, pi03039, pi03040, pi03041, pi03042, pi03043, pi03044, pi03045, pi03046, pi03047, pi03048, pi03049, pi03050, pi03051, pi03052, pi03053, pi03054, pi03055, pi03056, pi03057, pi03058, pi03059, pi03060, pi03061, pi03062, pi03063, pi03064, pi03065, pi03066, pi03067, pi03068, pi03069, pi03070, pi03071, pi03072, pi03073, pi03074, pi03075, pi03076, pi03077, pi03078, pi03079, pi03080, pi03081, pi03082, pi03083, pi03084, pi03085, pi03086, pi03087, pi03088, pi03089, pi03090, pi03091, pi03092, pi03093, pi03094, pi03095, pi03096, pi03097, pi03098, pi03099, pi03100, pi03101, pi03102, pi03103, pi03104, pi03105, pi03106, pi03107, pi03108, pi03109, pi03110, pi03111, pi03112, pi03113, pi03114, pi03115, pi03116, pi03117, pi03118, pi03119, pi03120, pi03121, pi03122, pi03123, pi03124, pi03125, pi03126, pi03127, pi03128, pi03129, pi03130, pi03131, pi03132, pi03133, pi03134, pi03135, pi03136, pi03137, pi03138, pi03139, pi03140, pi03141, pi03142, pi03143, pi03144, pi03145, pi03146, pi03147, pi03148, pi03149, pi03150, pi03151, pi03152, pi03153, pi03154, pi03155, pi03156, pi03157, pi03158, pi03159, pi03160, pi03161, pi03162, pi03163, pi03164, pi03165, pi03166, pi03167, pi03168, pi03169, pi03170, pi03171, pi03172, pi03173, pi03174, pi03175, pi03176, pi03177, pi03178, pi03179, pi03180, pi03181, pi03182, pi03183, pi03184, pi03185, pi03186, pi03187, pi03188, pi03189, pi03190, pi03191, pi03192, pi03193, pi03194, pi03195, pi03196, pi03197, pi03198, pi03199, pi03200, pi03201, pi03202, pi03203, pi03204, pi03205, pi03206, pi03207, pi03208, pi03209, pi03210, pi03211, pi03212, pi03213, pi03214, pi03215, pi03216, pi03217, pi03218, pi03219, pi03220, pi03221, pi03222, pi03223, pi03224, pi03225, pi03226, pi03227, pi03228, pi03229, pi03230, pi03231, pi03232, pi03233, pi03234, pi03235, pi03236, pi03237, pi03238, pi03239, pi03240, pi03241, pi03242, pi03243, pi03244, pi03245, pi03246, pi03247, pi03248, pi03249, pi03250, pi03251, pi03252, pi03253, pi03254, pi03255, pi03256, pi03257, pi03258, pi03259, pi03260, pi03261, pi03262, pi03263, pi03264, pi03265, pi03266, pi03267, pi03268, pi03269, pi03270, pi03271, pi03272, pi03273, pi03274, pi03275, pi03276, pi03277, pi03278, pi03279, pi03280, pi03281, pi03282, pi03283, pi03284, pi03285, pi03286, pi03287, pi03288, pi03289, pi03290, pi03291, pi03292, pi03293, pi03294, pi03295, pi03296, pi03297, pi03298, pi03299, pi03300, pi03301, pi03302, pi03303, pi03304, pi03305, pi03306, pi03307, pi03308, pi03309, pi03310, pi03311, pi03312, pi03313, pi03314, pi03315, pi03316, pi03317, pi03318, pi03319, pi03320, pi03321, pi03322, pi03323, pi03324, pi03325, pi03326, pi03327, pi03328, pi03329, pi03330, pi03331, pi03332, pi03333, pi03334, pi03335, pi03336, pi03337, pi03338, pi03339, pi03340, pi03341, pi03342, pi03343, pi03344, pi03345, pi03346, pi03347, pi03348, pi03349, pi03350, pi03351, pi03352, pi03353, pi03354, pi03355, pi03356, pi03357, pi03358, pi03359, pi03360, pi03361, pi03362, pi03363, pi03364, pi03365, pi03366, pi03367, pi03368, pi03369, pi03370, pi03371, pi03372, pi03373, pi03374, pi03375, pi03376, pi03377, pi03378, pi03379, pi03380, pi03381, pi03382, pi03383, pi03384, pi03385, pi03386, pi03387, pi03388, pi03389, pi03390, pi03391, pi03392, pi03393, pi03394, pi03395, pi03396, pi03397, pi03398, pi03399, pi03400, pi03401, pi03402, pi03403, pi03404, pi03405, pi03406, pi03407, pi03408, pi03409, pi03410, pi03411, pi03412, pi03413, pi03414, pi03415, pi03416, pi03417, pi03418, pi03419, pi03420, pi03421, pi03422, pi03423, pi03424, pi03425, pi03426, pi03427, pi03428, pi03429, pi03430, pi03431, pi03432, pi03433, pi03434, pi03435, pi03436, pi03437, pi03438, pi03439, pi03440, pi03441, pi03442, pi03443, pi03444, pi03445, pi03446, pi03447, pi03448, pi03449, pi03450, pi03451, pi03452, pi03453, pi03454, pi03455, pi03456, pi03457, pi03458, pi03459, pi03460, pi03461, pi03462, pi03463, pi03464, pi03465, pi03466, pi03467, pi03468, pi03469, pi03470, pi03471, pi03472, pi03473, pi03474, pi03475, pi03476, pi03477, pi03478, pi03479, pi03480, pi03481, pi03482, pi03483, pi03484, pi03485, pi03486, pi03487, pi03488, pi03489, pi03490, pi03491, pi03492, pi03493, pi03494, pi03495, pi03496, pi03497, pi03498, pi03499, pi03500, pi03501, pi03502, pi03503, pi03504, pi03505, pi03506, pi03507, pi03508, pi03509, pi03510, pi03511, pi03512, pi03513, pi03514, pi03515, pi03516, pi03517, pi03518, pi03519, pi03520, pi03521, pi03522, pi03523, pi03524, pi03525, pi03526, pi03527, pi03528, pi03529, pi03530, pi03531, pi03532, pi03533, pi03534, pi03535, pi03536, pi03537, pi03538, pi03539, pi03540, pi03541, pi03542, pi03543, pi03544, pi03545, pi03546, pi03547, pi03548, pi03549, pi03550, pi03551, pi03552, pi03553, pi03554, pi03555, pi03556, pi03557, pi03558, pi03559, pi03560, pi03561, pi03562, pi03563, pi03564, pi03565, pi03566, pi03567, pi03568, pi03569, pi03570, pi03571, pi03572, pi03573, pi03574, pi03575, pi03576, pi03577, pi03578, pi03579, pi03580, pi03581, pi03582, pi03583, pi03584, pi03585, pi03586, pi03587, pi03588, pi03589, pi03590, pi03591, pi03592, pi03593, pi03594, pi03595, pi03596, pi03597, pi03598, pi03599, pi03600, pi03601, pi03602, pi03603, pi03604, pi03605, pi03606, pi03607, pi03608, pi03609, pi03610, pi03611, pi03612, pi03613, pi03614, pi03615, pi03616, pi03617, pi03618, pi03619, pi03620, pi03621, pi03622, pi03623, pi03624, pi03625, pi03626, pi03627, pi03628, pi03629, pi03630, pi03631, pi03632, pi03633, pi03634, pi03635, pi03636, pi03637, pi03638, pi03639, pi03640, pi03641, pi03642, pi03643, pi03644, pi03645, pi03646, pi03647, pi03648, pi03649, pi03650, pi03651, pi03652, pi03653, pi03654, pi03655, pi03656, pi03657, pi03658, pi03659, pi03660, pi03661, pi03662, pi03663, pi03664, pi03665, pi03666, pi03667, pi03668, pi03669, pi03670, pi03671, pi03672, pi03673, pi03674, pi03675, pi03676, pi03677, pi03678, pi03679, pi03680, pi03681, pi03682, pi03683, pi03684, pi03685, pi03686, pi03687, pi03688, pi03689, pi03690, pi03691, pi03692, pi03693, pi03694, pi03695, pi03696, pi03697, pi03698, pi03699, pi03700, pi03701, pi03702, pi03703, pi03704, pi03705, pi03706, pi03707, pi03708, pi03709, pi03710, pi03711, pi03712, pi03713, pi03714, pi03715, pi03716, pi03717, pi03718, pi03719, pi03720, pi03721, pi03722, pi03723, pi03724, pi03725, pi03726, pi03727, pi03728, pi03729, pi03730, pi03731, pi03732, pi03733, pi03734, pi03735, pi03736, pi03737, pi03738, pi03739, pi03740, pi03741, pi03742, pi03743, pi03744, pi03745, pi03746, pi03747, pi03748, pi03749, pi03750, pi03751, pi03752, pi03753, pi03754, pi03755, pi03756, pi03757, pi03758, pi03759, pi03760, pi03761, pi03762, pi03763, pi03764, pi03765, pi03766, pi03767, pi03768, pi03769, pi03770, pi03771, pi03772, pi03773, pi03774, pi03775, pi03776, pi03777, pi03778, pi03779, pi03780, pi03781, pi03782, pi03783, pi03784, pi03785, pi03786, pi03787, pi03788, pi03789, pi03790, pi03791, pi03792, pi03793, pi03794, pi03795, pi03796, pi03797, pi03798, pi03799, pi03800, pi03801, pi03802, pi03803, pi03804, pi03805, pi03806, pi03807, pi03808, pi03809, pi03810, pi03811, pi03812, pi03813, pi03814, pi03815, pi03816, pi03817, pi03818, pi03819, pi03820, pi03821, pi03822, pi03823, pi03824, pi03825, pi03826, pi03827, pi03828, pi03829, pi03830, pi03831, pi03832, pi03833, pi03834, pi03835, pi03836, pi03837, pi03838, pi03839, pi03840, pi03841, pi03842, pi03843, pi03844, pi03845, pi03846, pi03847, pi03848, pi03849, pi03850, pi03851, pi03852, pi03853, pi03854, pi03855, pi03856, pi03857, pi03858, pi03859, pi03860, pi03861, pi03862, pi03863, pi03864, pi03865, pi03866, pi03867, pi03868, pi03869, pi03870, pi03871, pi03872, pi03873, pi03874, pi03875, pi03876, pi03877, pi03878, pi03879, pi03880, pi03881, pi03882, pi03883, pi03884, pi03885, pi03886, pi03887, pi03888, pi03889, pi03890, pi03891, pi03892, pi03893, pi03894, pi03895, pi03896, pi03897, pi03898, pi03899, pi03900, pi03901, pi03902, pi03903, pi03904, pi03905, pi03906, pi03907, pi03908, pi03909, pi03910, pi03911, pi03912, pi03913, pi03914, pi03915, pi03916, pi03917, pi03918, pi03919, pi03920, pi03921, pi03922, pi03923, pi03924, pi03925, pi03926, pi03927, pi03928, pi03929, pi03930, pi03931, pi03932, pi03933, pi03934, pi03935, pi03936, pi03937, pi03938, pi03939, pi03940, pi03941, pi03942, pi03943, pi03944, pi03945, pi03946, pi03947, pi03948, pi03949, pi03950, pi03951, pi03952, pi03953, pi03954, pi03955, pi03956, pi03957, pi03958, pi03959, pi03960, pi03961, pi03962, pi03963, pi03964, pi03965, pi03966, pi03967, pi03968, pi03969, pi03970, pi03971, pi03972, pi03973, pi03974, pi03975, pi03976, pi03977, pi03978, pi03979, pi03980, pi03981, pi03982, pi03983, pi03984, pi03985, pi03986, pi03987, pi03988, pi03989, pi03990, pi03991, pi03992, pi03993, pi03994, pi03995, pi03996, pi03997, pi03998, pi03999, pi04000, pi04001, pi04002, pi04003, pi04004, pi04005, pi04006, pi04007, pi04008, pi04009, pi04010, pi04011, pi04012, pi04013, pi04014, pi04015, pi04016, pi04017, pi04018, pi04019, pi04020, pi04021, pi04022, pi04023, pi04024, pi04025, pi04026, pi04027, pi04028, pi04029, pi04030, pi04031, pi04032, pi04033, pi04034, pi04035, pi04036, pi04037, pi04038, pi04039, pi04040, pi04041, pi04042, pi04043, pi04044, pi04045, pi04046, pi04047, pi04048, pi04049, pi04050, pi04051, pi04052, pi04053, pi04054, pi04055, pi04056, pi04057, pi04058, pi04059, pi04060, pi04061, pi04062, pi04063, pi04064, pi04065, pi04066, pi04067, pi04068, pi04069, pi04070, pi04071, pi04072, pi04073, pi04074, pi04075, pi04076, pi04077, pi04078, pi04079, pi04080, pi04081, pi04082, pi04083, pi04084, pi04085, pi04086, pi04087, pi04088, pi04089, pi04090, pi04091, pi04092, pi04093, pi04094, pi04095, pi04096, pi04097, pi04098, pi04099, pi04100, pi04101, pi04102, pi04103, pi04104, pi04105, pi04106, pi04107, pi04108, pi04109, pi04110, pi04111, pi04112, pi04113, pi04114, pi04115, pi04116, pi04117, pi04118, pi04119, pi04120, pi04121, pi04122, pi04123, pi04124, pi04125, pi04126, pi04127, pi04128, pi04129, pi04130, pi04131, pi04132, pi04133, pi04134, pi04135, pi04136, pi04137, pi04138, pi04139, pi04140, pi04141, pi04142, pi04143, pi04144, pi04145, pi04146, pi04147, pi04148, pi04149, pi04150, pi04151, pi04152, pi04153, pi04154, pi04155, pi04156, pi04157, pi04158, pi04159, pi04160, pi04161, pi04162, pi04163, pi04164, pi04165, pi04166, pi04167, pi04168, pi04169, pi04170, pi04171, pi04172, pi04173, pi04174, pi04175, pi04176, pi04177, pi04178, pi04179, pi04180, pi04181, pi04182, pi04183, pi04184, pi04185, pi04186, pi04187, pi04188, pi04189, pi04190, pi04191, pi04192, pi04193, pi04194, pi04195, pi04196, pi04197, pi04198, pi04199, pi04200, pi04201, pi04202, pi04203, pi04204, pi04205, pi04206, pi04207, pi04208, pi04209, pi04210, pi04211, pi04212, pi04213, pi04214, pi04215, pi04216, pi04217, pi04218, pi04219, pi04220, pi04221, pi04222, pi04223, pi04224, pi04225, pi04226, pi04227, pi04228, pi04229, pi04230, pi04231, pi04232, pi04233, pi04234, pi04235, pi04236, pi04237, pi04238, pi04239, pi04240, pi04241, pi04242, pi04243, pi04244, pi04245, pi04246, pi04247, pi04248, pi04249, pi04250, pi04251, pi04252, pi04253, pi04254, pi04255, pi04256, pi04257, pi04258, pi04259, pi04260, pi04261, pi04262, pi04263, pi04264, pi04265, pi04266, pi04267, pi04268, pi04269, pi04270, pi04271, pi04272, pi04273, pi04274, pi04275, pi04276, pi04277, pi04278, pi04279, pi04280, pi04281, pi04282, pi04283, pi04284, pi04285, pi04286, pi04287, pi04288, pi04289, pi04290, pi04291, pi04292, pi04293, pi04294, pi04295, pi04296, pi04297, pi04298, pi04299, pi04300, pi04301, pi04302, pi04303, pi04304, pi04305, pi04306, pi04307, pi04308, pi04309, pi04310, pi04311, pi04312, pi04313, pi04314, pi04315, pi04316, pi04317, pi04318, pi04319, pi04320, pi04321, pi04322, pi04323, pi04324, pi04325, pi04326, pi04327, pi04328, pi04329, pi04330, pi04331, pi04332, pi04333, pi04334, pi04335, pi04336, pi04337, pi04338, pi04339, pi04340, pi04341, pi04342, pi04343, pi04344, pi04345, pi04346, pi04347, pi04348, pi04349, pi04350, pi04351, pi04352, pi04353, pi04354, pi04355, pi04356, pi04357, pi04358, pi04359, pi04360, pi04361, pi04362, pi04363, pi04364, pi04365, pi04366, pi04367, pi04368, pi04369, pi04370, pi04371, pi04372, pi04373, pi04374, pi04375, pi04376, pi04377, pi04378, pi04379, pi04380, pi04381, pi04382, pi04383, pi04384, pi04385, pi04386, pi04387, pi04388, pi04389, pi04390, pi04391, pi04392, pi04393, pi04394, pi04395, pi04396, pi04397, pi04398, pi04399, pi04400, pi04401, pi04402, pi04403, pi04404, pi04405, pi04406, pi04407, pi04408, pi04409, pi04410, pi04411, pi04412, pi04413, pi04414, pi04415, pi04416, pi04417, pi04418, pi04419, pi04420, pi04421, pi04422, pi04423, pi04424, pi04425, pi04426, pi04427, pi04428, pi04429, pi04430, pi04431, pi04432, pi04433, pi04434, pi04435, pi04436, pi04437, pi04438, pi04439, pi04440, pi04441, pi04442, pi04443, pi04444, pi04445, pi04446, pi04447, pi04448, pi04449, pi04450, pi04451, pi04452, pi04453, pi04454, pi04455, pi04456, pi04457, pi04458, pi04459, pi04460, pi04461, pi04462, pi04463, pi04464, pi04465, pi04466, pi04467, pi04468, pi04469, pi04470, pi04471, pi04472, pi04473, pi04474, pi04475, pi04476, pi04477, pi04478, pi04479, pi04480, pi04481, pi04482, pi04483, pi04484, pi04485, pi04486, pi04487, pi04488, pi04489, pi04490, pi04491, pi04492, pi04493, pi04494, pi04495, pi04496, pi04497, pi04498, pi04499, pi04500, pi04501, pi04502, pi04503, pi04504, pi04505, pi04506, pi04507, pi04508, pi04509, pi04510, pi04511, pi04512, pi04513, pi04514, pi04515, pi04516, pi04517, pi04518, pi04519, pi04520, pi04521, pi04522, pi04523, pi04524, pi04525, pi04526, pi04527, pi04528, pi04529, pi04530, pi04531, pi04532, pi04533, pi04534, pi04535, pi04536, pi04537, pi04538, pi04539, pi04540, pi04541, pi04542, pi04543, pi04544, pi04545, pi04546, pi04547, pi04548, pi04549, pi04550, pi04551, pi04552, pi04553, pi04554, pi04555, pi04556, pi04557, pi04558, pi04559, pi04560, pi04561, pi04562, pi04563, pi04564, pi04565, pi04566, pi04567, pi04568, pi04569, pi04570, pi04571, pi04572, pi04573, pi04574, pi04575, pi04576, pi04577, pi04578, pi04579, pi04580, pi04581, pi04582, pi04583, pi04584, pi04585, pi04586, pi04587, pi04588, pi04589, pi04590, pi04591, pi04592, pi04593, pi04594, pi04595, pi04596, pi04597, pi04598, pi04599, pi04600, pi04601, pi04602, pi04603, pi04604, pi04605, pi04606, pi04607, pi04608, pi04609, pi04610, pi04611, pi04612, pi04613, pi04614, pi04615, pi04616, pi04617, pi04618, pi04619, pi04620, pi04621, pi04622, pi04623, pi04624, pi04625, pi04626, pi04627, pi04628, pi04629, pi04630, pi04631, pi04632, pi04633, pi04634, pi04635, pi04636, pi04637, pi04638, pi04639, pi04640, pi04641, pi04642, pi04643, pi04644, pi04645, pi04646, pi04647, pi04648, pi04649, pi04650, pi04651, pi04652, pi04653, pi04654, pi04655, pi04656, pi04657, pi04658, pi04659, pi04660, pi04661, pi04662, pi04663, pi04664, pi04665, pi04666, pi04667, pi04668, pi04669, pi04670, pi04671, pi04672, pi04673, pi04674, pi04675, pi04676, pi04677, pi04678, pi04679, pi04680, pi04681, pi04682, pi04683, pi04684, pi04685, pi04686, pi04687, pi04688, pi04689, pi04690, pi04691, pi04692, pi04693, pi04694, pi04695, pi04696, pi04697, pi04698, pi04699, pi04700, pi04701, pi04702, pi04703, pi04704, pi04705, pi04706, pi04707, pi04708, pi04709, pi04710, pi04711, pi04712, pi04713, pi04714, pi04715, pi04716, pi04717, pi04718, pi04719, pi04720, pi04721, pi04722, pi04723, pi04724, pi04725, pi04726, pi04727, pi04728, pi04729, pi04730, pi04731, pi04732, pi04733, pi04734, pi04735, pi04736, pi04737, pi04738, pi04739, pi04740, pi04741, pi04742, pi04743, pi04744, pi04745, pi04746, pi04747, pi04748, pi04749, pi04750, pi04751, pi04752, pi04753, pi04754, pi04755, pi04756, pi04757, pi04758, pi04759, pi04760, pi04761, pi04762, pi04763, pi04764, pi04765, pi04766, pi04767, pi04768, pi04769, pi04770, pi04771, pi04772, pi04773, pi04774, pi04775, pi04776, pi04777, pi04778, pi04779, pi04780, pi04781, pi04782, pi04783, pi04784, pi04785, pi04786, pi04787, pi04788, pi04789, pi04790, pi04791, pi04792, pi04793, pi04794, pi04795, pi04796, pi04797, pi04798, pi04799, pi04800, pi04801, pi04802, pi04803, pi04804, pi04805, pi04806, pi04807, pi04808, pi04809, pi04810, pi04811, pi04812, pi04813, pi04814, pi04815, pi04816, pi04817, pi04818, pi04819, pi04820, pi04821, pi04822, pi04823, pi04824, pi04825, pi04826, pi04827, pi04828, pi04829, pi04830, pi04831, pi04832, pi04833, pi04834, pi04835, pi04836, pi04837, pi04838, pi04839, pi04840, pi04841, pi04842, pi04843, pi04844, pi04845, pi04846, pi04847, pi04848, pi04849, pi04850, pi04851, pi04852, pi04853, pi04854, pi04855, pi04856, pi04857, pi04858, pi04859, pi04860, pi04861, pi04862, pi04863, pi04864, pi04865, pi04866, pi04867, pi04868, pi04869, pi04870, pi04871, pi04872, pi04873, pi04874, pi04875, pi04876, pi04877, pi04878, pi04879, pi04880, pi04881, pi04882, pi04883, pi04884, pi04885, pi04886, pi04887, pi04888, pi04889, pi04890, pi04891, pi04892, pi04893, pi04894, pi04895, pi04896, pi04897, pi04898, pi04899, pi04900, pi04901, pi04902, pi04903, pi04904, pi04905, pi04906, pi04907, pi04908, pi04909, pi04910, pi04911, pi04912, pi04913, pi04914, pi04915, pi04916, pi04917, pi04918, pi04919, pi04920, pi04921, pi04922, pi04923, pi04924, pi04925, pi04926, pi04927, pi04928, pi04929, pi04930, pi04931, pi04932, pi04933, pi04934, pi04935, pi04936, pi04937, pi04938, pi04939, pi04940, pi04941, pi04942, pi04943, pi04944, pi04945, pi04946, pi04947, pi04948, pi04949, pi04950, pi04951, pi04952, pi04953, pi04954, pi04955, pi04956, pi04957, pi04958, pi04959, pi04960, pi04961, pi04962, pi04963, pi04964, pi04965, pi04966, pi04967, pi04968, pi04969, pi04970, pi04971, pi04972, pi04973, pi04974, pi04975, pi04976, pi04977, pi04978, pi04979, pi04980, pi04981, pi04982, pi04983, pi04984, pi04985, pi04986, pi04987, pi04988, pi04989, pi04990, pi04991, pi04992, pi04993, pi04994, pi04995, pi04996, pi04997, pi04998, pi04999, pi05000, pi05001, pi05002, pi05003, pi05004, pi05005, pi05006, pi05007, pi05008, pi05009, pi05010, pi05011, pi05012, pi05013, pi05014, pi05015, pi05016, pi05017, pi05018, pi05019, pi05020, pi05021, pi05022, pi05023, pi05024, pi05025, pi05026, pi05027, pi05028, pi05029, pi05030, pi05031, pi05032, pi05033, pi05034, pi05035, pi05036, pi05037, pi05038, pi05039, pi05040, pi05041, pi05042, pi05043, pi05044, pi05045, pi05046, pi05047, pi05048, pi05049, pi05050, pi05051, pi05052, pi05053, pi05054, pi05055, pi05056, pi05057, pi05058, pi05059, pi05060, pi05061, pi05062, pi05063, pi05064, pi05065, pi05066, pi05067, pi05068, pi05069, pi05070, pi05071, pi05072, pi05073, pi05074, pi05075, pi05076, pi05077, pi05078, pi05079, pi05080, pi05081, pi05082, pi05083, pi05084, pi05085, pi05086, pi05087, pi05088, pi05089, pi05090, pi05091, pi05092, pi05093, pi05094, pi05095, pi05096, pi05097, pi05098, pi05099, pi05100, pi05101, pi05102, pi05103, pi05104, pi05105, pi05106, pi05107, pi05108, pi05109, pi05110, pi05111, pi05112, pi05113, pi05114, pi05115, pi05116, pi05117, pi05118, pi05119, pi05120, pi05121, pi05122, pi05123, pi05124, pi05125, pi05126, pi05127, pi05128, pi05129, pi05130, pi05131, pi05132, pi05133, pi05134, pi05135, pi05136, pi05137, pi05138, pi05139, pi05140, pi05141, pi05142, pi05143, pi05144, pi05145, pi05146, pi05147, pi05148, pi05149, pi05150, pi05151, pi05152, pi05153, pi05154, pi05155, pi05156, pi05157, pi05158, pi05159, pi05160, pi05161, pi05162, pi05163, pi05164, pi05165, pi05166, pi05167, pi05168, pi05169, pi05170, pi05171, pi05172, pi05173, pi05174, pi05175, pi05176, pi05177, pi05178, pi05179, pi05180, pi05181, pi05182, pi05183, pi05184, pi05185, pi05186, pi05187, pi05188, pi05189, pi05190, pi05191, pi05192, pi05193, pi05194, pi05195, pi05196, pi05197, pi05198, pi05199, pi05200, pi05201, pi05202, pi05203, pi05204, pi05205, pi05206, pi05207, pi05208, pi05209, pi05210, pi05211, pi05212, pi05213, pi05214, pi05215, pi05216, pi05217, pi05218, pi05219, pi05220, pi05221, pi05222, pi05223, pi05224, pi05225, pi05226, pi05227, pi05228, pi05229, pi05230, pi05231, pi05232, pi05233, pi05234, pi05235, pi05236, pi05237, pi05238, pi05239, pi05240, pi05241, pi05242, pi05243, pi05244, pi05245, pi05246, pi05247, pi05248, pi05249, pi05250, pi05251, pi05252, pi05253, pi05254, pi05255, pi05256, pi05257, pi05258, pi05259, pi05260, pi05261, pi05262, pi05263, pi05264, pi05265, pi05266, pi05267, pi05268, pi05269, pi05270, pi05271, pi05272, pi05273, pi05274, pi05275, pi05276, pi05277, pi05278, pi05279, pi05280, pi05281, pi05282, pi05283, pi05284, pi05285, pi05286, pi05287, pi05288, pi05289, pi05290, pi05291, pi05292, pi05293, pi05294, pi05295, pi05296, pi05297, pi05298, pi05299, pi05300, pi05301, pi05302, pi05303, pi05304, pi05305, pi05306, pi05307, pi05308, pi05309, pi05310, pi05311, pi05312, pi05313, pi05314, pi05315, pi05316, pi05317, pi05318, pi05319, pi05320, pi05321, pi05322, pi05323, pi05324, pi05325, pi05326, pi05327, pi05328, pi05329, pi05330, pi05331, pi05332, pi05333, pi05334, pi05335, pi05336, pi05337, pi05338, pi05339, pi05340, pi05341, pi05342, pi05343, pi05344, pi05345, pi05346, pi05347, pi05348, pi05349, pi05350, pi05351, pi05352, pi05353, pi05354, pi05355, pi05356, pi05357, pi05358, pi05359, pi05360, pi05361, pi05362, pi05363, pi05364, pi05365, pi05366, pi05367, pi05368, pi05369, pi05370, pi05371, pi05372, pi05373, pi05374, pi05375, pi05376, pi05377, pi05378, pi05379, pi05380, pi05381, pi05382, pi05383, pi05384, pi05385, pi05386, pi05387, pi05388, pi05389, pi05390, pi05391, pi05392, pi05393, pi05394, pi05395, pi05396, pi05397, pi05398, pi05399, pi05400, pi05401, pi05402, pi05403, pi05404, pi05405, pi05406, pi05407, pi05408, pi05409, pi05410, pi05411, pi05412, pi05413, pi05414, pi05415, pi05416, pi05417, pi05418, pi05419, pi05420, pi05421, pi05422, pi05423, pi05424, pi05425, pi05426, pi05427, pi05428, pi05429, pi05430, pi05431, pi05432, pi05433, pi05434, pi05435, pi05436, pi05437, pi05438, pi05439, pi05440, pi05441, pi05442, pi05443, pi05444, pi05445, pi05446, pi05447, pi05448, pi05449, pi05450, pi05451, pi05452, pi05453, pi05454, pi05455, pi05456, pi05457, pi05458, pi05459, pi05460, pi05461, pi05462, pi05463, pi05464, pi05465, pi05466, pi05467, pi05468, pi05469, pi05470, pi05471, pi05472, pi05473, pi05474, pi05475, pi05476, pi05477, pi05478, pi05479, pi05480, pi05481, pi05482, pi05483, pi05484, pi05485, pi05486, pi05487, pi05488, pi05489, pi05490, pi05491, pi05492, pi05493, pi05494, pi05495, pi05496, pi05497, pi05498, pi05499, pi05500, pi05501, pi05502, pi05503, pi05504, pi05505, pi05506, pi05507, pi05508, pi05509, pi05510, pi05511, pi05512, pi05513, pi05514, pi05515, pi05516, pi05517, pi05518, pi05519, pi05520, pi05521, pi05522, pi05523, pi05524, pi05525, pi05526, pi05527, pi05528, pi05529, pi05530, pi05531, pi05532, pi05533, pi05534, pi05535, pi05536, pi05537, pi05538, pi05539, pi05540, pi05541, pi05542, pi05543, pi05544, pi05545, pi05546, pi05547, pi05548, pi05549, pi05550, pi05551, pi05552, pi05553, pi05554, pi05555, pi05556, pi05557, pi05558, pi05559, pi05560, pi05561, pi05562, pi05563, pi05564, pi05565, pi05566, pi05567, pi05568, pi05569, pi05570, pi05571, pi05572, pi05573, pi05574, pi05575, pi05576, pi05577, pi05578, pi05579, pi05580, pi05581, pi05582, pi05583, pi05584, pi05585, pi05586, pi05587, pi05588, pi05589, pi05590, pi05591, pi05592, pi05593, pi05594, pi05595, pi05596, pi05597, pi05598, pi05599, pi05600, pi05601, pi05602, pi05603, pi05604, pi05605, pi05606, pi05607, pi05608, pi05609, pi05610, pi05611, pi05612, pi05613, pi05614, pi05615, pi05616, pi05617, pi05618, pi05619, pi05620, pi05621, pi05622, pi05623, pi05624, pi05625, pi05626, pi05627, pi05628, pi05629, pi05630, pi05631, pi05632, pi05633, pi05634, pi05635, pi05636, pi05637, pi05638, pi05639, pi05640, pi05641, pi05642, pi05643, pi05644, pi05645, pi05646, pi05647, pi05648, pi05649, pi05650, pi05651, pi05652, pi05653, pi05654, pi05655, pi05656, pi05657, pi05658, pi05659, pi05660, pi05661, pi05662, pi05663, pi05664, pi05665, pi05666, pi05667, pi05668, pi05669, pi05670, pi05671, pi05672, pi05673, pi05674, pi05675, pi05676, pi05677, pi05678, pi05679, pi05680, pi05681, pi05682, pi05683, pi05684, pi05685, pi05686, pi05687, pi05688, pi05689, pi05690, pi05691, pi05692, pi05693, pi05694, pi05695, pi05696, pi05697, pi05698, pi05699, pi05700, pi05701, pi05702, pi05703, pi05704, pi05705, pi05706, pi05707, pi05708, pi05709, pi05710, pi05711, pi05712, pi05713, pi05714, pi05715, pi05716, pi05717, pi05718, pi05719, pi05720, pi05721, pi05722, pi05723, pi05724, pi05725, pi05726, pi05727, pi05728, pi05729, pi05730, pi05731, pi05732, pi05733, pi05734, pi05735, pi05736, pi05737, pi05738, pi05739, pi05740, pi05741, pi05742, pi05743, pi05744, pi05745, pi05746, pi05747, pi05748, pi05749, pi05750, pi05751, pi05752, pi05753, pi05754, pi05755, pi05756, pi05757, pi05758, pi05759, pi05760, pi05761, pi05762, pi05763, pi05764, pi05765, pi05766, pi05767, pi05768, pi05769, pi05770, pi05771, pi05772, pi05773, pi05774, pi05775, pi05776, pi05777, pi05778, pi05779, pi05780, pi05781, pi05782, pi05783, pi05784, pi05785, pi05786, pi05787, pi05788, pi05789, pi05790, pi05791, pi05792, pi05793, pi05794, pi05795, pi05796, pi05797, pi05798, pi05799, pi05800, pi05801, pi05802, pi05803, pi05804, pi05805, pi05806, pi05807, pi05808, pi05809, pi05810, pi05811, pi05812, pi05813, pi05814, pi05815, pi05816, pi05817, pi05818, pi05819, pi05820, pi05821, pi05822, pi05823, pi05824, pi05825, pi05826, pi05827, pi05828, pi05829, pi05830, pi05831, pi05832, pi05833, pi05834, pi05835, pi05836, pi05837, pi05838, pi05839, pi05840, pi05841, pi05842, pi05843, pi05844, pi05845, pi05846, pi05847, pi05848, pi05849, pi05850, pi05851, pi05852, pi05853, pi05854, pi05855, pi05856, pi05857, pi05858, pi05859, pi05860, pi05861, pi05862, pi05863, pi05864, pi05865, pi05866, pi05867, pi05868, pi05869, pi05870, pi05871, pi05872, pi05873, pi05874, pi05875, pi05876, pi05877, pi05878, pi05879, pi05880, pi05881, pi05882, pi05883, pi05884, pi05885, pi05886, pi05887, pi05888, pi05889, pi05890, pi05891, pi05892, pi05893, pi05894, pi05895, pi05896, pi05897, pi05898, pi05899, pi05900, pi05901, pi05902, pi05903, pi05904, pi05905, pi05906, pi05907, pi05908, pi05909, pi05910, pi05911, pi05912, pi05913, pi05914, pi05915, pi05916, pi05917, pi05918, pi05919, pi05920, pi05921, pi05922, pi05923, pi05924, pi05925, pi05926, pi05927, pi05928, pi05929, pi05930, pi05931, pi05932, pi05933, pi05934, pi05935, pi05936, pi05937, pi05938, pi05939, pi05940, pi05941, pi05942, pi05943, pi05944, pi05945, pi05946, pi05947, pi05948, pi05949, pi05950, pi05951, pi05952, pi05953, pi05954, pi05955, pi05956, pi05957, pi05958, pi05959, pi05960, pi05961, pi05962, pi05963, pi05964, pi05965, pi05966, pi05967, pi05968, pi05969, pi05970, pi05971, pi05972, pi05973, pi05974, pi05975, pi05976, pi05977, pi05978, pi05979, pi05980, pi05981, pi05982, pi05983, pi05984, pi05985, pi05986, pi05987, pi05988, pi05989, pi05990, pi05991, pi05992, pi05993, pi05994, pi05995, pi05996, pi05997, pi05998, pi05999, pi06000, pi06001, pi06002, pi06003, pi06004, pi06005, pi06006, pi06007, pi06008, pi06009, pi06010, pi06011, pi06012, pi06013, pi06014, pi06015, pi06016, pi06017, pi06018, pi06019, pi06020, pi06021, pi06022, pi06023, pi06024, pi06025, pi06026, pi06027, pi06028, pi06029, pi06030, pi06031, pi06032, pi06033, pi06034, pi06035, pi06036, pi06037, pi06038, pi06039, pi06040, pi06041, pi06042, pi06043, pi06044, pi06045, pi06046, pi06047, pi06048, pi06049, pi06050, pi06051, pi06052, pi06053, pi06054, pi06055, pi06056, pi06057, pi06058, pi06059, pi06060, pi06061, pi06062, pi06063, pi06064, pi06065, pi06066, pi06067, pi06068, pi06069, pi06070, pi06071, pi06072, pi06073, pi06074, pi06075, pi06076, pi06077, pi06078, pi06079, pi06080, pi06081, pi06082, pi06083, pi06084, pi06085, pi06086, pi06087, pi06088, pi06089, pi06090, pi06091, pi06092, pi06093, pi06094, pi06095, pi06096, pi06097, pi06098, pi06099, pi06100, pi06101, pi06102, pi06103, pi06104, pi06105, pi06106, pi06107, pi06108, pi06109, pi06110, pi06111, pi06112, pi06113, pi06114, pi06115, pi06116, pi06117, pi06118, pi06119, pi06120, pi06121, pi06122, pi06123, pi06124, pi06125, pi06126, pi06127, pi06128, pi06129, pi06130, pi06131, pi06132, pi06133, pi06134, pi06135, pi06136, pi06137, pi06138, pi06139, pi06140, pi06141, pi06142, pi06143, pi06144, pi06145, pi06146, pi06147, pi06148, pi06149, pi06150, pi06151, pi06152, pi06153, pi06154, pi06155, pi06156, pi06157, pi06158, pi06159, pi06160, pi06161, pi06162, pi06163, pi06164, pi06165, pi06166, pi06167, pi06168, pi06169, pi06170, pi06171, pi06172, pi06173, pi06174, pi06175, pi06176, pi06177, pi06178, pi06179, pi06180, pi06181, pi06182, pi06183, pi06184, pi06185, pi06186, pi06187, pi06188, pi06189, pi06190, pi06191, pi06192, pi06193, pi06194, pi06195, pi06196, pi06197, pi06198, pi06199, pi06200, pi06201, pi06202, pi06203, pi06204, pi06205, pi06206, pi06207, pi06208, pi06209, pi06210, pi06211, pi06212, pi06213, pi06214, pi06215, pi06216, pi06217, pi06218, pi06219, pi06220, pi06221, pi06222, pi06223, pi06224, pi06225, pi06226, pi06227, pi06228, pi06229, pi06230, pi06231, pi06232, pi06233, pi06234, pi06235, pi06236, pi06237, pi06238, pi06239, pi06240, pi06241, pi06242, pi06243, pi06244, pi06245, pi06246, pi06247, pi06248, pi06249, pi06250, pi06251, pi06252, pi06253, pi06254, pi06255, pi06256, pi06257, pi06258, pi06259, pi06260, pi06261, pi06262, pi06263, pi06264, pi06265, pi06266, pi06267, pi06268, pi06269, pi06270, pi06271, pi06272, pi06273, pi06274, pi06275, pi06276, pi06277, pi06278, pi06279, pi06280, pi06281, pi06282, pi06283, pi06284, pi06285, pi06286, pi06287, pi06288, pi06289, pi06290, pi06291, pi06292, pi06293, pi06294, pi06295, pi06296, pi06297, pi06298, pi06299, pi06300, pi06301, pi06302, pi06303, pi06304, pi06305, pi06306, pi06307, pi06308, pi06309, pi06310, pi06311, pi06312, pi06313, pi06314, pi06315, pi06316, pi06317, pi06318, pi06319, pi06320, pi06321, pi06322, pi06323, pi06324, pi06325, pi06326, pi06327, pi06328, pi06329, pi06330, pi06331, pi06332, pi06333, pi06334, pi06335, pi06336, pi06337, pi06338, pi06339, pi06340, pi06341, pi06342, pi06343, pi06344, pi06345, pi06346, pi06347, pi06348, pi06349, pi06350, pi06351, pi06352, pi06353, pi06354, pi06355, pi06356, pi06357, pi06358, pi06359, pi06360, pi06361, pi06362, pi06363, pi06364, pi06365, pi06366, pi06367, pi06368, pi06369, pi06370, pi06371, pi06372, pi06373, pi06374, pi06375, pi06376, pi06377, pi06378, pi06379, pi06380, pi06381, pi06382, pi06383, pi06384, pi06385, pi06386, pi06387, pi06388, pi06389, pi06390, pi06391, pi06392, pi06393, pi06394, pi06395, pi06396, pi06397, pi06398, pi06399, pi06400, pi06401, pi06402, pi06403, pi06404, pi06405, pi06406, pi06407, pi06408, pi06409, pi06410, pi06411, pi06412, pi06413, pi06414, pi06415, pi06416, pi06417, pi06418, pi06419, pi06420, pi06421, pi06422, pi06423, pi06424, pi06425, pi06426, pi06427, pi06428, pi06429, pi06430, pi06431, pi06432, pi06433, pi06434, pi06435, pi06436, pi06437, pi06438, pi06439, pi06440, pi06441, pi06442, pi06443, pi06444, pi06445, pi06446, pi06447, pi06448, pi06449, pi06450, pi06451, pi06452, pi06453, pi06454, pi06455, pi06456, pi06457, pi06458, pi06459, pi06460, pi06461, pi06462, pi06463, pi06464, pi06465, pi06466, pi06467, pi06468, pi06469, pi06470, pi06471, pi06472, pi06473, pi06474, pi06475, pi06476, pi06477, pi06478, pi06479, pi06480, pi06481, pi06482, pi06483, pi06484, pi06485, pi06486, pi06487, pi06488, pi06489, pi06490, pi06491, pi06492, pi06493, pi06494, pi06495, pi06496, pi06497, pi06498, pi06499, pi06500, pi06501, pi06502, pi06503, pi06504, pi06505, pi06506, pi06507, pi06508, pi06509, pi06510, pi06511, pi06512, pi06513, pi06514, pi06515, pi06516, pi06517, pi06518, pi06519, pi06520, pi06521, pi06522, pi06523, pi06524, pi06525, pi06526, pi06527, pi06528, pi06529, pi06530, pi06531, pi06532, pi06533, pi06534, pi06535, pi06536, pi06537, pi06538, pi06539, pi06540, pi06541, pi06542, pi06543, pi06544, pi06545, pi06546, pi06547, pi06548, pi06549, pi06550, pi06551, pi06552, pi06553, pi06554, pi06555, pi06556, pi06557, pi06558, pi06559, pi06560, pi06561, pi06562, pi06563, pi06564, pi06565, pi06566, pi06567, pi06568, pi06569, pi06570, pi06571, pi06572, pi06573, pi06574, pi06575, pi06576, pi06577, pi06578, pi06579, pi06580, pi06581, pi06582, pi06583, pi06584, pi06585, pi06586, pi06587, pi06588, pi06589, pi06590, pi06591, pi06592, pi06593, pi06594, pi06595, pi06596, pi06597, pi06598, pi06599, pi06600, pi06601, pi06602, pi06603, pi06604, pi06605, pi06606, pi06607, pi06608, pi06609, pi06610, pi06611, pi06612, pi06613, pi06614, pi06615, pi06616, pi06617, pi06618, pi06619, pi06620, pi06621, pi06622, pi06623, pi06624, pi06625, pi06626, pi06627, pi06628, pi06629, pi06630, pi06631, pi06632, pi06633, pi06634, pi06635, pi06636, pi06637, pi06638, pi06639, pi06640, pi06641, pi06642, pi06643, pi06644, pi06645, pi06646, pi06647, pi06648, pi06649, pi06650, pi06651, pi06652, pi06653, pi06654, pi06655, pi06656, pi06657, pi06658, pi06659, pi06660, pi06661, pi06662, pi06663, pi06664, pi06665, pi06666, pi06667, pi06668, pi06669, pi06670, pi06671, pi06672, pi06673, pi06674, pi06675, pi06676, pi06677, pi06678, pi06679, pi06680, pi06681, pi06682, pi06683, pi06684, pi06685, pi06686, pi06687, pi06688, pi06689, pi06690, pi06691, pi06692, pi06693, pi06694, pi06695, pi06696, pi06697, pi06698, pi06699, pi06700, pi06701, pi06702, pi06703, pi06704, pi06705, pi06706, pi06707, pi06708, pi06709, pi06710, pi06711, pi06712, pi06713, pi06714, pi06715, pi06716, pi06717, pi06718, pi06719, pi06720, pi06721, pi06722, pi06723, pi06724, pi06725, pi06726, pi06727, pi06728, pi06729, pi06730, pi06731, pi06732, pi06733, pi06734, pi06735, pi06736, pi06737, pi06738, pi06739, pi06740, pi06741, pi06742, pi06743, pi06744, pi06745, pi06746, pi06747, pi06748, pi06749, pi06750, pi06751, pi06752, pi06753, pi06754, pi06755, pi06756, pi06757, pi06758, pi06759, pi06760, pi06761, pi06762, pi06763, pi06764, pi06765, pi06766, pi06767, pi06768, pi06769, pi06770, pi06771, pi06772, pi06773, pi06774, pi06775, pi06776, pi06777, pi06778, pi06779, pi06780, pi06781, pi06782, pi06783, pi06784, pi06785, pi06786, pi06787, pi06788, pi06789, pi06790, pi06791, pi06792, pi06793, pi06794, pi06795, pi06796, pi06797, pi06798, pi06799, pi06800, pi06801, pi06802, pi06803, pi06804, pi06805, pi06806, pi06807, pi06808, pi06809, pi06810, pi06811, pi06812, pi06813, pi06814, pi06815, pi06816, pi06817, pi06818, pi06819, pi06820, pi06821, pi06822, pi06823, pi06824, pi06825, pi06826, pi06827, pi06828, pi06829, pi06830, pi06831, pi06832, pi06833, pi06834, pi06835, pi06836, pi06837, pi06838, pi06839, pi06840, pi06841, pi06842, pi06843, pi06844, pi06845, pi06846, pi06847, pi06848, pi06849, pi06850, pi06851, pi06852, pi06853, pi06854, pi06855, pi06856, pi06857, pi06858, pi06859, pi06860, pi06861, pi06862, pi06863, pi06864, pi06865, pi06866, pi06867, pi06868, pi06869, pi06870, pi06871, pi06872, pi06873, pi06874, pi06875, pi06876, pi06877, pi06878, pi06879, pi06880, pi06881, pi06882, pi06883, pi06884, pi06885, pi06886, pi06887, pi06888, pi06889, pi06890, pi06891, pi06892, pi06893, pi06894, pi06895, pi06896, pi06897, pi06898, pi06899, pi06900, pi06901, pi06902, pi06903, pi06904, pi06905, pi06906, pi06907, pi06908, pi06909, pi06910, pi06911, pi06912, pi06913, pi06914, pi06915, pi06916, pi06917, pi06918, pi06919, pi06920, pi06921, pi06922, pi06923, pi06924, pi06925, pi06926, pi06927, pi06928, pi06929, pi06930, pi06931, pi06932, pi06933, pi06934, pi06935, pi06936, pi06937, pi06938, pi06939, pi06940, pi06941, pi06942, pi06943, pi06944, pi06945, pi06946, pi06947, pi06948, pi06949, pi06950, pi06951, pi06952, pi06953, pi06954, pi06955, pi06956, pi06957, pi06958, pi06959, pi06960, pi06961, pi06962, pi06963, pi06964, pi06965, pi06966, pi06967, pi06968, pi06969, pi06970, pi06971, pi06972, pi06973, pi06974, pi06975, pi06976, pi06977, pi06978, pi06979, pi06980, pi06981, pi06982, pi06983, pi06984, pi06985, pi06986, pi06987, pi06988, pi06989, pi06990, pi06991, pi06992, pi06993, pi06994, pi06995, pi06996, pi06997, pi06998, pi06999, pi07000, pi07001, pi07002, pi07003, pi07004, pi07005, pi07006, pi07007, pi07008, pi07009, pi07010, pi07011, pi07012, pi07013, pi07014, pi07015, pi07016, pi07017, pi07018, pi07019, pi07020, pi07021, pi07022, pi07023, pi07024, pi07025, pi07026, pi07027, pi07028, pi07029, pi07030, pi07031, pi07032, pi07033, pi07034, pi07035, pi07036, pi07037, pi07038, pi07039, pi07040, pi07041, pi07042, pi07043, pi07044, pi07045, pi07046, pi07047, pi07048, pi07049, pi07050, pi07051, pi07052, pi07053, pi07054, pi07055, pi07056, pi07057, pi07058, pi07059, pi07060, pi07061, pi07062, pi07063, pi07064, pi07065, pi07066, pi07067, pi07068, pi07069, pi07070, pi07071, pi07072, pi07073, pi07074, pi07075, pi07076, pi07077, pi07078, pi07079, pi07080, pi07081, pi07082, pi07083, pi07084, pi07085, pi07086, pi07087, pi07088, pi07089, pi07090, pi07091, pi07092, pi07093, pi07094, pi07095, pi07096, pi07097, pi07098, pi07099, pi07100, pi07101, pi07102, pi07103, pi07104, pi07105, pi07106, pi07107, pi07108, pi07109, pi07110, pi07111, pi07112, pi07113, pi07114, pi07115, pi07116, pi07117, pi07118, pi07119, pi07120, pi07121, pi07122, pi07123, pi07124, pi07125, pi07126, pi07127, pi07128, pi07129, pi07130, pi07131, pi07132, pi07133, pi07134, pi07135, pi07136, pi07137, pi07138, pi07139, pi07140, pi07141, pi07142, pi07143, pi07144, pi07145, pi07146, pi07147, pi07148, pi07149, pi07150, pi07151, pi07152, pi07153, pi07154, pi07155, pi07156, pi07157, pi07158, pi07159, pi07160, pi07161, pi07162, pi07163, pi07164, pi07165, pi07166, pi07167, pi07168, pi07169, pi07170, pi07171, pi07172, pi07173, pi07174, pi07175, pi07176, pi07177, pi07178, pi07179, pi07180, pi07181, pi07182, pi07183, pi07184, pi07185, pi07186, pi07187, pi07188, pi07189, pi07190, pi07191, pi07192, pi07193, pi07194, pi07195, pi07196, pi07197, pi07198, pi07199, pi07200, pi07201, pi07202, pi07203, pi07204, pi07205, pi07206, pi07207, pi07208, pi07209, pi07210, pi07211, pi07212, pi07213, pi07214, pi07215, pi07216, pi07217, pi07218, pi07219, pi07220, pi07221, pi07222, pi07223, pi07224, pi07225, pi07226, pi07227, pi07228, pi07229, pi07230, pi07231, pi07232, pi07233, pi07234, pi07235, pi07236, pi07237, pi07238, pi07239, pi07240, pi07241, pi07242, pi07243, pi07244, pi07245, pi07246, pi07247, pi07248, pi07249, pi07250, pi07251, pi07252, pi07253, pi07254, pi07255, pi07256, pi07257, pi07258, pi07259, pi07260, pi07261, pi07262, pi07263, pi07264, pi07265, pi07266, pi07267, pi07268, pi07269, pi07270, pi07271, pi07272, pi07273, pi07274, pi07275, pi07276, pi07277, pi07278, pi07279, pi07280, pi07281, pi07282, pi07283, pi07284, pi07285, pi07286, pi07287, pi07288, pi07289, pi07290, pi07291, pi07292, pi07293, pi07294, pi07295, pi07296, pi07297, pi07298, pi07299, pi07300, pi07301, pi07302, pi07303, pi07304, pi07305, pi07306, pi07307, pi07308, pi07309, pi07310, pi07311, pi07312, pi07313, pi07314, pi07315, pi07316, pi07317, pi07318, pi07319, pi07320, pi07321, pi07322, pi07323, pi07324, pi07325, pi07326, pi07327, pi07328, pi07329, pi07330, pi07331, pi07332, pi07333, pi07334, pi07335, pi07336, pi07337, pi07338, pi07339, pi07340, pi07341, pi07342, pi07343, pi07344, pi07345, pi07346, pi07347, pi07348, pi07349, pi07350, pi07351, pi07352, pi07353, pi07354, pi07355, pi07356, pi07357, pi07358, pi07359, pi07360, pi07361, pi07362, pi07363, pi07364, pi07365, pi07366, pi07367, pi07368, pi07369, pi07370, pi07371, pi07372, pi07373, pi07374, pi07375, pi07376, pi07377, pi07378, pi07379, pi07380, pi07381, pi07382, pi07383, pi07384, pi07385, pi07386, pi07387, pi07388, pi07389, pi07390, pi07391, pi07392, pi07393, pi07394, pi07395, pi07396, pi07397, pi07398, pi07399, pi07400, pi07401, pi07402, pi07403, pi07404, pi07405, pi07406, pi07407, pi07408, pi07409, pi07410, pi07411, pi07412, pi07413, pi07414, pi07415, pi07416, pi07417, pi07418, pi07419, pi07420, pi07421, pi07422, pi07423, pi07424, pi07425, pi07426, pi07427, pi07428, pi07429, pi07430, pi07431, pi07432, pi07433, pi07434, pi07435, pi07436, pi07437, pi07438, pi07439, pi07440, pi07441, pi07442, pi07443, pi07444, pi07445, pi07446, pi07447, pi07448, pi07449, pi07450, pi07451, pi07452, pi07453, pi07454, pi07455, pi07456, pi07457, pi07458, pi07459, pi07460, pi07461, pi07462, pi07463, pi07464, pi07465, pi07466, pi07467, pi07468, pi07469, pi07470, pi07471, pi07472, pi07473, pi07474, pi07475, pi07476, pi07477, pi07478, pi07479, pi07480, pi07481, pi07482, pi07483, pi07484, pi07485, pi07486, pi07487, pi07488, pi07489, pi07490, pi07491, pi07492, pi07493, pi07494, pi07495, pi07496, pi07497, pi07498, pi07499, pi07500, pi07501, pi07502, pi07503, pi07504, pi07505, pi07506, pi07507, pi07508, pi07509, pi07510, pi07511, pi07512, pi07513, pi07514, pi07515, pi07516, pi07517, pi07518, pi07519, pi07520, pi07521, pi07522, pi07523, pi07524, pi07525, pi07526, pi07527, pi07528, pi07529, pi07530, pi07531, pi07532, pi07533, pi07534, pi07535, pi07536, pi07537, pi07538, pi07539, pi07540, pi07541, pi07542, pi07543, pi07544, pi07545, pi07546, pi07547, pi07548, pi07549, pi07550, pi07551, pi07552, pi07553, pi07554, pi07555, pi07556, pi07557, pi07558, pi07559, pi07560, pi07561, pi07562, pi07563, pi07564, pi07565, pi07566, pi07567, pi07568, pi07569, pi07570, pi07571, pi07572, pi07573, pi07574, pi07575, pi07576, pi07577, pi07578, pi07579, pi07580, pi07581, pi07582, pi07583, pi07584, pi07585, pi07586, pi07587, pi07588, pi07589, pi07590, pi07591, pi07592, pi07593, pi07594, pi07595, pi07596, pi07597, pi07598, pi07599, pi07600, pi07601, pi07602, pi07603, pi07604, pi07605, pi07606, pi07607, pi07608, pi07609, pi07610, pi07611, pi07612, pi07613, pi07614, pi07615, pi07616, pi07617, pi07618, pi07619, pi07620, pi07621, pi07622, pi07623, pi07624, pi07625, pi07626, pi07627, pi07628, pi07629, pi07630, pi07631, pi07632, pi07633, pi07634, pi07635, pi07636, pi07637, pi07638, pi07639, pi07640, pi07641, pi07642, pi07643, pi07644, pi07645, pi07646, pi07647, pi07648, pi07649, pi07650, pi07651, pi07652, pi07653, pi07654, pi07655, pi07656, pi07657, pi07658, pi07659, pi07660, pi07661, pi07662, pi07663, pi07664, pi07665, pi07666, pi07667, pi07668, pi07669, pi07670, pi07671, pi07672, pi07673, pi07674, pi07675, pi07676, pi07677, pi07678, pi07679, pi07680, pi07681, pi07682, pi07683, pi07684, pi07685, pi07686, pi07687, pi07688, pi07689, pi07690, pi07691, pi07692, pi07693, pi07694, pi07695, pi07696, pi07697, pi07698, pi07699, pi07700, pi07701, pi07702, pi07703, pi07704, pi07705, pi07706, pi07707, pi07708, pi07709, pi07710, pi07711, pi07712, pi07713, pi07714, pi07715, pi07716, pi07717, pi07718, pi07719, pi07720, pi07721, pi07722, pi07723, pi07724, pi07725, pi07726, pi07727, pi07728, pi07729, pi07730, pi07731, pi07732, pi07733, pi07734, pi07735, pi07736, pi07737, pi07738, pi07739, pi07740, pi07741, pi07742, pi07743, pi07744, pi07745, pi07746, pi07747, pi07748, pi07749, pi07750, pi07751, pi07752, pi07753, pi07754, pi07755, pi07756, pi07757, pi07758, pi07759, pi07760, pi07761, pi07762, pi07763, pi07764, pi07765, pi07766, pi07767, pi07768, pi07769, pi07770, pi07771, pi07772, pi07773, pi07774, pi07775, pi07776, pi07777, pi07778, pi07779, pi07780, pi07781, pi07782, pi07783, pi07784, pi07785, pi07786, pi07787, pi07788, pi07789, pi07790, pi07791, pi07792, pi07793, pi07794, pi07795, pi07796, pi07797, pi07798, pi07799, pi07800, pi07801, pi07802, pi07803, pi07804, pi07805, pi07806, pi07807, pi07808, pi07809, pi07810, pi07811, pi07812, pi07813, pi07814, pi07815, pi07816, pi07817, pi07818, pi07819, pi07820, pi07821, pi07822, pi07823, pi07824, pi07825, pi07826, pi07827, pi07828, pi07829, pi07830, pi07831, pi07832, pi07833, pi07834, pi07835, pi07836, pi07837, pi07838, pi07839, pi07840, pi07841, pi07842, pi07843, pi07844, pi07845, pi07846, pi07847, pi07848, pi07849, pi07850, pi07851, pi07852, pi07853, pi07854, pi07855, pi07856, pi07857, pi07858, pi07859, pi07860, pi07861, pi07862, pi07863, pi07864, pi07865, pi07866, pi07867, pi07868, pi07869, pi07870, pi07871, pi07872, pi07873, pi07874, pi07875, pi07876, pi07877, pi07878, pi07879, pi07880, pi07881, pi07882, pi07883, pi07884, pi07885, pi07886, pi07887, pi07888, pi07889, pi07890, pi07891, pi07892, pi07893, pi07894, pi07895, pi07896, pi07897, pi07898, pi07899, pi07900, pi07901, pi07902, pi07903, pi07904, pi07905, pi07906, pi07907, pi07908, pi07909, pi07910, pi07911, pi07912, pi07913, pi07914, pi07915, pi07916, pi07917, pi07918, pi07919, pi07920, pi07921, pi07922, pi07923, pi07924, pi07925, pi07926, pi07927, pi07928, pi07929, pi07930, pi07931, pi07932, pi07933, pi07934, pi07935, pi07936, pi07937, pi07938, pi07939, pi07940, pi07941, pi07942, pi07943, pi07944, pi07945, pi07946, pi07947, pi07948, pi07949, pi07950, pi07951, pi07952, pi07953, pi07954, pi07955, pi07956, pi07957, pi07958, pi07959, pi07960, pi07961, pi07962, pi07963, pi07964, pi07965, pi07966, pi07967, pi07968, pi07969, pi07970, pi07971, pi07972, pi07973, pi07974, pi07975, pi07976, pi07977, pi07978, pi07979, pi07980, pi07981, pi07982, pi07983, pi07984, pi07985, pi07986, pi07987, pi07988, pi07989, pi07990, pi07991, pi07992, pi07993, pi07994, pi07995, pi07996, pi07997, pi07998, pi07999, pi08000, pi08001, pi08002, pi08003, pi08004, pi08005, pi08006, pi08007, pi08008, pi08009, pi08010, pi08011, pi08012, pi08013, pi08014, pi08015, pi08016, pi08017, pi08018, pi08019, pi08020, pi08021, pi08022, pi08023, pi08024, pi08025, pi08026, pi08027, pi08028, pi08029, pi08030, pi08031, pi08032, pi08033, pi08034, pi08035, pi08036, pi08037, pi08038, pi08039, pi08040, pi08041, pi08042, pi08043, pi08044, pi08045, pi08046, pi08047, pi08048, pi08049, pi08050, pi08051, pi08052, pi08053, pi08054, pi08055, pi08056, pi08057, pi08058, pi08059, pi08060, pi08061, pi08062, pi08063, pi08064, pi08065, pi08066, pi08067, pi08068, pi08069, pi08070, pi08071, pi08072, pi08073, pi08074, pi08075, pi08076, pi08077, pi08078, pi08079, pi08080, pi08081, pi08082, pi08083, pi08084, pi08085, pi08086, pi08087, pi08088, pi08089, pi08090, pi08091, pi08092, pi08093, pi08094, pi08095, pi08096, pi08097, pi08098, pi08099, pi08100, pi08101, pi08102, pi08103, pi08104, pi08105, pi08106, pi08107, pi08108, pi08109, pi08110, pi08111, pi08112, pi08113, pi08114, pi08115, pi08116, pi08117, pi08118, pi08119, pi08120, pi08121, pi08122, pi08123, pi08124, pi08125, pi08126, pi08127, pi08128, pi08129, pi08130, pi08131, pi08132, pi08133, pi08134, pi08135, pi08136, pi08137, pi08138, pi08139, pi08140, pi08141, pi08142, pi08143, pi08144, pi08145, pi08146, pi08147, pi08148, pi08149, pi08150, pi08151, pi08152, pi08153, pi08154, pi08155, pi08156, pi08157, pi08158, pi08159, pi08160, pi08161, pi08162, pi08163, pi08164, pi08165, pi08166, pi08167, pi08168, pi08169, pi08170, pi08171, pi08172, pi08173, pi08174, pi08175, pi08176, pi08177, pi08178, pi08179, pi08180, pi08181, pi08182, pi08183, pi08184, pi08185, pi08186, pi08187, pi08188, pi08189, pi08190, pi08191, pi08192, pi08193, pi08194, pi08195, pi08196, pi08197, pi08198, pi08199, pi08200, pi08201, pi08202, pi08203, pi08204, pi08205, pi08206, pi08207, pi08208, pi08209, pi08210, pi08211, pi08212, pi08213, pi08214, pi08215, pi08216, pi08217, pi08218, pi08219, pi08220, pi08221, pi08222, pi08223, pi08224, pi08225, pi08226, pi08227, pi08228, pi08229, pi08230, pi08231, pi08232, pi08233, pi08234, pi08235, pi08236, pi08237, pi08238, pi08239, pi08240, pi08241, pi08242, pi08243, pi08244, pi08245, pi08246, pi08247, pi08248, pi08249, pi08250, pi08251, pi08252, pi08253, pi08254, pi08255, pi08256, pi08257, pi08258, pi08259, pi08260, pi08261, pi08262, pi08263, pi08264, pi08265, pi08266, pi08267, pi08268, pi08269, pi08270, pi08271, pi08272, pi08273, pi08274, pi08275, pi08276, pi08277, pi08278, pi08279, pi08280, pi08281, pi08282, pi08283, pi08284, pi08285, pi08286, pi08287, pi08288, pi08289, pi08290, pi08291, pi08292, pi08293, pi08294, pi08295, pi08296, pi08297, pi08298, pi08299, pi08300, pi08301, pi08302, pi08303, pi08304, pi08305, pi08306, pi08307, pi08308, pi08309, pi08310, pi08311, pi08312, pi08313, pi08314, pi08315, pi08316, pi08317, pi08318, pi08319, pi08320, pi08321, pi08322, pi08323, pi08324, pi08325, pi08326, pi08327, pi08328, pi08329, pi08330, pi08331, pi08332, pi08333, pi08334, pi08335, pi08336, pi08337, pi08338, pi08339, pi08340, pi08341, pi08342, pi08343, pi08344, pi08345, pi08346, pi08347, pi08348, pi08349, pi08350, pi08351, pi08352, pi08353, pi08354, pi08355, pi08356, pi08357, pi08358, pi08359, pi08360, pi08361, pi08362, pi08363, pi08364, pi08365, pi08366, pi08367, pi08368, pi08369, pi08370, pi08371, pi08372, pi08373, pi08374, pi08375, pi08376, pi08377, pi08378, pi08379, pi08380, pi08381, pi08382, pi08383, pi08384, pi08385, pi08386, pi08387, pi08388, pi08389, pi08390, pi08391, pi08392, pi08393, pi08394, pi08395, pi08396, pi08397, pi08398, pi08399, pi08400, pi08401, pi08402, pi08403, pi08404, pi08405, pi08406, pi08407, pi08408, pi08409, pi08410, pi08411, pi08412, pi08413, pi08414, pi08415, pi08416, pi08417, pi08418, pi08419, pi08420, pi08421, pi08422, pi08423, pi08424, pi08425, pi08426, pi08427, pi08428, pi08429, pi08430, pi08431, pi08432, pi08433, pi08434, pi08435, pi08436, pi08437, pi08438, pi08439, pi08440, pi08441, pi08442, pi08443, pi08444, pi08445, pi08446, pi08447, pi08448, pi08449, pi08450, pi08451, pi08452, pi08453, pi08454, pi08455, pi08456, pi08457, pi08458, pi08459, pi08460, pi08461, pi08462, pi08463, pi08464, pi08465, pi08466, pi08467, pi08468, pi08469, pi08470, pi08471, pi08472, pi08473, pi08474, pi08475, pi08476, pi08477, pi08478, pi08479, pi08480, pi08481, pi08482, pi08483, pi08484, pi08485, pi08486, pi08487, pi08488, pi08489, pi08490, pi08491, pi08492, pi08493, pi08494, pi08495, pi08496, pi08497, pi08498, pi08499, pi08500, pi08501, pi08502, pi08503, pi08504, pi08505, pi08506, pi08507, pi08508, pi08509, pi08510, pi08511, pi08512, pi08513, pi08514, pi08515, pi08516, pi08517, pi08518, pi08519, pi08520, pi08521, pi08522, pi08523, pi08524, pi08525, pi08526, pi08527, pi08528, pi08529, pi08530, pi08531, pi08532, pi08533, pi08534, pi08535, pi08536, pi08537, pi08538, pi08539, pi08540, pi08541, pi08542, pi08543, pi08544, pi08545, pi08546, pi08547, pi08548, pi08549, pi08550, pi08551, pi08552, pi08553, pi08554, pi08555, pi08556, pi08557, pi08558, pi08559, pi08560, pi08561, pi08562, pi08563, pi08564, pi08565, pi08566, pi08567, pi08568, pi08569, pi08570, pi08571, pi08572, pi08573, pi08574, pi08575, pi08576, pi08577, pi08578, pi08579, pi08580, pi08581, pi08582, pi08583, pi08584, pi08585, pi08586, pi08587, pi08588, pi08589, pi08590, pi08591, pi08592, pi08593, pi08594, pi08595, pi08596, pi08597, pi08598, pi08599, pi08600, pi08601, pi08602, pi08603, pi08604, pi08605, pi08606, pi08607, pi08608, pi08609, pi08610, pi08611, pi08612, pi08613, pi08614, pi08615, pi08616, pi08617, pi08618, pi08619, pi08620, pi08621, pi08622, pi08623, pi08624, pi08625, pi08626, pi08627, pi08628, pi08629, pi08630, pi08631, pi08632, pi08633, pi08634, pi08635, pi08636, pi08637, pi08638, pi08639, pi08640, pi08641, pi08642, pi08643, pi08644, pi08645, pi08646, pi08647, pi08648, pi08649, pi08650, pi08651, pi08652, pi08653, pi08654, pi08655, pi08656, pi08657, pi08658, pi08659, pi08660, pi08661, pi08662, pi08663, pi08664, pi08665, pi08666, pi08667, pi08668, pi08669, pi08670, pi08671, pi08672, pi08673, pi08674, pi08675, pi08676, pi08677, pi08678, pi08679, pi08680, pi08681, pi08682, pi08683, pi08684, pi08685, pi08686, pi08687, pi08688, pi08689, pi08690, pi08691, pi08692, pi08693, pi08694, pi08695, pi08696, pi08697, pi08698, pi08699, pi08700, pi08701, pi08702, pi08703, pi08704, pi08705, pi08706, pi08707, pi08708, pi08709, pi08710, pi08711, pi08712, pi08713, pi08714, pi08715, pi08716, pi08717, pi08718, pi08719, pi08720, pi08721, pi08722, pi08723, pi08724, pi08725, pi08726, pi08727, pi08728, pi08729, pi08730, pi08731, pi08732, pi08733, pi08734, pi08735, pi08736, pi08737, pi08738, pi08739, pi08740, pi08741, pi08742, pi08743, pi08744, pi08745, pi08746, pi08747, pi08748, pi08749, pi08750, pi08751, pi08752, pi08753, pi08754, pi08755, pi08756, pi08757, pi08758, pi08759, pi08760, pi08761, pi08762, pi08763, pi08764, pi08765, pi08766, pi08767, pi08768, pi08769, pi08770, pi08771, pi08772, pi08773, pi08774, pi08775, pi08776, pi08777, pi08778, pi08779, pi08780, pi08781, pi08782, pi08783, pi08784, pi08785, pi08786, pi08787, pi08788, pi08789, pi08790, pi08791, pi08792, pi08793, pi08794, pi08795, pi08796, pi08797, pi08798, pi08799, pi08800, pi08801, pi08802, pi08803, pi08804, pi08805, pi08806, pi08807, pi08808, pi08809, pi08810, pi08811, pi08812, pi08813, pi08814, pi08815, pi08816, pi08817, pi08818, pi08819, pi08820, pi08821, pi08822, pi08823, pi08824, pi08825, pi08826, pi08827, pi08828, pi08829, pi08830, pi08831, pi08832, pi08833, pi08834, pi08835, pi08836, pi08837, pi08838, pi08839, pi08840, pi08841, pi08842, pi08843, pi08844, pi08845, pi08846, pi08847, pi08848, pi08849, pi08850, pi08851, pi08852, pi08853, pi08854, pi08855, pi08856, pi08857, pi08858, pi08859, pi08860, pi08861, pi08862, pi08863, pi08864, pi08865, pi08866, pi08867, pi08868, pi08869, pi08870, pi08871, pi08872, pi08873, pi08874, pi08875, pi08876, pi08877, pi08878, pi08879, pi08880, pi08881, pi08882, pi08883, pi08884, pi08885, pi08886, pi08887, pi08888, pi08889, pi08890, pi08891, pi08892, pi08893, pi08894, pi08895, pi08896, pi08897, pi08898, pi08899, pi08900, pi08901, pi08902, pi08903, pi08904, pi08905, pi08906, pi08907, pi08908, pi08909, pi08910, pi08911, pi08912, pi08913, pi08914, pi08915, pi08916, pi08917, pi08918, pi08919, pi08920, pi08921, pi08922, pi08923, pi08924, pi08925, pi08926, pi08927, pi08928, pi08929, pi08930, pi08931, pi08932, pi08933, pi08934, pi08935, pi08936, pi08937, pi08938, pi08939, pi08940, pi08941, pi08942, pi08943, pi08944, pi08945, pi08946, pi08947, pi08948, pi08949, pi08950, pi08951, pi08952, pi08953, pi08954, pi08955, pi08956, pi08957, pi08958, pi08959, pi08960, pi08961, pi08962, pi08963, pi08964, pi08965, pi08966, pi08967, pi08968, pi08969, pi08970, pi08971, pi08972, pi08973, pi08974, pi08975, pi08976, pi08977, pi08978, pi08979, pi08980, pi08981, pi08982, pi08983, pi08984, pi08985, pi08986, pi08987, pi08988, pi08989, pi08990, pi08991, pi08992, pi08993, pi08994, pi08995, pi08996, pi08997, pi08998, pi08999, pi09000, pi09001, pi09002, pi09003, pi09004, pi09005, pi09006, pi09007, pi09008, pi09009, pi09010, pi09011, pi09012, pi09013, pi09014, pi09015, pi09016, pi09017, pi09018, pi09019, pi09020, pi09021, pi09022, pi09023, pi09024, pi09025, pi09026, pi09027, pi09028, pi09029, pi09030, pi09031, pi09032, pi09033, pi09034, pi09035, pi09036, pi09037, pi09038, pi09039, pi09040, pi09041, pi09042, pi09043, pi09044, pi09045, pi09046, pi09047, pi09048, pi09049, pi09050, pi09051, pi09052, pi09053, pi09054, pi09055, pi09056, pi09057, pi09058, pi09059, pi09060, pi09061, pi09062, pi09063, pi09064, pi09065, pi09066, pi09067, pi09068, pi09069, pi09070, pi09071, pi09072, pi09073, pi09074, pi09075, pi09076, pi09077, pi09078, pi09079, pi09080, pi09081, pi09082, pi09083, pi09084, pi09085, pi09086, pi09087, pi09088, pi09089, pi09090, pi09091, pi09092, pi09093, pi09094, pi09095, pi09096, pi09097, pi09098, pi09099, pi09100, pi09101, pi09102, pi09103, pi09104, pi09105, pi09106, pi09107, pi09108, pi09109, pi09110, pi09111, pi09112, pi09113, pi09114, pi09115, pi09116, pi09117, pi09118, pi09119, pi09120, pi09121, pi09122, pi09123, pi09124, pi09125, pi09126, pi09127, pi09128, pi09129, pi09130, pi09131, pi09132, pi09133, pi09134, pi09135, pi09136, pi09137, pi09138, pi09139, pi09140, pi09141, pi09142, pi09143, pi09144, pi09145, pi09146, pi09147, pi09148, pi09149, pi09150, pi09151, pi09152, pi09153, pi09154, pi09155, pi09156, pi09157, pi09158, pi09159, pi09160, pi09161, pi09162, pi09163, pi09164, pi09165, pi09166, pi09167, pi09168, pi09169, pi09170, pi09171, pi09172, pi09173, pi09174, pi09175, pi09176, pi09177, pi09178, pi09179, pi09180, pi09181, pi09182, pi09183, pi09184, pi09185, pi09186, pi09187, pi09188, pi09189, pi09190, pi09191, pi09192, pi09193, pi09194, pi09195, pi09196, pi09197, pi09198, pi09199, pi09200, pi09201, pi09202, pi09203, pi09204, pi09205, pi09206, pi09207, pi09208, pi09209, pi09210, pi09211, pi09212, pi09213, pi09214, pi09215, pi09216, pi09217, pi09218, pi09219, pi09220, pi09221, pi09222, pi09223, pi09224, pi09225, pi09226, pi09227, pi09228, pi09229, pi09230, pi09231, pi09232, pi09233, pi09234, pi09235, pi09236, pi09237, pi09238, pi09239, pi09240, pi09241, pi09242, pi09243, pi09244, pi09245, pi09246, pi09247, pi09248, pi09249, pi09250, pi09251, pi09252, pi09253, pi09254, pi09255, pi09256, pi09257, pi09258, pi09259, pi09260, pi09261, pi09262, pi09263, pi09264, pi09265, pi09266, pi09267, pi09268, pi09269, pi09270, pi09271, pi09272, pi09273, pi09274, pi09275, pi09276, pi09277, pi09278, pi09279, pi09280, pi09281, pi09282, pi09283, pi09284, pi09285, pi09286, pi09287, pi09288, pi09289, pi09290, pi09291, pi09292, pi09293, pi09294, pi09295, pi09296, pi09297, pi09298, pi09299, pi09300, pi09301, pi09302, pi09303, pi09304, pi09305, pi09306, pi09307, pi09308, pi09309, pi09310, pi09311, pi09312, pi09313, pi09314, pi09315, pi09316, pi09317, pi09318, pi09319, pi09320, pi09321, pi09322, pi09323, pi09324, pi09325, pi09326, pi09327, pi09328, pi09329, pi09330, pi09331, pi09332, pi09333, pi09334, pi09335, pi09336, pi09337, pi09338, pi09339, pi09340, pi09341, pi09342, pi09343, pi09344, pi09345, pi09346, pi09347, pi09348, pi09349, pi09350, pi09351, pi09352, pi09353, pi09354, pi09355, pi09356, pi09357, pi09358, pi09359, pi09360, pi09361, pi09362, pi09363, pi09364, pi09365, pi09366, pi09367, pi09368, pi09369, pi09370, pi09371, pi09372, pi09373, pi09374, pi09375, pi09376, pi09377, pi09378, pi09379, pi09380, pi09381, pi09382, pi09383, pi09384, pi09385, pi09386, pi09387, pi09388, pi09389, pi09390, pi09391, pi09392, pi09393, pi09394, pi09395, pi09396, pi09397, pi09398, pi09399, pi09400, pi09401, pi09402, pi09403, pi09404, pi09405, pi09406, pi09407, pi09408, pi09409, pi09410, pi09411, pi09412, pi09413, pi09414, pi09415, pi09416, pi09417, pi09418, pi09419, pi09420, pi09421, pi09422, pi09423, pi09424, pi09425, pi09426, pi09427, pi09428, pi09429, pi09430, pi09431, pi09432, pi09433, pi09434, pi09435, pi09436, pi09437, pi09438, pi09439, pi09440, pi09441, pi09442, pi09443, pi09444, pi09445, pi09446, pi09447, pi09448, pi09449, pi09450, pi09451, pi09452, pi09453, pi09454, pi09455, pi09456, pi09457, pi09458, pi09459, pi09460, pi09461, pi09462, pi09463, pi09464, pi09465, pi09466, pi09467, pi09468, pi09469, pi09470, pi09471, pi09472, pi09473, pi09474, pi09475, pi09476, pi09477, pi09478, pi09479, pi09480, pi09481, pi09482, pi09483, pi09484, pi09485, pi09486, pi09487, pi09488, pi09489, pi09490, pi09491, pi09492, pi09493, pi09494, pi09495, pi09496, pi09497, pi09498, pi09499, pi09500, pi09501, pi09502, pi09503, pi09504, pi09505, pi09506, pi09507, pi09508, pi09509, pi09510, pi09511, pi09512, pi09513, pi09514, pi09515, pi09516, pi09517, pi09518, pi09519, pi09520, pi09521, pi09522, pi09523, pi09524, pi09525, pi09526, pi09527, pi09528, pi09529, pi09530, pi09531, pi09532, pi09533, pi09534, pi09535, pi09536, pi09537, pi09538, pi09539, pi09540, pi09541, pi09542, pi09543, pi09544, pi09545, pi09546, pi09547, pi09548, pi09549, pi09550, pi09551, pi09552, pi09553, pi09554, pi09555, pi09556, pi09557, pi09558, pi09559, pi09560, pi09561, pi09562, pi09563, pi09564, pi09565, pi09566, pi09567, pi09568, pi09569, pi09570, pi09571, pi09572, pi09573, pi09574, pi09575, pi09576, pi09577, pi09578, pi09579, pi09580, pi09581, pi09582, pi09583, pi09584, pi09585, pi09586, pi09587, pi09588, pi09589, pi09590, pi09591, pi09592, pi09593, pi09594, pi09595, pi09596, pi09597, pi09598, pi09599, pi09600, pi09601, pi09602, pi09603, pi09604, pi09605, pi09606, pi09607, pi09608, pi09609, pi09610, pi09611, pi09612, pi09613, pi09614, pi09615, pi09616, pi09617, pi09618, pi09619, pi09620, pi09621, pi09622, pi09623, pi09624, pi09625, pi09626, pi09627, pi09628, pi09629, pi09630, pi09631, pi09632, pi09633, pi09634, pi09635, pi09636, pi09637, pi09638, pi09639, pi09640, pi09641, pi09642, pi09643, pi09644, pi09645, pi09646, pi09647, pi09648, pi09649, pi09650, pi09651, pi09652, pi09653, pi09654, pi09655, pi09656, pi09657, pi09658, pi09659, pi09660, pi09661, pi09662, pi09663, pi09664, pi09665, pi09666, pi09667, pi09668, pi09669, pi09670, pi09671, pi09672, pi09673, pi09674, pi09675, pi09676, pi09677, pi09678, pi09679, pi09680, pi09681, pi09682, pi09683, pi09684, pi09685, pi09686, pi09687, pi09688, pi09689, pi09690, pi09691, pi09692, pi09693, pi09694, pi09695, pi09696, pi09697, pi09698, pi09699, pi09700, pi09701, pi09702, pi09703, pi09704, pi09705, pi09706, pi09707, pi09708, pi09709, pi09710, pi09711, pi09712, pi09713, pi09714, pi09715, pi09716, pi09717, pi09718, pi09719, pi09720, pi09721, pi09722, pi09723, pi09724, pi09725, pi09726, pi09727, pi09728, pi09729, pi09730, pi09731, pi09732, pi09733, pi09734, pi09735, pi09736, pi09737, pi09738, pi09739, pi09740, pi09741, pi09742, pi09743, pi09744, pi09745, pi09746, pi09747, pi09748, pi09749, pi09750, pi09751, pi09752, pi09753, pi09754, pi09755, pi09756, pi09757, pi09758, pi09759, pi09760, pi09761, pi09762, pi09763, pi09764, pi09765, pi09766, pi09767, pi09768, pi09769, pi09770, pi09771, pi09772, pi09773, pi09774, pi09775, pi09776, pi09777, pi09778, pi09779, pi09780, pi09781, pi09782, pi09783, pi09784, pi09785, pi09786, pi09787, pi09788, pi09789, pi09790, pi09791, pi09792, pi09793, pi09794, pi09795, pi09796, pi09797, pi09798, pi09799, pi09800, pi09801, pi09802, pi09803, pi09804, pi09805, pi09806, pi09807, pi09808, pi09809, pi09810, pi09811, pi09812, pi09813, pi09814, pi09815, pi09816, pi09817, pi09818, pi09819, pi09820, pi09821, pi09822, pi09823, pi09824, pi09825, pi09826, pi09827, pi09828, pi09829, pi09830, pi09831, pi09832, pi09833, pi09834, pi09835, pi09836, pi09837, pi09838, pi09839, pi09840, pi09841, pi09842, pi09843, pi09844, pi09845, pi09846, pi09847, pi09848, pi09849, pi09850, pi09851, pi09852, pi09853, pi09854, pi09855, pi09856, pi09857, pi09858, pi09859, pi09860, pi09861, pi09862, pi09863, pi09864, pi09865, pi09866, pi09867, pi09868, pi09869, pi09870, pi09871, pi09872, pi09873, pi09874, pi09875, pi09876, pi09877, pi09878, pi09879, pi09880, pi09881, pi09882, pi09883, pi09884, pi09885, pi09886, pi09887, pi09888, pi09889, pi09890, pi09891, pi09892, pi09893, pi09894, pi09895, pi09896, pi09897, pi09898, pi09899, pi09900, pi09901, pi09902, pi09903, pi09904, pi09905, pi09906, pi09907, pi09908, pi09909, pi09910, pi09911, pi09912, pi09913, pi09914, pi09915, pi09916, pi09917, pi09918, pi09919, pi09920, pi09921, pi09922, pi09923, pi09924, pi09925, pi09926, pi09927, pi09928, pi09929, pi09930, pi09931, pi09932, pi09933, pi09934, pi09935, pi09936, pi09937, pi09938, pi09939, pi09940, pi09941, pi09942, pi09943, pi09944, pi09945, pi09946, pi09947, pi09948, pi09949, pi09950, pi09951, pi09952, pi09953, pi09954, pi09955, pi09956, pi09957, pi09958, pi09959, pi09960, pi09961, pi09962, pi09963, pi09964, pi09965, pi09966, pi09967, pi09968, pi09969, pi09970, pi09971, pi09972, pi09973, pi09974, pi09975, pi09976, pi09977, pi09978, pi09979, pi09980, pi09981, pi09982, pi09983, pi09984, pi09985, pi09986, pi09987, pi09988, pi09989, pi09990, pi09991, pi09992, pi09993, pi09994, pi09995, pi09996, pi09997, pi09998, pi09999, pi10000, pi10001, pi10002, pi10003, pi10004, pi10005, pi10006, pi10007, pi10008, pi10009, pi10010, pi10011, pi10012, pi10013, pi10014, pi10015, pi10016, pi10017, pi10018, pi10019, pi10020, pi10021, pi10022, pi10023, pi10024, pi10025, pi10026, pi10027, pi10028, pi10029, pi10030, pi10031, pi10032, pi10033, pi10034, pi10035, pi10036, pi10037, pi10038, pi10039, pi10040, pi10041, pi10042, pi10043, pi10044, pi10045, pi10046, pi10047, pi10048, pi10049, pi10050, pi10051, pi10052, pi10053, pi10054, pi10055, pi10056, pi10057, pi10058, pi10059, pi10060, pi10061, pi10062, pi10063, pi10064, pi10065, pi10066, pi10067, pi10068, pi10069, pi10070, pi10071, pi10072, pi10073, pi10074, pi10075, pi10076, pi10077, pi10078, pi10079, pi10080, pi10081, pi10082, pi10083, pi10084, pi10085, pi10086, pi10087, pi10088, pi10089, pi10090, pi10091, pi10092, pi10093, pi10094, pi10095, pi10096, pi10097, pi10098, pi10099, pi10100, pi10101, pi10102, pi10103, pi10104, pi10105, pi10106, pi10107, pi10108, pi10109, pi10110, pi10111, pi10112, pi10113, pi10114, pi10115, pi10116, pi10117, pi10118, pi10119, pi10120, pi10121, pi10122, pi10123, pi10124, pi10125, pi10126, pi10127, pi10128, pi10129, pi10130, pi10131, pi10132, pi10133, pi10134, pi10135, pi10136, pi10137, pi10138, pi10139, pi10140, pi10141, pi10142, pi10143, pi10144, pi10145, pi10146, pi10147, pi10148, pi10149, pi10150, pi10151, pi10152, pi10153, pi10154, pi10155, pi10156, pi10157, pi10158, pi10159, pi10160, pi10161, pi10162, pi10163, pi10164, pi10165, pi10166, pi10167, pi10168, pi10169, pi10170, pi10171, pi10172, pi10173, pi10174, pi10175, pi10176, pi10177, pi10178, pi10179, pi10180, pi10181, pi10182, pi10183, pi10184, pi10185, pi10186, pi10187, pi10188, pi10189, pi10190, pi10191, pi10192, pi10193, pi10194, pi10195, pi10196, pi10197, pi10198, pi10199, pi10200, pi10201, pi10202, pi10203, pi10204, pi10205, pi10206, pi10207, pi10208, pi10209, pi10210, pi10211, pi10212, pi10213, pi10214, pi10215, pi10216, pi10217, pi10218, pi10219, pi10220, pi10221, pi10222, pi10223, pi10224, pi10225, pi10226, pi10227, pi10228, pi10229, pi10230, pi10231, pi10232, pi10233, pi10234, pi10235, pi10236, pi10237, pi10238, pi10239, pi10240, pi10241, pi10242, pi10243, pi10244, pi10245, pi10246, pi10247, pi10248, pi10249, pi10250, pi10251, pi10252, pi10253, pi10254, pi10255, pi10256, pi10257, pi10258, pi10259, pi10260, pi10261, pi10262, pi10263, pi10264, pi10265, pi10266, pi10267, pi10268, pi10269, pi10270, pi10271, pi10272, pi10273, pi10274, pi10275, pi10276, pi10277, pi10278, pi10279, pi10280, pi10281, pi10282, pi10283, pi10284, pi10285, pi10286, pi10287, pi10288, pi10289, pi10290, pi10291, pi10292, pi10293, pi10294, pi10295, pi10296, pi10297, pi10298, pi10299, pi10300, pi10301, pi10302, pi10303, pi10304, pi10305, pi10306, pi10307, pi10308, pi10309, pi10310, pi10311, pi10312, pi10313, pi10314, pi10315, pi10316, pi10317, pi10318, pi10319, pi10320, pi10321, pi10322, pi10323, pi10324, pi10325, pi10326, pi10327, pi10328, pi10329, pi10330, pi10331, pi10332, pi10333, pi10334, pi10335, pi10336, pi10337, pi10338, pi10339, pi10340, pi10341, pi10342, pi10343, pi10344, pi10345, pi10346, pi10347, pi10348, pi10349, pi10350, pi10351, pi10352, pi10353, pi10354, pi10355, pi10356, pi10357, pi10358, pi10359, pi10360, pi10361, pi10362, pi10363, pi10364, pi10365, pi10366, pi10367, pi10368, pi10369, pi10370, pi10371, pi10372, pi10373, pi10374, pi10375, pi10376, pi10377, pi10378, pi10379, pi10380, pi10381, pi10382, pi10383, pi10384, pi10385, pi10386, pi10387, pi10388, pi10389, pi10390, pi10391, pi10392, pi10393, pi10394, pi10395, pi10396, pi10397, pi10398, pi10399, pi10400, pi10401, pi10402, pi10403, pi10404, pi10405, pi10406, pi10407, pi10408, pi10409, pi10410, pi10411, pi10412, pi10413, pi10414, pi10415, pi10416, pi10417, pi10418, pi10419, pi10420, pi10421, pi10422, pi10423, pi10424, pi10425, pi10426, pi10427, pi10428, pi10429, pi10430, pi10431, pi10432, pi10433, pi10434, pi10435, pi10436, pi10437, pi10438, pi10439, pi10440, pi10441, pi10442, pi10443, pi10444, pi10445, pi10446, pi10447, pi10448, pi10449, pi10450, pi10451, pi10452, pi10453, pi10454, pi10455, pi10456, pi10457, pi10458, pi10459, pi10460, pi10461, pi10462, pi10463, pi10464, pi10465, pi10466, pi10467, pi10468, pi10469, pi10470, pi10471, pi10472, pi10473, pi10474, pi10475, pi10476, pi10477, pi10478, pi10479, pi10480, pi10481, pi10482, pi10483, pi10484, pi10485, pi10486, pi10487, pi10488, pi10489, pi10490, pi10491, pi10492, pi10493, pi10494, pi10495, pi10496, pi10497, pi10498, pi10499, pi10500, pi10501, pi10502, pi10503, pi10504, pi10505, pi10506, pi10507, pi10508, pi10509, pi10510, pi10511, pi10512, pi10513, pi10514, pi10515, pi10516, pi10517, pi10518, pi10519, pi10520, pi10521, pi10522, pi10523, pi10524, pi10525, pi10526, pi10527, pi10528, pi10529, pi10530, pi10531, pi10532, pi10533, pi10534, pi10535, pi10536, pi10537, pi10538, pi10539, pi10540, pi10541, pi10542, pi10543, pi10544, pi10545, pi10546, pi10547, pi10548, pi10549, pi10550, pi10551, pi10552, pi10553, pi10554, pi10555, pi10556, pi10557, pi10558, pi10559, pi10560, pi10561, pi10562, pi10563, pi10564, pi10565, pi10566, pi10567, pi10568, pi10569, pi10570, pi10571, pi10572, pi10573, pi10574, pi10575, pi10576, pi10577, pi10578, pi10579, pi10580, pi10581, pi10582, pi10583, pi10584, pi10585, pi10586, pi10587, pi10588, pi10589, pi10590, pi10591, pi10592, pi10593, pi10594, pi10595, pi10596, pi10597, pi10598, pi10599, pi10600, pi10601, pi10602, pi10603, pi10604, pi10605, pi10606, pi10607, pi10608, pi10609, pi10610, pi10611, pi10612, pi10613, pi10614, pi10615, pi10616, pi10617, pi10618, pi10619, pi10620, pi10621, pi10622, pi10623, pi10624, pi10625, pi10626, pi10627, pi10628, pi10629, pi10630, pi10631, pi10632, pi10633, pi10634, pi10635, pi10636, pi10637, pi10638, pi10639, pi10640, pi10641, pi10642, pi10643, pi10644, pi10645, pi10646, pi10647, pi10648, pi10649, pi10650, pi10651, pi10652, pi10653, pi10654, pi10655, pi10656, pi10657, pi10658, pi10659, pi10660, pi10661, pi10662, pi10663, pi10664, pi10665, pi10666, pi10667, pi10668, pi10669, pi10670, pi10671, 
            po00000, po00001, po00002, po00003, po00004, po00005, po00006, po00007, po00008, po00009, po00010, po00011, po00012, po00013, po00014, po00015, po00016, po00017, po00018, po00019, po00020, po00021, po00022, po00023, po00024, po00025, po00026, po00027, po00028, po00029, po00030, po00031, po00032, po00033, po00034, po00035, po00036, po00037, po00038, po00039, po00040, po00041, po00042, po00043, po00044, po00045, po00046, po00047, po00048, po00049, po00050, po00051, po00052, po00053, po00054, po00055, po00056, po00057, po00058, po00059, po00060, po00061, po00062, po00063, po00064, po00065, po00066, po00067, po00068, po00069, po00070, po00071, po00072, po00073, po00074, po00075, po00076, po00077, po00078, po00079, po00080, po00081, po00082, po00083, po00084, po00085, po00086, po00087, po00088, po00089, po00090, po00091, po00092, po00093, po00094, po00095, po00096, po00097, po00098, po00099, po00100, po00101, po00102, po00103, po00104, po00105, po00106, po00107, po00108, po00109, po00110, po00111, po00112, po00113, po00114, po00115, po00116, po00117, po00118, po00119, po00120, po00121, po00122, po00123, po00124, po00125, po00126, po00127, po00128, po00129, po00130, po00131, po00132, po00133, po00134, po00135, po00136, po00137, po00138, po00139, po00140, po00141, po00142, po00143, po00144, po00145, po00146, po00147, po00148, po00149, po00150, po00151, po00152, po00153, po00154, po00155, po00156, po00157, po00158, po00159, po00160, po00161, po00162, po00163, po00164, po00165, po00166, po00167, po00168, po00169, po00170, po00171, po00172, po00173, po00174, po00175, po00176, po00177, po00178, po00179, po00180, po00181, po00182, po00183, po00184, po00185, po00186, po00187, po00188, po00189, po00190, po00191, po00192, po00193, po00194, po00195, po00196, po00197, po00198, po00199, po00200, po00201, po00202, po00203, po00204, po00205, po00206, po00207, po00208, po00209, po00210, po00211, po00212, po00213, po00214, po00215, po00216, po00217, po00218, po00219, po00220, po00221, po00222, po00223, po00224, po00225, po00226, po00227, po00228, po00229, po00230, po00231, po00232, po00233, po00234, po00235, po00236, po00237, po00238, po00239, po00240, po00241, po00242, po00243, po00244, po00245, po00246, po00247, po00248, po00249, po00250, po00251, po00252, po00253, po00254, po00255, po00256, po00257, po00258, po00259, po00260, po00261, po00262, po00263, po00264, po00265, po00266, po00267, po00268, po00269, po00270, po00271, po00272, po00273, po00274, po00275, po00276, po00277, po00278, po00279, po00280, po00281, po00282, po00283, po00284, po00285, po00286, po00287, po00288, po00289, po00290, po00291, po00292, po00293, po00294, po00295, po00296, po00297, po00298, po00299, po00300, po00301, po00302, po00303, po00304, po00305, po00306, po00307, po00308, po00309, po00310, po00311, po00312, po00313, po00314, po00315, po00316, po00317, po00318, po00319, po00320, po00321, po00322, po00323, po00324, po00325, po00326, po00327, po00328, po00329, po00330, po00331, po00332, po00333, po00334, po00335, po00336, po00337, po00338, po00339, po00340, po00341, po00342, po00343, po00344, po00345, po00346, po00347, po00348, po00349, po00350, po00351, po00352, po00353, po00354, po00355, po00356, po00357, po00358, po00359, po00360, po00361, po00362, po00363, po00364, po00365, po00366, po00367, po00368, po00369, po00370, po00371, po00372, po00373, po00374, po00375, po00376, po00377, po00378, po00379, po00380, po00381, po00382, po00383, po00384, po00385, po00386, po00387, po00388, po00389, po00390, po00391, po00392, po00393, po00394, po00395, po00396, po00397, po00398, po00399, po00400, po00401, po00402, po00403, po00404, po00405, po00406, po00407, po00408, po00409, po00410, po00411, po00412, po00413, po00414, po00415, po00416, po00417, po00418, po00419, po00420, po00421, po00422, po00423, po00424, po00425, po00426, po00427, po00428, po00429, po00430, po00431, po00432, po00433, po00434, po00435, po00436, po00437, po00438, po00439, po00440, po00441, po00442, po00443, po00444, po00445, po00446, po00447, po00448, po00449, po00450, po00451, po00452, po00453, po00454, po00455, po00456, po00457, po00458, po00459, po00460, po00461, po00462, po00463, po00464, po00465, po00466, po00467, po00468, po00469, po00470, po00471, po00472, po00473, po00474, po00475, po00476, po00477, po00478, po00479, po00480, po00481, po00482, po00483, po00484, po00485, po00486, po00487, po00488, po00489, po00490, po00491, po00492, po00493, po00494, po00495, po00496, po00497, po00498, po00499, po00500, po00501, po00502, po00503, po00504, po00505, po00506, po00507, po00508, po00509, po00510, po00511, po00512, po00513, po00514, po00515, po00516, po00517, po00518, po00519, po00520, po00521, po00522, po00523, po00524, po00525, po00526, po00527, po00528, po00529, po00530, po00531, po00532, po00533, po00534, po00535, po00536, po00537, po00538, po00539, po00540, po00541, po00542, po00543, po00544, po00545, po00546, po00547, po00548, po00549, po00550, po00551, po00552, po00553, po00554, po00555, po00556, po00557, po00558, po00559, po00560, po00561, po00562, po00563, po00564, po00565, po00566, po00567, po00568, po00569, po00570, po00571, po00572, po00573, po00574, po00575, po00576, po00577, po00578, po00579, po00580, po00581, po00582, po00583, po00584, po00585, po00586, po00587, po00588, po00589, po00590, po00591, po00592, po00593, po00594, po00595, po00596, po00597, po00598, po00599, po00600, po00601, po00602, po00603, po00604, po00605, po00606, po00607, po00608, po00609, po00610, po00611, po00612, po00613, po00614, po00615, po00616, po00617, po00618, po00619, po00620, po00621, po00622, po00623, po00624, po00625, po00626, po00627, po00628, po00629, po00630, po00631, po00632, po00633, po00634, po00635, po00636, po00637, po00638, po00639, po00640, po00641, po00642, po00643, po00644, po00645, po00646, po00647, po00648, po00649, po00650, po00651, po00652, po00653, po00654, po00655, po00656, po00657, po00658, po00659, po00660, po00661, po00662, po00663, po00664, po00665, po00666, po00667, po00668, po00669, po00670, po00671, po00672, po00673, po00674, po00675, po00676, po00677, po00678, po00679, po00680, po00681, po00682, po00683, po00684, po00685, po00686, po00687, po00688, po00689, po00690, po00691, po00692, po00693, po00694, po00695, po00696, po00697, po00698, po00699, po00700, po00701, po00702, po00703, po00704, po00705, po00706, po00707, po00708, po00709, po00710, po00711, po00712, po00713, po00714, po00715, po00716, po00717, po00718, po00719, po00720, po00721, po00722, po00723, po00724, po00725, po00726, po00727, po00728, po00729, po00730, po00731, po00732, po00733, po00734, po00735, po00736, po00737, po00738, po00739, po00740, po00741, po00742, po00743, po00744, po00745, po00746, po00747, po00748, po00749, po00750, po00751, po00752, po00753, po00754, po00755, po00756, po00757, po00758, po00759, po00760, po00761, po00762, po00763, po00764, po00765, po00766, po00767, po00768, po00769, po00770, po00771, po00772, po00773, po00774, po00775, po00776, po00777, po00778, po00779, po00780, po00781, po00782, po00783, po00784, po00785, po00786, po00787, po00788, po00789, po00790, po00791, po00792, po00793, po00794, po00795, po00796, po00797, po00798, po00799, po00800, po00801, po00802, po00803, po00804, po00805, po00806, po00807, po00808, po00809, po00810, po00811, po00812, po00813, po00814, po00815, po00816, po00817, po00818, po00819, po00820, po00821, po00822, po00823, po00824, po00825, po00826, po00827, po00828, po00829, po00830, po00831, po00832, po00833, po00834, po00835, po00836, po00837, po00838, po00839, po00840, po00841, po00842, po00843, po00844, po00845, po00846, po00847, po00848, po00849, po00850, po00851, po00852, po00853, po00854, po00855, po00856, po00857, po00858, po00859, po00860, po00861, po00862, po00863, po00864, po00865, po00866, po00867, po00868, po00869, po00870, po00871, po00872, po00873, po00874, po00875, po00876, po00877, po00878, po00879, po00880, po00881, po00882, po00883, po00884, po00885, po00886, po00887, po00888, po00889, po00890, po00891, po00892, po00893, po00894, po00895, po00896, po00897, po00898, po00899, po00900, po00901, po00902, po00903, po00904, po00905, po00906, po00907, po00908, po00909, po00910, po00911, po00912, po00913, po00914, po00915, po00916, po00917, po00918, po00919, po00920, po00921, po00922, po00923, po00924, po00925, po00926, po00927, po00928, po00929, po00930, po00931, po00932, po00933, po00934, po00935, po00936, po00937, po00938, po00939, po00940, po00941, po00942, po00943, po00944, po00945, po00946, po00947, po00948, po00949, po00950, po00951, po00952, po00953, po00954, po00955, po00956, po00957, po00958, po00959, po00960, po00961, po00962, po00963, po00964, po00965, po00966, po00967, po00968, po00969, po00970, po00971, po00972, po00973, po00974, po00975, po00976, po00977, po00978, po00979, po00980, po00981, po00982, po00983, po00984, po00985, po00986, po00987, po00988, po00989, po00990, po00991, po00992, po00993, po00994, po00995, po00996, po00997, po00998, po00999, po01000, po01001, po01002, po01003, po01004, po01005, po01006, po01007, po01008, po01009, po01010, po01011, po01012, po01013, po01014, po01015, po01016, po01017, po01018, po01019, po01020, po01021, po01022, po01023, po01024, po01025, po01026, po01027, po01028, po01029, po01030, po01031, po01032, po01033, po01034, po01035, po01036, po01037, po01038, po01039, po01040, po01041, po01042, po01043, po01044, po01045, po01046, po01047, po01048, po01049, po01050, po01051, po01052, po01053, po01054, po01055, po01056, po01057, po01058, po01059, po01060, po01061, po01062, po01063, po01064, po01065, po01066, po01067, po01068, po01069, po01070, po01071, po01072, po01073, po01074, po01075, po01076, po01077, po01078, po01079, po01080, po01081, po01082, po01083, po01084, po01085, po01086, po01087, po01088, po01089, po01090, po01091, po01092, po01093, po01094, po01095, po01096, po01097, po01098, po01099, po01100, po01101, po01102, po01103, po01104, po01105, po01106, po01107, po01108, po01109, po01110, po01111, po01112, po01113, po01114, po01115, po01116, po01117, po01118, po01119, po01120, po01121, po01122, po01123, po01124, po01125, po01126, po01127, po01128, po01129, po01130, po01131, po01132, po01133, po01134, po01135, po01136, po01137, po01138, po01139, po01140, po01141, po01142, po01143, po01144, po01145, po01146, po01147, po01148, po01149, po01150, po01151, po01152, po01153, po01154, po01155, po01156, po01157, po01158, po01159, po01160, po01161, po01162, po01163, po01164, po01165, po01166, po01167, po01168, po01169, po01170, po01171, po01172, po01173, po01174, po01175, po01176, po01177, po01178, po01179, po01180, po01181, po01182, po01183, po01184, po01185, po01186, po01187, po01188, po01189, po01190, po01191, po01192, po01193, po01194, po01195, po01196, po01197, po01198, po01199, po01200, po01201, po01202, po01203, po01204, po01205, po01206, po01207, po01208, po01209, po01210, po01211, po01212, po01213, po01214, po01215, po01216, po01217, po01218, po01219, po01220, po01221, po01222, po01223, po01224, po01225, po01226, po01227, po01228, po01229, po01230, po01231, po01232, po01233, po01234, po01235, po01236, po01237, po01238, po01239, po01240, po01241, po01242, po01243, po01244, po01245, po01246, po01247, po01248, po01249, po01250, po01251, po01252, po01253, po01254, po01255, po01256, po01257, po01258, po01259, po01260, po01261, po01262, po01263, po01264, po01265, po01266, po01267, po01268, po01269, po01270, po01271, po01272, po01273, po01274, po01275, po01276, po01277, po01278, po01279, po01280, po01281, po01282, po01283, po01284, po01285, po01286, po01287, po01288, po01289, po01290, po01291, po01292, po01293, po01294, po01295, po01296, po01297, po01298, po01299, po01300, po01301, po01302, po01303, po01304, po01305, po01306, po01307, po01308, po01309, po01310, po01311, po01312, po01313, po01314, po01315, po01316, po01317, po01318, po01319, po01320, po01321, po01322, po01323, po01324, po01325, po01326, po01327, po01328, po01329, po01330, po01331, po01332, po01333, po01334, po01335, po01336, po01337, po01338, po01339, po01340, po01341, po01342, po01343, po01344, po01345, po01346, po01347, po01348, po01349, po01350, po01351, po01352, po01353, po01354, po01355, po01356, po01357, po01358, po01359, po01360, po01361, po01362, po01363, po01364, po01365, po01366, po01367, po01368, po01369, po01370, po01371, po01372, po01373, po01374, po01375, po01376, po01377, po01378, po01379, po01380, po01381, po01382, po01383, po01384, po01385, po01386, po01387, po01388, po01389, po01390, po01391, po01392, po01393, po01394, po01395, po01396, po01397, po01398, po01399, po01400, po01401, po01402, po01403, po01404, po01405, po01406, po01407, po01408, po01409, po01410, po01411, po01412, po01413, po01414, po01415, po01416, po01417, po01418, po01419, po01420, po01421, po01422, po01423, po01424, po01425, po01426, po01427, po01428, po01429, po01430, po01431, po01432, po01433, po01434, po01435, po01436, po01437, po01438, po01439, po01440, po01441, po01442, po01443, po01444, po01445, po01446, po01447, po01448, po01449, po01450, po01451, po01452, po01453, po01454, po01455, po01456, po01457, po01458, po01459, po01460, po01461, po01462, po01463, po01464, po01465, po01466, po01467, po01468, po01469, po01470, po01471, po01472, po01473, po01474, po01475, po01476, po01477, po01478, po01479, po01480, po01481, po01482, po01483, po01484, po01485, po01486, po01487, po01488, po01489, po01490, po01491, po01492, po01493, po01494, po01495, po01496, po01497, po01498, po01499, po01500, po01501, po01502, po01503, po01504, po01505, po01506, po01507, po01508, po01509, po01510, po01511, po01512, po01513, po01514, po01515, po01516, po01517, po01518, po01519, po01520, po01521, po01522, po01523, po01524, po01525, po01526, po01527, po01528, po01529, po01530, po01531, po01532, po01533, po01534, po01535, po01536, po01537, po01538, po01539, po01540, po01541, po01542, po01543, po01544, po01545, po01546, po01547, po01548, po01549, po01550, po01551, po01552, po01553, po01554, po01555, po01556, po01557, po01558, po01559, po01560, po01561, po01562, po01563, po01564, po01565, po01566, po01567, po01568, po01569, po01570, po01571, po01572, po01573, po01574, po01575, po01576, po01577, po01578, po01579, po01580, po01581, po01582, po01583, po01584, po01585, po01586, po01587, po01588, po01589, po01590, po01591, po01592, po01593, po01594, po01595, po01596, po01597, po01598, po01599, po01600, po01601, po01602, po01603, po01604, po01605, po01606, po01607, po01608, po01609, po01610, po01611, po01612, po01613, po01614, po01615, po01616, po01617, po01618, po01619, po01620, po01621, po01622, po01623, po01624, po01625, po01626, po01627, po01628, po01629, po01630, po01631, po01632, po01633, po01634, po01635, po01636, po01637, po01638, po01639, po01640, po01641, po01642, po01643, po01644, po01645, po01646, po01647, po01648, po01649, po01650, po01651, po01652, po01653, po01654, po01655, po01656, po01657, po01658, po01659, po01660, po01661, po01662, po01663, po01664, po01665, po01666, po01667, po01668, po01669, po01670, po01671, po01672, po01673, po01674, po01675, po01676, po01677, po01678, po01679, po01680, po01681, po01682, po01683, po01684, po01685, po01686, po01687, po01688, po01689, po01690, po01691, po01692, po01693, po01694, po01695, po01696, po01697, po01698, po01699, po01700, po01701, po01702, po01703, po01704, po01705, po01706, po01707, po01708, po01709, po01710, po01711, po01712, po01713, po01714, po01715, po01716, po01717, po01718, po01719, po01720, po01721, po01722, po01723, po01724, po01725, po01726, po01727, po01728, po01729, po01730, po01731, po01732, po01733, po01734, po01735, po01736, po01737, po01738, po01739, po01740, po01741, po01742, po01743, po01744, po01745, po01746, po01747, po01748, po01749, po01750, po01751, po01752, po01753, po01754, po01755, po01756, po01757, po01758, po01759, po01760, po01761, po01762, po01763, po01764, po01765, po01766, po01767, po01768, po01769, po01770, po01771, po01772, po01773, po01774, po01775, po01776, po01777, po01778, po01779, po01780, po01781, po01782, po01783, po01784, po01785, po01786, po01787, po01788, po01789, po01790, po01791, po01792, po01793, po01794, po01795, po01796, po01797, po01798, po01799, po01800, po01801, po01802, po01803, po01804, po01805, po01806, po01807, po01808, po01809, po01810, po01811, po01812, po01813, po01814, po01815, po01816, po01817, po01818, po01819, po01820, po01821, po01822, po01823, po01824, po01825, po01826, po01827, po01828, po01829, po01830, po01831, po01832, po01833, po01834, po01835, po01836, po01837, po01838, po01839, po01840, po01841, po01842, po01843, po01844, po01845, po01846, po01847, po01848, po01849, po01850, po01851, po01852, po01853, po01854, po01855, po01856, po01857, po01858, po01859, po01860, po01861, po01862, po01863, po01864, po01865, po01866, po01867, po01868, po01869, po01870, po01871, po01872, po01873, po01874, po01875, po01876, po01877, po01878, po01879, po01880, po01881, po01882, po01883, po01884, po01885, po01886, po01887, po01888, po01889, po01890, po01891, po01892, po01893, po01894, po01895, po01896, po01897, po01898, po01899, po01900, po01901, po01902, po01903, po01904, po01905, po01906, po01907, po01908, po01909, po01910, po01911, po01912, po01913, po01914, po01915, po01916, po01917, po01918, po01919, po01920, po01921, po01922, po01923, po01924, po01925, po01926, po01927, po01928, po01929, po01930, po01931, po01932, po01933, po01934, po01935, po01936, po01937, po01938, po01939, po01940, po01941, po01942, po01943, po01944, po01945, po01946, po01947, po01948, po01949, po01950, po01951, po01952, po01953, po01954, po01955, po01956, po01957, po01958, po01959, po01960, po01961, po01962, po01963, po01964, po01965, po01966, po01967, po01968, po01969, po01970, po01971, po01972, po01973, po01974, po01975, po01976, po01977, po01978, po01979, po01980, po01981, po01982, po01983, po01984, po01985, po01986, po01987, po01988, po01989, po01990, po01991, po01992, po01993, po01994, po01995, po01996, po01997, po01998, po01999, po02000, po02001, po02002, po02003, po02004, po02005, po02006, po02007, po02008, po02009, po02010, po02011, po02012, po02013, po02014, po02015, po02016, po02017, po02018, po02019, po02020, po02021, po02022, po02023, po02024, po02025, po02026, po02027, po02028, po02029, po02030, po02031, po02032, po02033, po02034, po02035, po02036, po02037, po02038, po02039, po02040, po02041, po02042, po02043, po02044, po02045, po02046, po02047, po02048, po02049, po02050, po02051, po02052, po02053, po02054, po02055, po02056, po02057, po02058, po02059, po02060, po02061, po02062, po02063, po02064, po02065, po02066, po02067, po02068, po02069, po02070, po02071, po02072, po02073, po02074, po02075, po02076, po02077, po02078, po02079, po02080, po02081, po02082, po02083, po02084, po02085, po02086, po02087, po02088, po02089, po02090, po02091, po02092, po02093, po02094, po02095, po02096, po02097, po02098, po02099, po02100, po02101, po02102, po02103, po02104, po02105, po02106, po02107, po02108, po02109, po02110, po02111, po02112, po02113, po02114, po02115, po02116, po02117, po02118, po02119, po02120, po02121, po02122, po02123, po02124, po02125, po02126, po02127, po02128, po02129, po02130, po02131, po02132, po02133, po02134, po02135, po02136, po02137, po02138, po02139, po02140, po02141, po02142, po02143, po02144, po02145, po02146, po02147, po02148, po02149, po02150, po02151, po02152, po02153, po02154, po02155, po02156, po02157, po02158, po02159, po02160, po02161, po02162, po02163, po02164, po02165, po02166, po02167, po02168, po02169, po02170, po02171, po02172, po02173, po02174, po02175, po02176, po02177, po02178, po02179, po02180, po02181, po02182, po02183, po02184, po02185, po02186, po02187, po02188, po02189, po02190, po02191, po02192, po02193, po02194, po02195, po02196, po02197, po02198, po02199, po02200, po02201, po02202, po02203, po02204, po02205, po02206, po02207, po02208, po02209, po02210, po02211, po02212, po02213, po02214, po02215, po02216, po02217, po02218, po02219, po02220, po02221, po02222, po02223, po02224, po02225, po02226, po02227, po02228, po02229, po02230, po02231, po02232, po02233, po02234, po02235, po02236, po02237, po02238, po02239, po02240, po02241, po02242, po02243, po02244, po02245, po02246, po02247, po02248, po02249, po02250, po02251, po02252, po02253, po02254, po02255, po02256, po02257, po02258, po02259, po02260, po02261, po02262, po02263, po02264, po02265, po02266, po02267, po02268, po02269, po02270, po02271, po02272, po02273, po02274, po02275, po02276, po02277, po02278, po02279, po02280, po02281, po02282, po02283, po02284, po02285, po02286, po02287, po02288, po02289, po02290, po02291, po02292, po02293, po02294, po02295, po02296, po02297, po02298, po02299, po02300, po02301, po02302, po02303, po02304, po02305, po02306, po02307, po02308, po02309, po02310, po02311, po02312, po02313, po02314, po02315, po02316, po02317, po02318, po02319, po02320, po02321, po02322, po02323, po02324, po02325, po02326, po02327, po02328, po02329, po02330, po02331, po02332, po02333, po02334, po02335, po02336, po02337, po02338, po02339, po02340, po02341, po02342, po02343, po02344, po02345, po02346, po02347, po02348, po02349, po02350, po02351, po02352, po02353, po02354, po02355, po02356, po02357, po02358, po02359, po02360, po02361, po02362, po02363, po02364, po02365, po02366, po02367, po02368, po02369, po02370, po02371, po02372, po02373, po02374, po02375, po02376, po02377, po02378, po02379, po02380, po02381, po02382, po02383, po02384, po02385, po02386, po02387, po02388, po02389, po02390, po02391, po02392, po02393, po02394, po02395, po02396, po02397, po02398, po02399, po02400, po02401, po02402, po02403, po02404, po02405, po02406, po02407, po02408, po02409, po02410, po02411, po02412, po02413, po02414, po02415, po02416, po02417, po02418, po02419, po02420, po02421, po02422, po02423, po02424, po02425, po02426, po02427, po02428, po02429, po02430, po02431, po02432, po02433, po02434, po02435, po02436, po02437, po02438, po02439, po02440, po02441, po02442, po02443, po02444, po02445, po02446, po02447, po02448, po02449, po02450, po02451, po02452, po02453, po02454, po02455, po02456, po02457, po02458, po02459, po02460, po02461, po02462, po02463, po02464, po02465, po02466, po02467, po02468, po02469, po02470, po02471, po02472, po02473, po02474, po02475, po02476, po02477, po02478, po02479, po02480, po02481, po02482, po02483, po02484, po02485, po02486, po02487, po02488, po02489, po02490, po02491, po02492, po02493, po02494, po02495, po02496, po02497, po02498, po02499, po02500, po02501, po02502, po02503, po02504, po02505, po02506, po02507, po02508, po02509, po02510, po02511, po02512, po02513, po02514, po02515, po02516, po02517, po02518, po02519, po02520, po02521, po02522, po02523, po02524, po02525, po02526, po02527, po02528, po02529, po02530, po02531, po02532, po02533, po02534, po02535, po02536, po02537, po02538, po02539, po02540, po02541, po02542, po02543, po02544, po02545, po02546, po02547, po02548, po02549, po02550, po02551, po02552, po02553, po02554, po02555, po02556, po02557, po02558, po02559, po02560, po02561, po02562, po02563, po02564, po02565, po02566, po02567, po02568, po02569, po02570, po02571, po02572, po02573, po02574, po02575, po02576, po02577, po02578, po02579, po02580, po02581, po02582, po02583, po02584, po02585, po02586, po02587, po02588, po02589, po02590, po02591, po02592, po02593, po02594, po02595, po02596, po02597, po02598, po02599, po02600, po02601, po02602, po02603, po02604, po02605, po02606, po02607, po02608, po02609, po02610, po02611, po02612, po02613, po02614, po02615, po02616, po02617, po02618, po02619, po02620, po02621, po02622, po02623, po02624, po02625, po02626, po02627, po02628, po02629, po02630, po02631, po02632, po02633, po02634, po02635, po02636, po02637, po02638, po02639, po02640, po02641, po02642, po02643, po02644, po02645, po02646, po02647, po02648, po02649, po02650, po02651, po02652, po02653, po02654, po02655, po02656, po02657, po02658, po02659, po02660, po02661, po02662, po02663, po02664, po02665, po02666, po02667, po02668, po02669, po02670, po02671, po02672, po02673, po02674, po02675, po02676, po02677, po02678, po02679, po02680, po02681, po02682, po02683, po02684, po02685, po02686, po02687, po02688, po02689, po02690, po02691, po02692, po02693, po02694, po02695, po02696, po02697, po02698, po02699, po02700, po02701, po02702, po02703, po02704, po02705, po02706, po02707, po02708, po02709, po02710, po02711, po02712, po02713, po02714, po02715, po02716, po02717, po02718, po02719, po02720, po02721, po02722, po02723, po02724, po02725, po02726, po02727, po02728, po02729, po02730, po02731, po02732, po02733, po02734, po02735, po02736, po02737, po02738, po02739, po02740, po02741, po02742, po02743, po02744, po02745, po02746, po02747, po02748, po02749, po02750, po02751, po02752, po02753, po02754, po02755, po02756, po02757, po02758, po02759, po02760, po02761, po02762, po02763, po02764, po02765, po02766, po02767, po02768, po02769, po02770, po02771, po02772, po02773, po02774, po02775, po02776, po02777, po02778, po02779, po02780, po02781, po02782, po02783, po02784, po02785, po02786, po02787, po02788, po02789, po02790, po02791, po02792, po02793, po02794, po02795, po02796, po02797, po02798, po02799, po02800, po02801, po02802, po02803, po02804, po02805, po02806, po02807, po02808, po02809, po02810, po02811, po02812, po02813, po02814, po02815, po02816, po02817, po02818, po02819, po02820, po02821, po02822, po02823, po02824, po02825, po02826, po02827, po02828, po02829, po02830, po02831, po02832, po02833, po02834, po02835, po02836, po02837, po02838, po02839, po02840, po02841, po02842, po02843, po02844, po02845, po02846, po02847, po02848, po02849, po02850, po02851, po02852, po02853, po02854, po02855, po02856, po02857, po02858, po02859, po02860, po02861, po02862, po02863, po02864, po02865, po02866, po02867, po02868, po02869, po02870, po02871, po02872, po02873, po02874, po02875, po02876, po02877, po02878, po02879, po02880, po02881, po02882, po02883, po02884, po02885, po02886, po02887, po02888, po02889, po02890, po02891, po02892, po02893, po02894, po02895, po02896, po02897, po02898, po02899, po02900, po02901, po02902, po02903, po02904, po02905, po02906, po02907, po02908, po02909, po02910, po02911, po02912, po02913, po02914, po02915, po02916, po02917, po02918, po02919, po02920, po02921, po02922, po02923, po02924, po02925, po02926, po02927, po02928, po02929, po02930, po02931, po02932, po02933, po02934, po02935, po02936, po02937, po02938, po02939, po02940, po02941, po02942, po02943, po02944, po02945, po02946, po02947, po02948, po02949, po02950, po02951, po02952, po02953, po02954, po02955, po02956, po02957, po02958, po02959, po02960, po02961, po02962, po02963, po02964, po02965, po02966, po02967, po02968, po02969, po02970, po02971, po02972, po02973, po02974, po02975, po02976, po02977, po02978, po02979, po02980, po02981, po02982, po02983, po02984, po02985, po02986, po02987, po02988, po02989, po02990, po02991, po02992, po02993, po02994, po02995, po02996, po02997, po02998, po02999, po03000, po03001, po03002, po03003, po03004, po03005, po03006, po03007, po03008, po03009, po03010, po03011, po03012, po03013, po03014, po03015, po03016, po03017, po03018, po03019, po03020, po03021, po03022, po03023, po03024, po03025, po03026, po03027, po03028, po03029, po03030, po03031, po03032, po03033, po03034, po03035, po03036, po03037, po03038, po03039, po03040, po03041, po03042, po03043, po03044, po03045, po03046, po03047, po03048, po03049, po03050, po03051, po03052, po03053, po03054, po03055, po03056, po03057, po03058, po03059, po03060, po03061, po03062, po03063, po03064, po03065, po03066, po03067, po03068, po03069, po03070, po03071, po03072, po03073, po03074, po03075, po03076, po03077, po03078, po03079, po03080, po03081, po03082, po03083, po03084, po03085, po03086, po03087, po03088, po03089, po03090, po03091, po03092, po03093, po03094, po03095, po03096, po03097, po03098, po03099, po03100, po03101, po03102, po03103, po03104, po03105, po03106, po03107, po03108, po03109, po03110, po03111, po03112, po03113, po03114, po03115, po03116, po03117, po03118, po03119, po03120, po03121, po03122, po03123, po03124, po03125, po03126, po03127, po03128, po03129, po03130, po03131, po03132, po03133, po03134, po03135, po03136, po03137, po03138, po03139, po03140, po03141, po03142, po03143, po03144, po03145, po03146, po03147, po03148, po03149, po03150, po03151, po03152, po03153, po03154, po03155, po03156, po03157, po03158, po03159, po03160, po03161, po03162, po03163, po03164, po03165, po03166, po03167, po03168, po03169, po03170, po03171, po03172, po03173, po03174, po03175, po03176, po03177, po03178, po03179, po03180, po03181, po03182, po03183, po03184, po03185, po03186, po03187, po03188, po03189, po03190, po03191, po03192, po03193, po03194, po03195, po03196, po03197, po03198, po03199, po03200, po03201, po03202, po03203, po03204, po03205, po03206, po03207, po03208, po03209, po03210, po03211, po03212, po03213, po03214, po03215, po03216, po03217, po03218, po03219, po03220, po03221, po03222, po03223, po03224, po03225, po03226, po03227, po03228, po03229, po03230, po03231, po03232, po03233, po03234, po03235, po03236, po03237, po03238, po03239, po03240, po03241, po03242, po03243, po03244, po03245, po03246, po03247, po03248, po03249, po03250, po03251, po03252, po03253, po03254, po03255, po03256, po03257, po03258, po03259, po03260, po03261, po03262, po03263, po03264, po03265, po03266, po03267, po03268, po03269, po03270, po03271, po03272, po03273, po03274, po03275, po03276, po03277, po03278, po03279, po03280, po03281, po03282, po03283, po03284, po03285, po03286, po03287, po03288, po03289, po03290, po03291, po03292, po03293, po03294, po03295, po03296, po03297, po03298, po03299, po03300, po03301, po03302, po03303, po03304, po03305, po03306, po03307, po03308, po03309, po03310, po03311, po03312, po03313, po03314, po03315, po03316, po03317, po03318, po03319, po03320, po03321, po03322, po03323, po03324, po03325, po03326, po03327, po03328, po03329, po03330, po03331, po03332, po03333, po03334, po03335, po03336, po03337, po03338, po03339, po03340, po03341, po03342, po03343, po03344, po03345, po03346, po03347, po03348, po03349, po03350, po03351, po03352, po03353, po03354, po03355, po03356, po03357, po03358, po03359, po03360, po03361, po03362, po03363, po03364, po03365, po03366, po03367, po03368, po03369, po03370, po03371, po03372, po03373, po03374, po03375, po03376, po03377, po03378, po03379, po03380, po03381, po03382, po03383, po03384, po03385, po03386, po03387, po03388, po03389, po03390, po03391, po03392, po03393, po03394, po03395, po03396, po03397, po03398, po03399, po03400, po03401, po03402, po03403, po03404, po03405, po03406, po03407, po03408, po03409, po03410, po03411, po03412, po03413, po03414, po03415, po03416, po03417, po03418, po03419, po03420, po03421, po03422, po03423, po03424, po03425, po03426, po03427, po03428, po03429, po03430, po03431, po03432, po03433, po03434, po03435, po03436, po03437, po03438, po03439, po03440, po03441, po03442, po03443, po03444, po03445, po03446, po03447, po03448, po03449, po03450, po03451, po03452, po03453, po03454, po03455, po03456, po03457, po03458, po03459, po03460, po03461, po03462, po03463, po03464, po03465, po03466, po03467, po03468, po03469, po03470, po03471, po03472, po03473, po03474, po03475, po03476, po03477, po03478, po03479, po03480, po03481, po03482, po03483, po03484, po03485, po03486, po03487, po03488, po03489, po03490, po03491, po03492, po03493, po03494, po03495, po03496, po03497, po03498, po03499, po03500, po03501, po03502, po03503, po03504, po03505, po03506, po03507, po03508, po03509, po03510, po03511, po03512, po03513, po03514, po03515, po03516, po03517, po03518, po03519, po03520, po03521, po03522, po03523, po03524, po03525, po03526, po03527, po03528, po03529, po03530, po03531, po03532, po03533, po03534, po03535, po03536, po03537, po03538, po03539, po03540, po03541, po03542, po03543, po03544, po03545, po03546, po03547, po03548, po03549, po03550, po03551, po03552, po03553, po03554, po03555, po03556, po03557, po03558, po03559, po03560, po03561, po03562, po03563, po03564, po03565, po03566, po03567, po03568, po03569, po03570, po03571, po03572, po03573, po03574, po03575, po03576, po03577, po03578, po03579, po03580, po03581, po03582, po03583, po03584, po03585, po03586, po03587, po03588, po03589, po03590, po03591, po03592, po03593, po03594, po03595, po03596, po03597, po03598, po03599, po03600, po03601, po03602, po03603, po03604, po03605, po03606, po03607, po03608, po03609, po03610, po03611, po03612, po03613, po03614, po03615, po03616, po03617, po03618, po03619, po03620, po03621, po03622, po03623, po03624, po03625, po03626, po03627, po03628, po03629, po03630, po03631, po03632, po03633, po03634, po03635, po03636, po03637, po03638, po03639, po03640, po03641, po03642, po03643, po03644, po03645, po03646, po03647, po03648, po03649, po03650, po03651, po03652, po03653, po03654, po03655, po03656, po03657, po03658, po03659, po03660, po03661, po03662, po03663, po03664, po03665, po03666, po03667, po03668, po03669, po03670, po03671, po03672, po03673, po03674, po03675, po03676, po03677, po03678, po03679, po03680, po03681, po03682, po03683, po03684, po03685, po03686, po03687, po03688, po03689, po03690, po03691, po03692, po03693, po03694, po03695, po03696, po03697, po03698, po03699, po03700, po03701, po03702, po03703, po03704, po03705, po03706, po03707, po03708, po03709, po03710, po03711, po03712, po03713, po03714, po03715, po03716, po03717, po03718, po03719, po03720, po03721, po03722, po03723, po03724, po03725, po03726, po03727, po03728, po03729, po03730, po03731, po03732, po03733, po03734, po03735, po03736, po03737, po03738, po03739, po03740, po03741, po03742, po03743, po03744, po03745, po03746, po03747, po03748, po03749, po03750, po03751, po03752, po03753, po03754, po03755, po03756, po03757, po03758, po03759, po03760, po03761, po03762, po03763, po03764, po03765, po03766, po03767, po03768, po03769, po03770, po03771, po03772, po03773, po03774, po03775, po03776, po03777, po03778, po03779, po03780, po03781, po03782, po03783, po03784, po03785, po03786, po03787, po03788, po03789, po03790, po03791, po03792, po03793, po03794, po03795, po03796, po03797, po03798, po03799, po03800, po03801, po03802, po03803, po03804, po03805, po03806, po03807, po03808, po03809, po03810, po03811, po03812, po03813, po03814, po03815, po03816, po03817, po03818, po03819, po03820, po03821, po03822, po03823, po03824, po03825, po03826, po03827, po03828, po03829, po03830, po03831, po03832, po03833, po03834, po03835, po03836, po03837, po03838, po03839, po03840, po03841, po03842, po03843, po03844, po03845, po03846, po03847, po03848, po03849, po03850, po03851, po03852, po03853, po03854, po03855, po03856, po03857, po03858, po03859, po03860, po03861, po03862, po03863, po03864, po03865, po03866, po03867, po03868, po03869, po03870, po03871, po03872, po03873, po03874, po03875, po03876, po03877, po03878, po03879, po03880, po03881, po03882, po03883, po03884, po03885, po03886, po03887, po03888, po03889, po03890, po03891, po03892, po03893, po03894, po03895, po03896, po03897, po03898, po03899, po03900, po03901, po03902, po03903, po03904, po03905, po03906, po03907, po03908, po03909, po03910, po03911, po03912, po03913, po03914, po03915, po03916, po03917, po03918, po03919, po03920, po03921, po03922, po03923, po03924, po03925, po03926, po03927, po03928, po03929, po03930, po03931, po03932, po03933, po03934, po03935, po03936, po03937, po03938, po03939, po03940, po03941, po03942, po03943, po03944, po03945, po03946, po03947, po03948, po03949, po03950, po03951, po03952, po03953, po03954, po03955, po03956, po03957, po03958, po03959, po03960, po03961, po03962, po03963, po03964, po03965, po03966, po03967, po03968, po03969, po03970, po03971, po03972, po03973, po03974, po03975, po03976, po03977, po03978, po03979, po03980, po03981, po03982, po03983, po03984, po03985, po03986, po03987, po03988, po03989, po03990, po03991, po03992, po03993, po03994, po03995, po03996, po03997, po03998, po03999, po04000, po04001, po04002, po04003, po04004, po04005, po04006, po04007, po04008, po04009, po04010, po04011, po04012, po04013, po04014, po04015, po04016, po04017, po04018, po04019, po04020, po04021, po04022, po04023, po04024, po04025, po04026, po04027, po04028, po04029, po04030, po04031, po04032, po04033, po04034, po04035, po04036, po04037, po04038, po04039, po04040, po04041, po04042, po04043, po04044, po04045, po04046, po04047, po04048, po04049, po04050, po04051, po04052, po04053, po04054, po04055, po04056, po04057, po04058, po04059, po04060, po04061, po04062, po04063, po04064, po04065, po04066, po04067, po04068, po04069, po04070, po04071, po04072, po04073, po04074, po04075, po04076, po04077, po04078, po04079, po04080, po04081, po04082, po04083, po04084, po04085, po04086, po04087, po04088, po04089, po04090, po04091, po04092, po04093, po04094, po04095, po04096, po04097, po04098, po04099, po04100, po04101, po04102, po04103, po04104, po04105, po04106, po04107, po04108, po04109, po04110, po04111, po04112, po04113, po04114, po04115, po04116, po04117, po04118, po04119, po04120, po04121, po04122, po04123, po04124, po04125, po04126, po04127, po04128, po04129, po04130, po04131, po04132, po04133, po04134, po04135, po04136, po04137, po04138, po04139, po04140, po04141, po04142, po04143, po04144, po04145, po04146, po04147, po04148, po04149, po04150, po04151, po04152, po04153, po04154, po04155, po04156, po04157, po04158, po04159, po04160, po04161, po04162, po04163, po04164, po04165, po04166, po04167, po04168, po04169, po04170, po04171, po04172, po04173, po04174, po04175, po04176, po04177, po04178, po04179, po04180, po04181, po04182, po04183, po04184, po04185, po04186, po04187, po04188, po04189, po04190, po04191, po04192, po04193, po04194, po04195, po04196, po04197, po04198, po04199, po04200, po04201, po04202, po04203, po04204, po04205, po04206, po04207, po04208, po04209, po04210, po04211, po04212, po04213, po04214, po04215, po04216, po04217, po04218, po04219, po04220, po04221, po04222, po04223, po04224, po04225, po04226, po04227, po04228, po04229, po04230, po04231, po04232, po04233, po04234, po04235, po04236, po04237, po04238, po04239, po04240, po04241, po04242, po04243, po04244, po04245, po04246, po04247, po04248, po04249, po04250, po04251, po04252, po04253, po04254, po04255, po04256, po04257, po04258, po04259, po04260, po04261, po04262, po04263, po04264, po04265, po04266, po04267, po04268, po04269, po04270, po04271, po04272, po04273, po04274, po04275, po04276, po04277, po04278, po04279, po04280, po04281, po04282, po04283, po04284, po04285, po04286, po04287, po04288, po04289, po04290, po04291, po04292, po04293, po04294, po04295, po04296, po04297, po04298, po04299, po04300, po04301, po04302, po04303, po04304, po04305, po04306, po04307, po04308, po04309, po04310, po04311, po04312, po04313, po04314, po04315, po04316, po04317, po04318, po04319, po04320, po04321, po04322, po04323, po04324, po04325, po04326, po04327, po04328, po04329, po04330, po04331, po04332, po04333, po04334, po04335, po04336, po04337, po04338, po04339, po04340, po04341, po04342, po04343, po04344, po04345, po04346, po04347, po04348, po04349, po04350, po04351, po04352, po04353, po04354, po04355, po04356, po04357, po04358, po04359, po04360, po04361, po04362, po04363, po04364, po04365, po04366, po04367, po04368, po04369, po04370, po04371, po04372, po04373, po04374, po04375, po04376, po04377, po04378, po04379, po04380, po04381, po04382, po04383, po04384, po04385, po04386, po04387, po04388, po04389, po04390, po04391, po04392, po04393, po04394, po04395, po04396, po04397, po04398, po04399, po04400, po04401, po04402, po04403, po04404, po04405, po04406, po04407, po04408, po04409, po04410, po04411, po04412, po04413, po04414, po04415, po04416, po04417, po04418, po04419, po04420, po04421, po04422, po04423, po04424, po04425, po04426, po04427, po04428, po04429, po04430, po04431, po04432, po04433, po04434, po04435, po04436, po04437, po04438, po04439, po04440, po04441, po04442, po04443, po04444, po04445, po04446, po04447, po04448, po04449, po04450, po04451, po04452, po04453, po04454, po04455, po04456, po04457, po04458, po04459, po04460, po04461, po04462, po04463, po04464, po04465, po04466, po04467, po04468, po04469, po04470, po04471, po04472, po04473, po04474, po04475, po04476, po04477, po04478, po04479, po04480, po04481, po04482, po04483, po04484, po04485, po04486, po04487, po04488, po04489, po04490, po04491, po04492, po04493, po04494, po04495, po04496, po04497, po04498, po04499, po04500, po04501, po04502, po04503, po04504, po04505, po04506, po04507, po04508, po04509, po04510, po04511, po04512, po04513, po04514, po04515, po04516, po04517, po04518, po04519, po04520, po04521, po04522, po04523, po04524, po04525, po04526, po04527, po04528, po04529, po04530, po04531, po04532, po04533, po04534, po04535, po04536, po04537, po04538, po04539, po04540, po04541, po04542, po04543, po04544, po04545, po04546, po04547, po04548, po04549, po04550, po04551, po04552, po04553, po04554, po04555, po04556, po04557, po04558, po04559, po04560, po04561, po04562, po04563, po04564, po04565, po04566, po04567, po04568, po04569, po04570, po04571, po04572, po04573, po04574, po04575, po04576, po04577, po04578, po04579, po04580, po04581, po04582, po04583, po04584, po04585, po04586, po04587, po04588, po04589, po04590, po04591, po04592, po04593, po04594, po04595, po04596, po04597, po04598, po04599, po04600, po04601, po04602, po04603, po04604, po04605, po04606, po04607, po04608, po04609, po04610, po04611, po04612, po04613, po04614, po04615, po04616, po04617, po04618, po04619, po04620, po04621, po04622, po04623, po04624, po04625, po04626, po04627, po04628, po04629, po04630, po04631, po04632, po04633, po04634, po04635, po04636, po04637, po04638, po04639, po04640, po04641, po04642, po04643, po04644, po04645, po04646, po04647, po04648, po04649, po04650, po04651, po04652, po04653, po04654, po04655, po04656, po04657, po04658, po04659, po04660, po04661, po04662, po04663, po04664, po04665, po04666, po04667, po04668, po04669, po04670, po04671, po04672, po04673, po04674, po04675, po04676, po04677, po04678, po04679, po04680, po04681, po04682, po04683, po04684, po04685, po04686, po04687, po04688, po04689, po04690, po04691, po04692, po04693, po04694, po04695, po04696, po04697, po04698, po04699, po04700, po04701, po04702, po04703, po04704, po04705, po04706, po04707, po04708, po04709, po04710, po04711, po04712, po04713, po04714, po04715, po04716, po04717, po04718, po04719, po04720, po04721, po04722, po04723, po04724, po04725, po04726, po04727, po04728, po04729, po04730, po04731, po04732, po04733, po04734, po04735, po04736, po04737, po04738, po04739, po04740, po04741, po04742, po04743, po04744, po04745, po04746, po04747, po04748, po04749, po04750, po04751, po04752, po04753, po04754, po04755, po04756, po04757, po04758, po04759, po04760, po04761, po04762, po04763, po04764, po04765, po04766, po04767, po04768, po04769, po04770, po04771, po04772, po04773, po04774, po04775, po04776, po04777, po04778, po04779, po04780, po04781, po04782, po04783, po04784, po04785, po04786, po04787, po04788, po04789, po04790, po04791, po04792, po04793, po04794, po04795, po04796, po04797, po04798, po04799, po04800, po04801, po04802, po04803, po04804, po04805, po04806, po04807, po04808, po04809, po04810, po04811, po04812, po04813, po04814, po04815, po04816, po04817, po04818, po04819, po04820, po04821, po04822, po04823, po04824, po04825, po04826, po04827, po04828, po04829, po04830, po04831, po04832, po04833, po04834, po04835, po04836, po04837, po04838, po04839, po04840, po04841, po04842, po04843, po04844, po04845, po04846, po04847, po04848, po04849, po04850, po04851, po04852, po04853, po04854, po04855, po04856, po04857, po04858, po04859, po04860, po04861, po04862, po04863, po04864, po04865, po04866, po04867, po04868, po04869, po04870, po04871, po04872, po04873, po04874, po04875, po04876, po04877, po04878, po04879, po04880, po04881, po04882, po04883, po04884, po04885, po04886, po04887, po04888, po04889, po04890, po04891, po04892, po04893, po04894, po04895, po04896, po04897, po04898, po04899, po04900, po04901, po04902, po04903, po04904, po04905, po04906, po04907, po04908, po04909, po04910, po04911, po04912, po04913, po04914, po04915, po04916, po04917, po04918, po04919, po04920, po04921, po04922, po04923, po04924, po04925, po04926, po04927, po04928, po04929, po04930, po04931, po04932, po04933, po04934, po04935, po04936, po04937, po04938, po04939, po04940, po04941, po04942, po04943, po04944, po04945, po04946, po04947, po04948, po04949, po04950, po04951, po04952, po04953, po04954, po04955, po04956, po04957, po04958, po04959, po04960, po04961, po04962, po04963, po04964, po04965, po04966, po04967, po04968, po04969, po04970, po04971, po04972, po04973, po04974, po04975, po04976, po04977, po04978, po04979, po04980, po04981, po04982, po04983, po04984, po04985, po04986, po04987, po04988, po04989, po04990, po04991, po04992, po04993, po04994, po04995, po04996, po04997, po04998, po04999, po05000, po05001, po05002, po05003, po05004, po05005, po05006, po05007, po05008, po05009, po05010, po05011, po05012, po05013, po05014, po05015, po05016, po05017, po05018, po05019, po05020, po05021, po05022, po05023, po05024, po05025, po05026, po05027, po05028, po05029, po05030, po05031, po05032, po05033, po05034, po05035, po05036, po05037, po05038, po05039, po05040, po05041, po05042, po05043, po05044, po05045, po05046, po05047, po05048, po05049, po05050, po05051, po05052, po05053, po05054, po05055, po05056, po05057, po05058, po05059, po05060, po05061, po05062, po05063, po05064, po05065, po05066, po05067, po05068, po05069, po05070, po05071, po05072, po05073, po05074, po05075, po05076, po05077, po05078, po05079, po05080, po05081, po05082, po05083, po05084, po05085, po05086, po05087, po05088, po05089, po05090, po05091, po05092, po05093, po05094, po05095, po05096, po05097, po05098, po05099, po05100, po05101, po05102, po05103, po05104, po05105, po05106, po05107, po05108, po05109, po05110, po05111, po05112, po05113, po05114, po05115, po05116, po05117, po05118, po05119, po05120, po05121, po05122, po05123, po05124, po05125, po05126, po05127, po05128, po05129, po05130, po05131, po05132, po05133, po05134, po05135, po05136, po05137, po05138, po05139, po05140, po05141, po05142, po05143, po05144, po05145, po05146, po05147, po05148, po05149, po05150, po05151, po05152, po05153, po05154, po05155, po05156, po05157, po05158, po05159, po05160, po05161, po05162, po05163, po05164, po05165, po05166, po05167, po05168, po05169, po05170, po05171, po05172, po05173, po05174, po05175, po05176, po05177, po05178, po05179, po05180, po05181, po05182, po05183, po05184, po05185, po05186, po05187, po05188, po05189, po05190, po05191, po05192, po05193, po05194, po05195, po05196, po05197, po05198, po05199, po05200, po05201, po05202, po05203, po05204, po05205, po05206, po05207, po05208, po05209, po05210, po05211, po05212, po05213, po05214, po05215, po05216, po05217, po05218, po05219, po05220, po05221, po05222, po05223, po05224, po05225, po05226, po05227, po05228, po05229, po05230, po05231, po05232, po05233, po05234, po05235, po05236, po05237, po05238, po05239, po05240, po05241, po05242, po05243, po05244, po05245, po05246, po05247, po05248, po05249, po05250, po05251, po05252, po05253, po05254, po05255, po05256, po05257, po05258, po05259, po05260, po05261, po05262, po05263, po05264, po05265, po05266, po05267, po05268, po05269, po05270, po05271, po05272, po05273, po05274, po05275, po05276, po05277, po05278, po05279, po05280, po05281, po05282, po05283, po05284, po05285, po05286, po05287, po05288, po05289, po05290, po05291, po05292, po05293, po05294, po05295, po05296, po05297, po05298, po05299, po05300, po05301, po05302, po05303, po05304, po05305, po05306, po05307, po05308, po05309, po05310, po05311, po05312, po05313, po05314, po05315, po05316, po05317, po05318, po05319, po05320, po05321, po05322, po05323, po05324, po05325, po05326, po05327, po05328, po05329, po05330, po05331, po05332, po05333, po05334, po05335, po05336, po05337, po05338, po05339, po05340, po05341, po05342, po05343, po05344, po05345, po05346, po05347, po05348, po05349, po05350, po05351, po05352, po05353, po05354, po05355, po05356, po05357, po05358, po05359, po05360, po05361, po05362, po05363, po05364, po05365, po05366, po05367, po05368, po05369, po05370, po05371, po05372, po05373, po05374, po05375, po05376, po05377, po05378, po05379, po05380, po05381, po05382, po05383, po05384, po05385, po05386, po05387, po05388, po05389, po05390, po05391, po05392, po05393, po05394, po05395, po05396, po05397, po05398, po05399, po05400, po05401, po05402, po05403, po05404, po05405, po05406, po05407, po05408, po05409, po05410, po05411, po05412, po05413, po05414, po05415, po05416, po05417, po05418, po05419, po05420, po05421, po05422, po05423, po05424, po05425, po05426, po05427, po05428, po05429, po05430, po05431, po05432, po05433, po05434, po05435, po05436, po05437, po05438, po05439, po05440, po05441, po05442, po05443, po05444, po05445, po05446, po05447, po05448, po05449, po05450, po05451, po05452, po05453, po05454, po05455, po05456, po05457, po05458, po05459, po05460, po05461, po05462, po05463, po05464, po05465, po05466, po05467, po05468, po05469, po05470, po05471, po05472, po05473, po05474, po05475, po05476, po05477, po05478, po05479, po05480, po05481, po05482, po05483, po05484, po05485, po05486, po05487, po05488, po05489, po05490, po05491, po05492, po05493, po05494, po05495, po05496, po05497, po05498, po05499, po05500, po05501, po05502, po05503, po05504, po05505, po05506, po05507, po05508, po05509, po05510, po05511, po05512, po05513, po05514, po05515, po05516, po05517, po05518, po05519, po05520, po05521, po05522, po05523, po05524, po05525, po05526, po05527, po05528, po05529, po05530, po05531, po05532, po05533, po05534, po05535, po05536, po05537, po05538, po05539, po05540, po05541, po05542, po05543, po05544, po05545, po05546, po05547, po05548, po05549, po05550, po05551, po05552, po05553, po05554, po05555, po05556, po05557, po05558, po05559, po05560, po05561, po05562, po05563, po05564, po05565, po05566, po05567, po05568, po05569, po05570, po05571, po05572, po05573, po05574, po05575, po05576, po05577, po05578, po05579, po05580, po05581, po05582, po05583, po05584, po05585, po05586, po05587, po05588, po05589, po05590, po05591, po05592, po05593, po05594, po05595, po05596, po05597, po05598, po05599, po05600, po05601, po05602, po05603, po05604, po05605, po05606, po05607, po05608, po05609, po05610, po05611, po05612, po05613, po05614, po05615, po05616, po05617, po05618, po05619, po05620, po05621, po05622, po05623, po05624, po05625, po05626, po05627, po05628, po05629, po05630, po05631, po05632, po05633, po05634, po05635, po05636, po05637, po05638, po05639, po05640, po05641, po05642, po05643, po05644, po05645, po05646, po05647, po05648, po05649, po05650, po05651, po05652, po05653, po05654, po05655, po05656, po05657, po05658, po05659, po05660, po05661, po05662, po05663, po05664, po05665, po05666, po05667, po05668, po05669, po05670, po05671, po05672, po05673, po05674, po05675, po05676, po05677, po05678, po05679, po05680, po05681, po05682, po05683, po05684, po05685, po05686, po05687, po05688, po05689, po05690, po05691, po05692, po05693, po05694, po05695, po05696, po05697, po05698, po05699, po05700, po05701, po05702, po05703, po05704, po05705, po05706, po05707, po05708, po05709, po05710, po05711, po05712, po05713, po05714, po05715, po05716, po05717, po05718, po05719, po05720, po05721, po05722, po05723, po05724, po05725, po05726, po05727, po05728, po05729, po05730, po05731, po05732, po05733, po05734, po05735, po05736, po05737, po05738, po05739, po05740, po05741, po05742, po05743, po05744, po05745, po05746, po05747, po05748, po05749, po05750, po05751, po05752, po05753, po05754, po05755, po05756, po05757, po05758, po05759, po05760, po05761, po05762, po05763, po05764, po05765, po05766, po05767, po05768, po05769, po05770, po05771, po05772, po05773, po05774, po05775, po05776, po05777, po05778, po05779, po05780, po05781, po05782, po05783, po05784, po05785, po05786, po05787, po05788, po05789, po05790, po05791, po05792, po05793, po05794, po05795, po05796, po05797, po05798, po05799, po05800, po05801, po05802, po05803, po05804, po05805, po05806, po05807, po05808, po05809, po05810, po05811, po05812, po05813, po05814, po05815, po05816, po05817, po05818, po05819, po05820, po05821, po05822, po05823, po05824, po05825, po05826, po05827, po05828, po05829, po05830, po05831, po05832, po05833, po05834, po05835, po05836, po05837, po05838, po05839, po05840, po05841, po05842, po05843, po05844, po05845, po05846, po05847, po05848, po05849, po05850, po05851, po05852, po05853, po05854, po05855, po05856, po05857, po05858, po05859, po05860, po05861, po05862, po05863, po05864, po05865, po05866, po05867, po05868, po05869, po05870, po05871, po05872, po05873, po05874, po05875, po05876, po05877, po05878, po05879, po05880, po05881, po05882, po05883, po05884, po05885, po05886, po05887, po05888, po05889, po05890, po05891, po05892, po05893, po05894, po05895, po05896, po05897, po05898, po05899, po05900, po05901, po05902, po05903, po05904, po05905, po05906, po05907, po05908, po05909, po05910, po05911, po05912, po05913, po05914, po05915, po05916, po05917, po05918, po05919, po05920, po05921, po05922, po05923, po05924, po05925, po05926, po05927, po05928, po05929, po05930, po05931, po05932, po05933, po05934, po05935, po05936, po05937, po05938, po05939, po05940, po05941, po05942, po05943, po05944, po05945, po05946, po05947, po05948, po05949, po05950, po05951, po05952, po05953, po05954, po05955, po05956, po05957, po05958, po05959, po05960, po05961, po05962, po05963, po05964, po05965, po05966, po05967, po05968, po05969, po05970, po05971, po05972, po05973, po05974, po05975, po05976, po05977, po05978, po05979, po05980, po05981, po05982, po05983, po05984, po05985, po05986, po05987, po05988, po05989, po05990, po05991, po05992, po05993, po05994, po05995, po05996, po05997, po05998, po05999, po06000, po06001, po06002, po06003, po06004, po06005, po06006, po06007, po06008, po06009, po06010, po06011, po06012, po06013, po06014, po06015, po06016, po06017, po06018, po06019, po06020, po06021, po06022, po06023, po06024, po06025, po06026, po06027, po06028, po06029, po06030, po06031, po06032, po06033, po06034, po06035, po06036, po06037, po06038, po06039, po06040, po06041, po06042, po06043, po06044, po06045, po06046, po06047, po06048, po06049, po06050, po06051, po06052, po06053, po06054, po06055, po06056, po06057, po06058, po06059, po06060, po06061, po06062, po06063, po06064, po06065, po06066, po06067, po06068, po06069, po06070, po06071, po06072, po06073, po06074, po06075, po06076, po06077, po06078, po06079, po06080, po06081, po06082, po06083, po06084, po06085, po06086, po06087, po06088, po06089, po06090, po06091, po06092, po06093, po06094, po06095, po06096, po06097, po06098, po06099, po06100, po06101, po06102, po06103, po06104, po06105, po06106, po06107, po06108, po06109, po06110, po06111, po06112, po06113, po06114, po06115, po06116, po06117, po06118, po06119, po06120, po06121, po06122, po06123, po06124, po06125, po06126, po06127, po06128, po06129, po06130, po06131, po06132, po06133, po06134, po06135, po06136, po06137, po06138, po06139, po06140, po06141, po06142, po06143, po06144, po06145, po06146, po06147, po06148, po06149, po06150, po06151, po06152, po06153, po06154, po06155, po06156, po06157, po06158, po06159, po06160, po06161, po06162, po06163, po06164, po06165, po06166, po06167, po06168, po06169, po06170, po06171, po06172, po06173, po06174, po06175, po06176, po06177, po06178, po06179, po06180, po06181, po06182, po06183, po06184, po06185, po06186, po06187, po06188, po06189, po06190, po06191, po06192, po06193, po06194, po06195, po06196, po06197, po06198, po06199, po06200, po06201, po06202, po06203, po06204, po06205, po06206, po06207, po06208, po06209, po06210, po06211, po06212, po06213, po06214, po06215, po06216, po06217, po06218, po06219, po06220, po06221, po06222, po06223, po06224, po06225, po06226, po06227, po06228, po06229, po06230, po06231, po06232, po06233, po06234, po06235, po06236, po06237, po06238, po06239, po06240, po06241, po06242, po06243, po06244, po06245, po06246, po06247, po06248, po06249, po06250, po06251, po06252, po06253, po06254, po06255, po06256, po06257, po06258, po06259, po06260, po06261, po06262, po06263, po06264, po06265, po06266, po06267, po06268, po06269, po06270, po06271, po06272, po06273, po06274, po06275, po06276, po06277, po06278, po06279, po06280, po06281, po06282, po06283, po06284, po06285, po06286, po06287, po06288, po06289, po06290, po06291, po06292, po06293, po06294, po06295, po06296, po06297, po06298, po06299, po06300, po06301, po06302, po06303, po06304, po06305, po06306, po06307, po06308, po06309, po06310, po06311, po06312, po06313, po06314, po06315, po06316, po06317, po06318, po06319, po06320, po06321, po06322, po06323, po06324, po06325, po06326, po06327, po06328, po06329, po06330, po06331, po06332, po06333, po06334, po06335, po06336, po06337, po06338, po06339, po06340, po06341, po06342, po06343, po06344, po06345, po06346, po06347, po06348, po06349, po06350, po06351, po06352, po06353, po06354, po06355, po06356, po06357, po06358, po06359, po06360, po06361, po06362, po06363, po06364, po06365, po06366, po06367, po06368, po06369, po06370, po06371, po06372, po06373, po06374, po06375, po06376, po06377, po06378, po06379, po06380, po06381, po06382, po06383, po06384, po06385, po06386, po06387, po06388, po06389, po06390, po06391, po06392, po06393, po06394, po06395, po06396, po06397, po06398, po06399, po06400, po06401, po06402, po06403, po06404, po06405, po06406, po06407, po06408, po06409, po06410, po06411, po06412, po06413, po06414, po06415, po06416, po06417, po06418, po06419, po06420, po06421, po06422, po06423, po06424, po06425, po06426, po06427, po06428, po06429, po06430, po06431, po06432, po06433, po06434, po06435, po06436, po06437, po06438, po06439, po06440, po06441, po06442, po06443, po06444, po06445, po06446, po06447, po06448, po06449, po06450, po06451, po06452, po06453, po06454, po06455, po06456, po06457, po06458, po06459, po06460, po06461, po06462, po06463, po06464, po06465, po06466, po06467, po06468, po06469, po06470, po06471, po06472, po06473, po06474, po06475, po06476, po06477, po06478, po06479, po06480, po06481, po06482, po06483, po06484, po06485, po06486, po06487, po06488, po06489, po06490, po06491, po06492, po06493, po06494, po06495, po06496, po06497, po06498, po06499, po06500, po06501, po06502, po06503, po06504, po06505, po06506, po06507, po06508, po06509, po06510, po06511, po06512, po06513, po06514, po06515, po06516, po06517, po06518, po06519, po06520, po06521, po06522, po06523, po06524, po06525, po06526, po06527, po06528, po06529, po06530, po06531, po06532, po06533, po06534, po06535, po06536, po06537, po06538, po06539, po06540, po06541, po06542, po06543, po06544, po06545, po06546, po06547, po06548, po06549, po06550, po06551, po06552, po06553, po06554, po06555, po06556, po06557, po06558, po06559, po06560, po06561, po06562, po06563, po06564, po06565, po06566, po06567, po06568, po06569, po06570, po06571, po06572, po06573, po06574, po06575, po06576, po06577, po06578, po06579, po06580, po06581, po06582, po06583, po06584, po06585, po06586, po06587, po06588, po06589, po06590, po06591, po06592, po06593, po06594, po06595, po06596, po06597, po06598, po06599, po06600, po06601, po06602, po06603, po06604, po06605, po06606, po06607, po06608, po06609, po06610, po06611, po06612, po06613, po06614, po06615, po06616, po06617, po06618, po06619, po06620, po06621, po06622, po06623, po06624, po06625, po06626, po06627, po06628, po06629, po06630, po06631, po06632, po06633, po06634, po06635, po06636, po06637, po06638, po06639, po06640, po06641, po06642, po06643, po06644, po06645, po06646, po06647, po06648, po06649, po06650, po06651, po06652, po06653, po06654, po06655, po06656, po06657, po06658, po06659, po06660, po06661, po06662, po06663, po06664, po06665, po06666, po06667, po06668, po06669, po06670, po06671, po06672, po06673, po06674, po06675, po06676, po06677, po06678, po06679, po06680, po06681, po06682, po06683, po06684, po06685, po06686, po06687, po06688, po06689, po06690, po06691, po06692, po06693, po06694, po06695, po06696, po06697, po06698, po06699, po06700, po06701, po06702, po06703, po06704, po06705, po06706, po06707, po06708, po06709, po06710, po06711, po06712, po06713, po06714, po06715, po06716, po06717, po06718, po06719, po06720, po06721, po06722, po06723, po06724, po06725, po06726, po06727, po06728, po06729, po06730, po06731, po06732, po06733, po06734, po06735, po06736, po06737, po06738, po06739, po06740, po06741, po06742, po06743, po06744, po06745, po06746, po06747, po06748, po06749, po06750, po06751, po06752, po06753, po06754, po06755, po06756, po06757, po06758, po06759, po06760, po06761, po06762, po06763, po06764, po06765, po06766, po06767, po06768, po06769, po06770, po06771, po06772, po06773, po06774, po06775, po06776, po06777, po06778, po06779, po06780, po06781, po06782, po06783, po06784, po06785, po06786, po06787, po06788, po06789, po06790, po06791, po06792, po06793, po06794, po06795, po06796, po06797, po06798, po06799, po06800, po06801, po06802, po06803, po06804, po06805, po06806, po06807, po06808, po06809, po06810, po06811, po06812, po06813, po06814, po06815, po06816, po06817, po06818, po06819, po06820, po06821, po06822, po06823, po06824, po06825, po06826, po06827, po06828, po06829, po06830, po06831, po06832, po06833, po06834, po06835, po06836, po06837, po06838, po06839, po06840, po06841, po06842, po06843, po06844, po06845, po06846, po06847, po06848, po06849, po06850, po06851, po06852, po06853, po06854, po06855, po06856, po06857, po06858, po06859, po06860, po06861, po06862, po06863, po06864, po06865, po06866, po06867, po06868, po06869, po06870, po06871, po06872, po06873, po06874, po06875, po06876, po06877, po06878, po06879, po06880, po06881, po06882, po06883, po06884, po06885, po06886, po06887, po06888, po06889, po06890, po06891, po06892, po06893, po06894, po06895, po06896, po06897, po06898, po06899, po06900, po06901, po06902, po06903, po06904, po06905, po06906, po06907, po06908, po06909, po06910, po06911, po06912, po06913, po06914, po06915, po06916, po06917, po06918, po06919, po06920, po06921, po06922, po06923, po06924, po06925, po06926, po06927, po06928, po06929, po06930, po06931, po06932, po06933, po06934, po06935, po06936, po06937, po06938, po06939, po06940, po06941, po06942, po06943, po06944, po06945, po06946, po06947, po06948, po06949, po06950, po06951, po06952, po06953, po06954, po06955, po06956, po06957, po06958, po06959, po06960, po06961, po06962, po06963, po06964, po06965, po06966, po06967, po06968, po06969, po06970, po06971, po06972, po06973, po06974, po06975, po06976, po06977, po06978, po06979, po06980, po06981, po06982, po06983, po06984, po06985, po06986, po06987, po06988, po06989, po06990, po06991, po06992, po06993, po06994, po06995, po06996, po06997, po06998, po06999, po07000, po07001, po07002, po07003, po07004, po07005, po07006, po07007, po07008, po07009, po07010, po07011, po07012, po07013, po07014, po07015, po07016, po07017, po07018, po07019, po07020, po07021, po07022, po07023, po07024, po07025, po07026, po07027, po07028, po07029, po07030, po07031, po07032, po07033, po07034, po07035, po07036, po07037, po07038, po07039, po07040, po07041, po07042, po07043, po07044, po07045, po07046, po07047, po07048, po07049, po07050, po07051, po07052, po07053, po07054, po07055, po07056, po07057, po07058, po07059, po07060, po07061, po07062, po07063, po07064, po07065, po07066, po07067, po07068, po07069, po07070, po07071, po07072, po07073, po07074, po07075, po07076, po07077, po07078, po07079, po07080, po07081, po07082, po07083, po07084, po07085, po07086, po07087, po07088, po07089, po07090, po07091, po07092, po07093, po07094, po07095, po07096, po07097, po07098, po07099, po07100, po07101, po07102, po07103, po07104, po07105, po07106, po07107, po07108, po07109, po07110, po07111, po07112, po07113, po07114, po07115, po07116, po07117, po07118, po07119, po07120, po07121, po07122, po07123, po07124, po07125, po07126, po07127, po07128, po07129, po07130, po07131, po07132, po07133, po07134, po07135, po07136, po07137, po07138, po07139, po07140, po07141, po07142, po07143, po07144, po07145, po07146, po07147, po07148, po07149, po07150, po07151, po07152, po07153, po07154, po07155, po07156, po07157, po07158, po07159, po07160, po07161, po07162, po07163, po07164, po07165, po07166, po07167, po07168, po07169, po07170, po07171, po07172, po07173, po07174, po07175, po07176, po07177, po07178, po07179, po07180, po07181, po07182, po07183, po07184, po07185, po07186, po07187, po07188, po07189, po07190, po07191, po07192, po07193, po07194, po07195, po07196, po07197, po07198, po07199, po07200, po07201, po07202, po07203, po07204, po07205, po07206, po07207, po07208, po07209, po07210, po07211, po07212, po07213, po07214, po07215, po07216, po07217, po07218, po07219, po07220, po07221, po07222, po07223, po07224, po07225, po07226, po07227, po07228, po07229, po07230, po07231, po07232, po07233, po07234, po07235, po07236, po07237, po07238, po07239, po07240, po07241, po07242, po07243, po07244, po07245, po07246, po07247, po07248, po07249, po07250, po07251, po07252, po07253, po07254, po07255, po07256, po07257, po07258, po07259, po07260, po07261, po07262, po07263, po07264, po07265, po07266, po07267, po07268, po07269, po07270, po07271, po07272, po07273, po07274, po07275, po07276, po07277, po07278, po07279, po07280, po07281, po07282, po07283, po07284, po07285, po07286, po07287, po07288, po07289, po07290, po07291, po07292, po07293, po07294, po07295, po07296, po07297, po07298, po07299, po07300, po07301, po07302, po07303, po07304, po07305, po07306, po07307, po07308, po07309, po07310, po07311, po07312, po07313, po07314, po07315, po07316, po07317, po07318, po07319, po07320, po07321, po07322, po07323, po07324, po07325, po07326, po07327, po07328, po07329, po07330, po07331, po07332, po07333, po07334, po07335, po07336, po07337, po07338, po07339, po07340, po07341, po07342, po07343, po07344, po07345, po07346, po07347, po07348, po07349, po07350, po07351, po07352, po07353, po07354, po07355, po07356, po07357, po07358, po07359, po07360, po07361, po07362, po07363, po07364, po07365, po07366, po07367, po07368, po07369, po07370, po07371, po07372, po07373, po07374, po07375, po07376, po07377, po07378, po07379, po07380, po07381, po07382, po07383, po07384, po07385, po07386, po07387, po07388, po07389, po07390, po07391, po07392, po07393, po07394, po07395, po07396, po07397, po07398, po07399, po07400, po07401, po07402, po07403, po07404, po07405, po07406, po07407, po07408, po07409, po07410, po07411, po07412, po07413, po07414, po07415, po07416, po07417, po07418, po07419, po07420, po07421, po07422, po07423, po07424, po07425, po07426, po07427, po07428, po07429, po07430, po07431, po07432, po07433, po07434, po07435, po07436, po07437, po07438, po07439, po07440, po07441, po07442, po07443, po07444, po07445, po07446, po07447, po07448, po07449, po07450, po07451, po07452, po07453, po07454, po07455, po07456, po07457, po07458, po07459, po07460, po07461, po07462, po07463, po07464, po07465, po07466, po07467, po07468, po07469, po07470, po07471, po07472, po07473, po07474, po07475, po07476, po07477, po07478, po07479, po07480, po07481, po07482, po07483, po07484, po07485, po07486, po07487, po07488, po07489, po07490, po07491, po07492, po07493, po07494, po07495, po07496, po07497, po07498, po07499, po07500, po07501, po07502, po07503, po07504, po07505, po07506, po07507, po07508, po07509, po07510, po07511, po07512, po07513, po07514, po07515, po07516, po07517, po07518, po07519, po07520, po07521, po07522, po07523, po07524, po07525, po07526, po07527, po07528, po07529, po07530, po07531, po07532, po07533, po07534, po07535, po07536, po07537, po07538, po07539, po07540, po07541, po07542, po07543, po07544, po07545, po07546, po07547, po07548, po07549, po07550, po07551, po07552, po07553, po07554, po07555, po07556, po07557, po07558, po07559, po07560, po07561, po07562, po07563, po07564, po07565, po07566, po07567, po07568, po07569, po07570, po07571, po07572, po07573, po07574, po07575, po07576, po07577, po07578, po07579, po07580, po07581, po07582, po07583, po07584, po07585, po07586, po07587, po07588, po07589, po07590, po07591, po07592, po07593, po07594, po07595, po07596, po07597, po07598, po07599, po07600, po07601, po07602, po07603, po07604, po07605, po07606, po07607, po07608, po07609, po07610, po07611, po07612, po07613, po07614, po07615, po07616, po07617, po07618, po07619, po07620, po07621, po07622, po07623, po07624, po07625, po07626, po07627, po07628, po07629, po07630, po07631, po07632, po07633, po07634, po07635, po07636, po07637, po07638, po07639, po07640, po07641, po07642, po07643, po07644, po07645, po07646, po07647, po07648, po07649, po07650, po07651, po07652, po07653, po07654, po07655, po07656, po07657, po07658, po07659, po07660, po07661, po07662, po07663, po07664, po07665, po07666, po07667, po07668, po07669, po07670, po07671, po07672, po07673, po07674, po07675, po07676, po07677, po07678, po07679, po07680, po07681, po07682, po07683, po07684, po07685, po07686, po07687, po07688, po07689, po07690, po07691, po07692, po07693, po07694, po07695, po07696, po07697, po07698, po07699, po07700, po07701, po07702, po07703, po07704, po07705, po07706, po07707, po07708, po07709, po07710, po07711, po07712, po07713, po07714, po07715, po07716, po07717, po07718, po07719, po07720, po07721, po07722, po07723, po07724, po07725, po07726, po07727, po07728, po07729, po07730, po07731, po07732, po07733, po07734, po07735, po07736, po07737, po07738, po07739, po07740, po07741, po07742, po07743, po07744, po07745, po07746, po07747, po07748, po07749, po07750, po07751, po07752, po07753, po07754, po07755, po07756, po07757, po07758, po07759, po07760, po07761, po07762, po07763, po07764, po07765, po07766, po07767, po07768, po07769, po07770, po07771, po07772, po07773, po07774, po07775, po07776, po07777, po07778, po07779, po07780, po07781, po07782, po07783, po07784, po07785, po07786, po07787, po07788, po07789, po07790, po07791, po07792, po07793, po07794, po07795, po07796, po07797, po07798, po07799, po07800, po07801, po07802, po07803, po07804, po07805, po07806, po07807, po07808, po07809, po07810, po07811, po07812, po07813, po07814, po07815, po07816, po07817, po07818, po07819, po07820, po07821, po07822, po07823, po07824, po07825, po07826, po07827, po07828, po07829, po07830, po07831, po07832, po07833, po07834, po07835, po07836, po07837, po07838, po07839, po07840, po07841, po07842, po07843, po07844, po07845, po07846, po07847, po07848, po07849, po07850, po07851, po07852, po07853, po07854, po07855, po07856, po07857, po07858, po07859, po07860, po07861, po07862, po07863, po07864, po07865, po07866, po07867, po07868, po07869, po07870, po07871, po07872, po07873, po07874, po07875, po07876, po07877, po07878, po07879, po07880, po07881, po07882, po07883, po07884, po07885, po07886, po07887, po07888, po07889, po07890, po07891, po07892, po07893, po07894, po07895, po07896, po07897, po07898, po07899, po07900, po07901, po07902, po07903, po07904, po07905, po07906, po07907, po07908, po07909, po07910, po07911, po07912, po07913, po07914, po07915, po07916, po07917, po07918, po07919, po07920, po07921, po07922, po07923, po07924, po07925, po07926, po07927, po07928, po07929, po07930, po07931, po07932, po07933, po07934, po07935, po07936, po07937, po07938, po07939, po07940, po07941, po07942, po07943, po07944, po07945, po07946, po07947, po07948, po07949, po07950, po07951, po07952, po07953, po07954, po07955, po07956, po07957, po07958, po07959, po07960, po07961, po07962, po07963, po07964, po07965, po07966, po07967, po07968, po07969, po07970, po07971, po07972, po07973, po07974, po07975, po07976, po07977, po07978, po07979, po07980, po07981, po07982, po07983, po07984, po07985, po07986, po07987, po07988, po07989, po07990, po07991, po07992, po07993, po07994, po07995, po07996, po07997, po07998, po07999, po08000, po08001, po08002, po08003, po08004, po08005, po08006, po08007, po08008, po08009, po08010, po08011, po08012, po08013, po08014, po08015, po08016, po08017, po08018, po08019, po08020, po08021, po08022, po08023, po08024, po08025, po08026, po08027, po08028, po08029, po08030, po08031, po08032, po08033, po08034, po08035, po08036, po08037, po08038, po08039, po08040, po08041, po08042, po08043, po08044, po08045, po08046, po08047, po08048, po08049, po08050, po08051, po08052, po08053, po08054, po08055, po08056, po08057, po08058, po08059, po08060, po08061, po08062, po08063, po08064, po08065, po08066, po08067, po08068, po08069, po08070, po08071, po08072, po08073, po08074, po08075, po08076, po08077, po08078, po08079, po08080, po08081, po08082, po08083, po08084, po08085, po08086, po08087, po08088, po08089, po08090, po08091, po08092, po08093, po08094, po08095, po08096, po08097, po08098, po08099, po08100, po08101, po08102, po08103, po08104, po08105, po08106, po08107, po08108, po08109, po08110, po08111, po08112, po08113, po08114, po08115, po08116, po08117, po08118, po08119, po08120, po08121, po08122, po08123, po08124, po08125, po08126, po08127, po08128, po08129, po08130, po08131, po08132, po08133, po08134, po08135, po08136, po08137, po08138, po08139, po08140, po08141, po08142, po08143, po08144, po08145, po08146, po08147, po08148, po08149, po08150, po08151, po08152, po08153, po08154, po08155, po08156, po08157, po08158, po08159, po08160, po08161, po08162, po08163, po08164, po08165, po08166, po08167, po08168, po08169, po08170, po08171, po08172, po08173, po08174, po08175, po08176, po08177, po08178, po08179, po08180, po08181, po08182, po08183, po08184, po08185, po08186, po08187, po08188, po08189, po08190, po08191, po08192, po08193, po08194, po08195, po08196, po08197, po08198, po08199, po08200, po08201, po08202, po08203, po08204, po08205, po08206, po08207, po08208, po08209, po08210, po08211, po08212, po08213, po08214, po08215, po08216, po08217, po08218, po08219, po08220, po08221, po08222, po08223, po08224, po08225, po08226, po08227, po08228, po08229, po08230, po08231, po08232, po08233, po08234, po08235, po08236, po08237, po08238, po08239, po08240, po08241, po08242, po08243, po08244, po08245, po08246, po08247, po08248, po08249, po08250, po08251, po08252, po08253, po08254, po08255, po08256, po08257, po08258, po08259, po08260, po08261, po08262, po08263, po08264, po08265, po08266, po08267, po08268, po08269, po08270, po08271, po08272, po08273, po08274, po08275, po08276, po08277, po08278, po08279, po08280, po08281, po08282, po08283, po08284, po08285, po08286, po08287, po08288, po08289, po08290, po08291, po08292, po08293, po08294, po08295, po08296, po08297, po08298, po08299, po08300, po08301, po08302, po08303, po08304, po08305, po08306, po08307, po08308, po08309, po08310, po08311, po08312, po08313, po08314, po08315, po08316, po08317, po08318, po08319, po08320, po08321, po08322, po08323, po08324, po08325, po08326, po08327, po08328, po08329, po08330, po08331, po08332, po08333, po08334, po08335, po08336, po08337, po08338, po08339, po08340, po08341, po08342, po08343, po08344, po08345, po08346, po08347, po08348, po08349, po08350, po08351, po08352, po08353, po08354, po08355, po08356, po08357, po08358, po08359, po08360, po08361, po08362, po08363, po08364, po08365, po08366, po08367, po08368, po08369, po08370, po08371, po08372, po08373, po08374, po08375, po08376, po08377, po08378, po08379, po08380, po08381, po08382, po08383, po08384, po08385, po08386, po08387, po08388, po08389, po08390, po08391, po08392, po08393, po08394, po08395, po08396, po08397, po08398, po08399, po08400, po08401, po08402, po08403, po08404, po08405, po08406, po08407, po08408, po08409, po08410, po08411, po08412, po08413, po08414, po08415, po08416, po08417, po08418, po08419, po08420, po08421, po08422, po08423, po08424, po08425, po08426, po08427, po08428, po08429, po08430, po08431, po08432, po08433, po08434, po08435, po08436, po08437, po08438, po08439, po08440, po08441, po08442, po08443, po08444, po08445, po08446, po08447, po08448, po08449, po08450, po08451, po08452, po08453, po08454, po08455, po08456, po08457, po08458, po08459, po08460, po08461, po08462, po08463, po08464, po08465, po08466, po08467, po08468, po08469, po08470, po08471, po08472, po08473, po08474, po08475, po08476, po08477, po08478, po08479, po08480, po08481, po08482, po08483, po08484, po08485, po08486, po08487, po08488, po08489, po08490, po08491, po08492, po08493, po08494, po08495, po08496, po08497, po08498, po08499, po08500, po08501, po08502, po08503, po08504, po08505, po08506, po08507, po08508, po08509, po08510, po08511, po08512, po08513, po08514, po08515, po08516, po08517, po08518, po08519, po08520, po08521, po08522, po08523, po08524, po08525, po08526, po08527, po08528, po08529, po08530, po08531, po08532, po08533, po08534, po08535, po08536, po08537, po08538, po08539, po08540, po08541, po08542, po08543, po08544, po08545, po08546, po08547, po08548, po08549, po08550, po08551, po08552, po08553, po08554, po08555, po08556, po08557, po08558, po08559, po08560, po08561, po08562, po08563, po08564, po08565, po08566, po08567, po08568, po08569, po08570, po08571, po08572, po08573, po08574, po08575, po08576, po08577, po08578, po08579, po08580, po08581, po08582, po08583, po08584, po08585, po08586, po08587, po08588, po08589, po08590, po08591, po08592, po08593, po08594, po08595, po08596, po08597, po08598, po08599, po08600, po08601, po08602, po08603, po08604, po08605, po08606, po08607, po08608, po08609, po08610, po08611, po08612, po08613, po08614, po08615, po08616, po08617, po08618, po08619, po08620, po08621, po08622, po08623, po08624, po08625, po08626, po08627, po08628, po08629, po08630, po08631, po08632, po08633, po08634, po08635, po08636, po08637, po08638, po08639, po08640, po08641, po08642, po08643, po08644, po08645, po08646, po08647, po08648, po08649, po08650, po08651, po08652, po08653, po08654, po08655, po08656, po08657, po08658, po08659, po08660, po08661, po08662, po08663, po08664, po08665, po08666, po08667, po08668, po08669, po08670, po08671, po08672, po08673, po08674, po08675, po08676, po08677, po08678, po08679, po08680, po08681, po08682, po08683, po08684, po08685, po08686, po08687, po08688, po08689, po08690, po08691, po08692, po08693, po08694, po08695, po08696, po08697, po08698, po08699, po08700, po08701, po08702, po08703, po08704, po08705, po08706, po08707, po08708, po08709, po08710, po08711, po08712, po08713, po08714, po08715, po08716, po08717, po08718, po08719, po08720, po08721, po08722, po08723, po08724, po08725, po08726, po08727, po08728, po08729, po08730, po08731, po08732, po08733, po08734, po08735, po08736, po08737, po08738, po08739, po08740, po08741, po08742, po08743, po08744, po08745, po08746, po08747, po08748, po08749, po08750, po08751, po08752, po08753, po08754, po08755, po08756, po08757, po08758, po08759, po08760, po08761, po08762, po08763, po08764, po08765, po08766, po08767, po08768, po08769, po08770, po08771, po08772, po08773, po08774, po08775, po08776, po08777, po08778, po08779, po08780, po08781, po08782, po08783, po08784, po08785, po08786, po08787, po08788, po08789, po08790, po08791, po08792, po08793, po08794, po08795, po08796, po08797, po08798, po08799, po08800, po08801, po08802, po08803, po08804, po08805, po08806, po08807, po08808, po08809, po08810, po08811, po08812, po08813, po08814, po08815, po08816, po08817, po08818, po08819, po08820, po08821, po08822, po08823, po08824, po08825, po08826, po08827, po08828, po08829, po08830, po08831, po08832, po08833, po08834, po08835, po08836, po08837, po08838, po08839, po08840, po08841, po08842, po08843, po08844, po08845, po08846, po08847, po08848, po08849, po08850, po08851, po08852, po08853, po08854, po08855, po08856, po08857, po08858, po08859, po08860, po08861, po08862, po08863, po08864, po08865, po08866, po08867, po08868, po08869, po08870, po08871, po08872, po08873, po08874, po08875, po08876, po08877, po08878, po08879, po08880, po08881, po08882, po08883, po08884, po08885, po08886, po08887, po08888, po08889, po08890, po08891, po08892, po08893, po08894, po08895, po08896, po08897, po08898, po08899, po08900, po08901, po08902, po08903, po08904, po08905, po08906, po08907, po08908, po08909, po08910, po08911, po08912, po08913, po08914, po08915, po08916, po08917, po08918, po08919, po08920, po08921, po08922, po08923, po08924, po08925, po08926, po08927, po08928, po08929, po08930, po08931, po08932, po08933, po08934, po08935, po08936, po08937, po08938, po08939, po08940, po08941, po08942, po08943, po08944, po08945, po08946, po08947, po08948, po08949, po08950, po08951, po08952, po08953, po08954, po08955, po08956, po08957, po08958, po08959, po08960, po08961, po08962, po08963, po08964, po08965, po08966, po08967, po08968, po08969, po08970, po08971, po08972, po08973, po08974, po08975, po08976, po08977, po08978, po08979, po08980, po08981, po08982, po08983, po08984, po08985, po08986, po08987, po08988, po08989, po08990, po08991, po08992, po08993, po08994, po08995, po08996, po08997, po08998, po08999, po09000, po09001, po09002, po09003, po09004, po09005, po09006, po09007, po09008, po09009, po09010, po09011, po09012, po09013, po09014, po09015, po09016, po09017, po09018, po09019, po09020, po09021, po09022, po09023, po09024, po09025, po09026, po09027, po09028, po09029, po09030, po09031, po09032, po09033, po09034, po09035, po09036, po09037, po09038, po09039, po09040, po09041, po09042, po09043, po09044, po09045, po09046, po09047, po09048, po09049, po09050, po09051, po09052, po09053, po09054, po09055, po09056, po09057, po09058, po09059, po09060, po09061, po09062, po09063, po09064, po09065, po09066, po09067, po09068, po09069, po09070, po09071, po09072, po09073, po09074, po09075, po09076, po09077, po09078, po09079, po09080, po09081, po09082, po09083, po09084, po09085, po09086, po09087, po09088, po09089, po09090, po09091, po09092, po09093, po09094, po09095, po09096, po09097, po09098, po09099, po09100, po09101, po09102, po09103, po09104, po09105, po09106, po09107, po09108, po09109, po09110, po09111, po09112, po09113, po09114, po09115, po09116, po09117, po09118, po09119, po09120, po09121, po09122, po09123, po09124, po09125, po09126, po09127, po09128, po09129, po09130, po09131, po09132, po09133, po09134, po09135, po09136, po09137, po09138, po09139, po09140, po09141, po09142, po09143, po09144, po09145, po09146, po09147, po09148, po09149, po09150, po09151, po09152, po09153, po09154, po09155, po09156, po09157, po09158, po09159, po09160, po09161, po09162, po09163, po09164, po09165, po09166, po09167, po09168, po09169, po09170, po09171, po09172, po09173, po09174, po09175, po09176, po09177, po09178, po09179, po09180, po09181, po09182, po09183, po09184, po09185, po09186, po09187, po09188, po09189, po09190, po09191, po09192, po09193, po09194, po09195, po09196, po09197, po09198, po09199, po09200, po09201, po09202, po09203, po09204, po09205, po09206, po09207, po09208, po09209, po09210, po09211, po09212, po09213, po09214, po09215, po09216, po09217, po09218, po09219, po09220, po09221, po09222, po09223, po09224, po09225, po09226, po09227, po09228, po09229, po09230, po09231, po09232, po09233, po09234, po09235, po09236, po09237, po09238, po09239, po09240, po09241, po09242, po09243, po09244, po09245, po09246, po09247, po09248, po09249, po09250, po09251, po09252, po09253, po09254, po09255, po09256, po09257, po09258, po09259, po09260, po09261, po09262, po09263, po09264, po09265, po09266, po09267, po09268, po09269, po09270, po09271, po09272, po09273, po09274, po09275, po09276, po09277, po09278, po09279, po09280, po09281, po09282, po09283, po09284, po09285, po09286, po09287, po09288, po09289, po09290, po09291, po09292, po09293, po09294, po09295, po09296, po09297, po09298, po09299, po09300, po09301, po09302, po09303, po09304, po09305, po09306, po09307, po09308, po09309, po09310, po09311, po09312, po09313, po09314, po09315, po09316, po09317, po09318, po09319, po09320, po09321, po09322, po09323, po09324, po09325, po09326, po09327, po09328, po09329, po09330, po09331, po09332, po09333, po09334, po09335, po09336, po09337, po09338, po09339, po09340, po09341, po09342, po09343, po09344, po09345, po09346, po09347, po09348, po09349, po09350, po09351, po09352, po09353, po09354, po09355, po09356, po09357, po09358, po09359, po09360, po09361, po09362, po09363, po09364, po09365, po09366, po09367, po09368, po09369, po09370, po09371, po09372, po09373, po09374, po09375, po09376, po09377, po09378, po09379, po09380, po09381, po09382, po09383, po09384, po09385, po09386, po09387, po09388, po09389, po09390, po09391, po09392, po09393, po09394, po09395, po09396, po09397, po09398, po09399, po09400, po09401, po09402, po09403, po09404, po09405, po09406, po09407, po09408, po09409, po09410, po09411, po09412, po09413, po09414, po09415, po09416, po09417, po09418, po09419, po09420, po09421, po09422, po09423, po09424, po09425, po09426, po09427, po09428, po09429, po09430, po09431, po09432, po09433, po09434, po09435, po09436, po09437, po09438, po09439, po09440, po09441, po09442, po09443, po09444, po09445, po09446, po09447, po09448, po09449, po09450, po09451, po09452, po09453, po09454, po09455, po09456, po09457, po09458, po09459, po09460, po09461, po09462, po09463, po09464, po09465, po09466, po09467, po09468, po09469, po09470, po09471, po09472, po09473, po09474, po09475, po09476, po09477, po09478, po09479, po09480, po09481, po09482, po09483, po09484, po09485, po09486, po09487, po09488, po09489, po09490, po09491, po09492, po09493, po09494, po09495, po09496, po09497, po09498, po09499, po09500, po09501, po09502, po09503, po09504, po09505, po09506, po09507, po09508, po09509, po09510, po09511, po09512, po09513, po09514, po09515, po09516, po09517, po09518, po09519, po09520, po09521, po09522, po09523, po09524, po09525, po09526, po09527, po09528, po09529, po09530, po09531, po09532, po09533, po09534, po09535, po09536, po09537, po09538, po09539, po09540, po09541, po09542, po09543, po09544, po09545, po09546, po09547, po09548, po09549, po09550, po09551, po09552, po09553, po09554, po09555, po09556, po09557, po09558, po09559, po09560, po09561, po09562, po09563, po09564, po09565, po09566, po09567, po09568, po09569, po09570, po09571, po09572, po09573, po09574, po09575, po09576, po09577, po09578, po09579, po09580, po09581, po09582, po09583, po09584, po09585, po09586, po09587, po09588, po09589, po09590, po09591, po09592, po09593, po09594, po09595, po09596, po09597, po09598, po09599, po09600, po09601, po09602, po09603, po09604, po09605, po09606, po09607, po09608, po09609, po09610, po09611, po09612, po09613, po09614, po09615, po09616, po09617, po09618, po09619, po09620, po09621, po09622, po09623, po09624, po09625, po09626, po09627, po09628, po09629, po09630, po09631, po09632, po09633, po09634, po09635, po09636, po09637, po09638, po09639, po09640, po09641, po09642, po09643, po09644, po09645, po09646, po09647, po09648, po09649, po09650, po09651, po09652, po09653, po09654, po09655, po09656, po09657, po09658, po09659, po09660, po09661, po09662, po09663, po09664, po09665, po09666, po09667, po09668, po09669, po09670, po09671, po09672, po09673, po09674, po09675, po09676, po09677, po09678, po09679, po09680, po09681, po09682, po09683, po09684, po09685, po09686, po09687, po09688, po09689, po09690, po09691, po09692, po09693, po09694, po09695, po09696, po09697, po09698, po09699, po09700, po09701, po09702, po09703, po09704, po09705, po09706, po09707, po09708, po09709, po09710, po09711, po09712, po09713, po09714, po09715, po09716, po09717, po09718, po09719, po09720, po09721, po09722, po09723, po09724, po09725, po09726, po09727, po09728, po09729, po09730, po09731, po09732, po09733, po09734, po09735, po09736, po09737, po09738, po09739, po09740, po09741, po09742, po09743, po09744, po09745, po09746, po09747, po09748, po09749, po09750, po09751, po09752, po09753, po09754, po09755, po09756, po09757, po09758, po09759, po09760, po09761, po09762, po09763, po09764, po09765, po09766, po09767, po09768, po09769, po09770, po09771, po09772, po09773, po09774, po09775, po09776, po09777, po09778, po09779, po09780, po09781, po09782, po09783, po09784, po09785, po09786, po09787, po09788, po09789, po09790, po09791, po09792, po09793, po09794, po09795, po09796, po09797, po09798, po09799, po09800, po09801, po09802, po09803, po09804, po09805, po09806, po09807, po09808, po09809, po09810, po09811, po09812, po09813, po09814, po09815, po09816, po09817, po09818, po09819, po09820, po09821, po09822, po09823, po09824, po09825, po09826, po09827, po09828, po09829, po09830, po09831, po09832, po09833, po09834, po09835, po09836, po09837, po09838, po09839, po09840, po09841, po09842, po09843, po09844, po09845, po09846, po09847, po09848, po09849, po09850, po09851, po09852, po09853, po09854, po09855, po09856, po09857, po09858, po09859, po09860, po09861, po09862, po09863, po09864, po09865, po09866, po09867, po09868, po09869, po09870, po09871, po09872, po09873, po09874, po09875, po09876, po09877, po09878, po09879, po09880, po09881, po09882, po09883, po09884, po09885, po09886, po09887, po09888, po09889, po09890, po09891, po09892, po09893, po09894, po09895, po09896, po09897, po09898, po09899, po09900, po09901, po09902, po09903, po09904, po09905, po09906, po09907, po09908, po09909, po09910, po09911, po09912, po09913, po09914, po09915, po09916, po09917, po09918, po09919, po09920, po09921, po09922, po09923, po09924, po09925, po09926, po09927, po09928, po09929, po09930, po09931, po09932, po09933, po09934, po09935, po09936, po09937, po09938, po09939, po09940, po09941, po09942, po09943, po09944, po09945, po09946, po09947, po09948, po09949, po09950, po09951, po09952, po09953, po09954, po09955, po09956, po09957, po09958, po09959, po09960, po09961, po09962, po09963, po09964, po09965, po09966, po09967, po09968, po09969, po09970, po09971, po09972, po09973, po09974, po09975, po09976, po09977, po09978, po09979, po09980, po09981, po09982, po09983, po09984, po09985, po09986, po09987, po09988, po09989, po09990, po09991, po09992, po09993, po09994, po09995, po09996, po09997, po09998, po09999, po10000, po10001, po10002, po10003, po10004, po10005, po10006, po10007, po10008, po10009, po10010, po10011, po10012, po10013, po10014, po10015, po10016, po10017, po10018, po10019, po10020, po10021, po10022, po10023, po10024, po10025, po10026, po10027, po10028, po10029, po10030, po10031, po10032, po10033, po10034, po10035, po10036, po10037, po10038, po10039, po10040, po10041, po10042, po10043, po10044, po10045, po10046, po10047, po10048, po10049, po10050, po10051, po10052, po10053, po10054, po10055, po10056, po10057, po10058, po10059, po10060, po10061, po10062, po10063, po10064, po10065, po10066, po10067, po10068, po10069, po10070, po10071, po10072, po10073, po10074, po10075, po10076, po10077, po10078, po10079, po10080, po10081, po10082, po10083, po10084, po10085, po10086, po10087, po10088, po10089, po10090, po10091, po10092, po10093, po10094, po10095, po10096, po10097, po10098, po10099, po10100, po10101, po10102, po10103, po10104, po10105, po10106, po10107, po10108, po10109, po10110, po10111, po10112, po10113, po10114, po10115, po10116, po10117, po10118, po10119, po10120, po10121, po10122, po10123, po10124, po10125, po10126, po10127, po10128, po10129, po10130, po10131, po10132, po10133, po10134, po10135, po10136, po10137, po10138, po10139, po10140, po10141, po10142, po10143, po10144, po10145, po10146, po10147, po10148, po10149, po10150, po10151, po10152, po10153, po10154, po10155, po10156, po10157, po10158, po10159, po10160, po10161, po10162, po10163, po10164, po10165, po10166, po10167, po10168, po10169, po10170, po10171, po10172, po10173, po10174, po10175, po10176, po10177, po10178, po10179, po10180, po10181, po10182, po10183, po10184, po10185, po10186, po10187, po10188, po10189, po10190, po10191, po10192, po10193, po10194, po10195, po10196, po10197, po10198, po10199, po10200, po10201, po10202, po10203, po10204, po10205, po10206, po10207, po10208, po10209, po10210, po10211, po10212, po10213, po10214, po10215, po10216, po10217, po10218, po10219, po10220, po10221, po10222, po10223, po10224, po10225, po10226, po10227, po10228, po10229, po10230, po10231, po10232, po10233, po10234, po10235, po10236, po10237, po10238, po10239, po10240, po10241, po10242, po10243, po10244, po10245, po10246, po10247, po10248, po10249, po10250, po10251, po10252, po10253, po10254, po10255, po10256, po10257, po10258, po10259, po10260, po10261, po10262, po10263, po10264, po10265, po10266, po10267, po10268, po10269, po10270, po10271, po10272, po10273, po10274, po10275, po10276, po10277, po10278, po10279, po10280, po10281, po10282, po10283, po10284, po10285, po10286, po10287, po10288, po10289, po10290, po10291, po10292, po10293, po10294, po10295, po10296, po10297, po10298, po10299, po10300, po10301, po10302, po10303, po10304, po10305, po10306, po10307, po10308, po10309, po10310, po10311, po10312, po10313, po10314, po10315, po10316, po10317, po10318, po10319, po10320, po10321, po10322, po10323, po10324, po10325, po10326, po10327, po10328, po10329, po10330, po10331, po10332, po10333, po10334, po10335, po10336, po10337, po10338, po10339, po10340, po10341, po10342, po10343, po10344, po10345, po10346, po10347, po10348, po10349, po10350, po10351, po10352, po10353, po10354, po10355, po10356, po10357, po10358, po10359, po10360, po10361, po10362, po10363, po10364, po10365, po10366, po10367, po10368, po10369, po10370, po10371, po10372, po10373, po10374, po10375, po10376, po10377, po10378, po10379, po10380, po10381, po10382, po10383, po10384, po10385, po10386, po10387, po10388, po10389, po10390, po10391, po10392, po10393, po10394, po10395, po10396, po10397, po10398, po10399, po10400, po10401, po10402, po10403, po10404, po10405, po10406, po10407, po10408, po10409, po10410, po10411, po10412, po10413, po10414, po10415, po10416, po10417, po10418, po10419, po10420, po10421, po10422, po10423, po10424, po10425, po10426, po10427, po10428, po10429, po10430, po10431, po10432, po10433, po10434, po10435, po10436, po10437, po10438, po10439, po10440, po10441, po10442, po10443, po10444, po10445, po10446, po10447, po10448, po10449, po10450, po10451, po10452, po10453, po10454, po10455, po10456, po10457, po10458, po10459, po10460, po10461, po10462, po10463, po10464, po10465, po10466, po10467, po10468, po10469, po10470, po10471, po10472, po10473, po10474, po10475, po10476, po10477, po10478, po10479, po10480, po10481, po10482, po10483, po10484, po10485, po10486, po10487, po10488, po10489, po10490, po10491, po10492, po10493, po10494, po10495, po10496, po10497, po10498, po10499, po10500, po10501, po10502, po10503, po10504, po10505, po10506, po10507, po10508, po10509, po10510, po10511, po10512, po10513, po10514, po10515, po10516, po10517, po10518, po10519, po10520, po10521, po10522, po10523, po10524, po10525, po10526, po10527, po10528, po10529, po10530, po10531, po10532, po10533, po10534, po10535, po10536, po10537, po10538, po10539, po10540, po10541, po10542, po10543, po10544, po10545, po10546, po10547, po10548, po10549, po10550, po10551, po10552, po10553, po10554, po10555, po10556, po10557, po10558, po10559, po10560, po10561, po10562, po10563, po10564, po10565, po10566, po10567, po10568, po10569, po10570, po10571, po10572, po10573, po10574, po10575, po10576, po10577, po10578, po10579, po10580, po10581, po10582, po10583, po10584, po10585, po10586, po10587, po10588, po10589, po10590, po10591, po10592, po10593, po10594, po10595, po10596, po10597, po10598, po10599, po10600, po10601, po10602, po10603, po10604, po10605, po10606, po10607, po10608, po10609, po10610, po10611, po10612, po10613, po10614, po10615, po10616, po10617, po10618, po10619, po10620, po10621, po10622, po10623, po10624, po10625, po10626, po10627, po10628, po10629, po10630, po10631, po10632, po10633, po10634, po10635, po10636, po10637, po10638, po10639, po10640, po10641, po10642, po10643, po10644, po10645, po10646, po10647, po10648, po10649, po10650, po10651, po10652, po10653, po10654, po10655, po10656, po10657, po10658, po10659, po10660, po10661, po10662, po10663, po10664, po10665, po10666, po10667, po10668, po10669, po10670, po10671, po10672, po10673, po10674, po10675, po10676, po10677, po10678, po10679, po10680, po10681, po10682, po10683, po10684, po10685, po10686, po10687, po10688, po10689, po10690, po10691, po10692, po10693, po10694, po10695);
input pi00000, pi00001, pi00002, pi00003, pi00004, pi00005, pi00006, pi00007, pi00008, pi00009, pi00010, pi00011, pi00012, pi00013, pi00014, pi00015, pi00016, pi00017, pi00018, pi00019, pi00020, pi00021, pi00022, pi00023, pi00024, pi00025, pi00026, pi00027, pi00028, pi00029, pi00030, pi00031, pi00032, pi00033, pi00034, pi00035, pi00036, pi00037, pi00038, pi00039, pi00040, pi00041, pi00042, pi00043, pi00044, pi00045, pi00046, pi00047, pi00048, pi00049, pi00050, pi00051, pi00052, pi00053, pi00054, pi00055, pi00056, pi00057, pi00058, pi00059, pi00060, pi00061, pi00062, pi00063, pi00064, pi00065, pi00066, pi00067, pi00068, pi00069, pi00070, pi00071, pi00072, pi00073, pi00074, pi00075, pi00076, pi00077, pi00078, pi00079, pi00080, pi00081, pi00082, pi00083, pi00084, pi00085, pi00086, pi00087, pi00088, pi00089, pi00090, pi00091, pi00092, pi00093, pi00094, pi00095, pi00096, pi00097, pi00098, pi00099, pi00100, pi00101, pi00102, pi00103, pi00104, pi00105, pi00106, pi00107, pi00108, pi00109, pi00110, pi00111, pi00112, pi00113, pi00114, pi00115, pi00116, pi00117, pi00118, pi00119, pi00120, pi00121, pi00122, pi00123, pi00124, pi00125, pi00126, pi00127, pi00128, pi00129, pi00130, pi00131, pi00132, pi00133, pi00134, pi00135, pi00136, pi00137, pi00138, pi00139, pi00140, pi00141, pi00142, pi00143, pi00144, pi00145, pi00146, pi00147, pi00148, pi00149, pi00150, pi00151, pi00152, pi00153, pi00154, pi00155, pi00156, pi00157, pi00158, pi00159, pi00160, pi00161, pi00162, pi00163, pi00164, pi00165, pi00166, pi00167, pi00168, pi00169, pi00170, pi00171, pi00172, pi00173, pi00174, pi00175, pi00176, pi00177, pi00178, pi00179, pi00180, pi00181, pi00182, pi00183, pi00184, pi00185, pi00186, pi00187, pi00188, pi00189, pi00190, pi00191, pi00192, pi00193, pi00194, pi00195, pi00196, pi00197, pi00198, pi00199, pi00200, pi00201, pi00202, pi00203, pi00204, pi00205, pi00206, pi00207, pi00208, pi00209, pi00210, pi00211, pi00212, pi00213, pi00214, pi00215, pi00216, pi00217, pi00218, pi00219, pi00220, pi00221, pi00222, pi00223, pi00224, pi00225, pi00226, pi00227, pi00228, pi00229, pi00230, pi00231, pi00232, pi00233, pi00234, pi00235, pi00236, pi00237, pi00238, pi00239, pi00240, pi00241, pi00242, pi00243, pi00244, pi00245, pi00246, pi00247, pi00248, pi00249, pi00250, pi00251, pi00252, pi00253, pi00254, pi00255, pi00256, pi00257, pi00258, pi00259, pi00260, pi00261, pi00262, pi00263, pi00264, pi00265, pi00266, pi00267, pi00268, pi00269, pi00270, pi00271, pi00272, pi00273, pi00274, pi00275, pi00276, pi00277, pi00278, pi00279, pi00280, pi00281, pi00282, pi00283, pi00284, pi00285, pi00286, pi00287, pi00288, pi00289, pi00290, pi00291, pi00292, pi00293, pi00294, pi00295, pi00296, pi00297, pi00298, pi00299, pi00300, pi00301, pi00302, pi00303, pi00304, pi00305, pi00306, pi00307, pi00308, pi00309, pi00310, pi00311, pi00312, pi00313, pi00314, pi00315, pi00316, pi00317, pi00318, pi00319, pi00320, pi00321, pi00322, pi00323, pi00324, pi00325, pi00326, pi00327, pi00328, pi00329, pi00330, pi00331, pi00332, pi00333, pi00334, pi00335, pi00336, pi00337, pi00338, pi00339, pi00340, pi00341, pi00342, pi00343, pi00344, pi00345, pi00346, pi00347, pi00348, pi00349, pi00350, pi00351, pi00352, pi00353, pi00354, pi00355, pi00356, pi00357, pi00358, pi00359, pi00360, pi00361, pi00362, pi00363, pi00364, pi00365, pi00366, pi00367, pi00368, pi00369, pi00370, pi00371, pi00372, pi00373, pi00374, pi00375, pi00376, pi00377, pi00378, pi00379, pi00380, pi00381, pi00382, pi00383, pi00384, pi00385, pi00386, pi00387, pi00388, pi00389, pi00390, pi00391, pi00392, pi00393, pi00394, pi00395, pi00396, pi00397, pi00398, pi00399, pi00400, pi00401, pi00402, pi00403, pi00404, pi00405, pi00406, pi00407, pi00408, pi00409, pi00410, pi00411, pi00412, pi00413, pi00414, pi00415, pi00416, pi00417, pi00418, pi00419, pi00420, pi00421, pi00422, pi00423, pi00424, pi00425, pi00426, pi00427, pi00428, pi00429, pi00430, pi00431, pi00432, pi00433, pi00434, pi00435, pi00436, pi00437, pi00438, pi00439, pi00440, pi00441, pi00442, pi00443, pi00444, pi00445, pi00446, pi00447, pi00448, pi00449, pi00450, pi00451, pi00452, pi00453, pi00454, pi00455, pi00456, pi00457, pi00458, pi00459, pi00460, pi00461, pi00462, pi00463, pi00464, pi00465, pi00466, pi00467, pi00468, pi00469, pi00470, pi00471, pi00472, pi00473, pi00474, pi00475, pi00476, pi00477, pi00478, pi00479, pi00480, pi00481, pi00482, pi00483, pi00484, pi00485, pi00486, pi00487, pi00488, pi00489, pi00490, pi00491, pi00492, pi00493, pi00494, pi00495, pi00496, pi00497, pi00498, pi00499, pi00500, pi00501, pi00502, pi00503, pi00504, pi00505, pi00506, pi00507, pi00508, pi00509, pi00510, pi00511, pi00512, pi00513, pi00514, pi00515, pi00516, pi00517, pi00518, pi00519, pi00520, pi00521, pi00522, pi00523, pi00524, pi00525, pi00526, pi00527, pi00528, pi00529, pi00530, pi00531, pi00532, pi00533, pi00534, pi00535, pi00536, pi00537, pi00538, pi00539, pi00540, pi00541, pi00542, pi00543, pi00544, pi00545, pi00546, pi00547, pi00548, pi00549, pi00550, pi00551, pi00552, pi00553, pi00554, pi00555, pi00556, pi00557, pi00558, pi00559, pi00560, pi00561, pi00562, pi00563, pi00564, pi00565, pi00566, pi00567, pi00568, pi00569, pi00570, pi00571, pi00572, pi00573, pi00574, pi00575, pi00576, pi00577, pi00578, pi00579, pi00580, pi00581, pi00582, pi00583, pi00584, pi00585, pi00586, pi00587, pi00588, pi00589, pi00590, pi00591, pi00592, pi00593, pi00594, pi00595, pi00596, pi00597, pi00598, pi00599, pi00600, pi00601, pi00602, pi00603, pi00604, pi00605, pi00606, pi00607, pi00608, pi00609, pi00610, pi00611, pi00612, pi00613, pi00614, pi00615, pi00616, pi00617, pi00618, pi00619, pi00620, pi00621, pi00622, pi00623, pi00624, pi00625, pi00626, pi00627, pi00628, pi00629, pi00630, pi00631, pi00632, pi00633, pi00634, pi00635, pi00636, pi00637, pi00638, pi00639, pi00640, pi00641, pi00642, pi00643, pi00644, pi00645, pi00646, pi00647, pi00648, pi00649, pi00650, pi00651, pi00652, pi00653, pi00654, pi00655, pi00656, pi00657, pi00658, pi00659, pi00660, pi00661, pi00662, pi00663, pi00664, pi00665, pi00666, pi00667, pi00668, pi00669, pi00670, pi00671, pi00672, pi00673, pi00674, pi00675, pi00676, pi00677, pi00678, pi00679, pi00680, pi00681, pi00682, pi00683, pi00684, pi00685, pi00686, pi00687, pi00688, pi00689, pi00690, pi00691, pi00692, pi00693, pi00694, pi00695, pi00696, pi00697, pi00698, pi00699, pi00700, pi00701, pi00702, pi00703, pi00704, pi00705, pi00706, pi00707, pi00708, pi00709, pi00710, pi00711, pi00712, pi00713, pi00714, pi00715, pi00716, pi00717, pi00718, pi00719, pi00720, pi00721, pi00722, pi00723, pi00724, pi00725, pi00726, pi00727, pi00728, pi00729, pi00730, pi00731, pi00732, pi00733, pi00734, pi00735, pi00736, pi00737, pi00738, pi00739, pi00740, pi00741, pi00742, pi00743, pi00744, pi00745, pi00746, pi00747, pi00748, pi00749, pi00750, pi00751, pi00752, pi00753, pi00754, pi00755, pi00756, pi00757, pi00758, pi00759, pi00760, pi00761, pi00762, pi00763, pi00764, pi00765, pi00766, pi00767, pi00768, pi00769, pi00770, pi00771, pi00772, pi00773, pi00774, pi00775, pi00776, pi00777, pi00778, pi00779, pi00780, pi00781, pi00782, pi00783, pi00784, pi00785, pi00786, pi00787, pi00788, pi00789, pi00790, pi00791, pi00792, pi00793, pi00794, pi00795, pi00796, pi00797, pi00798, pi00799, pi00800, pi00801, pi00802, pi00803, pi00804, pi00805, pi00806, pi00807, pi00808, pi00809, pi00810, pi00811, pi00812, pi00813, pi00814, pi00815, pi00816, pi00817, pi00818, pi00819, pi00820, pi00821, pi00822, pi00823, pi00824, pi00825, pi00826, pi00827, pi00828, pi00829, pi00830, pi00831, pi00832, pi00833, pi00834, pi00835, pi00836, pi00837, pi00838, pi00839, pi00840, pi00841, pi00842, pi00843, pi00844, pi00845, pi00846, pi00847, pi00848, pi00849, pi00850, pi00851, pi00852, pi00853, pi00854, pi00855, pi00856, pi00857, pi00858, pi00859, pi00860, pi00861, pi00862, pi00863, pi00864, pi00865, pi00866, pi00867, pi00868, pi00869, pi00870, pi00871, pi00872, pi00873, pi00874, pi00875, pi00876, pi00877, pi00878, pi00879, pi00880, pi00881, pi00882, pi00883, pi00884, pi00885, pi00886, pi00887, pi00888, pi00889, pi00890, pi00891, pi00892, pi00893, pi00894, pi00895, pi00896, pi00897, pi00898, pi00899, pi00900, pi00901, pi00902, pi00903, pi00904, pi00905, pi00906, pi00907, pi00908, pi00909, pi00910, pi00911, pi00912, pi00913, pi00914, pi00915, pi00916, pi00917, pi00918, pi00919, pi00920, pi00921, pi00922, pi00923, pi00924, pi00925, pi00926, pi00927, pi00928, pi00929, pi00930, pi00931, pi00932, pi00933, pi00934, pi00935, pi00936, pi00937, pi00938, pi00939, pi00940, pi00941, pi00942, pi00943, pi00944, pi00945, pi00946, pi00947, pi00948, pi00949, pi00950, pi00951, pi00952, pi00953, pi00954, pi00955, pi00956, pi00957, pi00958, pi00959, pi00960, pi00961, pi00962, pi00963, pi00964, pi00965, pi00966, pi00967, pi00968, pi00969, pi00970, pi00971, pi00972, pi00973, pi00974, pi00975, pi00976, pi00977, pi00978, pi00979, pi00980, pi00981, pi00982, pi00983, pi00984, pi00985, pi00986, pi00987, pi00988, pi00989, pi00990, pi00991, pi00992, pi00993, pi00994, pi00995, pi00996, pi00997, pi00998, pi00999, pi01000, pi01001, pi01002, pi01003, pi01004, pi01005, pi01006, pi01007, pi01008, pi01009, pi01010, pi01011, pi01012, pi01013, pi01014, pi01015, pi01016, pi01017, pi01018, pi01019, pi01020, pi01021, pi01022, pi01023, pi01024, pi01025, pi01026, pi01027, pi01028, pi01029, pi01030, pi01031, pi01032, pi01033, pi01034, pi01035, pi01036, pi01037, pi01038, pi01039, pi01040, pi01041, pi01042, pi01043, pi01044, pi01045, pi01046, pi01047, pi01048, pi01049, pi01050, pi01051, pi01052, pi01053, pi01054, pi01055, pi01056, pi01057, pi01058, pi01059, pi01060, pi01061, pi01062, pi01063, pi01064, pi01065, pi01066, pi01067, pi01068, pi01069, pi01070, pi01071, pi01072, pi01073, pi01074, pi01075, pi01076, pi01077, pi01078, pi01079, pi01080, pi01081, pi01082, pi01083, pi01084, pi01085, pi01086, pi01087, pi01088, pi01089, pi01090, pi01091, pi01092, pi01093, pi01094, pi01095, pi01096, pi01097, pi01098, pi01099, pi01100, pi01101, pi01102, pi01103, pi01104, pi01105, pi01106, pi01107, pi01108, pi01109, pi01110, pi01111, pi01112, pi01113, pi01114, pi01115, pi01116, pi01117, pi01118, pi01119, pi01120, pi01121, pi01122, pi01123, pi01124, pi01125, pi01126, pi01127, pi01128, pi01129, pi01130, pi01131, pi01132, pi01133, pi01134, pi01135, pi01136, pi01137, pi01138, pi01139, pi01140, pi01141, pi01142, pi01143, pi01144, pi01145, pi01146, pi01147, pi01148, pi01149, pi01150, pi01151, pi01152, pi01153, pi01154, pi01155, pi01156, pi01157, pi01158, pi01159, pi01160, pi01161, pi01162, pi01163, pi01164, pi01165, pi01166, pi01167, pi01168, pi01169, pi01170, pi01171, pi01172, pi01173, pi01174, pi01175, pi01176, pi01177, pi01178, pi01179, pi01180, pi01181, pi01182, pi01183, pi01184, pi01185, pi01186, pi01187, pi01188, pi01189, pi01190, pi01191, pi01192, pi01193, pi01194, pi01195, pi01196, pi01197, pi01198, pi01199, pi01200, pi01201, pi01202, pi01203, pi01204, pi01205, pi01206, pi01207, pi01208, pi01209, pi01210, pi01211, pi01212, pi01213, pi01214, pi01215, pi01216, pi01217, pi01218, pi01219, pi01220, pi01221, pi01222, pi01223, pi01224, pi01225, pi01226, pi01227, pi01228, pi01229, pi01230, pi01231, pi01232, pi01233, pi01234, pi01235, pi01236, pi01237, pi01238, pi01239, pi01240, pi01241, pi01242, pi01243, pi01244, pi01245, pi01246, pi01247, pi01248, pi01249, pi01250, pi01251, pi01252, pi01253, pi01254, pi01255, pi01256, pi01257, pi01258, pi01259, pi01260, pi01261, pi01262, pi01263, pi01264, pi01265, pi01266, pi01267, pi01268, pi01269, pi01270, pi01271, pi01272, pi01273, pi01274, pi01275, pi01276, pi01277, pi01278, pi01279, pi01280, pi01281, pi01282, pi01283, pi01284, pi01285, pi01286, pi01287, pi01288, pi01289, pi01290, pi01291, pi01292, pi01293, pi01294, pi01295, pi01296, pi01297, pi01298, pi01299, pi01300, pi01301, pi01302, pi01303, pi01304, pi01305, pi01306, pi01307, pi01308, pi01309, pi01310, pi01311, pi01312, pi01313, pi01314, pi01315, pi01316, pi01317, pi01318, pi01319, pi01320, pi01321, pi01322, pi01323, pi01324, pi01325, pi01326, pi01327, pi01328, pi01329, pi01330, pi01331, pi01332, pi01333, pi01334, pi01335, pi01336, pi01337, pi01338, pi01339, pi01340, pi01341, pi01342, pi01343, pi01344, pi01345, pi01346, pi01347, pi01348, pi01349, pi01350, pi01351, pi01352, pi01353, pi01354, pi01355, pi01356, pi01357, pi01358, pi01359, pi01360, pi01361, pi01362, pi01363, pi01364, pi01365, pi01366, pi01367, pi01368, pi01369, pi01370, pi01371, pi01372, pi01373, pi01374, pi01375, pi01376, pi01377, pi01378, pi01379, pi01380, pi01381, pi01382, pi01383, pi01384, pi01385, pi01386, pi01387, pi01388, pi01389, pi01390, pi01391, pi01392, pi01393, pi01394, pi01395, pi01396, pi01397, pi01398, pi01399, pi01400, pi01401, pi01402, pi01403, pi01404, pi01405, pi01406, pi01407, pi01408, pi01409, pi01410, pi01411, pi01412, pi01413, pi01414, pi01415, pi01416, pi01417, pi01418, pi01419, pi01420, pi01421, pi01422, pi01423, pi01424, pi01425, pi01426, pi01427, pi01428, pi01429, pi01430, pi01431, pi01432, pi01433, pi01434, pi01435, pi01436, pi01437, pi01438, pi01439, pi01440, pi01441, pi01442, pi01443, pi01444, pi01445, pi01446, pi01447, pi01448, pi01449, pi01450, pi01451, pi01452, pi01453, pi01454, pi01455, pi01456, pi01457, pi01458, pi01459, pi01460, pi01461, pi01462, pi01463, pi01464, pi01465, pi01466, pi01467, pi01468, pi01469, pi01470, pi01471, pi01472, pi01473, pi01474, pi01475, pi01476, pi01477, pi01478, pi01479, pi01480, pi01481, pi01482, pi01483, pi01484, pi01485, pi01486, pi01487, pi01488, pi01489, pi01490, pi01491, pi01492, pi01493, pi01494, pi01495, pi01496, pi01497, pi01498, pi01499, pi01500, pi01501, pi01502, pi01503, pi01504, pi01505, pi01506, pi01507, pi01508, pi01509, pi01510, pi01511, pi01512, pi01513, pi01514, pi01515, pi01516, pi01517, pi01518, pi01519, pi01520, pi01521, pi01522, pi01523, pi01524, pi01525, pi01526, pi01527, pi01528, pi01529, pi01530, pi01531, pi01532, pi01533, pi01534, pi01535, pi01536, pi01537, pi01538, pi01539, pi01540, pi01541, pi01542, pi01543, pi01544, pi01545, pi01546, pi01547, pi01548, pi01549, pi01550, pi01551, pi01552, pi01553, pi01554, pi01555, pi01556, pi01557, pi01558, pi01559, pi01560, pi01561, pi01562, pi01563, pi01564, pi01565, pi01566, pi01567, pi01568, pi01569, pi01570, pi01571, pi01572, pi01573, pi01574, pi01575, pi01576, pi01577, pi01578, pi01579, pi01580, pi01581, pi01582, pi01583, pi01584, pi01585, pi01586, pi01587, pi01588, pi01589, pi01590, pi01591, pi01592, pi01593, pi01594, pi01595, pi01596, pi01597, pi01598, pi01599, pi01600, pi01601, pi01602, pi01603, pi01604, pi01605, pi01606, pi01607, pi01608, pi01609, pi01610, pi01611, pi01612, pi01613, pi01614, pi01615, pi01616, pi01617, pi01618, pi01619, pi01620, pi01621, pi01622, pi01623, pi01624, pi01625, pi01626, pi01627, pi01628, pi01629, pi01630, pi01631, pi01632, pi01633, pi01634, pi01635, pi01636, pi01637, pi01638, pi01639, pi01640, pi01641, pi01642, pi01643, pi01644, pi01645, pi01646, pi01647, pi01648, pi01649, pi01650, pi01651, pi01652, pi01653, pi01654, pi01655, pi01656, pi01657, pi01658, pi01659, pi01660, pi01661, pi01662, pi01663, pi01664, pi01665, pi01666, pi01667, pi01668, pi01669, pi01670, pi01671, pi01672, pi01673, pi01674, pi01675, pi01676, pi01677, pi01678, pi01679, pi01680, pi01681, pi01682, pi01683, pi01684, pi01685, pi01686, pi01687, pi01688, pi01689, pi01690, pi01691, pi01692, pi01693, pi01694, pi01695, pi01696, pi01697, pi01698, pi01699, pi01700, pi01701, pi01702, pi01703, pi01704, pi01705, pi01706, pi01707, pi01708, pi01709, pi01710, pi01711, pi01712, pi01713, pi01714, pi01715, pi01716, pi01717, pi01718, pi01719, pi01720, pi01721, pi01722, pi01723, pi01724, pi01725, pi01726, pi01727, pi01728, pi01729, pi01730, pi01731, pi01732, pi01733, pi01734, pi01735, pi01736, pi01737, pi01738, pi01739, pi01740, pi01741, pi01742, pi01743, pi01744, pi01745, pi01746, pi01747, pi01748, pi01749, pi01750, pi01751, pi01752, pi01753, pi01754, pi01755, pi01756, pi01757, pi01758, pi01759, pi01760, pi01761, pi01762, pi01763, pi01764, pi01765, pi01766, pi01767, pi01768, pi01769, pi01770, pi01771, pi01772, pi01773, pi01774, pi01775, pi01776, pi01777, pi01778, pi01779, pi01780, pi01781, pi01782, pi01783, pi01784, pi01785, pi01786, pi01787, pi01788, pi01789, pi01790, pi01791, pi01792, pi01793, pi01794, pi01795, pi01796, pi01797, pi01798, pi01799, pi01800, pi01801, pi01802, pi01803, pi01804, pi01805, pi01806, pi01807, pi01808, pi01809, pi01810, pi01811, pi01812, pi01813, pi01814, pi01815, pi01816, pi01817, pi01818, pi01819, pi01820, pi01821, pi01822, pi01823, pi01824, pi01825, pi01826, pi01827, pi01828, pi01829, pi01830, pi01831, pi01832, pi01833, pi01834, pi01835, pi01836, pi01837, pi01838, pi01839, pi01840, pi01841, pi01842, pi01843, pi01844, pi01845, pi01846, pi01847, pi01848, pi01849, pi01850, pi01851, pi01852, pi01853, pi01854, pi01855, pi01856, pi01857, pi01858, pi01859, pi01860, pi01861, pi01862, pi01863, pi01864, pi01865, pi01866, pi01867, pi01868, pi01869, pi01870, pi01871, pi01872, pi01873, pi01874, pi01875, pi01876, pi01877, pi01878, pi01879, pi01880, pi01881, pi01882, pi01883, pi01884, pi01885, pi01886, pi01887, pi01888, pi01889, pi01890, pi01891, pi01892, pi01893, pi01894, pi01895, pi01896, pi01897, pi01898, pi01899, pi01900, pi01901, pi01902, pi01903, pi01904, pi01905, pi01906, pi01907, pi01908, pi01909, pi01910, pi01911, pi01912, pi01913, pi01914, pi01915, pi01916, pi01917, pi01918, pi01919, pi01920, pi01921, pi01922, pi01923, pi01924, pi01925, pi01926, pi01927, pi01928, pi01929, pi01930, pi01931, pi01932, pi01933, pi01934, pi01935, pi01936, pi01937, pi01938, pi01939, pi01940, pi01941, pi01942, pi01943, pi01944, pi01945, pi01946, pi01947, pi01948, pi01949, pi01950, pi01951, pi01952, pi01953, pi01954, pi01955, pi01956, pi01957, pi01958, pi01959, pi01960, pi01961, pi01962, pi01963, pi01964, pi01965, pi01966, pi01967, pi01968, pi01969, pi01970, pi01971, pi01972, pi01973, pi01974, pi01975, pi01976, pi01977, pi01978, pi01979, pi01980, pi01981, pi01982, pi01983, pi01984, pi01985, pi01986, pi01987, pi01988, pi01989, pi01990, pi01991, pi01992, pi01993, pi01994, pi01995, pi01996, pi01997, pi01998, pi01999, pi02000, pi02001, pi02002, pi02003, pi02004, pi02005, pi02006, pi02007, pi02008, pi02009, pi02010, pi02011, pi02012, pi02013, pi02014, pi02015, pi02016, pi02017, pi02018, pi02019, pi02020, pi02021, pi02022, pi02023, pi02024, pi02025, pi02026, pi02027, pi02028, pi02029, pi02030, pi02031, pi02032, pi02033, pi02034, pi02035, pi02036, pi02037, pi02038, pi02039, pi02040, pi02041, pi02042, pi02043, pi02044, pi02045, pi02046, pi02047, pi02048, pi02049, pi02050, pi02051, pi02052, pi02053, pi02054, pi02055, pi02056, pi02057, pi02058, pi02059, pi02060, pi02061, pi02062, pi02063, pi02064, pi02065, pi02066, pi02067, pi02068, pi02069, pi02070, pi02071, pi02072, pi02073, pi02074, pi02075, pi02076, pi02077, pi02078, pi02079, pi02080, pi02081, pi02082, pi02083, pi02084, pi02085, pi02086, pi02087, pi02088, pi02089, pi02090, pi02091, pi02092, pi02093, pi02094, pi02095, pi02096, pi02097, pi02098, pi02099, pi02100, pi02101, pi02102, pi02103, pi02104, pi02105, pi02106, pi02107, pi02108, pi02109, pi02110, pi02111, pi02112, pi02113, pi02114, pi02115, pi02116, pi02117, pi02118, pi02119, pi02120, pi02121, pi02122, pi02123, pi02124, pi02125, pi02126, pi02127, pi02128, pi02129, pi02130, pi02131, pi02132, pi02133, pi02134, pi02135, pi02136, pi02137, pi02138, pi02139, pi02140, pi02141, pi02142, pi02143, pi02144, pi02145, pi02146, pi02147, pi02148, pi02149, pi02150, pi02151, pi02152, pi02153, pi02154, pi02155, pi02156, pi02157, pi02158, pi02159, pi02160, pi02161, pi02162, pi02163, pi02164, pi02165, pi02166, pi02167, pi02168, pi02169, pi02170, pi02171, pi02172, pi02173, pi02174, pi02175, pi02176, pi02177, pi02178, pi02179, pi02180, pi02181, pi02182, pi02183, pi02184, pi02185, pi02186, pi02187, pi02188, pi02189, pi02190, pi02191, pi02192, pi02193, pi02194, pi02195, pi02196, pi02197, pi02198, pi02199, pi02200, pi02201, pi02202, pi02203, pi02204, pi02205, pi02206, pi02207, pi02208, pi02209, pi02210, pi02211, pi02212, pi02213, pi02214, pi02215, pi02216, pi02217, pi02218, pi02219, pi02220, pi02221, pi02222, pi02223, pi02224, pi02225, pi02226, pi02227, pi02228, pi02229, pi02230, pi02231, pi02232, pi02233, pi02234, pi02235, pi02236, pi02237, pi02238, pi02239, pi02240, pi02241, pi02242, pi02243, pi02244, pi02245, pi02246, pi02247, pi02248, pi02249, pi02250, pi02251, pi02252, pi02253, pi02254, pi02255, pi02256, pi02257, pi02258, pi02259, pi02260, pi02261, pi02262, pi02263, pi02264, pi02265, pi02266, pi02267, pi02268, pi02269, pi02270, pi02271, pi02272, pi02273, pi02274, pi02275, pi02276, pi02277, pi02278, pi02279, pi02280, pi02281, pi02282, pi02283, pi02284, pi02285, pi02286, pi02287, pi02288, pi02289, pi02290, pi02291, pi02292, pi02293, pi02294, pi02295, pi02296, pi02297, pi02298, pi02299, pi02300, pi02301, pi02302, pi02303, pi02304, pi02305, pi02306, pi02307, pi02308, pi02309, pi02310, pi02311, pi02312, pi02313, pi02314, pi02315, pi02316, pi02317, pi02318, pi02319, pi02320, pi02321, pi02322, pi02323, pi02324, pi02325, pi02326, pi02327, pi02328, pi02329, pi02330, pi02331, pi02332, pi02333, pi02334, pi02335, pi02336, pi02337, pi02338, pi02339, pi02340, pi02341, pi02342, pi02343, pi02344, pi02345, pi02346, pi02347, pi02348, pi02349, pi02350, pi02351, pi02352, pi02353, pi02354, pi02355, pi02356, pi02357, pi02358, pi02359, pi02360, pi02361, pi02362, pi02363, pi02364, pi02365, pi02366, pi02367, pi02368, pi02369, pi02370, pi02371, pi02372, pi02373, pi02374, pi02375, pi02376, pi02377, pi02378, pi02379, pi02380, pi02381, pi02382, pi02383, pi02384, pi02385, pi02386, pi02387, pi02388, pi02389, pi02390, pi02391, pi02392, pi02393, pi02394, pi02395, pi02396, pi02397, pi02398, pi02399, pi02400, pi02401, pi02402, pi02403, pi02404, pi02405, pi02406, pi02407, pi02408, pi02409, pi02410, pi02411, pi02412, pi02413, pi02414, pi02415, pi02416, pi02417, pi02418, pi02419, pi02420, pi02421, pi02422, pi02423, pi02424, pi02425, pi02426, pi02427, pi02428, pi02429, pi02430, pi02431, pi02432, pi02433, pi02434, pi02435, pi02436, pi02437, pi02438, pi02439, pi02440, pi02441, pi02442, pi02443, pi02444, pi02445, pi02446, pi02447, pi02448, pi02449, pi02450, pi02451, pi02452, pi02453, pi02454, pi02455, pi02456, pi02457, pi02458, pi02459, pi02460, pi02461, pi02462, pi02463, pi02464, pi02465, pi02466, pi02467, pi02468, pi02469, pi02470, pi02471, pi02472, pi02473, pi02474, pi02475, pi02476, pi02477, pi02478, pi02479, pi02480, pi02481, pi02482, pi02483, pi02484, pi02485, pi02486, pi02487, pi02488, pi02489, pi02490, pi02491, pi02492, pi02493, pi02494, pi02495, pi02496, pi02497, pi02498, pi02499, pi02500, pi02501, pi02502, pi02503, pi02504, pi02505, pi02506, pi02507, pi02508, pi02509, pi02510, pi02511, pi02512, pi02513, pi02514, pi02515, pi02516, pi02517, pi02518, pi02519, pi02520, pi02521, pi02522, pi02523, pi02524, pi02525, pi02526, pi02527, pi02528, pi02529, pi02530, pi02531, pi02532, pi02533, pi02534, pi02535, pi02536, pi02537, pi02538, pi02539, pi02540, pi02541, pi02542, pi02543, pi02544, pi02545, pi02546, pi02547, pi02548, pi02549, pi02550, pi02551, pi02552, pi02553, pi02554, pi02555, pi02556, pi02557, pi02558, pi02559, pi02560, pi02561, pi02562, pi02563, pi02564, pi02565, pi02566, pi02567, pi02568, pi02569, pi02570, pi02571, pi02572, pi02573, pi02574, pi02575, pi02576, pi02577, pi02578, pi02579, pi02580, pi02581, pi02582, pi02583, pi02584, pi02585, pi02586, pi02587, pi02588, pi02589, pi02590, pi02591, pi02592, pi02593, pi02594, pi02595, pi02596, pi02597, pi02598, pi02599, pi02600, pi02601, pi02602, pi02603, pi02604, pi02605, pi02606, pi02607, pi02608, pi02609, pi02610, pi02611, pi02612, pi02613, pi02614, pi02615, pi02616, pi02617, pi02618, pi02619, pi02620, pi02621, pi02622, pi02623, pi02624, pi02625, pi02626, pi02627, pi02628, pi02629, pi02630, pi02631, pi02632, pi02633, pi02634, pi02635, pi02636, pi02637, pi02638, pi02639, pi02640, pi02641, pi02642, pi02643, pi02644, pi02645, pi02646, pi02647, pi02648, pi02649, pi02650, pi02651, pi02652, pi02653, pi02654, pi02655, pi02656, pi02657, pi02658, pi02659, pi02660, pi02661, pi02662, pi02663, pi02664, pi02665, pi02666, pi02667, pi02668, pi02669, pi02670, pi02671, pi02672, pi02673, pi02674, pi02675, pi02676, pi02677, pi02678, pi02679, pi02680, pi02681, pi02682, pi02683, pi02684, pi02685, pi02686, pi02687, pi02688, pi02689, pi02690, pi02691, pi02692, pi02693, pi02694, pi02695, pi02696, pi02697, pi02698, pi02699, pi02700, pi02701, pi02702, pi02703, pi02704, pi02705, pi02706, pi02707, pi02708, pi02709, pi02710, pi02711, pi02712, pi02713, pi02714, pi02715, pi02716, pi02717, pi02718, pi02719, pi02720, pi02721, pi02722, pi02723, pi02724, pi02725, pi02726, pi02727, pi02728, pi02729, pi02730, pi02731, pi02732, pi02733, pi02734, pi02735, pi02736, pi02737, pi02738, pi02739, pi02740, pi02741, pi02742, pi02743, pi02744, pi02745, pi02746, pi02747, pi02748, pi02749, pi02750, pi02751, pi02752, pi02753, pi02754, pi02755, pi02756, pi02757, pi02758, pi02759, pi02760, pi02761, pi02762, pi02763, pi02764, pi02765, pi02766, pi02767, pi02768, pi02769, pi02770, pi02771, pi02772, pi02773, pi02774, pi02775, pi02776, pi02777, pi02778, pi02779, pi02780, pi02781, pi02782, pi02783, pi02784, pi02785, pi02786, pi02787, pi02788, pi02789, pi02790, pi02791, pi02792, pi02793, pi02794, pi02795, pi02796, pi02797, pi02798, pi02799, pi02800, pi02801, pi02802, pi02803, pi02804, pi02805, pi02806, pi02807, pi02808, pi02809, pi02810, pi02811, pi02812, pi02813, pi02814, pi02815, pi02816, pi02817, pi02818, pi02819, pi02820, pi02821, pi02822, pi02823, pi02824, pi02825, pi02826, pi02827, pi02828, pi02829, pi02830, pi02831, pi02832, pi02833, pi02834, pi02835, pi02836, pi02837, pi02838, pi02839, pi02840, pi02841, pi02842, pi02843, pi02844, pi02845, pi02846, pi02847, pi02848, pi02849, pi02850, pi02851, pi02852, pi02853, pi02854, pi02855, pi02856, pi02857, pi02858, pi02859, pi02860, pi02861, pi02862, pi02863, pi02864, pi02865, pi02866, pi02867, pi02868, pi02869, pi02870, pi02871, pi02872, pi02873, pi02874, pi02875, pi02876, pi02877, pi02878, pi02879, pi02880, pi02881, pi02882, pi02883, pi02884, pi02885, pi02886, pi02887, pi02888, pi02889, pi02890, pi02891, pi02892, pi02893, pi02894, pi02895, pi02896, pi02897, pi02898, pi02899, pi02900, pi02901, pi02902, pi02903, pi02904, pi02905, pi02906, pi02907, pi02908, pi02909, pi02910, pi02911, pi02912, pi02913, pi02914, pi02915, pi02916, pi02917, pi02918, pi02919, pi02920, pi02921, pi02922, pi02923, pi02924, pi02925, pi02926, pi02927, pi02928, pi02929, pi02930, pi02931, pi02932, pi02933, pi02934, pi02935, pi02936, pi02937, pi02938, pi02939, pi02940, pi02941, pi02942, pi02943, pi02944, pi02945, pi02946, pi02947, pi02948, pi02949, pi02950, pi02951, pi02952, pi02953, pi02954, pi02955, pi02956, pi02957, pi02958, pi02959, pi02960, pi02961, pi02962, pi02963, pi02964, pi02965, pi02966, pi02967, pi02968, pi02969, pi02970, pi02971, pi02972, pi02973, pi02974, pi02975, pi02976, pi02977, pi02978, pi02979, pi02980, pi02981, pi02982, pi02983, pi02984, pi02985, pi02986, pi02987, pi02988, pi02989, pi02990, pi02991, pi02992, pi02993, pi02994, pi02995, pi02996, pi02997, pi02998, pi02999, pi03000, pi03001, pi03002, pi03003, pi03004, pi03005, pi03006, pi03007, pi03008, pi03009, pi03010, pi03011, pi03012, pi03013, pi03014, pi03015, pi03016, pi03017, pi03018, pi03019, pi03020, pi03021, pi03022, pi03023, pi03024, pi03025, pi03026, pi03027, pi03028, pi03029, pi03030, pi03031, pi03032, pi03033, pi03034, pi03035, pi03036, pi03037, pi03038, pi03039, pi03040, pi03041, pi03042, pi03043, pi03044, pi03045, pi03046, pi03047, pi03048, pi03049, pi03050, pi03051, pi03052, pi03053, pi03054, pi03055, pi03056, pi03057, pi03058, pi03059, pi03060, pi03061, pi03062, pi03063, pi03064, pi03065, pi03066, pi03067, pi03068, pi03069, pi03070, pi03071, pi03072, pi03073, pi03074, pi03075, pi03076, pi03077, pi03078, pi03079, pi03080, pi03081, pi03082, pi03083, pi03084, pi03085, pi03086, pi03087, pi03088, pi03089, pi03090, pi03091, pi03092, pi03093, pi03094, pi03095, pi03096, pi03097, pi03098, pi03099, pi03100, pi03101, pi03102, pi03103, pi03104, pi03105, pi03106, pi03107, pi03108, pi03109, pi03110, pi03111, pi03112, pi03113, pi03114, pi03115, pi03116, pi03117, pi03118, pi03119, pi03120, pi03121, pi03122, pi03123, pi03124, pi03125, pi03126, pi03127, pi03128, pi03129, pi03130, pi03131, pi03132, pi03133, pi03134, pi03135, pi03136, pi03137, pi03138, pi03139, pi03140, pi03141, pi03142, pi03143, pi03144, pi03145, pi03146, pi03147, pi03148, pi03149, pi03150, pi03151, pi03152, pi03153, pi03154, pi03155, pi03156, pi03157, pi03158, pi03159, pi03160, pi03161, pi03162, pi03163, pi03164, pi03165, pi03166, pi03167, pi03168, pi03169, pi03170, pi03171, pi03172, pi03173, pi03174, pi03175, pi03176, pi03177, pi03178, pi03179, pi03180, pi03181, pi03182, pi03183, pi03184, pi03185, pi03186, pi03187, pi03188, pi03189, pi03190, pi03191, pi03192, pi03193, pi03194, pi03195, pi03196, pi03197, pi03198, pi03199, pi03200, pi03201, pi03202, pi03203, pi03204, pi03205, pi03206, pi03207, pi03208, pi03209, pi03210, pi03211, pi03212, pi03213, pi03214, pi03215, pi03216, pi03217, pi03218, pi03219, pi03220, pi03221, pi03222, pi03223, pi03224, pi03225, pi03226, pi03227, pi03228, pi03229, pi03230, pi03231, pi03232, pi03233, pi03234, pi03235, pi03236, pi03237, pi03238, pi03239, pi03240, pi03241, pi03242, pi03243, pi03244, pi03245, pi03246, pi03247, pi03248, pi03249, pi03250, pi03251, pi03252, pi03253, pi03254, pi03255, pi03256, pi03257, pi03258, pi03259, pi03260, pi03261, pi03262, pi03263, pi03264, pi03265, pi03266, pi03267, pi03268, pi03269, pi03270, pi03271, pi03272, pi03273, pi03274, pi03275, pi03276, pi03277, pi03278, pi03279, pi03280, pi03281, pi03282, pi03283, pi03284, pi03285, pi03286, pi03287, pi03288, pi03289, pi03290, pi03291, pi03292, pi03293, pi03294, pi03295, pi03296, pi03297, pi03298, pi03299, pi03300, pi03301, pi03302, pi03303, pi03304, pi03305, pi03306, pi03307, pi03308, pi03309, pi03310, pi03311, pi03312, pi03313, pi03314, pi03315, pi03316, pi03317, pi03318, pi03319, pi03320, pi03321, pi03322, pi03323, pi03324, pi03325, pi03326, pi03327, pi03328, pi03329, pi03330, pi03331, pi03332, pi03333, pi03334, pi03335, pi03336, pi03337, pi03338, pi03339, pi03340, pi03341, pi03342, pi03343, pi03344, pi03345, pi03346, pi03347, pi03348, pi03349, pi03350, pi03351, pi03352, pi03353, pi03354, pi03355, pi03356, pi03357, pi03358, pi03359, pi03360, pi03361, pi03362, pi03363, pi03364, pi03365, pi03366, pi03367, pi03368, pi03369, pi03370, pi03371, pi03372, pi03373, pi03374, pi03375, pi03376, pi03377, pi03378, pi03379, pi03380, pi03381, pi03382, pi03383, pi03384, pi03385, pi03386, pi03387, pi03388, pi03389, pi03390, pi03391, pi03392, pi03393, pi03394, pi03395, pi03396, pi03397, pi03398, pi03399, pi03400, pi03401, pi03402, pi03403, pi03404, pi03405, pi03406, pi03407, pi03408, pi03409, pi03410, pi03411, pi03412, pi03413, pi03414, pi03415, pi03416, pi03417, pi03418, pi03419, pi03420, pi03421, pi03422, pi03423, pi03424, pi03425, pi03426, pi03427, pi03428, pi03429, pi03430, pi03431, pi03432, pi03433, pi03434, pi03435, pi03436, pi03437, pi03438, pi03439, pi03440, pi03441, pi03442, pi03443, pi03444, pi03445, pi03446, pi03447, pi03448, pi03449, pi03450, pi03451, pi03452, pi03453, pi03454, pi03455, pi03456, pi03457, pi03458, pi03459, pi03460, pi03461, pi03462, pi03463, pi03464, pi03465, pi03466, pi03467, pi03468, pi03469, pi03470, pi03471, pi03472, pi03473, pi03474, pi03475, pi03476, pi03477, pi03478, pi03479, pi03480, pi03481, pi03482, pi03483, pi03484, pi03485, pi03486, pi03487, pi03488, pi03489, pi03490, pi03491, pi03492, pi03493, pi03494, pi03495, pi03496, pi03497, pi03498, pi03499, pi03500, pi03501, pi03502, pi03503, pi03504, pi03505, pi03506, pi03507, pi03508, pi03509, pi03510, pi03511, pi03512, pi03513, pi03514, pi03515, pi03516, pi03517, pi03518, pi03519, pi03520, pi03521, pi03522, pi03523, pi03524, pi03525, pi03526, pi03527, pi03528, pi03529, pi03530, pi03531, pi03532, pi03533, pi03534, pi03535, pi03536, pi03537, pi03538, pi03539, pi03540, pi03541, pi03542, pi03543, pi03544, pi03545, pi03546, pi03547, pi03548, pi03549, pi03550, pi03551, pi03552, pi03553, pi03554, pi03555, pi03556, pi03557, pi03558, pi03559, pi03560, pi03561, pi03562, pi03563, pi03564, pi03565, pi03566, pi03567, pi03568, pi03569, pi03570, pi03571, pi03572, pi03573, pi03574, pi03575, pi03576, pi03577, pi03578, pi03579, pi03580, pi03581, pi03582, pi03583, pi03584, pi03585, pi03586, pi03587, pi03588, pi03589, pi03590, pi03591, pi03592, pi03593, pi03594, pi03595, pi03596, pi03597, pi03598, pi03599, pi03600, pi03601, pi03602, pi03603, pi03604, pi03605, pi03606, pi03607, pi03608, pi03609, pi03610, pi03611, pi03612, pi03613, pi03614, pi03615, pi03616, pi03617, pi03618, pi03619, pi03620, pi03621, pi03622, pi03623, pi03624, pi03625, pi03626, pi03627, pi03628, pi03629, pi03630, pi03631, pi03632, pi03633, pi03634, pi03635, pi03636, pi03637, pi03638, pi03639, pi03640, pi03641, pi03642, pi03643, pi03644, pi03645, pi03646, pi03647, pi03648, pi03649, pi03650, pi03651, pi03652, pi03653, pi03654, pi03655, pi03656, pi03657, pi03658, pi03659, pi03660, pi03661, pi03662, pi03663, pi03664, pi03665, pi03666, pi03667, pi03668, pi03669, pi03670, pi03671, pi03672, pi03673, pi03674, pi03675, pi03676, pi03677, pi03678, pi03679, pi03680, pi03681, pi03682, pi03683, pi03684, pi03685, pi03686, pi03687, pi03688, pi03689, pi03690, pi03691, pi03692, pi03693, pi03694, pi03695, pi03696, pi03697, pi03698, pi03699, pi03700, pi03701, pi03702, pi03703, pi03704, pi03705, pi03706, pi03707, pi03708, pi03709, pi03710, pi03711, pi03712, pi03713, pi03714, pi03715, pi03716, pi03717, pi03718, pi03719, pi03720, pi03721, pi03722, pi03723, pi03724, pi03725, pi03726, pi03727, pi03728, pi03729, pi03730, pi03731, pi03732, pi03733, pi03734, pi03735, pi03736, pi03737, pi03738, pi03739, pi03740, pi03741, pi03742, pi03743, pi03744, pi03745, pi03746, pi03747, pi03748, pi03749, pi03750, pi03751, pi03752, pi03753, pi03754, pi03755, pi03756, pi03757, pi03758, pi03759, pi03760, pi03761, pi03762, pi03763, pi03764, pi03765, pi03766, pi03767, pi03768, pi03769, pi03770, pi03771, pi03772, pi03773, pi03774, pi03775, pi03776, pi03777, pi03778, pi03779, pi03780, pi03781, pi03782, pi03783, pi03784, pi03785, pi03786, pi03787, pi03788, pi03789, pi03790, pi03791, pi03792, pi03793, pi03794, pi03795, pi03796, pi03797, pi03798, pi03799, pi03800, pi03801, pi03802, pi03803, pi03804, pi03805, pi03806, pi03807, pi03808, pi03809, pi03810, pi03811, pi03812, pi03813, pi03814, pi03815, pi03816, pi03817, pi03818, pi03819, pi03820, pi03821, pi03822, pi03823, pi03824, pi03825, pi03826, pi03827, pi03828, pi03829, pi03830, pi03831, pi03832, pi03833, pi03834, pi03835, pi03836, pi03837, pi03838, pi03839, pi03840, pi03841, pi03842, pi03843, pi03844, pi03845, pi03846, pi03847, pi03848, pi03849, pi03850, pi03851, pi03852, pi03853, pi03854, pi03855, pi03856, pi03857, pi03858, pi03859, pi03860, pi03861, pi03862, pi03863, pi03864, pi03865, pi03866, pi03867, pi03868, pi03869, pi03870, pi03871, pi03872, pi03873, pi03874, pi03875, pi03876, pi03877, pi03878, pi03879, pi03880, pi03881, pi03882, pi03883, pi03884, pi03885, pi03886, pi03887, pi03888, pi03889, pi03890, pi03891, pi03892, pi03893, pi03894, pi03895, pi03896, pi03897, pi03898, pi03899, pi03900, pi03901, pi03902, pi03903, pi03904, pi03905, pi03906, pi03907, pi03908, pi03909, pi03910, pi03911, pi03912, pi03913, pi03914, pi03915, pi03916, pi03917, pi03918, pi03919, pi03920, pi03921, pi03922, pi03923, pi03924, pi03925, pi03926, pi03927, pi03928, pi03929, pi03930, pi03931, pi03932, pi03933, pi03934, pi03935, pi03936, pi03937, pi03938, pi03939, pi03940, pi03941, pi03942, pi03943, pi03944, pi03945, pi03946, pi03947, pi03948, pi03949, pi03950, pi03951, pi03952, pi03953, pi03954, pi03955, pi03956, pi03957, pi03958, pi03959, pi03960, pi03961, pi03962, pi03963, pi03964, pi03965, pi03966, pi03967, pi03968, pi03969, pi03970, pi03971, pi03972, pi03973, pi03974, pi03975, pi03976, pi03977, pi03978, pi03979, pi03980, pi03981, pi03982, pi03983, pi03984, pi03985, pi03986, pi03987, pi03988, pi03989, pi03990, pi03991, pi03992, pi03993, pi03994, pi03995, pi03996, pi03997, pi03998, pi03999, pi04000, pi04001, pi04002, pi04003, pi04004, pi04005, pi04006, pi04007, pi04008, pi04009, pi04010, pi04011, pi04012, pi04013, pi04014, pi04015, pi04016, pi04017, pi04018, pi04019, pi04020, pi04021, pi04022, pi04023, pi04024, pi04025, pi04026, pi04027, pi04028, pi04029, pi04030, pi04031, pi04032, pi04033, pi04034, pi04035, pi04036, pi04037, pi04038, pi04039, pi04040, pi04041, pi04042, pi04043, pi04044, pi04045, pi04046, pi04047, pi04048, pi04049, pi04050, pi04051, pi04052, pi04053, pi04054, pi04055, pi04056, pi04057, pi04058, pi04059, pi04060, pi04061, pi04062, pi04063, pi04064, pi04065, pi04066, pi04067, pi04068, pi04069, pi04070, pi04071, pi04072, pi04073, pi04074, pi04075, pi04076, pi04077, pi04078, pi04079, pi04080, pi04081, pi04082, pi04083, pi04084, pi04085, pi04086, pi04087, pi04088, pi04089, pi04090, pi04091, pi04092, pi04093, pi04094, pi04095, pi04096, pi04097, pi04098, pi04099, pi04100, pi04101, pi04102, pi04103, pi04104, pi04105, pi04106, pi04107, pi04108, pi04109, pi04110, pi04111, pi04112, pi04113, pi04114, pi04115, pi04116, pi04117, pi04118, pi04119, pi04120, pi04121, pi04122, pi04123, pi04124, pi04125, pi04126, pi04127, pi04128, pi04129, pi04130, pi04131, pi04132, pi04133, pi04134, pi04135, pi04136, pi04137, pi04138, pi04139, pi04140, pi04141, pi04142, pi04143, pi04144, pi04145, pi04146, pi04147, pi04148, pi04149, pi04150, pi04151, pi04152, pi04153, pi04154, pi04155, pi04156, pi04157, pi04158, pi04159, pi04160, pi04161, pi04162, pi04163, pi04164, pi04165, pi04166, pi04167, pi04168, pi04169, pi04170, pi04171, pi04172, pi04173, pi04174, pi04175, pi04176, pi04177, pi04178, pi04179, pi04180, pi04181, pi04182, pi04183, pi04184, pi04185, pi04186, pi04187, pi04188, pi04189, pi04190, pi04191, pi04192, pi04193, pi04194, pi04195, pi04196, pi04197, pi04198, pi04199, pi04200, pi04201, pi04202, pi04203, pi04204, pi04205, pi04206, pi04207, pi04208, pi04209, pi04210, pi04211, pi04212, pi04213, pi04214, pi04215, pi04216, pi04217, pi04218, pi04219, pi04220, pi04221, pi04222, pi04223, pi04224, pi04225, pi04226, pi04227, pi04228, pi04229, pi04230, pi04231, pi04232, pi04233, pi04234, pi04235, pi04236, pi04237, pi04238, pi04239, pi04240, pi04241, pi04242, pi04243, pi04244, pi04245, pi04246, pi04247, pi04248, pi04249, pi04250, pi04251, pi04252, pi04253, pi04254, pi04255, pi04256, pi04257, pi04258, pi04259, pi04260, pi04261, pi04262, pi04263, pi04264, pi04265, pi04266, pi04267, pi04268, pi04269, pi04270, pi04271, pi04272, pi04273, pi04274, pi04275, pi04276, pi04277, pi04278, pi04279, pi04280, pi04281, pi04282, pi04283, pi04284, pi04285, pi04286, pi04287, pi04288, pi04289, pi04290, pi04291, pi04292, pi04293, pi04294, pi04295, pi04296, pi04297, pi04298, pi04299, pi04300, pi04301, pi04302, pi04303, pi04304, pi04305, pi04306, pi04307, pi04308, pi04309, pi04310, pi04311, pi04312, pi04313, pi04314, pi04315, pi04316, pi04317, pi04318, pi04319, pi04320, pi04321, pi04322, pi04323, pi04324, pi04325, pi04326, pi04327, pi04328, pi04329, pi04330, pi04331, pi04332, pi04333, pi04334, pi04335, pi04336, pi04337, pi04338, pi04339, pi04340, pi04341, pi04342, pi04343, pi04344, pi04345, pi04346, pi04347, pi04348, pi04349, pi04350, pi04351, pi04352, pi04353, pi04354, pi04355, pi04356, pi04357, pi04358, pi04359, pi04360, pi04361, pi04362, pi04363, pi04364, pi04365, pi04366, pi04367, pi04368, pi04369, pi04370, pi04371, pi04372, pi04373, pi04374, pi04375, pi04376, pi04377, pi04378, pi04379, pi04380, pi04381, pi04382, pi04383, pi04384, pi04385, pi04386, pi04387, pi04388, pi04389, pi04390, pi04391, pi04392, pi04393, pi04394, pi04395, pi04396, pi04397, pi04398, pi04399, pi04400, pi04401, pi04402, pi04403, pi04404, pi04405, pi04406, pi04407, pi04408, pi04409, pi04410, pi04411, pi04412, pi04413, pi04414, pi04415, pi04416, pi04417, pi04418, pi04419, pi04420, pi04421, pi04422, pi04423, pi04424, pi04425, pi04426, pi04427, pi04428, pi04429, pi04430, pi04431, pi04432, pi04433, pi04434, pi04435, pi04436, pi04437, pi04438, pi04439, pi04440, pi04441, pi04442, pi04443, pi04444, pi04445, pi04446, pi04447, pi04448, pi04449, pi04450, pi04451, pi04452, pi04453, pi04454, pi04455, pi04456, pi04457, pi04458, pi04459, pi04460, pi04461, pi04462, pi04463, pi04464, pi04465, pi04466, pi04467, pi04468, pi04469, pi04470, pi04471, pi04472, pi04473, pi04474, pi04475, pi04476, pi04477, pi04478, pi04479, pi04480, pi04481, pi04482, pi04483, pi04484, pi04485, pi04486, pi04487, pi04488, pi04489, pi04490, pi04491, pi04492, pi04493, pi04494, pi04495, pi04496, pi04497, pi04498, pi04499, pi04500, pi04501, pi04502, pi04503, pi04504, pi04505, pi04506, pi04507, pi04508, pi04509, pi04510, pi04511, pi04512, pi04513, pi04514, pi04515, pi04516, pi04517, pi04518, pi04519, pi04520, pi04521, pi04522, pi04523, pi04524, pi04525, pi04526, pi04527, pi04528, pi04529, pi04530, pi04531, pi04532, pi04533, pi04534, pi04535, pi04536, pi04537, pi04538, pi04539, pi04540, pi04541, pi04542, pi04543, pi04544, pi04545, pi04546, pi04547, pi04548, pi04549, pi04550, pi04551, pi04552, pi04553, pi04554, pi04555, pi04556, pi04557, pi04558, pi04559, pi04560, pi04561, pi04562, pi04563, pi04564, pi04565, pi04566, pi04567, pi04568, pi04569, pi04570, pi04571, pi04572, pi04573, pi04574, pi04575, pi04576, pi04577, pi04578, pi04579, pi04580, pi04581, pi04582, pi04583, pi04584, pi04585, pi04586, pi04587, pi04588, pi04589, pi04590, pi04591, pi04592, pi04593, pi04594, pi04595, pi04596, pi04597, pi04598, pi04599, pi04600, pi04601, pi04602, pi04603, pi04604, pi04605, pi04606, pi04607, pi04608, pi04609, pi04610, pi04611, pi04612, pi04613, pi04614, pi04615, pi04616, pi04617, pi04618, pi04619, pi04620, pi04621, pi04622, pi04623, pi04624, pi04625, pi04626, pi04627, pi04628, pi04629, pi04630, pi04631, pi04632, pi04633, pi04634, pi04635, pi04636, pi04637, pi04638, pi04639, pi04640, pi04641, pi04642, pi04643, pi04644, pi04645, pi04646, pi04647, pi04648, pi04649, pi04650, pi04651, pi04652, pi04653, pi04654, pi04655, pi04656, pi04657, pi04658, pi04659, pi04660, pi04661, pi04662, pi04663, pi04664, pi04665, pi04666, pi04667, pi04668, pi04669, pi04670, pi04671, pi04672, pi04673, pi04674, pi04675, pi04676, pi04677, pi04678, pi04679, pi04680, pi04681, pi04682, pi04683, pi04684, pi04685, pi04686, pi04687, pi04688, pi04689, pi04690, pi04691, pi04692, pi04693, pi04694, pi04695, pi04696, pi04697, pi04698, pi04699, pi04700, pi04701, pi04702, pi04703, pi04704, pi04705, pi04706, pi04707, pi04708, pi04709, pi04710, pi04711, pi04712, pi04713, pi04714, pi04715, pi04716, pi04717, pi04718, pi04719, pi04720, pi04721, pi04722, pi04723, pi04724, pi04725, pi04726, pi04727, pi04728, pi04729, pi04730, pi04731, pi04732, pi04733, pi04734, pi04735, pi04736, pi04737, pi04738, pi04739, pi04740, pi04741, pi04742, pi04743, pi04744, pi04745, pi04746, pi04747, pi04748, pi04749, pi04750, pi04751, pi04752, pi04753, pi04754, pi04755, pi04756, pi04757, pi04758, pi04759, pi04760, pi04761, pi04762, pi04763, pi04764, pi04765, pi04766, pi04767, pi04768, pi04769, pi04770, pi04771, pi04772, pi04773, pi04774, pi04775, pi04776, pi04777, pi04778, pi04779, pi04780, pi04781, pi04782, pi04783, pi04784, pi04785, pi04786, pi04787, pi04788, pi04789, pi04790, pi04791, pi04792, pi04793, pi04794, pi04795, pi04796, pi04797, pi04798, pi04799, pi04800, pi04801, pi04802, pi04803, pi04804, pi04805, pi04806, pi04807, pi04808, pi04809, pi04810, pi04811, pi04812, pi04813, pi04814, pi04815, pi04816, pi04817, pi04818, pi04819, pi04820, pi04821, pi04822, pi04823, pi04824, pi04825, pi04826, pi04827, pi04828, pi04829, pi04830, pi04831, pi04832, pi04833, pi04834, pi04835, pi04836, pi04837, pi04838, pi04839, pi04840, pi04841, pi04842, pi04843, pi04844, pi04845, pi04846, pi04847, pi04848, pi04849, pi04850, pi04851, pi04852, pi04853, pi04854, pi04855, pi04856, pi04857, pi04858, pi04859, pi04860, pi04861, pi04862, pi04863, pi04864, pi04865, pi04866, pi04867, pi04868, pi04869, pi04870, pi04871, pi04872, pi04873, pi04874, pi04875, pi04876, pi04877, pi04878, pi04879, pi04880, pi04881, pi04882, pi04883, pi04884, pi04885, pi04886, pi04887, pi04888, pi04889, pi04890, pi04891, pi04892, pi04893, pi04894, pi04895, pi04896, pi04897, pi04898, pi04899, pi04900, pi04901, pi04902, pi04903, pi04904, pi04905, pi04906, pi04907, pi04908, pi04909, pi04910, pi04911, pi04912, pi04913, pi04914, pi04915, pi04916, pi04917, pi04918, pi04919, pi04920, pi04921, pi04922, pi04923, pi04924, pi04925, pi04926, pi04927, pi04928, pi04929, pi04930, pi04931, pi04932, pi04933, pi04934, pi04935, pi04936, pi04937, pi04938, pi04939, pi04940, pi04941, pi04942, pi04943, pi04944, pi04945, pi04946, pi04947, pi04948, pi04949, pi04950, pi04951, pi04952, pi04953, pi04954, pi04955, pi04956, pi04957, pi04958, pi04959, pi04960, pi04961, pi04962, pi04963, pi04964, pi04965, pi04966, pi04967, pi04968, pi04969, pi04970, pi04971, pi04972, pi04973, pi04974, pi04975, pi04976, pi04977, pi04978, pi04979, pi04980, pi04981, pi04982, pi04983, pi04984, pi04985, pi04986, pi04987, pi04988, pi04989, pi04990, pi04991, pi04992, pi04993, pi04994, pi04995, pi04996, pi04997, pi04998, pi04999, pi05000, pi05001, pi05002, pi05003, pi05004, pi05005, pi05006, pi05007, pi05008, pi05009, pi05010, pi05011, pi05012, pi05013, pi05014, pi05015, pi05016, pi05017, pi05018, pi05019, pi05020, pi05021, pi05022, pi05023, pi05024, pi05025, pi05026, pi05027, pi05028, pi05029, pi05030, pi05031, pi05032, pi05033, pi05034, pi05035, pi05036, pi05037, pi05038, pi05039, pi05040, pi05041, pi05042, pi05043, pi05044, pi05045, pi05046, pi05047, pi05048, pi05049, pi05050, pi05051, pi05052, pi05053, pi05054, pi05055, pi05056, pi05057, pi05058, pi05059, pi05060, pi05061, pi05062, pi05063, pi05064, pi05065, pi05066, pi05067, pi05068, pi05069, pi05070, pi05071, pi05072, pi05073, pi05074, pi05075, pi05076, pi05077, pi05078, pi05079, pi05080, pi05081, pi05082, pi05083, pi05084, pi05085, pi05086, pi05087, pi05088, pi05089, pi05090, pi05091, pi05092, pi05093, pi05094, pi05095, pi05096, pi05097, pi05098, pi05099, pi05100, pi05101, pi05102, pi05103, pi05104, pi05105, pi05106, pi05107, pi05108, pi05109, pi05110, pi05111, pi05112, pi05113, pi05114, pi05115, pi05116, pi05117, pi05118, pi05119, pi05120, pi05121, pi05122, pi05123, pi05124, pi05125, pi05126, pi05127, pi05128, pi05129, pi05130, pi05131, pi05132, pi05133, pi05134, pi05135, pi05136, pi05137, pi05138, pi05139, pi05140, pi05141, pi05142, pi05143, pi05144, pi05145, pi05146, pi05147, pi05148, pi05149, pi05150, pi05151, pi05152, pi05153, pi05154, pi05155, pi05156, pi05157, pi05158, pi05159, pi05160, pi05161, pi05162, pi05163, pi05164, pi05165, pi05166, pi05167, pi05168, pi05169, pi05170, pi05171, pi05172, pi05173, pi05174, pi05175, pi05176, pi05177, pi05178, pi05179, pi05180, pi05181, pi05182, pi05183, pi05184, pi05185, pi05186, pi05187, pi05188, pi05189, pi05190, pi05191, pi05192, pi05193, pi05194, pi05195, pi05196, pi05197, pi05198, pi05199, pi05200, pi05201, pi05202, pi05203, pi05204, pi05205, pi05206, pi05207, pi05208, pi05209, pi05210, pi05211, pi05212, pi05213, pi05214, pi05215, pi05216, pi05217, pi05218, pi05219, pi05220, pi05221, pi05222, pi05223, pi05224, pi05225, pi05226, pi05227, pi05228, pi05229, pi05230, pi05231, pi05232, pi05233, pi05234, pi05235, pi05236, pi05237, pi05238, pi05239, pi05240, pi05241, pi05242, pi05243, pi05244, pi05245, pi05246, pi05247, pi05248, pi05249, pi05250, pi05251, pi05252, pi05253, pi05254, pi05255, pi05256, pi05257, pi05258, pi05259, pi05260, pi05261, pi05262, pi05263, pi05264, pi05265, pi05266, pi05267, pi05268, pi05269, pi05270, pi05271, pi05272, pi05273, pi05274, pi05275, pi05276, pi05277, pi05278, pi05279, pi05280, pi05281, pi05282, pi05283, pi05284, pi05285, pi05286, pi05287, pi05288, pi05289, pi05290, pi05291, pi05292, pi05293, pi05294, pi05295, pi05296, pi05297, pi05298, pi05299, pi05300, pi05301, pi05302, pi05303, pi05304, pi05305, pi05306, pi05307, pi05308, pi05309, pi05310, pi05311, pi05312, pi05313, pi05314, pi05315, pi05316, pi05317, pi05318, pi05319, pi05320, pi05321, pi05322, pi05323, pi05324, pi05325, pi05326, pi05327, pi05328, pi05329, pi05330, pi05331, pi05332, pi05333, pi05334, pi05335, pi05336, pi05337, pi05338, pi05339, pi05340, pi05341, pi05342, pi05343, pi05344, pi05345, pi05346, pi05347, pi05348, pi05349, pi05350, pi05351, pi05352, pi05353, pi05354, pi05355, pi05356, pi05357, pi05358, pi05359, pi05360, pi05361, pi05362, pi05363, pi05364, pi05365, pi05366, pi05367, pi05368, pi05369, pi05370, pi05371, pi05372, pi05373, pi05374, pi05375, pi05376, pi05377, pi05378, pi05379, pi05380, pi05381, pi05382, pi05383, pi05384, pi05385, pi05386, pi05387, pi05388, pi05389, pi05390, pi05391, pi05392, pi05393, pi05394, pi05395, pi05396, pi05397, pi05398, pi05399, pi05400, pi05401, pi05402, pi05403, pi05404, pi05405, pi05406, pi05407, pi05408, pi05409, pi05410, pi05411, pi05412, pi05413, pi05414, pi05415, pi05416, pi05417, pi05418, pi05419, pi05420, pi05421, pi05422, pi05423, pi05424, pi05425, pi05426, pi05427, pi05428, pi05429, pi05430, pi05431, pi05432, pi05433, pi05434, pi05435, pi05436, pi05437, pi05438, pi05439, pi05440, pi05441, pi05442, pi05443, pi05444, pi05445, pi05446, pi05447, pi05448, pi05449, pi05450, pi05451, pi05452, pi05453, pi05454, pi05455, pi05456, pi05457, pi05458, pi05459, pi05460, pi05461, pi05462, pi05463, pi05464, pi05465, pi05466, pi05467, pi05468, pi05469, pi05470, pi05471, pi05472, pi05473, pi05474, pi05475, pi05476, pi05477, pi05478, pi05479, pi05480, pi05481, pi05482, pi05483, pi05484, pi05485, pi05486, pi05487, pi05488, pi05489, pi05490, pi05491, pi05492, pi05493, pi05494, pi05495, pi05496, pi05497, pi05498, pi05499, pi05500, pi05501, pi05502, pi05503, pi05504, pi05505, pi05506, pi05507, pi05508, pi05509, pi05510, pi05511, pi05512, pi05513, pi05514, pi05515, pi05516, pi05517, pi05518, pi05519, pi05520, pi05521, pi05522, pi05523, pi05524, pi05525, pi05526, pi05527, pi05528, pi05529, pi05530, pi05531, pi05532, pi05533, pi05534, pi05535, pi05536, pi05537, pi05538, pi05539, pi05540, pi05541, pi05542, pi05543, pi05544, pi05545, pi05546, pi05547, pi05548, pi05549, pi05550, pi05551, pi05552, pi05553, pi05554, pi05555, pi05556, pi05557, pi05558, pi05559, pi05560, pi05561, pi05562, pi05563, pi05564, pi05565, pi05566, pi05567, pi05568, pi05569, pi05570, pi05571, pi05572, pi05573, pi05574, pi05575, pi05576, pi05577, pi05578, pi05579, pi05580, pi05581, pi05582, pi05583, pi05584, pi05585, pi05586, pi05587, pi05588, pi05589, pi05590, pi05591, pi05592, pi05593, pi05594, pi05595, pi05596, pi05597, pi05598, pi05599, pi05600, pi05601, pi05602, pi05603, pi05604, pi05605, pi05606, pi05607, pi05608, pi05609, pi05610, pi05611, pi05612, pi05613, pi05614, pi05615, pi05616, pi05617, pi05618, pi05619, pi05620, pi05621, pi05622, pi05623, pi05624, pi05625, pi05626, pi05627, pi05628, pi05629, pi05630, pi05631, pi05632, pi05633, pi05634, pi05635, pi05636, pi05637, pi05638, pi05639, pi05640, pi05641, pi05642, pi05643, pi05644, pi05645, pi05646, pi05647, pi05648, pi05649, pi05650, pi05651, pi05652, pi05653, pi05654, pi05655, pi05656, pi05657, pi05658, pi05659, pi05660, pi05661, pi05662, pi05663, pi05664, pi05665, pi05666, pi05667, pi05668, pi05669, pi05670, pi05671, pi05672, pi05673, pi05674, pi05675, pi05676, pi05677, pi05678, pi05679, pi05680, pi05681, pi05682, pi05683, pi05684, pi05685, pi05686, pi05687, pi05688, pi05689, pi05690, pi05691, pi05692, pi05693, pi05694, pi05695, pi05696, pi05697, pi05698, pi05699, pi05700, pi05701, pi05702, pi05703, pi05704, pi05705, pi05706, pi05707, pi05708, pi05709, pi05710, pi05711, pi05712, pi05713, pi05714, pi05715, pi05716, pi05717, pi05718, pi05719, pi05720, pi05721, pi05722, pi05723, pi05724, pi05725, pi05726, pi05727, pi05728, pi05729, pi05730, pi05731, pi05732, pi05733, pi05734, pi05735, pi05736, pi05737, pi05738, pi05739, pi05740, pi05741, pi05742, pi05743, pi05744, pi05745, pi05746, pi05747, pi05748, pi05749, pi05750, pi05751, pi05752, pi05753, pi05754, pi05755, pi05756, pi05757, pi05758, pi05759, pi05760, pi05761, pi05762, pi05763, pi05764, pi05765, pi05766, pi05767, pi05768, pi05769, pi05770, pi05771, pi05772, pi05773, pi05774, pi05775, pi05776, pi05777, pi05778, pi05779, pi05780, pi05781, pi05782, pi05783, pi05784, pi05785, pi05786, pi05787, pi05788, pi05789, pi05790, pi05791, pi05792, pi05793, pi05794, pi05795, pi05796, pi05797, pi05798, pi05799, pi05800, pi05801, pi05802, pi05803, pi05804, pi05805, pi05806, pi05807, pi05808, pi05809, pi05810, pi05811, pi05812, pi05813, pi05814, pi05815, pi05816, pi05817, pi05818, pi05819, pi05820, pi05821, pi05822, pi05823, pi05824, pi05825, pi05826, pi05827, pi05828, pi05829, pi05830, pi05831, pi05832, pi05833, pi05834, pi05835, pi05836, pi05837, pi05838, pi05839, pi05840, pi05841, pi05842, pi05843, pi05844, pi05845, pi05846, pi05847, pi05848, pi05849, pi05850, pi05851, pi05852, pi05853, pi05854, pi05855, pi05856, pi05857, pi05858, pi05859, pi05860, pi05861, pi05862, pi05863, pi05864, pi05865, pi05866, pi05867, pi05868, pi05869, pi05870, pi05871, pi05872, pi05873, pi05874, pi05875, pi05876, pi05877, pi05878, pi05879, pi05880, pi05881, pi05882, pi05883, pi05884, pi05885, pi05886, pi05887, pi05888, pi05889, pi05890, pi05891, pi05892, pi05893, pi05894, pi05895, pi05896, pi05897, pi05898, pi05899, pi05900, pi05901, pi05902, pi05903, pi05904, pi05905, pi05906, pi05907, pi05908, pi05909, pi05910, pi05911, pi05912, pi05913, pi05914, pi05915, pi05916, pi05917, pi05918, pi05919, pi05920, pi05921, pi05922, pi05923, pi05924, pi05925, pi05926, pi05927, pi05928, pi05929, pi05930, pi05931, pi05932, pi05933, pi05934, pi05935, pi05936, pi05937, pi05938, pi05939, pi05940, pi05941, pi05942, pi05943, pi05944, pi05945, pi05946, pi05947, pi05948, pi05949, pi05950, pi05951, pi05952, pi05953, pi05954, pi05955, pi05956, pi05957, pi05958, pi05959, pi05960, pi05961, pi05962, pi05963, pi05964, pi05965, pi05966, pi05967, pi05968, pi05969, pi05970, pi05971, pi05972, pi05973, pi05974, pi05975, pi05976, pi05977, pi05978, pi05979, pi05980, pi05981, pi05982, pi05983, pi05984, pi05985, pi05986, pi05987, pi05988, pi05989, pi05990, pi05991, pi05992, pi05993, pi05994, pi05995, pi05996, pi05997, pi05998, pi05999, pi06000, pi06001, pi06002, pi06003, pi06004, pi06005, pi06006, pi06007, pi06008, pi06009, pi06010, pi06011, pi06012, pi06013, pi06014, pi06015, pi06016, pi06017, pi06018, pi06019, pi06020, pi06021, pi06022, pi06023, pi06024, pi06025, pi06026, pi06027, pi06028, pi06029, pi06030, pi06031, pi06032, pi06033, pi06034, pi06035, pi06036, pi06037, pi06038, pi06039, pi06040, pi06041, pi06042, pi06043, pi06044, pi06045, pi06046, pi06047, pi06048, pi06049, pi06050, pi06051, pi06052, pi06053, pi06054, pi06055, pi06056, pi06057, pi06058, pi06059, pi06060, pi06061, pi06062, pi06063, pi06064, pi06065, pi06066, pi06067, pi06068, pi06069, pi06070, pi06071, pi06072, pi06073, pi06074, pi06075, pi06076, pi06077, pi06078, pi06079, pi06080, pi06081, pi06082, pi06083, pi06084, pi06085, pi06086, pi06087, pi06088, pi06089, pi06090, pi06091, pi06092, pi06093, pi06094, pi06095, pi06096, pi06097, pi06098, pi06099, pi06100, pi06101, pi06102, pi06103, pi06104, pi06105, pi06106, pi06107, pi06108, pi06109, pi06110, pi06111, pi06112, pi06113, pi06114, pi06115, pi06116, pi06117, pi06118, pi06119, pi06120, pi06121, pi06122, pi06123, pi06124, pi06125, pi06126, pi06127, pi06128, pi06129, pi06130, pi06131, pi06132, pi06133, pi06134, pi06135, pi06136, pi06137, pi06138, pi06139, pi06140, pi06141, pi06142, pi06143, pi06144, pi06145, pi06146, pi06147, pi06148, pi06149, pi06150, pi06151, pi06152, pi06153, pi06154, pi06155, pi06156, pi06157, pi06158, pi06159, pi06160, pi06161, pi06162, pi06163, pi06164, pi06165, pi06166, pi06167, pi06168, pi06169, pi06170, pi06171, pi06172, pi06173, pi06174, pi06175, pi06176, pi06177, pi06178, pi06179, pi06180, pi06181, pi06182, pi06183, pi06184, pi06185, pi06186, pi06187, pi06188, pi06189, pi06190, pi06191, pi06192, pi06193, pi06194, pi06195, pi06196, pi06197, pi06198, pi06199, pi06200, pi06201, pi06202, pi06203, pi06204, pi06205, pi06206, pi06207, pi06208, pi06209, pi06210, pi06211, pi06212, pi06213, pi06214, pi06215, pi06216, pi06217, pi06218, pi06219, pi06220, pi06221, pi06222, pi06223, pi06224, pi06225, pi06226, pi06227, pi06228, pi06229, pi06230, pi06231, pi06232, pi06233, pi06234, pi06235, pi06236, pi06237, pi06238, pi06239, pi06240, pi06241, pi06242, pi06243, pi06244, pi06245, pi06246, pi06247, pi06248, pi06249, pi06250, pi06251, pi06252, pi06253, pi06254, pi06255, pi06256, pi06257, pi06258, pi06259, pi06260, pi06261, pi06262, pi06263, pi06264, pi06265, pi06266, pi06267, pi06268, pi06269, pi06270, pi06271, pi06272, pi06273, pi06274, pi06275, pi06276, pi06277, pi06278, pi06279, pi06280, pi06281, pi06282, pi06283, pi06284, pi06285, pi06286, pi06287, pi06288, pi06289, pi06290, pi06291, pi06292, pi06293, pi06294, pi06295, pi06296, pi06297, pi06298, pi06299, pi06300, pi06301, pi06302, pi06303, pi06304, pi06305, pi06306, pi06307, pi06308, pi06309, pi06310, pi06311, pi06312, pi06313, pi06314, pi06315, pi06316, pi06317, pi06318, pi06319, pi06320, pi06321, pi06322, pi06323, pi06324, pi06325, pi06326, pi06327, pi06328, pi06329, pi06330, pi06331, pi06332, pi06333, pi06334, pi06335, pi06336, pi06337, pi06338, pi06339, pi06340, pi06341, pi06342, pi06343, pi06344, pi06345, pi06346, pi06347, pi06348, pi06349, pi06350, pi06351, pi06352, pi06353, pi06354, pi06355, pi06356, pi06357, pi06358, pi06359, pi06360, pi06361, pi06362, pi06363, pi06364, pi06365, pi06366, pi06367, pi06368, pi06369, pi06370, pi06371, pi06372, pi06373, pi06374, pi06375, pi06376, pi06377, pi06378, pi06379, pi06380, pi06381, pi06382, pi06383, pi06384, pi06385, pi06386, pi06387, pi06388, pi06389, pi06390, pi06391, pi06392, pi06393, pi06394, pi06395, pi06396, pi06397, pi06398, pi06399, pi06400, pi06401, pi06402, pi06403, pi06404, pi06405, pi06406, pi06407, pi06408, pi06409, pi06410, pi06411, pi06412, pi06413, pi06414, pi06415, pi06416, pi06417, pi06418, pi06419, pi06420, pi06421, pi06422, pi06423, pi06424, pi06425, pi06426, pi06427, pi06428, pi06429, pi06430, pi06431, pi06432, pi06433, pi06434, pi06435, pi06436, pi06437, pi06438, pi06439, pi06440, pi06441, pi06442, pi06443, pi06444, pi06445, pi06446, pi06447, pi06448, pi06449, pi06450, pi06451, pi06452, pi06453, pi06454, pi06455, pi06456, pi06457, pi06458, pi06459, pi06460, pi06461, pi06462, pi06463, pi06464, pi06465, pi06466, pi06467, pi06468, pi06469, pi06470, pi06471, pi06472, pi06473, pi06474, pi06475, pi06476, pi06477, pi06478, pi06479, pi06480, pi06481, pi06482, pi06483, pi06484, pi06485, pi06486, pi06487, pi06488, pi06489, pi06490, pi06491, pi06492, pi06493, pi06494, pi06495, pi06496, pi06497, pi06498, pi06499, pi06500, pi06501, pi06502, pi06503, pi06504, pi06505, pi06506, pi06507, pi06508, pi06509, pi06510, pi06511, pi06512, pi06513, pi06514, pi06515, pi06516, pi06517, pi06518, pi06519, pi06520, pi06521, pi06522, pi06523, pi06524, pi06525, pi06526, pi06527, pi06528, pi06529, pi06530, pi06531, pi06532, pi06533, pi06534, pi06535, pi06536, pi06537, pi06538, pi06539, pi06540, pi06541, pi06542, pi06543, pi06544, pi06545, pi06546, pi06547, pi06548, pi06549, pi06550, pi06551, pi06552, pi06553, pi06554, pi06555, pi06556, pi06557, pi06558, pi06559, pi06560, pi06561, pi06562, pi06563, pi06564, pi06565, pi06566, pi06567, pi06568, pi06569, pi06570, pi06571, pi06572, pi06573, pi06574, pi06575, pi06576, pi06577, pi06578, pi06579, pi06580, pi06581, pi06582, pi06583, pi06584, pi06585, pi06586, pi06587, pi06588, pi06589, pi06590, pi06591, pi06592, pi06593, pi06594, pi06595, pi06596, pi06597, pi06598, pi06599, pi06600, pi06601, pi06602, pi06603, pi06604, pi06605, pi06606, pi06607, pi06608, pi06609, pi06610, pi06611, pi06612, pi06613, pi06614, pi06615, pi06616, pi06617, pi06618, pi06619, pi06620, pi06621, pi06622, pi06623, pi06624, pi06625, pi06626, pi06627, pi06628, pi06629, pi06630, pi06631, pi06632, pi06633, pi06634, pi06635, pi06636, pi06637, pi06638, pi06639, pi06640, pi06641, pi06642, pi06643, pi06644, pi06645, pi06646, pi06647, pi06648, pi06649, pi06650, pi06651, pi06652, pi06653, pi06654, pi06655, pi06656, pi06657, pi06658, pi06659, pi06660, pi06661, pi06662, pi06663, pi06664, pi06665, pi06666, pi06667, pi06668, pi06669, pi06670, pi06671, pi06672, pi06673, pi06674, pi06675, pi06676, pi06677, pi06678, pi06679, pi06680, pi06681, pi06682, pi06683, pi06684, pi06685, pi06686, pi06687, pi06688, pi06689, pi06690, pi06691, pi06692, pi06693, pi06694, pi06695, pi06696, pi06697, pi06698, pi06699, pi06700, pi06701, pi06702, pi06703, pi06704, pi06705, pi06706, pi06707, pi06708, pi06709, pi06710, pi06711, pi06712, pi06713, pi06714, pi06715, pi06716, pi06717, pi06718, pi06719, pi06720, pi06721, pi06722, pi06723, pi06724, pi06725, pi06726, pi06727, pi06728, pi06729, pi06730, pi06731, pi06732, pi06733, pi06734, pi06735, pi06736, pi06737, pi06738, pi06739, pi06740, pi06741, pi06742, pi06743, pi06744, pi06745, pi06746, pi06747, pi06748, pi06749, pi06750, pi06751, pi06752, pi06753, pi06754, pi06755, pi06756, pi06757, pi06758, pi06759, pi06760, pi06761, pi06762, pi06763, pi06764, pi06765, pi06766, pi06767, pi06768, pi06769, pi06770, pi06771, pi06772, pi06773, pi06774, pi06775, pi06776, pi06777, pi06778, pi06779, pi06780, pi06781, pi06782, pi06783, pi06784, pi06785, pi06786, pi06787, pi06788, pi06789, pi06790, pi06791, pi06792, pi06793, pi06794, pi06795, pi06796, pi06797, pi06798, pi06799, pi06800, pi06801, pi06802, pi06803, pi06804, pi06805, pi06806, pi06807, pi06808, pi06809, pi06810, pi06811, pi06812, pi06813, pi06814, pi06815, pi06816, pi06817, pi06818, pi06819, pi06820, pi06821, pi06822, pi06823, pi06824, pi06825, pi06826, pi06827, pi06828, pi06829, pi06830, pi06831, pi06832, pi06833, pi06834, pi06835, pi06836, pi06837, pi06838, pi06839, pi06840, pi06841, pi06842, pi06843, pi06844, pi06845, pi06846, pi06847, pi06848, pi06849, pi06850, pi06851, pi06852, pi06853, pi06854, pi06855, pi06856, pi06857, pi06858, pi06859, pi06860, pi06861, pi06862, pi06863, pi06864, pi06865, pi06866, pi06867, pi06868, pi06869, pi06870, pi06871, pi06872, pi06873, pi06874, pi06875, pi06876, pi06877, pi06878, pi06879, pi06880, pi06881, pi06882, pi06883, pi06884, pi06885, pi06886, pi06887, pi06888, pi06889, pi06890, pi06891, pi06892, pi06893, pi06894, pi06895, pi06896, pi06897, pi06898, pi06899, pi06900, pi06901, pi06902, pi06903, pi06904, pi06905, pi06906, pi06907, pi06908, pi06909, pi06910, pi06911, pi06912, pi06913, pi06914, pi06915, pi06916, pi06917, pi06918, pi06919, pi06920, pi06921, pi06922, pi06923, pi06924, pi06925, pi06926, pi06927, pi06928, pi06929, pi06930, pi06931, pi06932, pi06933, pi06934, pi06935, pi06936, pi06937, pi06938, pi06939, pi06940, pi06941, pi06942, pi06943, pi06944, pi06945, pi06946, pi06947, pi06948, pi06949, pi06950, pi06951, pi06952, pi06953, pi06954, pi06955, pi06956, pi06957, pi06958, pi06959, pi06960, pi06961, pi06962, pi06963, pi06964, pi06965, pi06966, pi06967, pi06968, pi06969, pi06970, pi06971, pi06972, pi06973, pi06974, pi06975, pi06976, pi06977, pi06978, pi06979, pi06980, pi06981, pi06982, pi06983, pi06984, pi06985, pi06986, pi06987, pi06988, pi06989, pi06990, pi06991, pi06992, pi06993, pi06994, pi06995, pi06996, pi06997, pi06998, pi06999, pi07000, pi07001, pi07002, pi07003, pi07004, pi07005, pi07006, pi07007, pi07008, pi07009, pi07010, pi07011, pi07012, pi07013, pi07014, pi07015, pi07016, pi07017, pi07018, pi07019, pi07020, pi07021, pi07022, pi07023, pi07024, pi07025, pi07026, pi07027, pi07028, pi07029, pi07030, pi07031, pi07032, pi07033, pi07034, pi07035, pi07036, pi07037, pi07038, pi07039, pi07040, pi07041, pi07042, pi07043, pi07044, pi07045, pi07046, pi07047, pi07048, pi07049, pi07050, pi07051, pi07052, pi07053, pi07054, pi07055, pi07056, pi07057, pi07058, pi07059, pi07060, pi07061, pi07062, pi07063, pi07064, pi07065, pi07066, pi07067, pi07068, pi07069, pi07070, pi07071, pi07072, pi07073, pi07074, pi07075, pi07076, pi07077, pi07078, pi07079, pi07080, pi07081, pi07082, pi07083, pi07084, pi07085, pi07086, pi07087, pi07088, pi07089, pi07090, pi07091, pi07092, pi07093, pi07094, pi07095, pi07096, pi07097, pi07098, pi07099, pi07100, pi07101, pi07102, pi07103, pi07104, pi07105, pi07106, pi07107, pi07108, pi07109, pi07110, pi07111, pi07112, pi07113, pi07114, pi07115, pi07116, pi07117, pi07118, pi07119, pi07120, pi07121, pi07122, pi07123, pi07124, pi07125, pi07126, pi07127, pi07128, pi07129, pi07130, pi07131, pi07132, pi07133, pi07134, pi07135, pi07136, pi07137, pi07138, pi07139, pi07140, pi07141, pi07142, pi07143, pi07144, pi07145, pi07146, pi07147, pi07148, pi07149, pi07150, pi07151, pi07152, pi07153, pi07154, pi07155, pi07156, pi07157, pi07158, pi07159, pi07160, pi07161, pi07162, pi07163, pi07164, pi07165, pi07166, pi07167, pi07168, pi07169, pi07170, pi07171, pi07172, pi07173, pi07174, pi07175, pi07176, pi07177, pi07178, pi07179, pi07180, pi07181, pi07182, pi07183, pi07184, pi07185, pi07186, pi07187, pi07188, pi07189, pi07190, pi07191, pi07192, pi07193, pi07194, pi07195, pi07196, pi07197, pi07198, pi07199, pi07200, pi07201, pi07202, pi07203, pi07204, pi07205, pi07206, pi07207, pi07208, pi07209, pi07210, pi07211, pi07212, pi07213, pi07214, pi07215, pi07216, pi07217, pi07218, pi07219, pi07220, pi07221, pi07222, pi07223, pi07224, pi07225, pi07226, pi07227, pi07228, pi07229, pi07230, pi07231, pi07232, pi07233, pi07234, pi07235, pi07236, pi07237, pi07238, pi07239, pi07240, pi07241, pi07242, pi07243, pi07244, pi07245, pi07246, pi07247, pi07248, pi07249, pi07250, pi07251, pi07252, pi07253, pi07254, pi07255, pi07256, pi07257, pi07258, pi07259, pi07260, pi07261, pi07262, pi07263, pi07264, pi07265, pi07266, pi07267, pi07268, pi07269, pi07270, pi07271, pi07272, pi07273, pi07274, pi07275, pi07276, pi07277, pi07278, pi07279, pi07280, pi07281, pi07282, pi07283, pi07284, pi07285, pi07286, pi07287, pi07288, pi07289, pi07290, pi07291, pi07292, pi07293, pi07294, pi07295, pi07296, pi07297, pi07298, pi07299, pi07300, pi07301, pi07302, pi07303, pi07304, pi07305, pi07306, pi07307, pi07308, pi07309, pi07310, pi07311, pi07312, pi07313, pi07314, pi07315, pi07316, pi07317, pi07318, pi07319, pi07320, pi07321, pi07322, pi07323, pi07324, pi07325, pi07326, pi07327, pi07328, pi07329, pi07330, pi07331, pi07332, pi07333, pi07334, pi07335, pi07336, pi07337, pi07338, pi07339, pi07340, pi07341, pi07342, pi07343, pi07344, pi07345, pi07346, pi07347, pi07348, pi07349, pi07350, pi07351, pi07352, pi07353, pi07354, pi07355, pi07356, pi07357, pi07358, pi07359, pi07360, pi07361, pi07362, pi07363, pi07364, pi07365, pi07366, pi07367, pi07368, pi07369, pi07370, pi07371, pi07372, pi07373, pi07374, pi07375, pi07376, pi07377, pi07378, pi07379, pi07380, pi07381, pi07382, pi07383, pi07384, pi07385, pi07386, pi07387, pi07388, pi07389, pi07390, pi07391, pi07392, pi07393, pi07394, pi07395, pi07396, pi07397, pi07398, pi07399, pi07400, pi07401, pi07402, pi07403, pi07404, pi07405, pi07406, pi07407, pi07408, pi07409, pi07410, pi07411, pi07412, pi07413, pi07414, pi07415, pi07416, pi07417, pi07418, pi07419, pi07420, pi07421, pi07422, pi07423, pi07424, pi07425, pi07426, pi07427, pi07428, pi07429, pi07430, pi07431, pi07432, pi07433, pi07434, pi07435, pi07436, pi07437, pi07438, pi07439, pi07440, pi07441, pi07442, pi07443, pi07444, pi07445, pi07446, pi07447, pi07448, pi07449, pi07450, pi07451, pi07452, pi07453, pi07454, pi07455, pi07456, pi07457, pi07458, pi07459, pi07460, pi07461, pi07462, pi07463, pi07464, pi07465, pi07466, pi07467, pi07468, pi07469, pi07470, pi07471, pi07472, pi07473, pi07474, pi07475, pi07476, pi07477, pi07478, pi07479, pi07480, pi07481, pi07482, pi07483, pi07484, pi07485, pi07486, pi07487, pi07488, pi07489, pi07490, pi07491, pi07492, pi07493, pi07494, pi07495, pi07496, pi07497, pi07498, pi07499, pi07500, pi07501, pi07502, pi07503, pi07504, pi07505, pi07506, pi07507, pi07508, pi07509, pi07510, pi07511, pi07512, pi07513, pi07514, pi07515, pi07516, pi07517, pi07518, pi07519, pi07520, pi07521, pi07522, pi07523, pi07524, pi07525, pi07526, pi07527, pi07528, pi07529, pi07530, pi07531, pi07532, pi07533, pi07534, pi07535, pi07536, pi07537, pi07538, pi07539, pi07540, pi07541, pi07542, pi07543, pi07544, pi07545, pi07546, pi07547, pi07548, pi07549, pi07550, pi07551, pi07552, pi07553, pi07554, pi07555, pi07556, pi07557, pi07558, pi07559, pi07560, pi07561, pi07562, pi07563, pi07564, pi07565, pi07566, pi07567, pi07568, pi07569, pi07570, pi07571, pi07572, pi07573, pi07574, pi07575, pi07576, pi07577, pi07578, pi07579, pi07580, pi07581, pi07582, pi07583, pi07584, pi07585, pi07586, pi07587, pi07588, pi07589, pi07590, pi07591, pi07592, pi07593, pi07594, pi07595, pi07596, pi07597, pi07598, pi07599, pi07600, pi07601, pi07602, pi07603, pi07604, pi07605, pi07606, pi07607, pi07608, pi07609, pi07610, pi07611, pi07612, pi07613, pi07614, pi07615, pi07616, pi07617, pi07618, pi07619, pi07620, pi07621, pi07622, pi07623, pi07624, pi07625, pi07626, pi07627, pi07628, pi07629, pi07630, pi07631, pi07632, pi07633, pi07634, pi07635, pi07636, pi07637, pi07638, pi07639, pi07640, pi07641, pi07642, pi07643, pi07644, pi07645, pi07646, pi07647, pi07648, pi07649, pi07650, pi07651, pi07652, pi07653, pi07654, pi07655, pi07656, pi07657, pi07658, pi07659, pi07660, pi07661, pi07662, pi07663, pi07664, pi07665, pi07666, pi07667, pi07668, pi07669, pi07670, pi07671, pi07672, pi07673, pi07674, pi07675, pi07676, pi07677, pi07678, pi07679, pi07680, pi07681, pi07682, pi07683, pi07684, pi07685, pi07686, pi07687, pi07688, pi07689, pi07690, pi07691, pi07692, pi07693, pi07694, pi07695, pi07696, pi07697, pi07698, pi07699, pi07700, pi07701, pi07702, pi07703, pi07704, pi07705, pi07706, pi07707, pi07708, pi07709, pi07710, pi07711, pi07712, pi07713, pi07714, pi07715, pi07716, pi07717, pi07718, pi07719, pi07720, pi07721, pi07722, pi07723, pi07724, pi07725, pi07726, pi07727, pi07728, pi07729, pi07730, pi07731, pi07732, pi07733, pi07734, pi07735, pi07736, pi07737, pi07738, pi07739, pi07740, pi07741, pi07742, pi07743, pi07744, pi07745, pi07746, pi07747, pi07748, pi07749, pi07750, pi07751, pi07752, pi07753, pi07754, pi07755, pi07756, pi07757, pi07758, pi07759, pi07760, pi07761, pi07762, pi07763, pi07764, pi07765, pi07766, pi07767, pi07768, pi07769, pi07770, pi07771, pi07772, pi07773, pi07774, pi07775, pi07776, pi07777, pi07778, pi07779, pi07780, pi07781, pi07782, pi07783, pi07784, pi07785, pi07786, pi07787, pi07788, pi07789, pi07790, pi07791, pi07792, pi07793, pi07794, pi07795, pi07796, pi07797, pi07798, pi07799, pi07800, pi07801, pi07802, pi07803, pi07804, pi07805, pi07806, pi07807, pi07808, pi07809, pi07810, pi07811, pi07812, pi07813, pi07814, pi07815, pi07816, pi07817, pi07818, pi07819, pi07820, pi07821, pi07822, pi07823, pi07824, pi07825, pi07826, pi07827, pi07828, pi07829, pi07830, pi07831, pi07832, pi07833, pi07834, pi07835, pi07836, pi07837, pi07838, pi07839, pi07840, pi07841, pi07842, pi07843, pi07844, pi07845, pi07846, pi07847, pi07848, pi07849, pi07850, pi07851, pi07852, pi07853, pi07854, pi07855, pi07856, pi07857, pi07858, pi07859, pi07860, pi07861, pi07862, pi07863, pi07864, pi07865, pi07866, pi07867, pi07868, pi07869, pi07870, pi07871, pi07872, pi07873, pi07874, pi07875, pi07876, pi07877, pi07878, pi07879, pi07880, pi07881, pi07882, pi07883, pi07884, pi07885, pi07886, pi07887, pi07888, pi07889, pi07890, pi07891, pi07892, pi07893, pi07894, pi07895, pi07896, pi07897, pi07898, pi07899, pi07900, pi07901, pi07902, pi07903, pi07904, pi07905, pi07906, pi07907, pi07908, pi07909, pi07910, pi07911, pi07912, pi07913, pi07914, pi07915, pi07916, pi07917, pi07918, pi07919, pi07920, pi07921, pi07922, pi07923, pi07924, pi07925, pi07926, pi07927, pi07928, pi07929, pi07930, pi07931, pi07932, pi07933, pi07934, pi07935, pi07936, pi07937, pi07938, pi07939, pi07940, pi07941, pi07942, pi07943, pi07944, pi07945, pi07946, pi07947, pi07948, pi07949, pi07950, pi07951, pi07952, pi07953, pi07954, pi07955, pi07956, pi07957, pi07958, pi07959, pi07960, pi07961, pi07962, pi07963, pi07964, pi07965, pi07966, pi07967, pi07968, pi07969, pi07970, pi07971, pi07972, pi07973, pi07974, pi07975, pi07976, pi07977, pi07978, pi07979, pi07980, pi07981, pi07982, pi07983, pi07984, pi07985, pi07986, pi07987, pi07988, pi07989, pi07990, pi07991, pi07992, pi07993, pi07994, pi07995, pi07996, pi07997, pi07998, pi07999, pi08000, pi08001, pi08002, pi08003, pi08004, pi08005, pi08006, pi08007, pi08008, pi08009, pi08010, pi08011, pi08012, pi08013, pi08014, pi08015, pi08016, pi08017, pi08018, pi08019, pi08020, pi08021, pi08022, pi08023, pi08024, pi08025, pi08026, pi08027, pi08028, pi08029, pi08030, pi08031, pi08032, pi08033, pi08034, pi08035, pi08036, pi08037, pi08038, pi08039, pi08040, pi08041, pi08042, pi08043, pi08044, pi08045, pi08046, pi08047, pi08048, pi08049, pi08050, pi08051, pi08052, pi08053, pi08054, pi08055, pi08056, pi08057, pi08058, pi08059, pi08060, pi08061, pi08062, pi08063, pi08064, pi08065, pi08066, pi08067, pi08068, pi08069, pi08070, pi08071, pi08072, pi08073, pi08074, pi08075, pi08076, pi08077, pi08078, pi08079, pi08080, pi08081, pi08082, pi08083, pi08084, pi08085, pi08086, pi08087, pi08088, pi08089, pi08090, pi08091, pi08092, pi08093, pi08094, pi08095, pi08096, pi08097, pi08098, pi08099, pi08100, pi08101, pi08102, pi08103, pi08104, pi08105, pi08106, pi08107, pi08108, pi08109, pi08110, pi08111, pi08112, pi08113, pi08114, pi08115, pi08116, pi08117, pi08118, pi08119, pi08120, pi08121, pi08122, pi08123, pi08124, pi08125, pi08126, pi08127, pi08128, pi08129, pi08130, pi08131, pi08132, pi08133, pi08134, pi08135, pi08136, pi08137, pi08138, pi08139, pi08140, pi08141, pi08142, pi08143, pi08144, pi08145, pi08146, pi08147, pi08148, pi08149, pi08150, pi08151, pi08152, pi08153, pi08154, pi08155, pi08156, pi08157, pi08158, pi08159, pi08160, pi08161, pi08162, pi08163, pi08164, pi08165, pi08166, pi08167, pi08168, pi08169, pi08170, pi08171, pi08172, pi08173, pi08174, pi08175, pi08176, pi08177, pi08178, pi08179, pi08180, pi08181, pi08182, pi08183, pi08184, pi08185, pi08186, pi08187, pi08188, pi08189, pi08190, pi08191, pi08192, pi08193, pi08194, pi08195, pi08196, pi08197, pi08198, pi08199, pi08200, pi08201, pi08202, pi08203, pi08204, pi08205, pi08206, pi08207, pi08208, pi08209, pi08210, pi08211, pi08212, pi08213, pi08214, pi08215, pi08216, pi08217, pi08218, pi08219, pi08220, pi08221, pi08222, pi08223, pi08224, pi08225, pi08226, pi08227, pi08228, pi08229, pi08230, pi08231, pi08232, pi08233, pi08234, pi08235, pi08236, pi08237, pi08238, pi08239, pi08240, pi08241, pi08242, pi08243, pi08244, pi08245, pi08246, pi08247, pi08248, pi08249, pi08250, pi08251, pi08252, pi08253, pi08254, pi08255, pi08256, pi08257, pi08258, pi08259, pi08260, pi08261, pi08262, pi08263, pi08264, pi08265, pi08266, pi08267, pi08268, pi08269, pi08270, pi08271, pi08272, pi08273, pi08274, pi08275, pi08276, pi08277, pi08278, pi08279, pi08280, pi08281, pi08282, pi08283, pi08284, pi08285, pi08286, pi08287, pi08288, pi08289, pi08290, pi08291, pi08292, pi08293, pi08294, pi08295, pi08296, pi08297, pi08298, pi08299, pi08300, pi08301, pi08302, pi08303, pi08304, pi08305, pi08306, pi08307, pi08308, pi08309, pi08310, pi08311, pi08312, pi08313, pi08314, pi08315, pi08316, pi08317, pi08318, pi08319, pi08320, pi08321, pi08322, pi08323, pi08324, pi08325, pi08326, pi08327, pi08328, pi08329, pi08330, pi08331, pi08332, pi08333, pi08334, pi08335, pi08336, pi08337, pi08338, pi08339, pi08340, pi08341, pi08342, pi08343, pi08344, pi08345, pi08346, pi08347, pi08348, pi08349, pi08350, pi08351, pi08352, pi08353, pi08354, pi08355, pi08356, pi08357, pi08358, pi08359, pi08360, pi08361, pi08362, pi08363, pi08364, pi08365, pi08366, pi08367, pi08368, pi08369, pi08370, pi08371, pi08372, pi08373, pi08374, pi08375, pi08376, pi08377, pi08378, pi08379, pi08380, pi08381, pi08382, pi08383, pi08384, pi08385, pi08386, pi08387, pi08388, pi08389, pi08390, pi08391, pi08392, pi08393, pi08394, pi08395, pi08396, pi08397, pi08398, pi08399, pi08400, pi08401, pi08402, pi08403, pi08404, pi08405, pi08406, pi08407, pi08408, pi08409, pi08410, pi08411, pi08412, pi08413, pi08414, pi08415, pi08416, pi08417, pi08418, pi08419, pi08420, pi08421, pi08422, pi08423, pi08424, pi08425, pi08426, pi08427, pi08428, pi08429, pi08430, pi08431, pi08432, pi08433, pi08434, pi08435, pi08436, pi08437, pi08438, pi08439, pi08440, pi08441, pi08442, pi08443, pi08444, pi08445, pi08446, pi08447, pi08448, pi08449, pi08450, pi08451, pi08452, pi08453, pi08454, pi08455, pi08456, pi08457, pi08458, pi08459, pi08460, pi08461, pi08462, pi08463, pi08464, pi08465, pi08466, pi08467, pi08468, pi08469, pi08470, pi08471, pi08472, pi08473, pi08474, pi08475, pi08476, pi08477, pi08478, pi08479, pi08480, pi08481, pi08482, pi08483, pi08484, pi08485, pi08486, pi08487, pi08488, pi08489, pi08490, pi08491, pi08492, pi08493, pi08494, pi08495, pi08496, pi08497, pi08498, pi08499, pi08500, pi08501, pi08502, pi08503, pi08504, pi08505, pi08506, pi08507, pi08508, pi08509, pi08510, pi08511, pi08512, pi08513, pi08514, pi08515, pi08516, pi08517, pi08518, pi08519, pi08520, pi08521, pi08522, pi08523, pi08524, pi08525, pi08526, pi08527, pi08528, pi08529, pi08530, pi08531, pi08532, pi08533, pi08534, pi08535, pi08536, pi08537, pi08538, pi08539, pi08540, pi08541, pi08542, pi08543, pi08544, pi08545, pi08546, pi08547, pi08548, pi08549, pi08550, pi08551, pi08552, pi08553, pi08554, pi08555, pi08556, pi08557, pi08558, pi08559, pi08560, pi08561, pi08562, pi08563, pi08564, pi08565, pi08566, pi08567, pi08568, pi08569, pi08570, pi08571, pi08572, pi08573, pi08574, pi08575, pi08576, pi08577, pi08578, pi08579, pi08580, pi08581, pi08582, pi08583, pi08584, pi08585, pi08586, pi08587, pi08588, pi08589, pi08590, pi08591, pi08592, pi08593, pi08594, pi08595, pi08596, pi08597, pi08598, pi08599, pi08600, pi08601, pi08602, pi08603, pi08604, pi08605, pi08606, pi08607, pi08608, pi08609, pi08610, pi08611, pi08612, pi08613, pi08614, pi08615, pi08616, pi08617, pi08618, pi08619, pi08620, pi08621, pi08622, pi08623, pi08624, pi08625, pi08626, pi08627, pi08628, pi08629, pi08630, pi08631, pi08632, pi08633, pi08634, pi08635, pi08636, pi08637, pi08638, pi08639, pi08640, pi08641, pi08642, pi08643, pi08644, pi08645, pi08646, pi08647, pi08648, pi08649, pi08650, pi08651, pi08652, pi08653, pi08654, pi08655, pi08656, pi08657, pi08658, pi08659, pi08660, pi08661, pi08662, pi08663, pi08664, pi08665, pi08666, pi08667, pi08668, pi08669, pi08670, pi08671, pi08672, pi08673, pi08674, pi08675, pi08676, pi08677, pi08678, pi08679, pi08680, pi08681, pi08682, pi08683, pi08684, pi08685, pi08686, pi08687, pi08688, pi08689, pi08690, pi08691, pi08692, pi08693, pi08694, pi08695, pi08696, pi08697, pi08698, pi08699, pi08700, pi08701, pi08702, pi08703, pi08704, pi08705, pi08706, pi08707, pi08708, pi08709, pi08710, pi08711, pi08712, pi08713, pi08714, pi08715, pi08716, pi08717, pi08718, pi08719, pi08720, pi08721, pi08722, pi08723, pi08724, pi08725, pi08726, pi08727, pi08728, pi08729, pi08730, pi08731, pi08732, pi08733, pi08734, pi08735, pi08736, pi08737, pi08738, pi08739, pi08740, pi08741, pi08742, pi08743, pi08744, pi08745, pi08746, pi08747, pi08748, pi08749, pi08750, pi08751, pi08752, pi08753, pi08754, pi08755, pi08756, pi08757, pi08758, pi08759, pi08760, pi08761, pi08762, pi08763, pi08764, pi08765, pi08766, pi08767, pi08768, pi08769, pi08770, pi08771, pi08772, pi08773, pi08774, pi08775, pi08776, pi08777, pi08778, pi08779, pi08780, pi08781, pi08782, pi08783, pi08784, pi08785, pi08786, pi08787, pi08788, pi08789, pi08790, pi08791, pi08792, pi08793, pi08794, pi08795, pi08796, pi08797, pi08798, pi08799, pi08800, pi08801, pi08802, pi08803, pi08804, pi08805, pi08806, pi08807, pi08808, pi08809, pi08810, pi08811, pi08812, pi08813, pi08814, pi08815, pi08816, pi08817, pi08818, pi08819, pi08820, pi08821, pi08822, pi08823, pi08824, pi08825, pi08826, pi08827, pi08828, pi08829, pi08830, pi08831, pi08832, pi08833, pi08834, pi08835, pi08836, pi08837, pi08838, pi08839, pi08840, pi08841, pi08842, pi08843, pi08844, pi08845, pi08846, pi08847, pi08848, pi08849, pi08850, pi08851, pi08852, pi08853, pi08854, pi08855, pi08856, pi08857, pi08858, pi08859, pi08860, pi08861, pi08862, pi08863, pi08864, pi08865, pi08866, pi08867, pi08868, pi08869, pi08870, pi08871, pi08872, pi08873, pi08874, pi08875, pi08876, pi08877, pi08878, pi08879, pi08880, pi08881, pi08882, pi08883, pi08884, pi08885, pi08886, pi08887, pi08888, pi08889, pi08890, pi08891, pi08892, pi08893, pi08894, pi08895, pi08896, pi08897, pi08898, pi08899, pi08900, pi08901, pi08902, pi08903, pi08904, pi08905, pi08906, pi08907, pi08908, pi08909, pi08910, pi08911, pi08912, pi08913, pi08914, pi08915, pi08916, pi08917, pi08918, pi08919, pi08920, pi08921, pi08922, pi08923, pi08924, pi08925, pi08926, pi08927, pi08928, pi08929, pi08930, pi08931, pi08932, pi08933, pi08934, pi08935, pi08936, pi08937, pi08938, pi08939, pi08940, pi08941, pi08942, pi08943, pi08944, pi08945, pi08946, pi08947, pi08948, pi08949, pi08950, pi08951, pi08952, pi08953, pi08954, pi08955, pi08956, pi08957, pi08958, pi08959, pi08960, pi08961, pi08962, pi08963, pi08964, pi08965, pi08966, pi08967, pi08968, pi08969, pi08970, pi08971, pi08972, pi08973, pi08974, pi08975, pi08976, pi08977, pi08978, pi08979, pi08980, pi08981, pi08982, pi08983, pi08984, pi08985, pi08986, pi08987, pi08988, pi08989, pi08990, pi08991, pi08992, pi08993, pi08994, pi08995, pi08996, pi08997, pi08998, pi08999, pi09000, pi09001, pi09002, pi09003, pi09004, pi09005, pi09006, pi09007, pi09008, pi09009, pi09010, pi09011, pi09012, pi09013, pi09014, pi09015, pi09016, pi09017, pi09018, pi09019, pi09020, pi09021, pi09022, pi09023, pi09024, pi09025, pi09026, pi09027, pi09028, pi09029, pi09030, pi09031, pi09032, pi09033, pi09034, pi09035, pi09036, pi09037, pi09038, pi09039, pi09040, pi09041, pi09042, pi09043, pi09044, pi09045, pi09046, pi09047, pi09048, pi09049, pi09050, pi09051, pi09052, pi09053, pi09054, pi09055, pi09056, pi09057, pi09058, pi09059, pi09060, pi09061, pi09062, pi09063, pi09064, pi09065, pi09066, pi09067, pi09068, pi09069, pi09070, pi09071, pi09072, pi09073, pi09074, pi09075, pi09076, pi09077, pi09078, pi09079, pi09080, pi09081, pi09082, pi09083, pi09084, pi09085, pi09086, pi09087, pi09088, pi09089, pi09090, pi09091, pi09092, pi09093, pi09094, pi09095, pi09096, pi09097, pi09098, pi09099, pi09100, pi09101, pi09102, pi09103, pi09104, pi09105, pi09106, pi09107, pi09108, pi09109, pi09110, pi09111, pi09112, pi09113, pi09114, pi09115, pi09116, pi09117, pi09118, pi09119, pi09120, pi09121, pi09122, pi09123, pi09124, pi09125, pi09126, pi09127, pi09128, pi09129, pi09130, pi09131, pi09132, pi09133, pi09134, pi09135, pi09136, pi09137, pi09138, pi09139, pi09140, pi09141, pi09142, pi09143, pi09144, pi09145, pi09146, pi09147, pi09148, pi09149, pi09150, pi09151, pi09152, pi09153, pi09154, pi09155, pi09156, pi09157, pi09158, pi09159, pi09160, pi09161, pi09162, pi09163, pi09164, pi09165, pi09166, pi09167, pi09168, pi09169, pi09170, pi09171, pi09172, pi09173, pi09174, pi09175, pi09176, pi09177, pi09178, pi09179, pi09180, pi09181, pi09182, pi09183, pi09184, pi09185, pi09186, pi09187, pi09188, pi09189, pi09190, pi09191, pi09192, pi09193, pi09194, pi09195, pi09196, pi09197, pi09198, pi09199, pi09200, pi09201, pi09202, pi09203, pi09204, pi09205, pi09206, pi09207, pi09208, pi09209, pi09210, pi09211, pi09212, pi09213, pi09214, pi09215, pi09216, pi09217, pi09218, pi09219, pi09220, pi09221, pi09222, pi09223, pi09224, pi09225, pi09226, pi09227, pi09228, pi09229, pi09230, pi09231, pi09232, pi09233, pi09234, pi09235, pi09236, pi09237, pi09238, pi09239, pi09240, pi09241, pi09242, pi09243, pi09244, pi09245, pi09246, pi09247, pi09248, pi09249, pi09250, pi09251, pi09252, pi09253, pi09254, pi09255, pi09256, pi09257, pi09258, pi09259, pi09260, pi09261, pi09262, pi09263, pi09264, pi09265, pi09266, pi09267, pi09268, pi09269, pi09270, pi09271, pi09272, pi09273, pi09274, pi09275, pi09276, pi09277, pi09278, pi09279, pi09280, pi09281, pi09282, pi09283, pi09284, pi09285, pi09286, pi09287, pi09288, pi09289, pi09290, pi09291, pi09292, pi09293, pi09294, pi09295, pi09296, pi09297, pi09298, pi09299, pi09300, pi09301, pi09302, pi09303, pi09304, pi09305, pi09306, pi09307, pi09308, pi09309, pi09310, pi09311, pi09312, pi09313, pi09314, pi09315, pi09316, pi09317, pi09318, pi09319, pi09320, pi09321, pi09322, pi09323, pi09324, pi09325, pi09326, pi09327, pi09328, pi09329, pi09330, pi09331, pi09332, pi09333, pi09334, pi09335, pi09336, pi09337, pi09338, pi09339, pi09340, pi09341, pi09342, pi09343, pi09344, pi09345, pi09346, pi09347, pi09348, pi09349, pi09350, pi09351, pi09352, pi09353, pi09354, pi09355, pi09356, pi09357, pi09358, pi09359, pi09360, pi09361, pi09362, pi09363, pi09364, pi09365, pi09366, pi09367, pi09368, pi09369, pi09370, pi09371, pi09372, pi09373, pi09374, pi09375, pi09376, pi09377, pi09378, pi09379, pi09380, pi09381, pi09382, pi09383, pi09384, pi09385, pi09386, pi09387, pi09388, pi09389, pi09390, pi09391, pi09392, pi09393, pi09394, pi09395, pi09396, pi09397, pi09398, pi09399, pi09400, pi09401, pi09402, pi09403, pi09404, pi09405, pi09406, pi09407, pi09408, pi09409, pi09410, pi09411, pi09412, pi09413, pi09414, pi09415, pi09416, pi09417, pi09418, pi09419, pi09420, pi09421, pi09422, pi09423, pi09424, pi09425, pi09426, pi09427, pi09428, pi09429, pi09430, pi09431, pi09432, pi09433, pi09434, pi09435, pi09436, pi09437, pi09438, pi09439, pi09440, pi09441, pi09442, pi09443, pi09444, pi09445, pi09446, pi09447, pi09448, pi09449, pi09450, pi09451, pi09452, pi09453, pi09454, pi09455, pi09456, pi09457, pi09458, pi09459, pi09460, pi09461, pi09462, pi09463, pi09464, pi09465, pi09466, pi09467, pi09468, pi09469, pi09470, pi09471, pi09472, pi09473, pi09474, pi09475, pi09476, pi09477, pi09478, pi09479, pi09480, pi09481, pi09482, pi09483, pi09484, pi09485, pi09486, pi09487, pi09488, pi09489, pi09490, pi09491, pi09492, pi09493, pi09494, pi09495, pi09496, pi09497, pi09498, pi09499, pi09500, pi09501, pi09502, pi09503, pi09504, pi09505, pi09506, pi09507, pi09508, pi09509, pi09510, pi09511, pi09512, pi09513, pi09514, pi09515, pi09516, pi09517, pi09518, pi09519, pi09520, pi09521, pi09522, pi09523, pi09524, pi09525, pi09526, pi09527, pi09528, pi09529, pi09530, pi09531, pi09532, pi09533, pi09534, pi09535, pi09536, pi09537, pi09538, pi09539, pi09540, pi09541, pi09542, pi09543, pi09544, pi09545, pi09546, pi09547, pi09548, pi09549, pi09550, pi09551, pi09552, pi09553, pi09554, pi09555, pi09556, pi09557, pi09558, pi09559, pi09560, pi09561, pi09562, pi09563, pi09564, pi09565, pi09566, pi09567, pi09568, pi09569, pi09570, pi09571, pi09572, pi09573, pi09574, pi09575, pi09576, pi09577, pi09578, pi09579, pi09580, pi09581, pi09582, pi09583, pi09584, pi09585, pi09586, pi09587, pi09588, pi09589, pi09590, pi09591, pi09592, pi09593, pi09594, pi09595, pi09596, pi09597, pi09598, pi09599, pi09600, pi09601, pi09602, pi09603, pi09604, pi09605, pi09606, pi09607, pi09608, pi09609, pi09610, pi09611, pi09612, pi09613, pi09614, pi09615, pi09616, pi09617, pi09618, pi09619, pi09620, pi09621, pi09622, pi09623, pi09624, pi09625, pi09626, pi09627, pi09628, pi09629, pi09630, pi09631, pi09632, pi09633, pi09634, pi09635, pi09636, pi09637, pi09638, pi09639, pi09640, pi09641, pi09642, pi09643, pi09644, pi09645, pi09646, pi09647, pi09648, pi09649, pi09650, pi09651, pi09652, pi09653, pi09654, pi09655, pi09656, pi09657, pi09658, pi09659, pi09660, pi09661, pi09662, pi09663, pi09664, pi09665, pi09666, pi09667, pi09668, pi09669, pi09670, pi09671, pi09672, pi09673, pi09674, pi09675, pi09676, pi09677, pi09678, pi09679, pi09680, pi09681, pi09682, pi09683, pi09684, pi09685, pi09686, pi09687, pi09688, pi09689, pi09690, pi09691, pi09692, pi09693, pi09694, pi09695, pi09696, pi09697, pi09698, pi09699, pi09700, pi09701, pi09702, pi09703, pi09704, pi09705, pi09706, pi09707, pi09708, pi09709, pi09710, pi09711, pi09712, pi09713, pi09714, pi09715, pi09716, pi09717, pi09718, pi09719, pi09720, pi09721, pi09722, pi09723, pi09724, pi09725, pi09726, pi09727, pi09728, pi09729, pi09730, pi09731, pi09732, pi09733, pi09734, pi09735, pi09736, pi09737, pi09738, pi09739, pi09740, pi09741, pi09742, pi09743, pi09744, pi09745, pi09746, pi09747, pi09748, pi09749, pi09750, pi09751, pi09752, pi09753, pi09754, pi09755, pi09756, pi09757, pi09758, pi09759, pi09760, pi09761, pi09762, pi09763, pi09764, pi09765, pi09766, pi09767, pi09768, pi09769, pi09770, pi09771, pi09772, pi09773, pi09774, pi09775, pi09776, pi09777, pi09778, pi09779, pi09780, pi09781, pi09782, pi09783, pi09784, pi09785, pi09786, pi09787, pi09788, pi09789, pi09790, pi09791, pi09792, pi09793, pi09794, pi09795, pi09796, pi09797, pi09798, pi09799, pi09800, pi09801, pi09802, pi09803, pi09804, pi09805, pi09806, pi09807, pi09808, pi09809, pi09810, pi09811, pi09812, pi09813, pi09814, pi09815, pi09816, pi09817, pi09818, pi09819, pi09820, pi09821, pi09822, pi09823, pi09824, pi09825, pi09826, pi09827, pi09828, pi09829, pi09830, pi09831, pi09832, pi09833, pi09834, pi09835, pi09836, pi09837, pi09838, pi09839, pi09840, pi09841, pi09842, pi09843, pi09844, pi09845, pi09846, pi09847, pi09848, pi09849, pi09850, pi09851, pi09852, pi09853, pi09854, pi09855, pi09856, pi09857, pi09858, pi09859, pi09860, pi09861, pi09862, pi09863, pi09864, pi09865, pi09866, pi09867, pi09868, pi09869, pi09870, pi09871, pi09872, pi09873, pi09874, pi09875, pi09876, pi09877, pi09878, pi09879, pi09880, pi09881, pi09882, pi09883, pi09884, pi09885, pi09886, pi09887, pi09888, pi09889, pi09890, pi09891, pi09892, pi09893, pi09894, pi09895, pi09896, pi09897, pi09898, pi09899, pi09900, pi09901, pi09902, pi09903, pi09904, pi09905, pi09906, pi09907, pi09908, pi09909, pi09910, pi09911, pi09912, pi09913, pi09914, pi09915, pi09916, pi09917, pi09918, pi09919, pi09920, pi09921, pi09922, pi09923, pi09924, pi09925, pi09926, pi09927, pi09928, pi09929, pi09930, pi09931, pi09932, pi09933, pi09934, pi09935, pi09936, pi09937, pi09938, pi09939, pi09940, pi09941, pi09942, pi09943, pi09944, pi09945, pi09946, pi09947, pi09948, pi09949, pi09950, pi09951, pi09952, pi09953, pi09954, pi09955, pi09956, pi09957, pi09958, pi09959, pi09960, pi09961, pi09962, pi09963, pi09964, pi09965, pi09966, pi09967, pi09968, pi09969, pi09970, pi09971, pi09972, pi09973, pi09974, pi09975, pi09976, pi09977, pi09978, pi09979, pi09980, pi09981, pi09982, pi09983, pi09984, pi09985, pi09986, pi09987, pi09988, pi09989, pi09990, pi09991, pi09992, pi09993, pi09994, pi09995, pi09996, pi09997, pi09998, pi09999, pi10000, pi10001, pi10002, pi10003, pi10004, pi10005, pi10006, pi10007, pi10008, pi10009, pi10010, pi10011, pi10012, pi10013, pi10014, pi10015, pi10016, pi10017, pi10018, pi10019, pi10020, pi10021, pi10022, pi10023, pi10024, pi10025, pi10026, pi10027, pi10028, pi10029, pi10030, pi10031, pi10032, pi10033, pi10034, pi10035, pi10036, pi10037, pi10038, pi10039, pi10040, pi10041, pi10042, pi10043, pi10044, pi10045, pi10046, pi10047, pi10048, pi10049, pi10050, pi10051, pi10052, pi10053, pi10054, pi10055, pi10056, pi10057, pi10058, pi10059, pi10060, pi10061, pi10062, pi10063, pi10064, pi10065, pi10066, pi10067, pi10068, pi10069, pi10070, pi10071, pi10072, pi10073, pi10074, pi10075, pi10076, pi10077, pi10078, pi10079, pi10080, pi10081, pi10082, pi10083, pi10084, pi10085, pi10086, pi10087, pi10088, pi10089, pi10090, pi10091, pi10092, pi10093, pi10094, pi10095, pi10096, pi10097, pi10098, pi10099, pi10100, pi10101, pi10102, pi10103, pi10104, pi10105, pi10106, pi10107, pi10108, pi10109, pi10110, pi10111, pi10112, pi10113, pi10114, pi10115, pi10116, pi10117, pi10118, pi10119, pi10120, pi10121, pi10122, pi10123, pi10124, pi10125, pi10126, pi10127, pi10128, pi10129, pi10130, pi10131, pi10132, pi10133, pi10134, pi10135, pi10136, pi10137, pi10138, pi10139, pi10140, pi10141, pi10142, pi10143, pi10144, pi10145, pi10146, pi10147, pi10148, pi10149, pi10150, pi10151, pi10152, pi10153, pi10154, pi10155, pi10156, pi10157, pi10158, pi10159, pi10160, pi10161, pi10162, pi10163, pi10164, pi10165, pi10166, pi10167, pi10168, pi10169, pi10170, pi10171, pi10172, pi10173, pi10174, pi10175, pi10176, pi10177, pi10178, pi10179, pi10180, pi10181, pi10182, pi10183, pi10184, pi10185, pi10186, pi10187, pi10188, pi10189, pi10190, pi10191, pi10192, pi10193, pi10194, pi10195, pi10196, pi10197, pi10198, pi10199, pi10200, pi10201, pi10202, pi10203, pi10204, pi10205, pi10206, pi10207, pi10208, pi10209, pi10210, pi10211, pi10212, pi10213, pi10214, pi10215, pi10216, pi10217, pi10218, pi10219, pi10220, pi10221, pi10222, pi10223, pi10224, pi10225, pi10226, pi10227, pi10228, pi10229, pi10230, pi10231, pi10232, pi10233, pi10234, pi10235, pi10236, pi10237, pi10238, pi10239, pi10240, pi10241, pi10242, pi10243, pi10244, pi10245, pi10246, pi10247, pi10248, pi10249, pi10250, pi10251, pi10252, pi10253, pi10254, pi10255, pi10256, pi10257, pi10258, pi10259, pi10260, pi10261, pi10262, pi10263, pi10264, pi10265, pi10266, pi10267, pi10268, pi10269, pi10270, pi10271, pi10272, pi10273, pi10274, pi10275, pi10276, pi10277, pi10278, pi10279, pi10280, pi10281, pi10282, pi10283, pi10284, pi10285, pi10286, pi10287, pi10288, pi10289, pi10290, pi10291, pi10292, pi10293, pi10294, pi10295, pi10296, pi10297, pi10298, pi10299, pi10300, pi10301, pi10302, pi10303, pi10304, pi10305, pi10306, pi10307, pi10308, pi10309, pi10310, pi10311, pi10312, pi10313, pi10314, pi10315, pi10316, pi10317, pi10318, pi10319, pi10320, pi10321, pi10322, pi10323, pi10324, pi10325, pi10326, pi10327, pi10328, pi10329, pi10330, pi10331, pi10332, pi10333, pi10334, pi10335, pi10336, pi10337, pi10338, pi10339, pi10340, pi10341, pi10342, pi10343, pi10344, pi10345, pi10346, pi10347, pi10348, pi10349, pi10350, pi10351, pi10352, pi10353, pi10354, pi10355, pi10356, pi10357, pi10358, pi10359, pi10360, pi10361, pi10362, pi10363, pi10364, pi10365, pi10366, pi10367, pi10368, pi10369, pi10370, pi10371, pi10372, pi10373, pi10374, pi10375, pi10376, pi10377, pi10378, pi10379, pi10380, pi10381, pi10382, pi10383, pi10384, pi10385, pi10386, pi10387, pi10388, pi10389, pi10390, pi10391, pi10392, pi10393, pi10394, pi10395, pi10396, pi10397, pi10398, pi10399, pi10400, pi10401, pi10402, pi10403, pi10404, pi10405, pi10406, pi10407, pi10408, pi10409, pi10410, pi10411, pi10412, pi10413, pi10414, pi10415, pi10416, pi10417, pi10418, pi10419, pi10420, pi10421, pi10422, pi10423, pi10424, pi10425, pi10426, pi10427, pi10428, pi10429, pi10430, pi10431, pi10432, pi10433, pi10434, pi10435, pi10436, pi10437, pi10438, pi10439, pi10440, pi10441, pi10442, pi10443, pi10444, pi10445, pi10446, pi10447, pi10448, pi10449, pi10450, pi10451, pi10452, pi10453, pi10454, pi10455, pi10456, pi10457, pi10458, pi10459, pi10460, pi10461, pi10462, pi10463, pi10464, pi10465, pi10466, pi10467, pi10468, pi10469, pi10470, pi10471, pi10472, pi10473, pi10474, pi10475, pi10476, pi10477, pi10478, pi10479, pi10480, pi10481, pi10482, pi10483, pi10484, pi10485, pi10486, pi10487, pi10488, pi10489, pi10490, pi10491, pi10492, pi10493, pi10494, pi10495, pi10496, pi10497, pi10498, pi10499, pi10500, pi10501, pi10502, pi10503, pi10504, pi10505, pi10506, pi10507, pi10508, pi10509, pi10510, pi10511, pi10512, pi10513, pi10514, pi10515, pi10516, pi10517, pi10518, pi10519, pi10520, pi10521, pi10522, pi10523, pi10524, pi10525, pi10526, pi10527, pi10528, pi10529, pi10530, pi10531, pi10532, pi10533, pi10534, pi10535, pi10536, pi10537, pi10538, pi10539, pi10540, pi10541, pi10542, pi10543, pi10544, pi10545, pi10546, pi10547, pi10548, pi10549, pi10550, pi10551, pi10552, pi10553, pi10554, pi10555, pi10556, pi10557, pi10558, pi10559, pi10560, pi10561, pi10562, pi10563, pi10564, pi10565, pi10566, pi10567, pi10568, pi10569, pi10570, pi10571, pi10572, pi10573, pi10574, pi10575, pi10576, pi10577, pi10578, pi10579, pi10580, pi10581, pi10582, pi10583, pi10584, pi10585, pi10586, pi10587, pi10588, pi10589, pi10590, pi10591, pi10592, pi10593, pi10594, pi10595, pi10596, pi10597, pi10598, pi10599, pi10600, pi10601, pi10602, pi10603, pi10604, pi10605, pi10606, pi10607, pi10608, pi10609, pi10610, pi10611, pi10612, pi10613, pi10614, pi10615, pi10616, pi10617, pi10618, pi10619, pi10620, pi10621, pi10622, pi10623, pi10624, pi10625, pi10626, pi10627, pi10628, pi10629, pi10630, pi10631, pi10632, pi10633, pi10634, pi10635, pi10636, pi10637, pi10638, pi10639, pi10640, pi10641, pi10642, pi10643, pi10644, pi10645, pi10646, pi10647, pi10648, pi10649, pi10650, pi10651, pi10652, pi10653, pi10654, pi10655, pi10656, pi10657, pi10658, pi10659, pi10660, pi10661, pi10662, pi10663, pi10664, pi10665, pi10666, pi10667, pi10668, pi10669, pi10670, pi10671;
output po00000, po00001, po00002, po00003, po00004, po00005, po00006, po00007, po00008, po00009, po00010, po00011, po00012, po00013, po00014, po00015, po00016, po00017, po00018, po00019, po00020, po00021, po00022, po00023, po00024, po00025, po00026, po00027, po00028, po00029, po00030, po00031, po00032, po00033, po00034, po00035, po00036, po00037, po00038, po00039, po00040, po00041, po00042, po00043, po00044, po00045, po00046, po00047, po00048, po00049, po00050, po00051, po00052, po00053, po00054, po00055, po00056, po00057, po00058, po00059, po00060, po00061, po00062, po00063, po00064, po00065, po00066, po00067, po00068, po00069, po00070, po00071, po00072, po00073, po00074, po00075, po00076, po00077, po00078, po00079, po00080, po00081, po00082, po00083, po00084, po00085, po00086, po00087, po00088, po00089, po00090, po00091, po00092, po00093, po00094, po00095, po00096, po00097, po00098, po00099, po00100, po00101, po00102, po00103, po00104, po00105, po00106, po00107, po00108, po00109, po00110, po00111, po00112, po00113, po00114, po00115, po00116, po00117, po00118, po00119, po00120, po00121, po00122, po00123, po00124, po00125, po00126, po00127, po00128, po00129, po00130, po00131, po00132, po00133, po00134, po00135, po00136, po00137, po00138, po00139, po00140, po00141, po00142, po00143, po00144, po00145, po00146, po00147, po00148, po00149, po00150, po00151, po00152, po00153, po00154, po00155, po00156, po00157, po00158, po00159, po00160, po00161, po00162, po00163, po00164, po00165, po00166, po00167, po00168, po00169, po00170, po00171, po00172, po00173, po00174, po00175, po00176, po00177, po00178, po00179, po00180, po00181, po00182, po00183, po00184, po00185, po00186, po00187, po00188, po00189, po00190, po00191, po00192, po00193, po00194, po00195, po00196, po00197, po00198, po00199, po00200, po00201, po00202, po00203, po00204, po00205, po00206, po00207, po00208, po00209, po00210, po00211, po00212, po00213, po00214, po00215, po00216, po00217, po00218, po00219, po00220, po00221, po00222, po00223, po00224, po00225, po00226, po00227, po00228, po00229, po00230, po00231, po00232, po00233, po00234, po00235, po00236, po00237, po00238, po00239, po00240, po00241, po00242, po00243, po00244, po00245, po00246, po00247, po00248, po00249, po00250, po00251, po00252, po00253, po00254, po00255, po00256, po00257, po00258, po00259, po00260, po00261, po00262, po00263, po00264, po00265, po00266, po00267, po00268, po00269, po00270, po00271, po00272, po00273, po00274, po00275, po00276, po00277, po00278, po00279, po00280, po00281, po00282, po00283, po00284, po00285, po00286, po00287, po00288, po00289, po00290, po00291, po00292, po00293, po00294, po00295, po00296, po00297, po00298, po00299, po00300, po00301, po00302, po00303, po00304, po00305, po00306, po00307, po00308, po00309, po00310, po00311, po00312, po00313, po00314, po00315, po00316, po00317, po00318, po00319, po00320, po00321, po00322, po00323, po00324, po00325, po00326, po00327, po00328, po00329, po00330, po00331, po00332, po00333, po00334, po00335, po00336, po00337, po00338, po00339, po00340, po00341, po00342, po00343, po00344, po00345, po00346, po00347, po00348, po00349, po00350, po00351, po00352, po00353, po00354, po00355, po00356, po00357, po00358, po00359, po00360, po00361, po00362, po00363, po00364, po00365, po00366, po00367, po00368, po00369, po00370, po00371, po00372, po00373, po00374, po00375, po00376, po00377, po00378, po00379, po00380, po00381, po00382, po00383, po00384, po00385, po00386, po00387, po00388, po00389, po00390, po00391, po00392, po00393, po00394, po00395, po00396, po00397, po00398, po00399, po00400, po00401, po00402, po00403, po00404, po00405, po00406, po00407, po00408, po00409, po00410, po00411, po00412, po00413, po00414, po00415, po00416, po00417, po00418, po00419, po00420, po00421, po00422, po00423, po00424, po00425, po00426, po00427, po00428, po00429, po00430, po00431, po00432, po00433, po00434, po00435, po00436, po00437, po00438, po00439, po00440, po00441, po00442, po00443, po00444, po00445, po00446, po00447, po00448, po00449, po00450, po00451, po00452, po00453, po00454, po00455, po00456, po00457, po00458, po00459, po00460, po00461, po00462, po00463, po00464, po00465, po00466, po00467, po00468, po00469, po00470, po00471, po00472, po00473, po00474, po00475, po00476, po00477, po00478, po00479, po00480, po00481, po00482, po00483, po00484, po00485, po00486, po00487, po00488, po00489, po00490, po00491, po00492, po00493, po00494, po00495, po00496, po00497, po00498, po00499, po00500, po00501, po00502, po00503, po00504, po00505, po00506, po00507, po00508, po00509, po00510, po00511, po00512, po00513, po00514, po00515, po00516, po00517, po00518, po00519, po00520, po00521, po00522, po00523, po00524, po00525, po00526, po00527, po00528, po00529, po00530, po00531, po00532, po00533, po00534, po00535, po00536, po00537, po00538, po00539, po00540, po00541, po00542, po00543, po00544, po00545, po00546, po00547, po00548, po00549, po00550, po00551, po00552, po00553, po00554, po00555, po00556, po00557, po00558, po00559, po00560, po00561, po00562, po00563, po00564, po00565, po00566, po00567, po00568, po00569, po00570, po00571, po00572, po00573, po00574, po00575, po00576, po00577, po00578, po00579, po00580, po00581, po00582, po00583, po00584, po00585, po00586, po00587, po00588, po00589, po00590, po00591, po00592, po00593, po00594, po00595, po00596, po00597, po00598, po00599, po00600, po00601, po00602, po00603, po00604, po00605, po00606, po00607, po00608, po00609, po00610, po00611, po00612, po00613, po00614, po00615, po00616, po00617, po00618, po00619, po00620, po00621, po00622, po00623, po00624, po00625, po00626, po00627, po00628, po00629, po00630, po00631, po00632, po00633, po00634, po00635, po00636, po00637, po00638, po00639, po00640, po00641, po00642, po00643, po00644, po00645, po00646, po00647, po00648, po00649, po00650, po00651, po00652, po00653, po00654, po00655, po00656, po00657, po00658, po00659, po00660, po00661, po00662, po00663, po00664, po00665, po00666, po00667, po00668, po00669, po00670, po00671, po00672, po00673, po00674, po00675, po00676, po00677, po00678, po00679, po00680, po00681, po00682, po00683, po00684, po00685, po00686, po00687, po00688, po00689, po00690, po00691, po00692, po00693, po00694, po00695, po00696, po00697, po00698, po00699, po00700, po00701, po00702, po00703, po00704, po00705, po00706, po00707, po00708, po00709, po00710, po00711, po00712, po00713, po00714, po00715, po00716, po00717, po00718, po00719, po00720, po00721, po00722, po00723, po00724, po00725, po00726, po00727, po00728, po00729, po00730, po00731, po00732, po00733, po00734, po00735, po00736, po00737, po00738, po00739, po00740, po00741, po00742, po00743, po00744, po00745, po00746, po00747, po00748, po00749, po00750, po00751, po00752, po00753, po00754, po00755, po00756, po00757, po00758, po00759, po00760, po00761, po00762, po00763, po00764, po00765, po00766, po00767, po00768, po00769, po00770, po00771, po00772, po00773, po00774, po00775, po00776, po00777, po00778, po00779, po00780, po00781, po00782, po00783, po00784, po00785, po00786, po00787, po00788, po00789, po00790, po00791, po00792, po00793, po00794, po00795, po00796, po00797, po00798, po00799, po00800, po00801, po00802, po00803, po00804, po00805, po00806, po00807, po00808, po00809, po00810, po00811, po00812, po00813, po00814, po00815, po00816, po00817, po00818, po00819, po00820, po00821, po00822, po00823, po00824, po00825, po00826, po00827, po00828, po00829, po00830, po00831, po00832, po00833, po00834, po00835, po00836, po00837, po00838, po00839, po00840, po00841, po00842, po00843, po00844, po00845, po00846, po00847, po00848, po00849, po00850, po00851, po00852, po00853, po00854, po00855, po00856, po00857, po00858, po00859, po00860, po00861, po00862, po00863, po00864, po00865, po00866, po00867, po00868, po00869, po00870, po00871, po00872, po00873, po00874, po00875, po00876, po00877, po00878, po00879, po00880, po00881, po00882, po00883, po00884, po00885, po00886, po00887, po00888, po00889, po00890, po00891, po00892, po00893, po00894, po00895, po00896, po00897, po00898, po00899, po00900, po00901, po00902, po00903, po00904, po00905, po00906, po00907, po00908, po00909, po00910, po00911, po00912, po00913, po00914, po00915, po00916, po00917, po00918, po00919, po00920, po00921, po00922, po00923, po00924, po00925, po00926, po00927, po00928, po00929, po00930, po00931, po00932, po00933, po00934, po00935, po00936, po00937, po00938, po00939, po00940, po00941, po00942, po00943, po00944, po00945, po00946, po00947, po00948, po00949, po00950, po00951, po00952, po00953, po00954, po00955, po00956, po00957, po00958, po00959, po00960, po00961, po00962, po00963, po00964, po00965, po00966, po00967, po00968, po00969, po00970, po00971, po00972, po00973, po00974, po00975, po00976, po00977, po00978, po00979, po00980, po00981, po00982, po00983, po00984, po00985, po00986, po00987, po00988, po00989, po00990, po00991, po00992, po00993, po00994, po00995, po00996, po00997, po00998, po00999, po01000, po01001, po01002, po01003, po01004, po01005, po01006, po01007, po01008, po01009, po01010, po01011, po01012, po01013, po01014, po01015, po01016, po01017, po01018, po01019, po01020, po01021, po01022, po01023, po01024, po01025, po01026, po01027, po01028, po01029, po01030, po01031, po01032, po01033, po01034, po01035, po01036, po01037, po01038, po01039, po01040, po01041, po01042, po01043, po01044, po01045, po01046, po01047, po01048, po01049, po01050, po01051, po01052, po01053, po01054, po01055, po01056, po01057, po01058, po01059, po01060, po01061, po01062, po01063, po01064, po01065, po01066, po01067, po01068, po01069, po01070, po01071, po01072, po01073, po01074, po01075, po01076, po01077, po01078, po01079, po01080, po01081, po01082, po01083, po01084, po01085, po01086, po01087, po01088, po01089, po01090, po01091, po01092, po01093, po01094, po01095, po01096, po01097, po01098, po01099, po01100, po01101, po01102, po01103, po01104, po01105, po01106, po01107, po01108, po01109, po01110, po01111, po01112, po01113, po01114, po01115, po01116, po01117, po01118, po01119, po01120, po01121, po01122, po01123, po01124, po01125, po01126, po01127, po01128, po01129, po01130, po01131, po01132, po01133, po01134, po01135, po01136, po01137, po01138, po01139, po01140, po01141, po01142, po01143, po01144, po01145, po01146, po01147, po01148, po01149, po01150, po01151, po01152, po01153, po01154, po01155, po01156, po01157, po01158, po01159, po01160, po01161, po01162, po01163, po01164, po01165, po01166, po01167, po01168, po01169, po01170, po01171, po01172, po01173, po01174, po01175, po01176, po01177, po01178, po01179, po01180, po01181, po01182, po01183, po01184, po01185, po01186, po01187, po01188, po01189, po01190, po01191, po01192, po01193, po01194, po01195, po01196, po01197, po01198, po01199, po01200, po01201, po01202, po01203, po01204, po01205, po01206, po01207, po01208, po01209, po01210, po01211, po01212, po01213, po01214, po01215, po01216, po01217, po01218, po01219, po01220, po01221, po01222, po01223, po01224, po01225, po01226, po01227, po01228, po01229, po01230, po01231, po01232, po01233, po01234, po01235, po01236, po01237, po01238, po01239, po01240, po01241, po01242, po01243, po01244, po01245, po01246, po01247, po01248, po01249, po01250, po01251, po01252, po01253, po01254, po01255, po01256, po01257, po01258, po01259, po01260, po01261, po01262, po01263, po01264, po01265, po01266, po01267, po01268, po01269, po01270, po01271, po01272, po01273, po01274, po01275, po01276, po01277, po01278, po01279, po01280, po01281, po01282, po01283, po01284, po01285, po01286, po01287, po01288, po01289, po01290, po01291, po01292, po01293, po01294, po01295, po01296, po01297, po01298, po01299, po01300, po01301, po01302, po01303, po01304, po01305, po01306, po01307, po01308, po01309, po01310, po01311, po01312, po01313, po01314, po01315, po01316, po01317, po01318, po01319, po01320, po01321, po01322, po01323, po01324, po01325, po01326, po01327, po01328, po01329, po01330, po01331, po01332, po01333, po01334, po01335, po01336, po01337, po01338, po01339, po01340, po01341, po01342, po01343, po01344, po01345, po01346, po01347, po01348, po01349, po01350, po01351, po01352, po01353, po01354, po01355, po01356, po01357, po01358, po01359, po01360, po01361, po01362, po01363, po01364, po01365, po01366, po01367, po01368, po01369, po01370, po01371, po01372, po01373, po01374, po01375, po01376, po01377, po01378, po01379, po01380, po01381, po01382, po01383, po01384, po01385, po01386, po01387, po01388, po01389, po01390, po01391, po01392, po01393, po01394, po01395, po01396, po01397, po01398, po01399, po01400, po01401, po01402, po01403, po01404, po01405, po01406, po01407, po01408, po01409, po01410, po01411, po01412, po01413, po01414, po01415, po01416, po01417, po01418, po01419, po01420, po01421, po01422, po01423, po01424, po01425, po01426, po01427, po01428, po01429, po01430, po01431, po01432, po01433, po01434, po01435, po01436, po01437, po01438, po01439, po01440, po01441, po01442, po01443, po01444, po01445, po01446, po01447, po01448, po01449, po01450, po01451, po01452, po01453, po01454, po01455, po01456, po01457, po01458, po01459, po01460, po01461, po01462, po01463, po01464, po01465, po01466, po01467, po01468, po01469, po01470, po01471, po01472, po01473, po01474, po01475, po01476, po01477, po01478, po01479, po01480, po01481, po01482, po01483, po01484, po01485, po01486, po01487, po01488, po01489, po01490, po01491, po01492, po01493, po01494, po01495, po01496, po01497, po01498, po01499, po01500, po01501, po01502, po01503, po01504, po01505, po01506, po01507, po01508, po01509, po01510, po01511, po01512, po01513, po01514, po01515, po01516, po01517, po01518, po01519, po01520, po01521, po01522, po01523, po01524, po01525, po01526, po01527, po01528, po01529, po01530, po01531, po01532, po01533, po01534, po01535, po01536, po01537, po01538, po01539, po01540, po01541, po01542, po01543, po01544, po01545, po01546, po01547, po01548, po01549, po01550, po01551, po01552, po01553, po01554, po01555, po01556, po01557, po01558, po01559, po01560, po01561, po01562, po01563, po01564, po01565, po01566, po01567, po01568, po01569, po01570, po01571, po01572, po01573, po01574, po01575, po01576, po01577, po01578, po01579, po01580, po01581, po01582, po01583, po01584, po01585, po01586, po01587, po01588, po01589, po01590, po01591, po01592, po01593, po01594, po01595, po01596, po01597, po01598, po01599, po01600, po01601, po01602, po01603, po01604, po01605, po01606, po01607, po01608, po01609, po01610, po01611, po01612, po01613, po01614, po01615, po01616, po01617, po01618, po01619, po01620, po01621, po01622, po01623, po01624, po01625, po01626, po01627, po01628, po01629, po01630, po01631, po01632, po01633, po01634, po01635, po01636, po01637, po01638, po01639, po01640, po01641, po01642, po01643, po01644, po01645, po01646, po01647, po01648, po01649, po01650, po01651, po01652, po01653, po01654, po01655, po01656, po01657, po01658, po01659, po01660, po01661, po01662, po01663, po01664, po01665, po01666, po01667, po01668, po01669, po01670, po01671, po01672, po01673, po01674, po01675, po01676, po01677, po01678, po01679, po01680, po01681, po01682, po01683, po01684, po01685, po01686, po01687, po01688, po01689, po01690, po01691, po01692, po01693, po01694, po01695, po01696, po01697, po01698, po01699, po01700, po01701, po01702, po01703, po01704, po01705, po01706, po01707, po01708, po01709, po01710, po01711, po01712, po01713, po01714, po01715, po01716, po01717, po01718, po01719, po01720, po01721, po01722, po01723, po01724, po01725, po01726, po01727, po01728, po01729, po01730, po01731, po01732, po01733, po01734, po01735, po01736, po01737, po01738, po01739, po01740, po01741, po01742, po01743, po01744, po01745, po01746, po01747, po01748, po01749, po01750, po01751, po01752, po01753, po01754, po01755, po01756, po01757, po01758, po01759, po01760, po01761, po01762, po01763, po01764, po01765, po01766, po01767, po01768, po01769, po01770, po01771, po01772, po01773, po01774, po01775, po01776, po01777, po01778, po01779, po01780, po01781, po01782, po01783, po01784, po01785, po01786, po01787, po01788, po01789, po01790, po01791, po01792, po01793, po01794, po01795, po01796, po01797, po01798, po01799, po01800, po01801, po01802, po01803, po01804, po01805, po01806, po01807, po01808, po01809, po01810, po01811, po01812, po01813, po01814, po01815, po01816, po01817, po01818, po01819, po01820, po01821, po01822, po01823, po01824, po01825, po01826, po01827, po01828, po01829, po01830, po01831, po01832, po01833, po01834, po01835, po01836, po01837, po01838, po01839, po01840, po01841, po01842, po01843, po01844, po01845, po01846, po01847, po01848, po01849, po01850, po01851, po01852, po01853, po01854, po01855, po01856, po01857, po01858, po01859, po01860, po01861, po01862, po01863, po01864, po01865, po01866, po01867, po01868, po01869, po01870, po01871, po01872, po01873, po01874, po01875, po01876, po01877, po01878, po01879, po01880, po01881, po01882, po01883, po01884, po01885, po01886, po01887, po01888, po01889, po01890, po01891, po01892, po01893, po01894, po01895, po01896, po01897, po01898, po01899, po01900, po01901, po01902, po01903, po01904, po01905, po01906, po01907, po01908, po01909, po01910, po01911, po01912, po01913, po01914, po01915, po01916, po01917, po01918, po01919, po01920, po01921, po01922, po01923, po01924, po01925, po01926, po01927, po01928, po01929, po01930, po01931, po01932, po01933, po01934, po01935, po01936, po01937, po01938, po01939, po01940, po01941, po01942, po01943, po01944, po01945, po01946, po01947, po01948, po01949, po01950, po01951, po01952, po01953, po01954, po01955, po01956, po01957, po01958, po01959, po01960, po01961, po01962, po01963, po01964, po01965, po01966, po01967, po01968, po01969, po01970, po01971, po01972, po01973, po01974, po01975, po01976, po01977, po01978, po01979, po01980, po01981, po01982, po01983, po01984, po01985, po01986, po01987, po01988, po01989, po01990, po01991, po01992, po01993, po01994, po01995, po01996, po01997, po01998, po01999, po02000, po02001, po02002, po02003, po02004, po02005, po02006, po02007, po02008, po02009, po02010, po02011, po02012, po02013, po02014, po02015, po02016, po02017, po02018, po02019, po02020, po02021, po02022, po02023, po02024, po02025, po02026, po02027, po02028, po02029, po02030, po02031, po02032, po02033, po02034, po02035, po02036, po02037, po02038, po02039, po02040, po02041, po02042, po02043, po02044, po02045, po02046, po02047, po02048, po02049, po02050, po02051, po02052, po02053, po02054, po02055, po02056, po02057, po02058, po02059, po02060, po02061, po02062, po02063, po02064, po02065, po02066, po02067, po02068, po02069, po02070, po02071, po02072, po02073, po02074, po02075, po02076, po02077, po02078, po02079, po02080, po02081, po02082, po02083, po02084, po02085, po02086, po02087, po02088, po02089, po02090, po02091, po02092, po02093, po02094, po02095, po02096, po02097, po02098, po02099, po02100, po02101, po02102, po02103, po02104, po02105, po02106, po02107, po02108, po02109, po02110, po02111, po02112, po02113, po02114, po02115, po02116, po02117, po02118, po02119, po02120, po02121, po02122, po02123, po02124, po02125, po02126, po02127, po02128, po02129, po02130, po02131, po02132, po02133, po02134, po02135, po02136, po02137, po02138, po02139, po02140, po02141, po02142, po02143, po02144, po02145, po02146, po02147, po02148, po02149, po02150, po02151, po02152, po02153, po02154, po02155, po02156, po02157, po02158, po02159, po02160, po02161, po02162, po02163, po02164, po02165, po02166, po02167, po02168, po02169, po02170, po02171, po02172, po02173, po02174, po02175, po02176, po02177, po02178, po02179, po02180, po02181, po02182, po02183, po02184, po02185, po02186, po02187, po02188, po02189, po02190, po02191, po02192, po02193, po02194, po02195, po02196, po02197, po02198, po02199, po02200, po02201, po02202, po02203, po02204, po02205, po02206, po02207, po02208, po02209, po02210, po02211, po02212, po02213, po02214, po02215, po02216, po02217, po02218, po02219, po02220, po02221, po02222, po02223, po02224, po02225, po02226, po02227, po02228, po02229, po02230, po02231, po02232, po02233, po02234, po02235, po02236, po02237, po02238, po02239, po02240, po02241, po02242, po02243, po02244, po02245, po02246, po02247, po02248, po02249, po02250, po02251, po02252, po02253, po02254, po02255, po02256, po02257, po02258, po02259, po02260, po02261, po02262, po02263, po02264, po02265, po02266, po02267, po02268, po02269, po02270, po02271, po02272, po02273, po02274, po02275, po02276, po02277, po02278, po02279, po02280, po02281, po02282, po02283, po02284, po02285, po02286, po02287, po02288, po02289, po02290, po02291, po02292, po02293, po02294, po02295, po02296, po02297, po02298, po02299, po02300, po02301, po02302, po02303, po02304, po02305, po02306, po02307, po02308, po02309, po02310, po02311, po02312, po02313, po02314, po02315, po02316, po02317, po02318, po02319, po02320, po02321, po02322, po02323, po02324, po02325, po02326, po02327, po02328, po02329, po02330, po02331, po02332, po02333, po02334, po02335, po02336, po02337, po02338, po02339, po02340, po02341, po02342, po02343, po02344, po02345, po02346, po02347, po02348, po02349, po02350, po02351, po02352, po02353, po02354, po02355, po02356, po02357, po02358, po02359, po02360, po02361, po02362, po02363, po02364, po02365, po02366, po02367, po02368, po02369, po02370, po02371, po02372, po02373, po02374, po02375, po02376, po02377, po02378, po02379, po02380, po02381, po02382, po02383, po02384, po02385, po02386, po02387, po02388, po02389, po02390, po02391, po02392, po02393, po02394, po02395, po02396, po02397, po02398, po02399, po02400, po02401, po02402, po02403, po02404, po02405, po02406, po02407, po02408, po02409, po02410, po02411, po02412, po02413, po02414, po02415, po02416, po02417, po02418, po02419, po02420, po02421, po02422, po02423, po02424, po02425, po02426, po02427, po02428, po02429, po02430, po02431, po02432, po02433, po02434, po02435, po02436, po02437, po02438, po02439, po02440, po02441, po02442, po02443, po02444, po02445, po02446, po02447, po02448, po02449, po02450, po02451, po02452, po02453, po02454, po02455, po02456, po02457, po02458, po02459, po02460, po02461, po02462, po02463, po02464, po02465, po02466, po02467, po02468, po02469, po02470, po02471, po02472, po02473, po02474, po02475, po02476, po02477, po02478, po02479, po02480, po02481, po02482, po02483, po02484, po02485, po02486, po02487, po02488, po02489, po02490, po02491, po02492, po02493, po02494, po02495, po02496, po02497, po02498, po02499, po02500, po02501, po02502, po02503, po02504, po02505, po02506, po02507, po02508, po02509, po02510, po02511, po02512, po02513, po02514, po02515, po02516, po02517, po02518, po02519, po02520, po02521, po02522, po02523, po02524, po02525, po02526, po02527, po02528, po02529, po02530, po02531, po02532, po02533, po02534, po02535, po02536, po02537, po02538, po02539, po02540, po02541, po02542, po02543, po02544, po02545, po02546, po02547, po02548, po02549, po02550, po02551, po02552, po02553, po02554, po02555, po02556, po02557, po02558, po02559, po02560, po02561, po02562, po02563, po02564, po02565, po02566, po02567, po02568, po02569, po02570, po02571, po02572, po02573, po02574, po02575, po02576, po02577, po02578, po02579, po02580, po02581, po02582, po02583, po02584, po02585, po02586, po02587, po02588, po02589, po02590, po02591, po02592, po02593, po02594, po02595, po02596, po02597, po02598, po02599, po02600, po02601, po02602, po02603, po02604, po02605, po02606, po02607, po02608, po02609, po02610, po02611, po02612, po02613, po02614, po02615, po02616, po02617, po02618, po02619, po02620, po02621, po02622, po02623, po02624, po02625, po02626, po02627, po02628, po02629, po02630, po02631, po02632, po02633, po02634, po02635, po02636, po02637, po02638, po02639, po02640, po02641, po02642, po02643, po02644, po02645, po02646, po02647, po02648, po02649, po02650, po02651, po02652, po02653, po02654, po02655, po02656, po02657, po02658, po02659, po02660, po02661, po02662, po02663, po02664, po02665, po02666, po02667, po02668, po02669, po02670, po02671, po02672, po02673, po02674, po02675, po02676, po02677, po02678, po02679, po02680, po02681, po02682, po02683, po02684, po02685, po02686, po02687, po02688, po02689, po02690, po02691, po02692, po02693, po02694, po02695, po02696, po02697, po02698, po02699, po02700, po02701, po02702, po02703, po02704, po02705, po02706, po02707, po02708, po02709, po02710, po02711, po02712, po02713, po02714, po02715, po02716, po02717, po02718, po02719, po02720, po02721, po02722, po02723, po02724, po02725, po02726, po02727, po02728, po02729, po02730, po02731, po02732, po02733, po02734, po02735, po02736, po02737, po02738, po02739, po02740, po02741, po02742, po02743, po02744, po02745, po02746, po02747, po02748, po02749, po02750, po02751, po02752, po02753, po02754, po02755, po02756, po02757, po02758, po02759, po02760, po02761, po02762, po02763, po02764, po02765, po02766, po02767, po02768, po02769, po02770, po02771, po02772, po02773, po02774, po02775, po02776, po02777, po02778, po02779, po02780, po02781, po02782, po02783, po02784, po02785, po02786, po02787, po02788, po02789, po02790, po02791, po02792, po02793, po02794, po02795, po02796, po02797, po02798, po02799, po02800, po02801, po02802, po02803, po02804, po02805, po02806, po02807, po02808, po02809, po02810, po02811, po02812, po02813, po02814, po02815, po02816, po02817, po02818, po02819, po02820, po02821, po02822, po02823, po02824, po02825, po02826, po02827, po02828, po02829, po02830, po02831, po02832, po02833, po02834, po02835, po02836, po02837, po02838, po02839, po02840, po02841, po02842, po02843, po02844, po02845, po02846, po02847, po02848, po02849, po02850, po02851, po02852, po02853, po02854, po02855, po02856, po02857, po02858, po02859, po02860, po02861, po02862, po02863, po02864, po02865, po02866, po02867, po02868, po02869, po02870, po02871, po02872, po02873, po02874, po02875, po02876, po02877, po02878, po02879, po02880, po02881, po02882, po02883, po02884, po02885, po02886, po02887, po02888, po02889, po02890, po02891, po02892, po02893, po02894, po02895, po02896, po02897, po02898, po02899, po02900, po02901, po02902, po02903, po02904, po02905, po02906, po02907, po02908, po02909, po02910, po02911, po02912, po02913, po02914, po02915, po02916, po02917, po02918, po02919, po02920, po02921, po02922, po02923, po02924, po02925, po02926, po02927, po02928, po02929, po02930, po02931, po02932, po02933, po02934, po02935, po02936, po02937, po02938, po02939, po02940, po02941, po02942, po02943, po02944, po02945, po02946, po02947, po02948, po02949, po02950, po02951, po02952, po02953, po02954, po02955, po02956, po02957, po02958, po02959, po02960, po02961, po02962, po02963, po02964, po02965, po02966, po02967, po02968, po02969, po02970, po02971, po02972, po02973, po02974, po02975, po02976, po02977, po02978, po02979, po02980, po02981, po02982, po02983, po02984, po02985, po02986, po02987, po02988, po02989, po02990, po02991, po02992, po02993, po02994, po02995, po02996, po02997, po02998, po02999, po03000, po03001, po03002, po03003, po03004, po03005, po03006, po03007, po03008, po03009, po03010, po03011, po03012, po03013, po03014, po03015, po03016, po03017, po03018, po03019, po03020, po03021, po03022, po03023, po03024, po03025, po03026, po03027, po03028, po03029, po03030, po03031, po03032, po03033, po03034, po03035, po03036, po03037, po03038, po03039, po03040, po03041, po03042, po03043, po03044, po03045, po03046, po03047, po03048, po03049, po03050, po03051, po03052, po03053, po03054, po03055, po03056, po03057, po03058, po03059, po03060, po03061, po03062, po03063, po03064, po03065, po03066, po03067, po03068, po03069, po03070, po03071, po03072, po03073, po03074, po03075, po03076, po03077, po03078, po03079, po03080, po03081, po03082, po03083, po03084, po03085, po03086, po03087, po03088, po03089, po03090, po03091, po03092, po03093, po03094, po03095, po03096, po03097, po03098, po03099, po03100, po03101, po03102, po03103, po03104, po03105, po03106, po03107, po03108, po03109, po03110, po03111, po03112, po03113, po03114, po03115, po03116, po03117, po03118, po03119, po03120, po03121, po03122, po03123, po03124, po03125, po03126, po03127, po03128, po03129, po03130, po03131, po03132, po03133, po03134, po03135, po03136, po03137, po03138, po03139, po03140, po03141, po03142, po03143, po03144, po03145, po03146, po03147, po03148, po03149, po03150, po03151, po03152, po03153, po03154, po03155, po03156, po03157, po03158, po03159, po03160, po03161, po03162, po03163, po03164, po03165, po03166, po03167, po03168, po03169, po03170, po03171, po03172, po03173, po03174, po03175, po03176, po03177, po03178, po03179, po03180, po03181, po03182, po03183, po03184, po03185, po03186, po03187, po03188, po03189, po03190, po03191, po03192, po03193, po03194, po03195, po03196, po03197, po03198, po03199, po03200, po03201, po03202, po03203, po03204, po03205, po03206, po03207, po03208, po03209, po03210, po03211, po03212, po03213, po03214, po03215, po03216, po03217, po03218, po03219, po03220, po03221, po03222, po03223, po03224, po03225, po03226, po03227, po03228, po03229, po03230, po03231, po03232, po03233, po03234, po03235, po03236, po03237, po03238, po03239, po03240, po03241, po03242, po03243, po03244, po03245, po03246, po03247, po03248, po03249, po03250, po03251, po03252, po03253, po03254, po03255, po03256, po03257, po03258, po03259, po03260, po03261, po03262, po03263, po03264, po03265, po03266, po03267, po03268, po03269, po03270, po03271, po03272, po03273, po03274, po03275, po03276, po03277, po03278, po03279, po03280, po03281, po03282, po03283, po03284, po03285, po03286, po03287, po03288, po03289, po03290, po03291, po03292, po03293, po03294, po03295, po03296, po03297, po03298, po03299, po03300, po03301, po03302, po03303, po03304, po03305, po03306, po03307, po03308, po03309, po03310, po03311, po03312, po03313, po03314, po03315, po03316, po03317, po03318, po03319, po03320, po03321, po03322, po03323, po03324, po03325, po03326, po03327, po03328, po03329, po03330, po03331, po03332, po03333, po03334, po03335, po03336, po03337, po03338, po03339, po03340, po03341, po03342, po03343, po03344, po03345, po03346, po03347, po03348, po03349, po03350, po03351, po03352, po03353, po03354, po03355, po03356, po03357, po03358, po03359, po03360, po03361, po03362, po03363, po03364, po03365, po03366, po03367, po03368, po03369, po03370, po03371, po03372, po03373, po03374, po03375, po03376, po03377, po03378, po03379, po03380, po03381, po03382, po03383, po03384, po03385, po03386, po03387, po03388, po03389, po03390, po03391, po03392, po03393, po03394, po03395, po03396, po03397, po03398, po03399, po03400, po03401, po03402, po03403, po03404, po03405, po03406, po03407, po03408, po03409, po03410, po03411, po03412, po03413, po03414, po03415, po03416, po03417, po03418, po03419, po03420, po03421, po03422, po03423, po03424, po03425, po03426, po03427, po03428, po03429, po03430, po03431, po03432, po03433, po03434, po03435, po03436, po03437, po03438, po03439, po03440, po03441, po03442, po03443, po03444, po03445, po03446, po03447, po03448, po03449, po03450, po03451, po03452, po03453, po03454, po03455, po03456, po03457, po03458, po03459, po03460, po03461, po03462, po03463, po03464, po03465, po03466, po03467, po03468, po03469, po03470, po03471, po03472, po03473, po03474, po03475, po03476, po03477, po03478, po03479, po03480, po03481, po03482, po03483, po03484, po03485, po03486, po03487, po03488, po03489, po03490, po03491, po03492, po03493, po03494, po03495, po03496, po03497, po03498, po03499, po03500, po03501, po03502, po03503, po03504, po03505, po03506, po03507, po03508, po03509, po03510, po03511, po03512, po03513, po03514, po03515, po03516, po03517, po03518, po03519, po03520, po03521, po03522, po03523, po03524, po03525, po03526, po03527, po03528, po03529, po03530, po03531, po03532, po03533, po03534, po03535, po03536, po03537, po03538, po03539, po03540, po03541, po03542, po03543, po03544, po03545, po03546, po03547, po03548, po03549, po03550, po03551, po03552, po03553, po03554, po03555, po03556, po03557, po03558, po03559, po03560, po03561, po03562, po03563, po03564, po03565, po03566, po03567, po03568, po03569, po03570, po03571, po03572, po03573, po03574, po03575, po03576, po03577, po03578, po03579, po03580, po03581, po03582, po03583, po03584, po03585, po03586, po03587, po03588, po03589, po03590, po03591, po03592, po03593, po03594, po03595, po03596, po03597, po03598, po03599, po03600, po03601, po03602, po03603, po03604, po03605, po03606, po03607, po03608, po03609, po03610, po03611, po03612, po03613, po03614, po03615, po03616, po03617, po03618, po03619, po03620, po03621, po03622, po03623, po03624, po03625, po03626, po03627, po03628, po03629, po03630, po03631, po03632, po03633, po03634, po03635, po03636, po03637, po03638, po03639, po03640, po03641, po03642, po03643, po03644, po03645, po03646, po03647, po03648, po03649, po03650, po03651, po03652, po03653, po03654, po03655, po03656, po03657, po03658, po03659, po03660, po03661, po03662, po03663, po03664, po03665, po03666, po03667, po03668, po03669, po03670, po03671, po03672, po03673, po03674, po03675, po03676, po03677, po03678, po03679, po03680, po03681, po03682, po03683, po03684, po03685, po03686, po03687, po03688, po03689, po03690, po03691, po03692, po03693, po03694, po03695, po03696, po03697, po03698, po03699, po03700, po03701, po03702, po03703, po03704, po03705, po03706, po03707, po03708, po03709, po03710, po03711, po03712, po03713, po03714, po03715, po03716, po03717, po03718, po03719, po03720, po03721, po03722, po03723, po03724, po03725, po03726, po03727, po03728, po03729, po03730, po03731, po03732, po03733, po03734, po03735, po03736, po03737, po03738, po03739, po03740, po03741, po03742, po03743, po03744, po03745, po03746, po03747, po03748, po03749, po03750, po03751, po03752, po03753, po03754, po03755, po03756, po03757, po03758, po03759, po03760, po03761, po03762, po03763, po03764, po03765, po03766, po03767, po03768, po03769, po03770, po03771, po03772, po03773, po03774, po03775, po03776, po03777, po03778, po03779, po03780, po03781, po03782, po03783, po03784, po03785, po03786, po03787, po03788, po03789, po03790, po03791, po03792, po03793, po03794, po03795, po03796, po03797, po03798, po03799, po03800, po03801, po03802, po03803, po03804, po03805, po03806, po03807, po03808, po03809, po03810, po03811, po03812, po03813, po03814, po03815, po03816, po03817, po03818, po03819, po03820, po03821, po03822, po03823, po03824, po03825, po03826, po03827, po03828, po03829, po03830, po03831, po03832, po03833, po03834, po03835, po03836, po03837, po03838, po03839, po03840, po03841, po03842, po03843, po03844, po03845, po03846, po03847, po03848, po03849, po03850, po03851, po03852, po03853, po03854, po03855, po03856, po03857, po03858, po03859, po03860, po03861, po03862, po03863, po03864, po03865, po03866, po03867, po03868, po03869, po03870, po03871, po03872, po03873, po03874, po03875, po03876, po03877, po03878, po03879, po03880, po03881, po03882, po03883, po03884, po03885, po03886, po03887, po03888, po03889, po03890, po03891, po03892, po03893, po03894, po03895, po03896, po03897, po03898, po03899, po03900, po03901, po03902, po03903, po03904, po03905, po03906, po03907, po03908, po03909, po03910, po03911, po03912, po03913, po03914, po03915, po03916, po03917, po03918, po03919, po03920, po03921, po03922, po03923, po03924, po03925, po03926, po03927, po03928, po03929, po03930, po03931, po03932, po03933, po03934, po03935, po03936, po03937, po03938, po03939, po03940, po03941, po03942, po03943, po03944, po03945, po03946, po03947, po03948, po03949, po03950, po03951, po03952, po03953, po03954, po03955, po03956, po03957, po03958, po03959, po03960, po03961, po03962, po03963, po03964, po03965, po03966, po03967, po03968, po03969, po03970, po03971, po03972, po03973, po03974, po03975, po03976, po03977, po03978, po03979, po03980, po03981, po03982, po03983, po03984, po03985, po03986, po03987, po03988, po03989, po03990, po03991, po03992, po03993, po03994, po03995, po03996, po03997, po03998, po03999, po04000, po04001, po04002, po04003, po04004, po04005, po04006, po04007, po04008, po04009, po04010, po04011, po04012, po04013, po04014, po04015, po04016, po04017, po04018, po04019, po04020, po04021, po04022, po04023, po04024, po04025, po04026, po04027, po04028, po04029, po04030, po04031, po04032, po04033, po04034, po04035, po04036, po04037, po04038, po04039, po04040, po04041, po04042, po04043, po04044, po04045, po04046, po04047, po04048, po04049, po04050, po04051, po04052, po04053, po04054, po04055, po04056, po04057, po04058, po04059, po04060, po04061, po04062, po04063, po04064, po04065, po04066, po04067, po04068, po04069, po04070, po04071, po04072, po04073, po04074, po04075, po04076, po04077, po04078, po04079, po04080, po04081, po04082, po04083, po04084, po04085, po04086, po04087, po04088, po04089, po04090, po04091, po04092, po04093, po04094, po04095, po04096, po04097, po04098, po04099, po04100, po04101, po04102, po04103, po04104, po04105, po04106, po04107, po04108, po04109, po04110, po04111, po04112, po04113, po04114, po04115, po04116, po04117, po04118, po04119, po04120, po04121, po04122, po04123, po04124, po04125, po04126, po04127, po04128, po04129, po04130, po04131, po04132, po04133, po04134, po04135, po04136, po04137, po04138, po04139, po04140, po04141, po04142, po04143, po04144, po04145, po04146, po04147, po04148, po04149, po04150, po04151, po04152, po04153, po04154, po04155, po04156, po04157, po04158, po04159, po04160, po04161, po04162, po04163, po04164, po04165, po04166, po04167, po04168, po04169, po04170, po04171, po04172, po04173, po04174, po04175, po04176, po04177, po04178, po04179, po04180, po04181, po04182, po04183, po04184, po04185, po04186, po04187, po04188, po04189, po04190, po04191, po04192, po04193, po04194, po04195, po04196, po04197, po04198, po04199, po04200, po04201, po04202, po04203, po04204, po04205, po04206, po04207, po04208, po04209, po04210, po04211, po04212, po04213, po04214, po04215, po04216, po04217, po04218, po04219, po04220, po04221, po04222, po04223, po04224, po04225, po04226, po04227, po04228, po04229, po04230, po04231, po04232, po04233, po04234, po04235, po04236, po04237, po04238, po04239, po04240, po04241, po04242, po04243, po04244, po04245, po04246, po04247, po04248, po04249, po04250, po04251, po04252, po04253, po04254, po04255, po04256, po04257, po04258, po04259, po04260, po04261, po04262, po04263, po04264, po04265, po04266, po04267, po04268, po04269, po04270, po04271, po04272, po04273, po04274, po04275, po04276, po04277, po04278, po04279, po04280, po04281, po04282, po04283, po04284, po04285, po04286, po04287, po04288, po04289, po04290, po04291, po04292, po04293, po04294, po04295, po04296, po04297, po04298, po04299, po04300, po04301, po04302, po04303, po04304, po04305, po04306, po04307, po04308, po04309, po04310, po04311, po04312, po04313, po04314, po04315, po04316, po04317, po04318, po04319, po04320, po04321, po04322, po04323, po04324, po04325, po04326, po04327, po04328, po04329, po04330, po04331, po04332, po04333, po04334, po04335, po04336, po04337, po04338, po04339, po04340, po04341, po04342, po04343, po04344, po04345, po04346, po04347, po04348, po04349, po04350, po04351, po04352, po04353, po04354, po04355, po04356, po04357, po04358, po04359, po04360, po04361, po04362, po04363, po04364, po04365, po04366, po04367, po04368, po04369, po04370, po04371, po04372, po04373, po04374, po04375, po04376, po04377, po04378, po04379, po04380, po04381, po04382, po04383, po04384, po04385, po04386, po04387, po04388, po04389, po04390, po04391, po04392, po04393, po04394, po04395, po04396, po04397, po04398, po04399, po04400, po04401, po04402, po04403, po04404, po04405, po04406, po04407, po04408, po04409, po04410, po04411, po04412, po04413, po04414, po04415, po04416, po04417, po04418, po04419, po04420, po04421, po04422, po04423, po04424, po04425, po04426, po04427, po04428, po04429, po04430, po04431, po04432, po04433, po04434, po04435, po04436, po04437, po04438, po04439, po04440, po04441, po04442, po04443, po04444, po04445, po04446, po04447, po04448, po04449, po04450, po04451, po04452, po04453, po04454, po04455, po04456, po04457, po04458, po04459, po04460, po04461, po04462, po04463, po04464, po04465, po04466, po04467, po04468, po04469, po04470, po04471, po04472, po04473, po04474, po04475, po04476, po04477, po04478, po04479, po04480, po04481, po04482, po04483, po04484, po04485, po04486, po04487, po04488, po04489, po04490, po04491, po04492, po04493, po04494, po04495, po04496, po04497, po04498, po04499, po04500, po04501, po04502, po04503, po04504, po04505, po04506, po04507, po04508, po04509, po04510, po04511, po04512, po04513, po04514, po04515, po04516, po04517, po04518, po04519, po04520, po04521, po04522, po04523, po04524, po04525, po04526, po04527, po04528, po04529, po04530, po04531, po04532, po04533, po04534, po04535, po04536, po04537, po04538, po04539, po04540, po04541, po04542, po04543, po04544, po04545, po04546, po04547, po04548, po04549, po04550, po04551, po04552, po04553, po04554, po04555, po04556, po04557, po04558, po04559, po04560, po04561, po04562, po04563, po04564, po04565, po04566, po04567, po04568, po04569, po04570, po04571, po04572, po04573, po04574, po04575, po04576, po04577, po04578, po04579, po04580, po04581, po04582, po04583, po04584, po04585, po04586, po04587, po04588, po04589, po04590, po04591, po04592, po04593, po04594, po04595, po04596, po04597, po04598, po04599, po04600, po04601, po04602, po04603, po04604, po04605, po04606, po04607, po04608, po04609, po04610, po04611, po04612, po04613, po04614, po04615, po04616, po04617, po04618, po04619, po04620, po04621, po04622, po04623, po04624, po04625, po04626, po04627, po04628, po04629, po04630, po04631, po04632, po04633, po04634, po04635, po04636, po04637, po04638, po04639, po04640, po04641, po04642, po04643, po04644, po04645, po04646, po04647, po04648, po04649, po04650, po04651, po04652, po04653, po04654, po04655, po04656, po04657, po04658, po04659, po04660, po04661, po04662, po04663, po04664, po04665, po04666, po04667, po04668, po04669, po04670, po04671, po04672, po04673, po04674, po04675, po04676, po04677, po04678, po04679, po04680, po04681, po04682, po04683, po04684, po04685, po04686, po04687, po04688, po04689, po04690, po04691, po04692, po04693, po04694, po04695, po04696, po04697, po04698, po04699, po04700, po04701, po04702, po04703, po04704, po04705, po04706, po04707, po04708, po04709, po04710, po04711, po04712, po04713, po04714, po04715, po04716, po04717, po04718, po04719, po04720, po04721, po04722, po04723, po04724, po04725, po04726, po04727, po04728, po04729, po04730, po04731, po04732, po04733, po04734, po04735, po04736, po04737, po04738, po04739, po04740, po04741, po04742, po04743, po04744, po04745, po04746, po04747, po04748, po04749, po04750, po04751, po04752, po04753, po04754, po04755, po04756, po04757, po04758, po04759, po04760, po04761, po04762, po04763, po04764, po04765, po04766, po04767, po04768, po04769, po04770, po04771, po04772, po04773, po04774, po04775, po04776, po04777, po04778, po04779, po04780, po04781, po04782, po04783, po04784, po04785, po04786, po04787, po04788, po04789, po04790, po04791, po04792, po04793, po04794, po04795, po04796, po04797, po04798, po04799, po04800, po04801, po04802, po04803, po04804, po04805, po04806, po04807, po04808, po04809, po04810, po04811, po04812, po04813, po04814, po04815, po04816, po04817, po04818, po04819, po04820, po04821, po04822, po04823, po04824, po04825, po04826, po04827, po04828, po04829, po04830, po04831, po04832, po04833, po04834, po04835, po04836, po04837, po04838, po04839, po04840, po04841, po04842, po04843, po04844, po04845, po04846, po04847, po04848, po04849, po04850, po04851, po04852, po04853, po04854, po04855, po04856, po04857, po04858, po04859, po04860, po04861, po04862, po04863, po04864, po04865, po04866, po04867, po04868, po04869, po04870, po04871, po04872, po04873, po04874, po04875, po04876, po04877, po04878, po04879, po04880, po04881, po04882, po04883, po04884, po04885, po04886, po04887, po04888, po04889, po04890, po04891, po04892, po04893, po04894, po04895, po04896, po04897, po04898, po04899, po04900, po04901, po04902, po04903, po04904, po04905, po04906, po04907, po04908, po04909, po04910, po04911, po04912, po04913, po04914, po04915, po04916, po04917, po04918, po04919, po04920, po04921, po04922, po04923, po04924, po04925, po04926, po04927, po04928, po04929, po04930, po04931, po04932, po04933, po04934, po04935, po04936, po04937, po04938, po04939, po04940, po04941, po04942, po04943, po04944, po04945, po04946, po04947, po04948, po04949, po04950, po04951, po04952, po04953, po04954, po04955, po04956, po04957, po04958, po04959, po04960, po04961, po04962, po04963, po04964, po04965, po04966, po04967, po04968, po04969, po04970, po04971, po04972, po04973, po04974, po04975, po04976, po04977, po04978, po04979, po04980, po04981, po04982, po04983, po04984, po04985, po04986, po04987, po04988, po04989, po04990, po04991, po04992, po04993, po04994, po04995, po04996, po04997, po04998, po04999, po05000, po05001, po05002, po05003, po05004, po05005, po05006, po05007, po05008, po05009, po05010, po05011, po05012, po05013, po05014, po05015, po05016, po05017, po05018, po05019, po05020, po05021, po05022, po05023, po05024, po05025, po05026, po05027, po05028, po05029, po05030, po05031, po05032, po05033, po05034, po05035, po05036, po05037, po05038, po05039, po05040, po05041, po05042, po05043, po05044, po05045, po05046, po05047, po05048, po05049, po05050, po05051, po05052, po05053, po05054, po05055, po05056, po05057, po05058, po05059, po05060, po05061, po05062, po05063, po05064, po05065, po05066, po05067, po05068, po05069, po05070, po05071, po05072, po05073, po05074, po05075, po05076, po05077, po05078, po05079, po05080, po05081, po05082, po05083, po05084, po05085, po05086, po05087, po05088, po05089, po05090, po05091, po05092, po05093, po05094, po05095, po05096, po05097, po05098, po05099, po05100, po05101, po05102, po05103, po05104, po05105, po05106, po05107, po05108, po05109, po05110, po05111, po05112, po05113, po05114, po05115, po05116, po05117, po05118, po05119, po05120, po05121, po05122, po05123, po05124, po05125, po05126, po05127, po05128, po05129, po05130, po05131, po05132, po05133, po05134, po05135, po05136, po05137, po05138, po05139, po05140, po05141, po05142, po05143, po05144, po05145, po05146, po05147, po05148, po05149, po05150, po05151, po05152, po05153, po05154, po05155, po05156, po05157, po05158, po05159, po05160, po05161, po05162, po05163, po05164, po05165, po05166, po05167, po05168, po05169, po05170, po05171, po05172, po05173, po05174, po05175, po05176, po05177, po05178, po05179, po05180, po05181, po05182, po05183, po05184, po05185, po05186, po05187, po05188, po05189, po05190, po05191, po05192, po05193, po05194, po05195, po05196, po05197, po05198, po05199, po05200, po05201, po05202, po05203, po05204, po05205, po05206, po05207, po05208, po05209, po05210, po05211, po05212, po05213, po05214, po05215, po05216, po05217, po05218, po05219, po05220, po05221, po05222, po05223, po05224, po05225, po05226, po05227, po05228, po05229, po05230, po05231, po05232, po05233, po05234, po05235, po05236, po05237, po05238, po05239, po05240, po05241, po05242, po05243, po05244, po05245, po05246, po05247, po05248, po05249, po05250, po05251, po05252, po05253, po05254, po05255, po05256, po05257, po05258, po05259, po05260, po05261, po05262, po05263, po05264, po05265, po05266, po05267, po05268, po05269, po05270, po05271, po05272, po05273, po05274, po05275, po05276, po05277, po05278, po05279, po05280, po05281, po05282, po05283, po05284, po05285, po05286, po05287, po05288, po05289, po05290, po05291, po05292, po05293, po05294, po05295, po05296, po05297, po05298, po05299, po05300, po05301, po05302, po05303, po05304, po05305, po05306, po05307, po05308, po05309, po05310, po05311, po05312, po05313, po05314, po05315, po05316, po05317, po05318, po05319, po05320, po05321, po05322, po05323, po05324, po05325, po05326, po05327, po05328, po05329, po05330, po05331, po05332, po05333, po05334, po05335, po05336, po05337, po05338, po05339, po05340, po05341, po05342, po05343, po05344, po05345, po05346, po05347, po05348, po05349, po05350, po05351, po05352, po05353, po05354, po05355, po05356, po05357, po05358, po05359, po05360, po05361, po05362, po05363, po05364, po05365, po05366, po05367, po05368, po05369, po05370, po05371, po05372, po05373, po05374, po05375, po05376, po05377, po05378, po05379, po05380, po05381, po05382, po05383, po05384, po05385, po05386, po05387, po05388, po05389, po05390, po05391, po05392, po05393, po05394, po05395, po05396, po05397, po05398, po05399, po05400, po05401, po05402, po05403, po05404, po05405, po05406, po05407, po05408, po05409, po05410, po05411, po05412, po05413, po05414, po05415, po05416, po05417, po05418, po05419, po05420, po05421, po05422, po05423, po05424, po05425, po05426, po05427, po05428, po05429, po05430, po05431, po05432, po05433, po05434, po05435, po05436, po05437, po05438, po05439, po05440, po05441, po05442, po05443, po05444, po05445, po05446, po05447, po05448, po05449, po05450, po05451, po05452, po05453, po05454, po05455, po05456, po05457, po05458, po05459, po05460, po05461, po05462, po05463, po05464, po05465, po05466, po05467, po05468, po05469, po05470, po05471, po05472, po05473, po05474, po05475, po05476, po05477, po05478, po05479, po05480, po05481, po05482, po05483, po05484, po05485, po05486, po05487, po05488, po05489, po05490, po05491, po05492, po05493, po05494, po05495, po05496, po05497, po05498, po05499, po05500, po05501, po05502, po05503, po05504, po05505, po05506, po05507, po05508, po05509, po05510, po05511, po05512, po05513, po05514, po05515, po05516, po05517, po05518, po05519, po05520, po05521, po05522, po05523, po05524, po05525, po05526, po05527, po05528, po05529, po05530, po05531, po05532, po05533, po05534, po05535, po05536, po05537, po05538, po05539, po05540, po05541, po05542, po05543, po05544, po05545, po05546, po05547, po05548, po05549, po05550, po05551, po05552, po05553, po05554, po05555, po05556, po05557, po05558, po05559, po05560, po05561, po05562, po05563, po05564, po05565, po05566, po05567, po05568, po05569, po05570, po05571, po05572, po05573, po05574, po05575, po05576, po05577, po05578, po05579, po05580, po05581, po05582, po05583, po05584, po05585, po05586, po05587, po05588, po05589, po05590, po05591, po05592, po05593, po05594, po05595, po05596, po05597, po05598, po05599, po05600, po05601, po05602, po05603, po05604, po05605, po05606, po05607, po05608, po05609, po05610, po05611, po05612, po05613, po05614, po05615, po05616, po05617, po05618, po05619, po05620, po05621, po05622, po05623, po05624, po05625, po05626, po05627, po05628, po05629, po05630, po05631, po05632, po05633, po05634, po05635, po05636, po05637, po05638, po05639, po05640, po05641, po05642, po05643, po05644, po05645, po05646, po05647, po05648, po05649, po05650, po05651, po05652, po05653, po05654, po05655, po05656, po05657, po05658, po05659, po05660, po05661, po05662, po05663, po05664, po05665, po05666, po05667, po05668, po05669, po05670, po05671, po05672, po05673, po05674, po05675, po05676, po05677, po05678, po05679, po05680, po05681, po05682, po05683, po05684, po05685, po05686, po05687, po05688, po05689, po05690, po05691, po05692, po05693, po05694, po05695, po05696, po05697, po05698, po05699, po05700, po05701, po05702, po05703, po05704, po05705, po05706, po05707, po05708, po05709, po05710, po05711, po05712, po05713, po05714, po05715, po05716, po05717, po05718, po05719, po05720, po05721, po05722, po05723, po05724, po05725, po05726, po05727, po05728, po05729, po05730, po05731, po05732, po05733, po05734, po05735, po05736, po05737, po05738, po05739, po05740, po05741, po05742, po05743, po05744, po05745, po05746, po05747, po05748, po05749, po05750, po05751, po05752, po05753, po05754, po05755, po05756, po05757, po05758, po05759, po05760, po05761, po05762, po05763, po05764, po05765, po05766, po05767, po05768, po05769, po05770, po05771, po05772, po05773, po05774, po05775, po05776, po05777, po05778, po05779, po05780, po05781, po05782, po05783, po05784, po05785, po05786, po05787, po05788, po05789, po05790, po05791, po05792, po05793, po05794, po05795, po05796, po05797, po05798, po05799, po05800, po05801, po05802, po05803, po05804, po05805, po05806, po05807, po05808, po05809, po05810, po05811, po05812, po05813, po05814, po05815, po05816, po05817, po05818, po05819, po05820, po05821, po05822, po05823, po05824, po05825, po05826, po05827, po05828, po05829, po05830, po05831, po05832, po05833, po05834, po05835, po05836, po05837, po05838, po05839, po05840, po05841, po05842, po05843, po05844, po05845, po05846, po05847, po05848, po05849, po05850, po05851, po05852, po05853, po05854, po05855, po05856, po05857, po05858, po05859, po05860, po05861, po05862, po05863, po05864, po05865, po05866, po05867, po05868, po05869, po05870, po05871, po05872, po05873, po05874, po05875, po05876, po05877, po05878, po05879, po05880, po05881, po05882, po05883, po05884, po05885, po05886, po05887, po05888, po05889, po05890, po05891, po05892, po05893, po05894, po05895, po05896, po05897, po05898, po05899, po05900, po05901, po05902, po05903, po05904, po05905, po05906, po05907, po05908, po05909, po05910, po05911, po05912, po05913, po05914, po05915, po05916, po05917, po05918, po05919, po05920, po05921, po05922, po05923, po05924, po05925, po05926, po05927, po05928, po05929, po05930, po05931, po05932, po05933, po05934, po05935, po05936, po05937, po05938, po05939, po05940, po05941, po05942, po05943, po05944, po05945, po05946, po05947, po05948, po05949, po05950, po05951, po05952, po05953, po05954, po05955, po05956, po05957, po05958, po05959, po05960, po05961, po05962, po05963, po05964, po05965, po05966, po05967, po05968, po05969, po05970, po05971, po05972, po05973, po05974, po05975, po05976, po05977, po05978, po05979, po05980, po05981, po05982, po05983, po05984, po05985, po05986, po05987, po05988, po05989, po05990, po05991, po05992, po05993, po05994, po05995, po05996, po05997, po05998, po05999, po06000, po06001, po06002, po06003, po06004, po06005, po06006, po06007, po06008, po06009, po06010, po06011, po06012, po06013, po06014, po06015, po06016, po06017, po06018, po06019, po06020, po06021, po06022, po06023, po06024, po06025, po06026, po06027, po06028, po06029, po06030, po06031, po06032, po06033, po06034, po06035, po06036, po06037, po06038, po06039, po06040, po06041, po06042, po06043, po06044, po06045, po06046, po06047, po06048, po06049, po06050, po06051, po06052, po06053, po06054, po06055, po06056, po06057, po06058, po06059, po06060, po06061, po06062, po06063, po06064, po06065, po06066, po06067, po06068, po06069, po06070, po06071, po06072, po06073, po06074, po06075, po06076, po06077, po06078, po06079, po06080, po06081, po06082, po06083, po06084, po06085, po06086, po06087, po06088, po06089, po06090, po06091, po06092, po06093, po06094, po06095, po06096, po06097, po06098, po06099, po06100, po06101, po06102, po06103, po06104, po06105, po06106, po06107, po06108, po06109, po06110, po06111, po06112, po06113, po06114, po06115, po06116, po06117, po06118, po06119, po06120, po06121, po06122, po06123, po06124, po06125, po06126, po06127, po06128, po06129, po06130, po06131, po06132, po06133, po06134, po06135, po06136, po06137, po06138, po06139, po06140, po06141, po06142, po06143, po06144, po06145, po06146, po06147, po06148, po06149, po06150, po06151, po06152, po06153, po06154, po06155, po06156, po06157, po06158, po06159, po06160, po06161, po06162, po06163, po06164, po06165, po06166, po06167, po06168, po06169, po06170, po06171, po06172, po06173, po06174, po06175, po06176, po06177, po06178, po06179, po06180, po06181, po06182, po06183, po06184, po06185, po06186, po06187, po06188, po06189, po06190, po06191, po06192, po06193, po06194, po06195, po06196, po06197, po06198, po06199, po06200, po06201, po06202, po06203, po06204, po06205, po06206, po06207, po06208, po06209, po06210, po06211, po06212, po06213, po06214, po06215, po06216, po06217, po06218, po06219, po06220, po06221, po06222, po06223, po06224, po06225, po06226, po06227, po06228, po06229, po06230, po06231, po06232, po06233, po06234, po06235, po06236, po06237, po06238, po06239, po06240, po06241, po06242, po06243, po06244, po06245, po06246, po06247, po06248, po06249, po06250, po06251, po06252, po06253, po06254, po06255, po06256, po06257, po06258, po06259, po06260, po06261, po06262, po06263, po06264, po06265, po06266, po06267, po06268, po06269, po06270, po06271, po06272, po06273, po06274, po06275, po06276, po06277, po06278, po06279, po06280, po06281, po06282, po06283, po06284, po06285, po06286, po06287, po06288, po06289, po06290, po06291, po06292, po06293, po06294, po06295, po06296, po06297, po06298, po06299, po06300, po06301, po06302, po06303, po06304, po06305, po06306, po06307, po06308, po06309, po06310, po06311, po06312, po06313, po06314, po06315, po06316, po06317, po06318, po06319, po06320, po06321, po06322, po06323, po06324, po06325, po06326, po06327, po06328, po06329, po06330, po06331, po06332, po06333, po06334, po06335, po06336, po06337, po06338, po06339, po06340, po06341, po06342, po06343, po06344, po06345, po06346, po06347, po06348, po06349, po06350, po06351, po06352, po06353, po06354, po06355, po06356, po06357, po06358, po06359, po06360, po06361, po06362, po06363, po06364, po06365, po06366, po06367, po06368, po06369, po06370, po06371, po06372, po06373, po06374, po06375, po06376, po06377, po06378, po06379, po06380, po06381, po06382, po06383, po06384, po06385, po06386, po06387, po06388, po06389, po06390, po06391, po06392, po06393, po06394, po06395, po06396, po06397, po06398, po06399, po06400, po06401, po06402, po06403, po06404, po06405, po06406, po06407, po06408, po06409, po06410, po06411, po06412, po06413, po06414, po06415, po06416, po06417, po06418, po06419, po06420, po06421, po06422, po06423, po06424, po06425, po06426, po06427, po06428, po06429, po06430, po06431, po06432, po06433, po06434, po06435, po06436, po06437, po06438, po06439, po06440, po06441, po06442, po06443, po06444, po06445, po06446, po06447, po06448, po06449, po06450, po06451, po06452, po06453, po06454, po06455, po06456, po06457, po06458, po06459, po06460, po06461, po06462, po06463, po06464, po06465, po06466, po06467, po06468, po06469, po06470, po06471, po06472, po06473, po06474, po06475, po06476, po06477, po06478, po06479, po06480, po06481, po06482, po06483, po06484, po06485, po06486, po06487, po06488, po06489, po06490, po06491, po06492, po06493, po06494, po06495, po06496, po06497, po06498, po06499, po06500, po06501, po06502, po06503, po06504, po06505, po06506, po06507, po06508, po06509, po06510, po06511, po06512, po06513, po06514, po06515, po06516, po06517, po06518, po06519, po06520, po06521, po06522, po06523, po06524, po06525, po06526, po06527, po06528, po06529, po06530, po06531, po06532, po06533, po06534, po06535, po06536, po06537, po06538, po06539, po06540, po06541, po06542, po06543, po06544, po06545, po06546, po06547, po06548, po06549, po06550, po06551, po06552, po06553, po06554, po06555, po06556, po06557, po06558, po06559, po06560, po06561, po06562, po06563, po06564, po06565, po06566, po06567, po06568, po06569, po06570, po06571, po06572, po06573, po06574, po06575, po06576, po06577, po06578, po06579, po06580, po06581, po06582, po06583, po06584, po06585, po06586, po06587, po06588, po06589, po06590, po06591, po06592, po06593, po06594, po06595, po06596, po06597, po06598, po06599, po06600, po06601, po06602, po06603, po06604, po06605, po06606, po06607, po06608, po06609, po06610, po06611, po06612, po06613, po06614, po06615, po06616, po06617, po06618, po06619, po06620, po06621, po06622, po06623, po06624, po06625, po06626, po06627, po06628, po06629, po06630, po06631, po06632, po06633, po06634, po06635, po06636, po06637, po06638, po06639, po06640, po06641, po06642, po06643, po06644, po06645, po06646, po06647, po06648, po06649, po06650, po06651, po06652, po06653, po06654, po06655, po06656, po06657, po06658, po06659, po06660, po06661, po06662, po06663, po06664, po06665, po06666, po06667, po06668, po06669, po06670, po06671, po06672, po06673, po06674, po06675, po06676, po06677, po06678, po06679, po06680, po06681, po06682, po06683, po06684, po06685, po06686, po06687, po06688, po06689, po06690, po06691, po06692, po06693, po06694, po06695, po06696, po06697, po06698, po06699, po06700, po06701, po06702, po06703, po06704, po06705, po06706, po06707, po06708, po06709, po06710, po06711, po06712, po06713, po06714, po06715, po06716, po06717, po06718, po06719, po06720, po06721, po06722, po06723, po06724, po06725, po06726, po06727, po06728, po06729, po06730, po06731, po06732, po06733, po06734, po06735, po06736, po06737, po06738, po06739, po06740, po06741, po06742, po06743, po06744, po06745, po06746, po06747, po06748, po06749, po06750, po06751, po06752, po06753, po06754, po06755, po06756, po06757, po06758, po06759, po06760, po06761, po06762, po06763, po06764, po06765, po06766, po06767, po06768, po06769, po06770, po06771, po06772, po06773, po06774, po06775, po06776, po06777, po06778, po06779, po06780, po06781, po06782, po06783, po06784, po06785, po06786, po06787, po06788, po06789, po06790, po06791, po06792, po06793, po06794, po06795, po06796, po06797, po06798, po06799, po06800, po06801, po06802, po06803, po06804, po06805, po06806, po06807, po06808, po06809, po06810, po06811, po06812, po06813, po06814, po06815, po06816, po06817, po06818, po06819, po06820, po06821, po06822, po06823, po06824, po06825, po06826, po06827, po06828, po06829, po06830, po06831, po06832, po06833, po06834, po06835, po06836, po06837, po06838, po06839, po06840, po06841, po06842, po06843, po06844, po06845, po06846, po06847, po06848, po06849, po06850, po06851, po06852, po06853, po06854, po06855, po06856, po06857, po06858, po06859, po06860, po06861, po06862, po06863, po06864, po06865, po06866, po06867, po06868, po06869, po06870, po06871, po06872, po06873, po06874, po06875, po06876, po06877, po06878, po06879, po06880, po06881, po06882, po06883, po06884, po06885, po06886, po06887, po06888, po06889, po06890, po06891, po06892, po06893, po06894, po06895, po06896, po06897, po06898, po06899, po06900, po06901, po06902, po06903, po06904, po06905, po06906, po06907, po06908, po06909, po06910, po06911, po06912, po06913, po06914, po06915, po06916, po06917, po06918, po06919, po06920, po06921, po06922, po06923, po06924, po06925, po06926, po06927, po06928, po06929, po06930, po06931, po06932, po06933, po06934, po06935, po06936, po06937, po06938, po06939, po06940, po06941, po06942, po06943, po06944, po06945, po06946, po06947, po06948, po06949, po06950, po06951, po06952, po06953, po06954, po06955, po06956, po06957, po06958, po06959, po06960, po06961, po06962, po06963, po06964, po06965, po06966, po06967, po06968, po06969, po06970, po06971, po06972, po06973, po06974, po06975, po06976, po06977, po06978, po06979, po06980, po06981, po06982, po06983, po06984, po06985, po06986, po06987, po06988, po06989, po06990, po06991, po06992, po06993, po06994, po06995, po06996, po06997, po06998, po06999, po07000, po07001, po07002, po07003, po07004, po07005, po07006, po07007, po07008, po07009, po07010, po07011, po07012, po07013, po07014, po07015, po07016, po07017, po07018, po07019, po07020, po07021, po07022, po07023, po07024, po07025, po07026, po07027, po07028, po07029, po07030, po07031, po07032, po07033, po07034, po07035, po07036, po07037, po07038, po07039, po07040, po07041, po07042, po07043, po07044, po07045, po07046, po07047, po07048, po07049, po07050, po07051, po07052, po07053, po07054, po07055, po07056, po07057, po07058, po07059, po07060, po07061, po07062, po07063, po07064, po07065, po07066, po07067, po07068, po07069, po07070, po07071, po07072, po07073, po07074, po07075, po07076, po07077, po07078, po07079, po07080, po07081, po07082, po07083, po07084, po07085, po07086, po07087, po07088, po07089, po07090, po07091, po07092, po07093, po07094, po07095, po07096, po07097, po07098, po07099, po07100, po07101, po07102, po07103, po07104, po07105, po07106, po07107, po07108, po07109, po07110, po07111, po07112, po07113, po07114, po07115, po07116, po07117, po07118, po07119, po07120, po07121, po07122, po07123, po07124, po07125, po07126, po07127, po07128, po07129, po07130, po07131, po07132, po07133, po07134, po07135, po07136, po07137, po07138, po07139, po07140, po07141, po07142, po07143, po07144, po07145, po07146, po07147, po07148, po07149, po07150, po07151, po07152, po07153, po07154, po07155, po07156, po07157, po07158, po07159, po07160, po07161, po07162, po07163, po07164, po07165, po07166, po07167, po07168, po07169, po07170, po07171, po07172, po07173, po07174, po07175, po07176, po07177, po07178, po07179, po07180, po07181, po07182, po07183, po07184, po07185, po07186, po07187, po07188, po07189, po07190, po07191, po07192, po07193, po07194, po07195, po07196, po07197, po07198, po07199, po07200, po07201, po07202, po07203, po07204, po07205, po07206, po07207, po07208, po07209, po07210, po07211, po07212, po07213, po07214, po07215, po07216, po07217, po07218, po07219, po07220, po07221, po07222, po07223, po07224, po07225, po07226, po07227, po07228, po07229, po07230, po07231, po07232, po07233, po07234, po07235, po07236, po07237, po07238, po07239, po07240, po07241, po07242, po07243, po07244, po07245, po07246, po07247, po07248, po07249, po07250, po07251, po07252, po07253, po07254, po07255, po07256, po07257, po07258, po07259, po07260, po07261, po07262, po07263, po07264, po07265, po07266, po07267, po07268, po07269, po07270, po07271, po07272, po07273, po07274, po07275, po07276, po07277, po07278, po07279, po07280, po07281, po07282, po07283, po07284, po07285, po07286, po07287, po07288, po07289, po07290, po07291, po07292, po07293, po07294, po07295, po07296, po07297, po07298, po07299, po07300, po07301, po07302, po07303, po07304, po07305, po07306, po07307, po07308, po07309, po07310, po07311, po07312, po07313, po07314, po07315, po07316, po07317, po07318, po07319, po07320, po07321, po07322, po07323, po07324, po07325, po07326, po07327, po07328, po07329, po07330, po07331, po07332, po07333, po07334, po07335, po07336, po07337, po07338, po07339, po07340, po07341, po07342, po07343, po07344, po07345, po07346, po07347, po07348, po07349, po07350, po07351, po07352, po07353, po07354, po07355, po07356, po07357, po07358, po07359, po07360, po07361, po07362, po07363, po07364, po07365, po07366, po07367, po07368, po07369, po07370, po07371, po07372, po07373, po07374, po07375, po07376, po07377, po07378, po07379, po07380, po07381, po07382, po07383, po07384, po07385, po07386, po07387, po07388, po07389, po07390, po07391, po07392, po07393, po07394, po07395, po07396, po07397, po07398, po07399, po07400, po07401, po07402, po07403, po07404, po07405, po07406, po07407, po07408, po07409, po07410, po07411, po07412, po07413, po07414, po07415, po07416, po07417, po07418, po07419, po07420, po07421, po07422, po07423, po07424, po07425, po07426, po07427, po07428, po07429, po07430, po07431, po07432, po07433, po07434, po07435, po07436, po07437, po07438, po07439, po07440, po07441, po07442, po07443, po07444, po07445, po07446, po07447, po07448, po07449, po07450, po07451, po07452, po07453, po07454, po07455, po07456, po07457, po07458, po07459, po07460, po07461, po07462, po07463, po07464, po07465, po07466, po07467, po07468, po07469, po07470, po07471, po07472, po07473, po07474, po07475, po07476, po07477, po07478, po07479, po07480, po07481, po07482, po07483, po07484, po07485, po07486, po07487, po07488, po07489, po07490, po07491, po07492, po07493, po07494, po07495, po07496, po07497, po07498, po07499, po07500, po07501, po07502, po07503, po07504, po07505, po07506, po07507, po07508, po07509, po07510, po07511, po07512, po07513, po07514, po07515, po07516, po07517, po07518, po07519, po07520, po07521, po07522, po07523, po07524, po07525, po07526, po07527, po07528, po07529, po07530, po07531, po07532, po07533, po07534, po07535, po07536, po07537, po07538, po07539, po07540, po07541, po07542, po07543, po07544, po07545, po07546, po07547, po07548, po07549, po07550, po07551, po07552, po07553, po07554, po07555, po07556, po07557, po07558, po07559, po07560, po07561, po07562, po07563, po07564, po07565, po07566, po07567, po07568, po07569, po07570, po07571, po07572, po07573, po07574, po07575, po07576, po07577, po07578, po07579, po07580, po07581, po07582, po07583, po07584, po07585, po07586, po07587, po07588, po07589, po07590, po07591, po07592, po07593, po07594, po07595, po07596, po07597, po07598, po07599, po07600, po07601, po07602, po07603, po07604, po07605, po07606, po07607, po07608, po07609, po07610, po07611, po07612, po07613, po07614, po07615, po07616, po07617, po07618, po07619, po07620, po07621, po07622, po07623, po07624, po07625, po07626, po07627, po07628, po07629, po07630, po07631, po07632, po07633, po07634, po07635, po07636, po07637, po07638, po07639, po07640, po07641, po07642, po07643, po07644, po07645, po07646, po07647, po07648, po07649, po07650, po07651, po07652, po07653, po07654, po07655, po07656, po07657, po07658, po07659, po07660, po07661, po07662, po07663, po07664, po07665, po07666, po07667, po07668, po07669, po07670, po07671, po07672, po07673, po07674, po07675, po07676, po07677, po07678, po07679, po07680, po07681, po07682, po07683, po07684, po07685, po07686, po07687, po07688, po07689, po07690, po07691, po07692, po07693, po07694, po07695, po07696, po07697, po07698, po07699, po07700, po07701, po07702, po07703, po07704, po07705, po07706, po07707, po07708, po07709, po07710, po07711, po07712, po07713, po07714, po07715, po07716, po07717, po07718, po07719, po07720, po07721, po07722, po07723, po07724, po07725, po07726, po07727, po07728, po07729, po07730, po07731, po07732, po07733, po07734, po07735, po07736, po07737, po07738, po07739, po07740, po07741, po07742, po07743, po07744, po07745, po07746, po07747, po07748, po07749, po07750, po07751, po07752, po07753, po07754, po07755, po07756, po07757, po07758, po07759, po07760, po07761, po07762, po07763, po07764, po07765, po07766, po07767, po07768, po07769, po07770, po07771, po07772, po07773, po07774, po07775, po07776, po07777, po07778, po07779, po07780, po07781, po07782, po07783, po07784, po07785, po07786, po07787, po07788, po07789, po07790, po07791, po07792, po07793, po07794, po07795, po07796, po07797, po07798, po07799, po07800, po07801, po07802, po07803, po07804, po07805, po07806, po07807, po07808, po07809, po07810, po07811, po07812, po07813, po07814, po07815, po07816, po07817, po07818, po07819, po07820, po07821, po07822, po07823, po07824, po07825, po07826, po07827, po07828, po07829, po07830, po07831, po07832, po07833, po07834, po07835, po07836, po07837, po07838, po07839, po07840, po07841, po07842, po07843, po07844, po07845, po07846, po07847, po07848, po07849, po07850, po07851, po07852, po07853, po07854, po07855, po07856, po07857, po07858, po07859, po07860, po07861, po07862, po07863, po07864, po07865, po07866, po07867, po07868, po07869, po07870, po07871, po07872, po07873, po07874, po07875, po07876, po07877, po07878, po07879, po07880, po07881, po07882, po07883, po07884, po07885, po07886, po07887, po07888, po07889, po07890, po07891, po07892, po07893, po07894, po07895, po07896, po07897, po07898, po07899, po07900, po07901, po07902, po07903, po07904, po07905, po07906, po07907, po07908, po07909, po07910, po07911, po07912, po07913, po07914, po07915, po07916, po07917, po07918, po07919, po07920, po07921, po07922, po07923, po07924, po07925, po07926, po07927, po07928, po07929, po07930, po07931, po07932, po07933, po07934, po07935, po07936, po07937, po07938, po07939, po07940, po07941, po07942, po07943, po07944, po07945, po07946, po07947, po07948, po07949, po07950, po07951, po07952, po07953, po07954, po07955, po07956, po07957, po07958, po07959, po07960, po07961, po07962, po07963, po07964, po07965, po07966, po07967, po07968, po07969, po07970, po07971, po07972, po07973, po07974, po07975, po07976, po07977, po07978, po07979, po07980, po07981, po07982, po07983, po07984, po07985, po07986, po07987, po07988, po07989, po07990, po07991, po07992, po07993, po07994, po07995, po07996, po07997, po07998, po07999, po08000, po08001, po08002, po08003, po08004, po08005, po08006, po08007, po08008, po08009, po08010, po08011, po08012, po08013, po08014, po08015, po08016, po08017, po08018, po08019, po08020, po08021, po08022, po08023, po08024, po08025, po08026, po08027, po08028, po08029, po08030, po08031, po08032, po08033, po08034, po08035, po08036, po08037, po08038, po08039, po08040, po08041, po08042, po08043, po08044, po08045, po08046, po08047, po08048, po08049, po08050, po08051, po08052, po08053, po08054, po08055, po08056, po08057, po08058, po08059, po08060, po08061, po08062, po08063, po08064, po08065, po08066, po08067, po08068, po08069, po08070, po08071, po08072, po08073, po08074, po08075, po08076, po08077, po08078, po08079, po08080, po08081, po08082, po08083, po08084, po08085, po08086, po08087, po08088, po08089, po08090, po08091, po08092, po08093, po08094, po08095, po08096, po08097, po08098, po08099, po08100, po08101, po08102, po08103, po08104, po08105, po08106, po08107, po08108, po08109, po08110, po08111, po08112, po08113, po08114, po08115, po08116, po08117, po08118, po08119, po08120, po08121, po08122, po08123, po08124, po08125, po08126, po08127, po08128, po08129, po08130, po08131, po08132, po08133, po08134, po08135, po08136, po08137, po08138, po08139, po08140, po08141, po08142, po08143, po08144, po08145, po08146, po08147, po08148, po08149, po08150, po08151, po08152, po08153, po08154, po08155, po08156, po08157, po08158, po08159, po08160, po08161, po08162, po08163, po08164, po08165, po08166, po08167, po08168, po08169, po08170, po08171, po08172, po08173, po08174, po08175, po08176, po08177, po08178, po08179, po08180, po08181, po08182, po08183, po08184, po08185, po08186, po08187, po08188, po08189, po08190, po08191, po08192, po08193, po08194, po08195, po08196, po08197, po08198, po08199, po08200, po08201, po08202, po08203, po08204, po08205, po08206, po08207, po08208, po08209, po08210, po08211, po08212, po08213, po08214, po08215, po08216, po08217, po08218, po08219, po08220, po08221, po08222, po08223, po08224, po08225, po08226, po08227, po08228, po08229, po08230, po08231, po08232, po08233, po08234, po08235, po08236, po08237, po08238, po08239, po08240, po08241, po08242, po08243, po08244, po08245, po08246, po08247, po08248, po08249, po08250, po08251, po08252, po08253, po08254, po08255, po08256, po08257, po08258, po08259, po08260, po08261, po08262, po08263, po08264, po08265, po08266, po08267, po08268, po08269, po08270, po08271, po08272, po08273, po08274, po08275, po08276, po08277, po08278, po08279, po08280, po08281, po08282, po08283, po08284, po08285, po08286, po08287, po08288, po08289, po08290, po08291, po08292, po08293, po08294, po08295, po08296, po08297, po08298, po08299, po08300, po08301, po08302, po08303, po08304, po08305, po08306, po08307, po08308, po08309, po08310, po08311, po08312, po08313, po08314, po08315, po08316, po08317, po08318, po08319, po08320, po08321, po08322, po08323, po08324, po08325, po08326, po08327, po08328, po08329, po08330, po08331, po08332, po08333, po08334, po08335, po08336, po08337, po08338, po08339, po08340, po08341, po08342, po08343, po08344, po08345, po08346, po08347, po08348, po08349, po08350, po08351, po08352, po08353, po08354, po08355, po08356, po08357, po08358, po08359, po08360, po08361, po08362, po08363, po08364, po08365, po08366, po08367, po08368, po08369, po08370, po08371, po08372, po08373, po08374, po08375, po08376, po08377, po08378, po08379, po08380, po08381, po08382, po08383, po08384, po08385, po08386, po08387, po08388, po08389, po08390, po08391, po08392, po08393, po08394, po08395, po08396, po08397, po08398, po08399, po08400, po08401, po08402, po08403, po08404, po08405, po08406, po08407, po08408, po08409, po08410, po08411, po08412, po08413, po08414, po08415, po08416, po08417, po08418, po08419, po08420, po08421, po08422, po08423, po08424, po08425, po08426, po08427, po08428, po08429, po08430, po08431, po08432, po08433, po08434, po08435, po08436, po08437, po08438, po08439, po08440, po08441, po08442, po08443, po08444, po08445, po08446, po08447, po08448, po08449, po08450, po08451, po08452, po08453, po08454, po08455, po08456, po08457, po08458, po08459, po08460, po08461, po08462, po08463, po08464, po08465, po08466, po08467, po08468, po08469, po08470, po08471, po08472, po08473, po08474, po08475, po08476, po08477, po08478, po08479, po08480, po08481, po08482, po08483, po08484, po08485, po08486, po08487, po08488, po08489, po08490, po08491, po08492, po08493, po08494, po08495, po08496, po08497, po08498, po08499, po08500, po08501, po08502, po08503, po08504, po08505, po08506, po08507, po08508, po08509, po08510, po08511, po08512, po08513, po08514, po08515, po08516, po08517, po08518, po08519, po08520, po08521, po08522, po08523, po08524, po08525, po08526, po08527, po08528, po08529, po08530, po08531, po08532, po08533, po08534, po08535, po08536, po08537, po08538, po08539, po08540, po08541, po08542, po08543, po08544, po08545, po08546, po08547, po08548, po08549, po08550, po08551, po08552, po08553, po08554, po08555, po08556, po08557, po08558, po08559, po08560, po08561, po08562, po08563, po08564, po08565, po08566, po08567, po08568, po08569, po08570, po08571, po08572, po08573, po08574, po08575, po08576, po08577, po08578, po08579, po08580, po08581, po08582, po08583, po08584, po08585, po08586, po08587, po08588, po08589, po08590, po08591, po08592, po08593, po08594, po08595, po08596, po08597, po08598, po08599, po08600, po08601, po08602, po08603, po08604, po08605, po08606, po08607, po08608, po08609, po08610, po08611, po08612, po08613, po08614, po08615, po08616, po08617, po08618, po08619, po08620, po08621, po08622, po08623, po08624, po08625, po08626, po08627, po08628, po08629, po08630, po08631, po08632, po08633, po08634, po08635, po08636, po08637, po08638, po08639, po08640, po08641, po08642, po08643, po08644, po08645, po08646, po08647, po08648, po08649, po08650, po08651, po08652, po08653, po08654, po08655, po08656, po08657, po08658, po08659, po08660, po08661, po08662, po08663, po08664, po08665, po08666, po08667, po08668, po08669, po08670, po08671, po08672, po08673, po08674, po08675, po08676, po08677, po08678, po08679, po08680, po08681, po08682, po08683, po08684, po08685, po08686, po08687, po08688, po08689, po08690, po08691, po08692, po08693, po08694, po08695, po08696, po08697, po08698, po08699, po08700, po08701, po08702, po08703, po08704, po08705, po08706, po08707, po08708, po08709, po08710, po08711, po08712, po08713, po08714, po08715, po08716, po08717, po08718, po08719, po08720, po08721, po08722, po08723, po08724, po08725, po08726, po08727, po08728, po08729, po08730, po08731, po08732, po08733, po08734, po08735, po08736, po08737, po08738, po08739, po08740, po08741, po08742, po08743, po08744, po08745, po08746, po08747, po08748, po08749, po08750, po08751, po08752, po08753, po08754, po08755, po08756, po08757, po08758, po08759, po08760, po08761, po08762, po08763, po08764, po08765, po08766, po08767, po08768, po08769, po08770, po08771, po08772, po08773, po08774, po08775, po08776, po08777, po08778, po08779, po08780, po08781, po08782, po08783, po08784, po08785, po08786, po08787, po08788, po08789, po08790, po08791, po08792, po08793, po08794, po08795, po08796, po08797, po08798, po08799, po08800, po08801, po08802, po08803, po08804, po08805, po08806, po08807, po08808, po08809, po08810, po08811, po08812, po08813, po08814, po08815, po08816, po08817, po08818, po08819, po08820, po08821, po08822, po08823, po08824, po08825, po08826, po08827, po08828, po08829, po08830, po08831, po08832, po08833, po08834, po08835, po08836, po08837, po08838, po08839, po08840, po08841, po08842, po08843, po08844, po08845, po08846, po08847, po08848, po08849, po08850, po08851, po08852, po08853, po08854, po08855, po08856, po08857, po08858, po08859, po08860, po08861, po08862, po08863, po08864, po08865, po08866, po08867, po08868, po08869, po08870, po08871, po08872, po08873, po08874, po08875, po08876, po08877, po08878, po08879, po08880, po08881, po08882, po08883, po08884, po08885, po08886, po08887, po08888, po08889, po08890, po08891, po08892, po08893, po08894, po08895, po08896, po08897, po08898, po08899, po08900, po08901, po08902, po08903, po08904, po08905, po08906, po08907, po08908, po08909, po08910, po08911, po08912, po08913, po08914, po08915, po08916, po08917, po08918, po08919, po08920, po08921, po08922, po08923, po08924, po08925, po08926, po08927, po08928, po08929, po08930, po08931, po08932, po08933, po08934, po08935, po08936, po08937, po08938, po08939, po08940, po08941, po08942, po08943, po08944, po08945, po08946, po08947, po08948, po08949, po08950, po08951, po08952, po08953, po08954, po08955, po08956, po08957, po08958, po08959, po08960, po08961, po08962, po08963, po08964, po08965, po08966, po08967, po08968, po08969, po08970, po08971, po08972, po08973, po08974, po08975, po08976, po08977, po08978, po08979, po08980, po08981, po08982, po08983, po08984, po08985, po08986, po08987, po08988, po08989, po08990, po08991, po08992, po08993, po08994, po08995, po08996, po08997, po08998, po08999, po09000, po09001, po09002, po09003, po09004, po09005, po09006, po09007, po09008, po09009, po09010, po09011, po09012, po09013, po09014, po09015, po09016, po09017, po09018, po09019, po09020, po09021, po09022, po09023, po09024, po09025, po09026, po09027, po09028, po09029, po09030, po09031, po09032, po09033, po09034, po09035, po09036, po09037, po09038, po09039, po09040, po09041, po09042, po09043, po09044, po09045, po09046, po09047, po09048, po09049, po09050, po09051, po09052, po09053, po09054, po09055, po09056, po09057, po09058, po09059, po09060, po09061, po09062, po09063, po09064, po09065, po09066, po09067, po09068, po09069, po09070, po09071, po09072, po09073, po09074, po09075, po09076, po09077, po09078, po09079, po09080, po09081, po09082, po09083, po09084, po09085, po09086, po09087, po09088, po09089, po09090, po09091, po09092, po09093, po09094, po09095, po09096, po09097, po09098, po09099, po09100, po09101, po09102, po09103, po09104, po09105, po09106, po09107, po09108, po09109, po09110, po09111, po09112, po09113, po09114, po09115, po09116, po09117, po09118, po09119, po09120, po09121, po09122, po09123, po09124, po09125, po09126, po09127, po09128, po09129, po09130, po09131, po09132, po09133, po09134, po09135, po09136, po09137, po09138, po09139, po09140, po09141, po09142, po09143, po09144, po09145, po09146, po09147, po09148, po09149, po09150, po09151, po09152, po09153, po09154, po09155, po09156, po09157, po09158, po09159, po09160, po09161, po09162, po09163, po09164, po09165, po09166, po09167, po09168, po09169, po09170, po09171, po09172, po09173, po09174, po09175, po09176, po09177, po09178, po09179, po09180, po09181, po09182, po09183, po09184, po09185, po09186, po09187, po09188, po09189, po09190, po09191, po09192, po09193, po09194, po09195, po09196, po09197, po09198, po09199, po09200, po09201, po09202, po09203, po09204, po09205, po09206, po09207, po09208, po09209, po09210, po09211, po09212, po09213, po09214, po09215, po09216, po09217, po09218, po09219, po09220, po09221, po09222, po09223, po09224, po09225, po09226, po09227, po09228, po09229, po09230, po09231, po09232, po09233, po09234, po09235, po09236, po09237, po09238, po09239, po09240, po09241, po09242, po09243, po09244, po09245, po09246, po09247, po09248, po09249, po09250, po09251, po09252, po09253, po09254, po09255, po09256, po09257, po09258, po09259, po09260, po09261, po09262, po09263, po09264, po09265, po09266, po09267, po09268, po09269, po09270, po09271, po09272, po09273, po09274, po09275, po09276, po09277, po09278, po09279, po09280, po09281, po09282, po09283, po09284, po09285, po09286, po09287, po09288, po09289, po09290, po09291, po09292, po09293, po09294, po09295, po09296, po09297, po09298, po09299, po09300, po09301, po09302, po09303, po09304, po09305, po09306, po09307, po09308, po09309, po09310, po09311, po09312, po09313, po09314, po09315, po09316, po09317, po09318, po09319, po09320, po09321, po09322, po09323, po09324, po09325, po09326, po09327, po09328, po09329, po09330, po09331, po09332, po09333, po09334, po09335, po09336, po09337, po09338, po09339, po09340, po09341, po09342, po09343, po09344, po09345, po09346, po09347, po09348, po09349, po09350, po09351, po09352, po09353, po09354, po09355, po09356, po09357, po09358, po09359, po09360, po09361, po09362, po09363, po09364, po09365, po09366, po09367, po09368, po09369, po09370, po09371, po09372, po09373, po09374, po09375, po09376, po09377, po09378, po09379, po09380, po09381, po09382, po09383, po09384, po09385, po09386, po09387, po09388, po09389, po09390, po09391, po09392, po09393, po09394, po09395, po09396, po09397, po09398, po09399, po09400, po09401, po09402, po09403, po09404, po09405, po09406, po09407, po09408, po09409, po09410, po09411, po09412, po09413, po09414, po09415, po09416, po09417, po09418, po09419, po09420, po09421, po09422, po09423, po09424, po09425, po09426, po09427, po09428, po09429, po09430, po09431, po09432, po09433, po09434, po09435, po09436, po09437, po09438, po09439, po09440, po09441, po09442, po09443, po09444, po09445, po09446, po09447, po09448, po09449, po09450, po09451, po09452, po09453, po09454, po09455, po09456, po09457, po09458, po09459, po09460, po09461, po09462, po09463, po09464, po09465, po09466, po09467, po09468, po09469, po09470, po09471, po09472, po09473, po09474, po09475, po09476, po09477, po09478, po09479, po09480, po09481, po09482, po09483, po09484, po09485, po09486, po09487, po09488, po09489, po09490, po09491, po09492, po09493, po09494, po09495, po09496, po09497, po09498, po09499, po09500, po09501, po09502, po09503, po09504, po09505, po09506, po09507, po09508, po09509, po09510, po09511, po09512, po09513, po09514, po09515, po09516, po09517, po09518, po09519, po09520, po09521, po09522, po09523, po09524, po09525, po09526, po09527, po09528, po09529, po09530, po09531, po09532, po09533, po09534, po09535, po09536, po09537, po09538, po09539, po09540, po09541, po09542, po09543, po09544, po09545, po09546, po09547, po09548, po09549, po09550, po09551, po09552, po09553, po09554, po09555, po09556, po09557, po09558, po09559, po09560, po09561, po09562, po09563, po09564, po09565, po09566, po09567, po09568, po09569, po09570, po09571, po09572, po09573, po09574, po09575, po09576, po09577, po09578, po09579, po09580, po09581, po09582, po09583, po09584, po09585, po09586, po09587, po09588, po09589, po09590, po09591, po09592, po09593, po09594, po09595, po09596, po09597, po09598, po09599, po09600, po09601, po09602, po09603, po09604, po09605, po09606, po09607, po09608, po09609, po09610, po09611, po09612, po09613, po09614, po09615, po09616, po09617, po09618, po09619, po09620, po09621, po09622, po09623, po09624, po09625, po09626, po09627, po09628, po09629, po09630, po09631, po09632, po09633, po09634, po09635, po09636, po09637, po09638, po09639, po09640, po09641, po09642, po09643, po09644, po09645, po09646, po09647, po09648, po09649, po09650, po09651, po09652, po09653, po09654, po09655, po09656, po09657, po09658, po09659, po09660, po09661, po09662, po09663, po09664, po09665, po09666, po09667, po09668, po09669, po09670, po09671, po09672, po09673, po09674, po09675, po09676, po09677, po09678, po09679, po09680, po09681, po09682, po09683, po09684, po09685, po09686, po09687, po09688, po09689, po09690, po09691, po09692, po09693, po09694, po09695, po09696, po09697, po09698, po09699, po09700, po09701, po09702, po09703, po09704, po09705, po09706, po09707, po09708, po09709, po09710, po09711, po09712, po09713, po09714, po09715, po09716, po09717, po09718, po09719, po09720, po09721, po09722, po09723, po09724, po09725, po09726, po09727, po09728, po09729, po09730, po09731, po09732, po09733, po09734, po09735, po09736, po09737, po09738, po09739, po09740, po09741, po09742, po09743, po09744, po09745, po09746, po09747, po09748, po09749, po09750, po09751, po09752, po09753, po09754, po09755, po09756, po09757, po09758, po09759, po09760, po09761, po09762, po09763, po09764, po09765, po09766, po09767, po09768, po09769, po09770, po09771, po09772, po09773, po09774, po09775, po09776, po09777, po09778, po09779, po09780, po09781, po09782, po09783, po09784, po09785, po09786, po09787, po09788, po09789, po09790, po09791, po09792, po09793, po09794, po09795, po09796, po09797, po09798, po09799, po09800, po09801, po09802, po09803, po09804, po09805, po09806, po09807, po09808, po09809, po09810, po09811, po09812, po09813, po09814, po09815, po09816, po09817, po09818, po09819, po09820, po09821, po09822, po09823, po09824, po09825, po09826, po09827, po09828, po09829, po09830, po09831, po09832, po09833, po09834, po09835, po09836, po09837, po09838, po09839, po09840, po09841, po09842, po09843, po09844, po09845, po09846, po09847, po09848, po09849, po09850, po09851, po09852, po09853, po09854, po09855, po09856, po09857, po09858, po09859, po09860, po09861, po09862, po09863, po09864, po09865, po09866, po09867, po09868, po09869, po09870, po09871, po09872, po09873, po09874, po09875, po09876, po09877, po09878, po09879, po09880, po09881, po09882, po09883, po09884, po09885, po09886, po09887, po09888, po09889, po09890, po09891, po09892, po09893, po09894, po09895, po09896, po09897, po09898, po09899, po09900, po09901, po09902, po09903, po09904, po09905, po09906, po09907, po09908, po09909, po09910, po09911, po09912, po09913, po09914, po09915, po09916, po09917, po09918, po09919, po09920, po09921, po09922, po09923, po09924, po09925, po09926, po09927, po09928, po09929, po09930, po09931, po09932, po09933, po09934, po09935, po09936, po09937, po09938, po09939, po09940, po09941, po09942, po09943, po09944, po09945, po09946, po09947, po09948, po09949, po09950, po09951, po09952, po09953, po09954, po09955, po09956, po09957, po09958, po09959, po09960, po09961, po09962, po09963, po09964, po09965, po09966, po09967, po09968, po09969, po09970, po09971, po09972, po09973, po09974, po09975, po09976, po09977, po09978, po09979, po09980, po09981, po09982, po09983, po09984, po09985, po09986, po09987, po09988, po09989, po09990, po09991, po09992, po09993, po09994, po09995, po09996, po09997, po09998, po09999, po10000, po10001, po10002, po10003, po10004, po10005, po10006, po10007, po10008, po10009, po10010, po10011, po10012, po10013, po10014, po10015, po10016, po10017, po10018, po10019, po10020, po10021, po10022, po10023, po10024, po10025, po10026, po10027, po10028, po10029, po10030, po10031, po10032, po10033, po10034, po10035, po10036, po10037, po10038, po10039, po10040, po10041, po10042, po10043, po10044, po10045, po10046, po10047, po10048, po10049, po10050, po10051, po10052, po10053, po10054, po10055, po10056, po10057, po10058, po10059, po10060, po10061, po10062, po10063, po10064, po10065, po10066, po10067, po10068, po10069, po10070, po10071, po10072, po10073, po10074, po10075, po10076, po10077, po10078, po10079, po10080, po10081, po10082, po10083, po10084, po10085, po10086, po10087, po10088, po10089, po10090, po10091, po10092, po10093, po10094, po10095, po10096, po10097, po10098, po10099, po10100, po10101, po10102, po10103, po10104, po10105, po10106, po10107, po10108, po10109, po10110, po10111, po10112, po10113, po10114, po10115, po10116, po10117, po10118, po10119, po10120, po10121, po10122, po10123, po10124, po10125, po10126, po10127, po10128, po10129, po10130, po10131, po10132, po10133, po10134, po10135, po10136, po10137, po10138, po10139, po10140, po10141, po10142, po10143, po10144, po10145, po10146, po10147, po10148, po10149, po10150, po10151, po10152, po10153, po10154, po10155, po10156, po10157, po10158, po10159, po10160, po10161, po10162, po10163, po10164, po10165, po10166, po10167, po10168, po10169, po10170, po10171, po10172, po10173, po10174, po10175, po10176, po10177, po10178, po10179, po10180, po10181, po10182, po10183, po10184, po10185, po10186, po10187, po10188, po10189, po10190, po10191, po10192, po10193, po10194, po10195, po10196, po10197, po10198, po10199, po10200, po10201, po10202, po10203, po10204, po10205, po10206, po10207, po10208, po10209, po10210, po10211, po10212, po10213, po10214, po10215, po10216, po10217, po10218, po10219, po10220, po10221, po10222, po10223, po10224, po10225, po10226, po10227, po10228, po10229, po10230, po10231, po10232, po10233, po10234, po10235, po10236, po10237, po10238, po10239, po10240, po10241, po10242, po10243, po10244, po10245, po10246, po10247, po10248, po10249, po10250, po10251, po10252, po10253, po10254, po10255, po10256, po10257, po10258, po10259, po10260, po10261, po10262, po10263, po10264, po10265, po10266, po10267, po10268, po10269, po10270, po10271, po10272, po10273, po10274, po10275, po10276, po10277, po10278, po10279, po10280, po10281, po10282, po10283, po10284, po10285, po10286, po10287, po10288, po10289, po10290, po10291, po10292, po10293, po10294, po10295, po10296, po10297, po10298, po10299, po10300, po10301, po10302, po10303, po10304, po10305, po10306, po10307, po10308, po10309, po10310, po10311, po10312, po10313, po10314, po10315, po10316, po10317, po10318, po10319, po10320, po10321, po10322, po10323, po10324, po10325, po10326, po10327, po10328, po10329, po10330, po10331, po10332, po10333, po10334, po10335, po10336, po10337, po10338, po10339, po10340, po10341, po10342, po10343, po10344, po10345, po10346, po10347, po10348, po10349, po10350, po10351, po10352, po10353, po10354, po10355, po10356, po10357, po10358, po10359, po10360, po10361, po10362, po10363, po10364, po10365, po10366, po10367, po10368, po10369, po10370, po10371, po10372, po10373, po10374, po10375, po10376, po10377, po10378, po10379, po10380, po10381, po10382, po10383, po10384, po10385, po10386, po10387, po10388, po10389, po10390, po10391, po10392, po10393, po10394, po10395, po10396, po10397, po10398, po10399, po10400, po10401, po10402, po10403, po10404, po10405, po10406, po10407, po10408, po10409, po10410, po10411, po10412, po10413, po10414, po10415, po10416, po10417, po10418, po10419, po10420, po10421, po10422, po10423, po10424, po10425, po10426, po10427, po10428, po10429, po10430, po10431, po10432, po10433, po10434, po10435, po10436, po10437, po10438, po10439, po10440, po10441, po10442, po10443, po10444, po10445, po10446, po10447, po10448, po10449, po10450, po10451, po10452, po10453, po10454, po10455, po10456, po10457, po10458, po10459, po10460, po10461, po10462, po10463, po10464, po10465, po10466, po10467, po10468, po10469, po10470, po10471, po10472, po10473, po10474, po10475, po10476, po10477, po10478, po10479, po10480, po10481, po10482, po10483, po10484, po10485, po10486, po10487, po10488, po10489, po10490, po10491, po10492, po10493, po10494, po10495, po10496, po10497, po10498, po10499, po10500, po10501, po10502, po10503, po10504, po10505, po10506, po10507, po10508, po10509, po10510, po10511, po10512, po10513, po10514, po10515, po10516, po10517, po10518, po10519, po10520, po10521, po10522, po10523, po10524, po10525, po10526, po10527, po10528, po10529, po10530, po10531, po10532, po10533, po10534, po10535, po10536, po10537, po10538, po10539, po10540, po10541, po10542, po10543, po10544, po10545, po10546, po10547, po10548, po10549, po10550, po10551, po10552, po10553, po10554, po10555, po10556, po10557, po10558, po10559, po10560, po10561, po10562, po10563, po10564, po10565, po10566, po10567, po10568, po10569, po10570, po10571, po10572, po10573, po10574, po10575, po10576, po10577, po10578, po10579, po10580, po10581, po10582, po10583, po10584, po10585, po10586, po10587, po10588, po10589, po10590, po10591, po10592, po10593, po10594, po10595, po10596, po10597, po10598, po10599, po10600, po10601, po10602, po10603, po10604, po10605, po10606, po10607, po10608, po10609, po10610, po10611, po10612, po10613, po10614, po10615, po10616, po10617, po10618, po10619, po10620, po10621, po10622, po10623, po10624, po10625, po10626, po10627, po10628, po10629, po10630, po10631, po10632, po10633, po10634, po10635, po10636, po10637, po10638, po10639, po10640, po10641, po10642, po10643, po10644, po10645, po10646, po10647, po10648, po10649, po10650, po10651, po10652, po10653, po10654, po10655, po10656, po10657, po10658, po10659, po10660, po10661, po10662, po10663, po10664, po10665, po10666, po10667, po10668, po10669, po10670, po10671, po10672, po10673, po10674, po10675, po10676, po10677, po10678, po10679, po10680, po10681, po10682, po10683, po10684, po10685, po10686, po10687, po10688, po10689, po10690, po10691, po10692, po10693, po10694, po10695;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835, w46836, w46837, w46838, w46839, w46840, w46841, w46842, w46843, w46844, w46845, w46846, w46847, w46848, w46849, w46850, w46851, w46852, w46853, w46854, w46855, w46856, w46857, w46858, w46859, w46860, w46861, w46862, w46863, w46864, w46865, w46866, w46867, w46868, w46869, w46870, w46871, w46872, w46873, w46874, w46875, w46876, w46877, w46878, w46879, w46880, w46881, w46882, w46883, w46884, w46885, w46886, w46887, w46888, w46889, w46890, w46891, w46892, w46893, w46894, w46895, w46896, w46897, w46898, w46899, w46900, w46901, w46902, w46903, w46904, w46905, w46906, w46907, w46908, w46909, w46910, w46911, w46912, w46913, w46914, w46915, w46916, w46917, w46918, w46919, w46920, w46921, w46922, w46923, w46924, w46925, w46926, w46927, w46928, w46929, w46930, w46931, w46932, w46933, w46934, w46935, w46936, w46937, w46938, w46939, w46940, w46941, w46942, w46943, w46944, w46945, w46946, w46947, w46948, w46949, w46950, w46951, w46952, w46953, w46954, w46955, w46956, w46957, w46958, w46959, w46960, w46961, w46962, w46963, w46964, w46965, w46966, w46967, w46968, w46969, w46970, w46971, w46972, w46973, w46974, w46975, w46976, w46977, w46978, w46979, w46980, w46981, w46982, w46983, w46984, w46985, w46986, w46987, w46988, w46989, w46990, w46991, w46992, w46993, w46994, w46995, w46996, w46997, w46998, w46999, w47000, w47001, w47002, w47003, w47004, w47005, w47006, w47007, w47008, w47009, w47010, w47011, w47012, w47013, w47014, w47015, w47016, w47017, w47018, w47019, w47020, w47021, w47022, w47023, w47024, w47025, w47026, w47027, w47028, w47029, w47030, w47031, w47032, w47033, w47034, w47035, w47036, w47037, w47038, w47039, w47040, w47041, w47042, w47043, w47044, w47045, w47046, w47047, w47048, w47049, w47050, w47051, w47052, w47053, w47054, w47055, w47056, w47057, w47058, w47059, w47060, w47061, w47062, w47063, w47064, w47065, w47066, w47067, w47068, w47069, w47070, w47071, w47072, w47073, w47074, w47075, w47076, w47077, w47078, w47079, w47080, w47081, w47082, w47083, w47084, w47085, w47086, w47087, w47088, w47089, w47090, w47091, w47092, w47093, w47094, w47095, w47096, w47097, w47098, w47099, w47100, w47101, w47102, w47103, w47104, w47105, w47106, w47107, w47108, w47109, w47110, w47111, w47112, w47113, w47114, w47115, w47116, w47117, w47118, w47119, w47120, w47121, w47122, w47123, w47124, w47125, w47126, w47127, w47128, w47129, w47130, w47131, w47132, w47133, w47134, w47135, w47136, w47137, w47138, w47139, w47140, w47141, w47142, w47143, w47144, w47145, w47146, w47147, w47148, w47149, w47150, w47151, w47152, w47153, w47154, w47155, w47156, w47157, w47158, w47159, w47160, w47161, w47162, w47163, w47164, w47165, w47166, w47167, w47168, w47169, w47170, w47171, w47172, w47173, w47174, w47175, w47176, w47177, w47178, w47179, w47180, w47181, w47182, w47183, w47184, w47185, w47186, w47187, w47188, w47189, w47190, w47191, w47192, w47193, w47194, w47195, w47196, w47197, w47198, w47199, w47200, w47201, w47202, w47203, w47204, w47205, w47206, w47207, w47208, w47209, w47210, w47211, w47212, w47213, w47214, w47215, w47216, w47217, w47218, w47219, w47220, w47221, w47222, w47223, w47224, w47225, w47226, w47227, w47228, w47229, w47230, w47231, w47232, w47233, w47234, w47235, w47236, w47237, w47238, w47239, w47240, w47241, w47242, w47243, w47244, w47245, w47246, w47247, w47248, w47249, w47250, w47251, w47252, w47253, w47254, w47255, w47256, w47257, w47258, w47259, w47260, w47261, w47262, w47263, w47264, w47265, w47266, w47267, w47268, w47269, w47270, w47271, w47272, w47273, w47274, w47275, w47276, w47277, w47278, w47279, w47280, w47281, w47282, w47283, w47284, w47285, w47286, w47287, w47288, w47289, w47290, w47291, w47292, w47293, w47294, w47295, w47296, w47297, w47298, w47299, w47300, w47301, w47302, w47303, w47304, w47305, w47306, w47307, w47308, w47309, w47310, w47311, w47312, w47313, w47314, w47315, w47316, w47317, w47318, w47319, w47320, w47321, w47322, w47323, w47324, w47325, w47326, w47327, w47328, w47329, w47330, w47331, w47332, w47333, w47334, w47335, w47336, w47337, w47338, w47339, w47340, w47341, w47342, w47343, w47344, w47345, w47346, w47347, w47348, w47349, w47350, w47351, w47352, w47353, w47354, w47355, w47356, w47357, w47358, w47359, w47360, w47361, w47362, w47363, w47364, w47365, w47366, w47367, w47368, w47369, w47370, w47371, w47372, w47373, w47374, w47375, w47376, w47377, w47378, w47379, w47380, w47381, w47382, w47383, w47384, w47385, w47386, w47387, w47388, w47389, w47390, w47391, w47392, w47393, w47394, w47395, w47396, w47397, w47398, w47399, w47400, w47401, w47402, w47403, w47404, w47405, w47406, w47407, w47408, w47409, w47410, w47411, w47412, w47413, w47414, w47415, w47416, w47417, w47418, w47419, w47420, w47421, w47422, w47423, w47424, w47425, w47426, w47427, w47428, w47429, w47430, w47431, w47432, w47433, w47434, w47435, w47436, w47437, w47438, w47439, w47440, w47441, w47442, w47443, w47444, w47445, w47446, w47447, w47448, w47449, w47450, w47451, w47452, w47453, w47454, w47455, w47456, w47457, w47458, w47459, w47460, w47461, w47462, w47463, w47464, w47465, w47466, w47467, w47468, w47469, w47470, w47471, w47472, w47473, w47474, w47475, w47476, w47477, w47478, w47479, w47480, w47481, w47482, w47483, w47484, w47485, w47486, w47487, w47488, w47489, w47490, w47491, w47492, w47493, w47494, w47495, w47496, w47497, w47498, w47499, w47500, w47501, w47502, w47503, w47504, w47505, w47506, w47507, w47508, w47509, w47510, w47511, w47512, w47513, w47514, w47515, w47516, w47517, w47518, w47519, w47520, w47521, w47522, w47523, w47524, w47525, w47526, w47527, w47528, w47529, w47530, w47531, w47532, w47533, w47534, w47535, w47536, w47537, w47538, w47539, w47540, w47541, w47542, w47543, w47544, w47545, w47546, w47547, w47548, w47549, w47550, w47551, w47552, w47553, w47554, w47555, w47556, w47557, w47558, w47559, w47560, w47561, w47562, w47563, w47564, w47565, w47566, w47567, w47568, w47569, w47570, w47571, w47572, w47573, w47574, w47575, w47576, w47577, w47578, w47579, w47580, w47581, w47582, w47583, w47584, w47585, w47586, w47587, w47588, w47589, w47590, w47591, w47592, w47593, w47594, w47595, w47596, w47597, w47598, w47599, w47600, w47601, w47602, w47603, w47604, w47605, w47606, w47607, w47608, w47609, w47610, w47611, w47612, w47613, w47614, w47615, w47616, w47617, w47618, w47619, w47620, w47621, w47622, w47623, w47624, w47625, w47626, w47627, w47628, w47629, w47630, w47631, w47632, w47633, w47634, w47635, w47636, w47637, w47638, w47639, w47640, w47641, w47642, w47643, w47644, w47645, w47646, w47647, w47648, w47649, w47650, w47651, w47652, w47653, w47654, w47655, w47656, w47657, w47658, w47659, w47660, w47661, w47662, w47663, w47664, w47665, w47666, w47667, w47668, w47669, w47670, w47671, w47672, w47673, w47674, w47675, w47676, w47677, w47678, w47679, w47680, w47681, w47682, w47683, w47684, w47685, w47686, w47687, w47688, w47689, w47690, w47691, w47692, w47693, w47694, w47695, w47696, w47697, w47698, w47699, w47700, w47701, w47702, w47703, w47704, w47705, w47706, w47707, w47708, w47709, w47710, w47711, w47712, w47713, w47714, w47715, w47716, w47717, w47718, w47719, w47720, w47721, w47722, w47723, w47724, w47725, w47726, w47727, w47728, w47729, w47730, w47731, w47732, w47733, w47734, w47735, w47736, w47737, w47738, w47739, w47740, w47741, w47742, w47743, w47744, w47745, w47746, w47747, w47748, w47749, w47750, w47751, w47752, w47753, w47754, w47755, w47756, w47757, w47758, w47759, w47760, w47761, w47762, w47763, w47764, w47765, w47766, w47767, w47768, w47769, w47770, w47771, w47772, w47773, w47774, w47775, w47776, w47777, w47778, w47779, w47780, w47781, w47782, w47783, w47784, w47785, w47786, w47787, w47788, w47789, w47790, w47791, w47792, w47793, w47794, w47795, w47796, w47797, w47798, w47799, w47800, w47801, w47802, w47803, w47804, w47805, w47806, w47807, w47808, w47809, w47810, w47811, w47812, w47813, w47814, w47815, w47816, w47817, w47818, w47819, w47820, w47821, w47822, w47823, w47824, w47825, w47826, w47827, w47828, w47829, w47830, w47831, w47832, w47833, w47834, w47835, w47836, w47837, w47838, w47839, w47840, w47841, w47842, w47843, w47844, w47845, w47846, w47847, w47848, w47849, w47850, w47851, w47852, w47853, w47854, w47855, w47856, w47857, w47858, w47859, w47860, w47861, w47862, w47863, w47864, w47865, w47866, w47867, w47868, w47869, w47870, w47871, w47872, w47873, w47874, w47875, w47876, w47877, w47878, w47879, w47880, w47881, w47882, w47883, w47884, w47885, w47886, w47887, w47888, w47889, w47890, w47891, w47892, w47893, w47894, w47895, w47896, w47897, w47898, w47899, w47900, w47901, w47902, w47903, w47904, w47905, w47906, w47907, w47908, w47909, w47910, w47911, w47912, w47913, w47914, w47915, w47916, w47917, w47918, w47919, w47920, w47921, w47922, w47923, w47924, w47925, w47926, w47927, w47928, w47929, w47930, w47931, w47932, w47933, w47934, w47935, w47936, w47937, w47938, w47939, w47940, w47941, w47942, w47943, w47944, w47945, w47946, w47947, w47948, w47949, w47950, w47951, w47952, w47953, w47954, w47955, w47956, w47957, w47958, w47959, w47960, w47961, w47962, w47963, w47964, w47965, w47966, w47967, w47968, w47969, w47970, w47971, w47972, w47973, w47974, w47975, w47976, w47977, w47978, w47979, w47980, w47981, w47982, w47983, w47984, w47985, w47986, w47987, w47988, w47989, w47990, w47991, w47992, w47993, w47994, w47995, w47996, w47997, w47998, w47999, w48000, w48001, w48002, w48003, w48004, w48005, w48006, w48007, w48008, w48009, w48010, w48011, w48012, w48013, w48014, w48015, w48016, w48017, w48018, w48019, w48020, w48021, w48022, w48023, w48024, w48025, w48026, w48027, w48028, w48029, w48030, w48031, w48032, w48033, w48034, w48035, w48036, w48037, w48038, w48039, w48040, w48041, w48042, w48043, w48044, w48045, w48046, w48047, w48048, w48049, w48050, w48051, w48052, w48053, w48054, w48055, w48056, w48057, w48058, w48059, w48060, w48061, w48062, w48063, w48064, w48065, w48066, w48067, w48068, w48069, w48070, w48071, w48072, w48073, w48074, w48075, w48076, w48077, w48078, w48079, w48080, w48081, w48082, w48083, w48084, w48085, w48086, w48087, w48088, w48089, w48090, w48091, w48092, w48093, w48094, w48095, w48096, w48097, w48098, w48099, w48100, w48101, w48102, w48103, w48104, w48105, w48106, w48107, w48108, w48109, w48110, w48111, w48112, w48113, w48114, w48115, w48116, w48117, w48118, w48119, w48120, w48121, w48122, w48123, w48124, w48125, w48126, w48127, w48128, w48129, w48130, w48131, w48132, w48133, w48134, w48135, w48136, w48137, w48138, w48139, w48140, w48141, w48142, w48143, w48144, w48145, w48146, w48147, w48148, w48149, w48150, w48151, w48152, w48153, w48154, w48155, w48156, w48157, w48158, w48159, w48160, w48161, w48162, w48163, w48164, w48165, w48166, w48167, w48168, w48169, w48170, w48171, w48172, w48173, w48174, w48175, w48176, w48177, w48178, w48179, w48180, w48181, w48182, w48183, w48184, w48185, w48186, w48187, w48188, w48189, w48190, w48191, w48192, w48193, w48194, w48195, w48196, w48197, w48198, w48199, w48200, w48201, w48202, w48203, w48204, w48205, w48206, w48207, w48208, w48209, w48210, w48211, w48212, w48213, w48214, w48215, w48216, w48217, w48218, w48219, w48220, w48221, w48222, w48223, w48224, w48225, w48226, w48227, w48228, w48229, w48230, w48231, w48232, w48233, w48234, w48235, w48236, w48237, w48238, w48239, w48240, w48241, w48242, w48243, w48244, w48245, w48246, w48247, w48248, w48249, w48250, w48251, w48252, w48253, w48254, w48255, w48256, w48257, w48258, w48259, w48260, w48261, w48262, w48263, w48264, w48265, w48266, w48267, w48268, w48269, w48270, w48271, w48272, w48273, w48274, w48275, w48276, w48277, w48278, w48279, w48280, w48281, w48282, w48283, w48284, w48285, w48286, w48287, w48288, w48289, w48290, w48291, w48292, w48293, w48294, w48295, w48296, w48297, w48298, w48299, w48300, w48301, w48302, w48303, w48304, w48305, w48306, w48307, w48308, w48309, w48310, w48311, w48312, w48313, w48314, w48315, w48316, w48317, w48318, w48319, w48320, w48321, w48322, w48323, w48324, w48325, w48326, w48327, w48328, w48329, w48330, w48331, w48332, w48333, w48334, w48335, w48336, w48337, w48338, w48339, w48340, w48341, w48342, w48343, w48344, w48345, w48346, w48347, w48348, w48349, w48350, w48351, w48352, w48353, w48354, w48355, w48356, w48357, w48358, w48359, w48360, w48361, w48362, w48363, w48364, w48365, w48366, w48367, w48368, w48369, w48370, w48371, w48372, w48373, w48374, w48375, w48376, w48377, w48378, w48379, w48380, w48381, w48382, w48383, w48384, w48385, w48386, w48387, w48388, w48389, w48390, w48391, w48392, w48393, w48394, w48395, w48396, w48397, w48398, w48399, w48400, w48401, w48402, w48403, w48404, w48405, w48406, w48407, w48408, w48409, w48410, w48411, w48412, w48413, w48414, w48415, w48416, w48417, w48418, w48419, w48420, w48421, w48422, w48423, w48424, w48425, w48426, w48427, w48428, w48429, w48430, w48431, w48432, w48433, w48434, w48435, w48436, w48437, w48438, w48439, w48440, w48441, w48442, w48443, w48444, w48445, w48446, w48447, w48448, w48449, w48450, w48451, w48452, w48453, w48454, w48455, w48456, w48457, w48458, w48459, w48460, w48461, w48462, w48463, w48464, w48465, w48466, w48467, w48468, w48469, w48470, w48471, w48472, w48473, w48474, w48475, w48476, w48477, w48478, w48479, w48480, w48481, w48482, w48483, w48484, w48485, w48486, w48487, w48488, w48489, w48490, w48491, w48492, w48493, w48494, w48495, w48496, w48497, w48498, w48499, w48500, w48501, w48502, w48503, w48504, w48505, w48506, w48507, w48508, w48509, w48510, w48511, w48512, w48513, w48514, w48515, w48516, w48517, w48518, w48519, w48520, w48521, w48522, w48523, w48524, w48525, w48526, w48527, w48528, w48529, w48530, w48531, w48532, w48533, w48534, w48535, w48536, w48537, w48538, w48539, w48540, w48541, w48542, w48543, w48544, w48545, w48546, w48547, w48548, w48549, w48550, w48551, w48552, w48553, w48554, w48555, w48556, w48557, w48558, w48559, w48560, w48561, w48562, w48563, w48564, w48565, w48566, w48567, w48568, w48569, w48570, w48571, w48572, w48573, w48574, w48575, w48576, w48577, w48578, w48579, w48580, w48581, w48582, w48583, w48584, w48585, w48586, w48587, w48588, w48589, w48590, w48591, w48592, w48593, w48594, w48595, w48596, w48597, w48598, w48599, w48600, w48601, w48602, w48603, w48604, w48605, w48606, w48607, w48608, w48609, w48610, w48611, w48612, w48613, w48614, w48615, w48616, w48617, w48618, w48619, w48620, w48621, w48622, w48623, w48624, w48625, w48626, w48627, w48628, w48629, w48630, w48631, w48632, w48633, w48634, w48635, w48636, w48637, w48638, w48639, w48640, w48641, w48642, w48643, w48644, w48645, w48646, w48647, w48648, w48649, w48650, w48651, w48652, w48653, w48654, w48655, w48656, w48657, w48658, w48659, w48660, w48661, w48662, w48663, w48664, w48665, w48666, w48667, w48668, w48669, w48670, w48671, w48672, w48673, w48674, w48675, w48676, w48677, w48678, w48679, w48680, w48681, w48682, w48683, w48684, w48685, w48686, w48687, w48688, w48689, w48690, w48691, w48692, w48693, w48694, w48695, w48696, w48697, w48698, w48699, w48700, w48701, w48702, w48703, w48704, w48705, w48706, w48707, w48708, w48709, w48710, w48711, w48712, w48713, w48714, w48715, w48716, w48717, w48718, w48719, w48720, w48721, w48722, w48723, w48724, w48725, w48726, w48727, w48728, w48729, w48730, w48731, w48732, w48733, w48734, w48735, w48736, w48737, w48738, w48739, w48740, w48741, w48742, w48743, w48744, w48745, w48746, w48747, w48748, w48749, w48750, w48751, w48752, w48753, w48754, w48755, w48756, w48757, w48758, w48759, w48760, w48761, w48762, w48763, w48764, w48765, w48766, w48767, w48768, w48769, w48770, w48771, w48772, w48773, w48774, w48775, w48776, w48777, w48778, w48779, w48780, w48781, w48782, w48783, w48784, w48785, w48786, w48787, w48788, w48789, w48790, w48791, w48792, w48793, w48794, w48795, w48796, w48797, w48798, w48799, w48800, w48801, w48802, w48803, w48804, w48805, w48806, w48807, w48808, w48809, w48810, w48811, w48812, w48813, w48814, w48815, w48816, w48817, w48818, w48819, w48820, w48821, w48822, w48823, w48824, w48825, w48826, w48827, w48828, w48829, w48830, w48831, w48832, w48833, w48834, w48835, w48836, w48837, w48838, w48839, w48840, w48841, w48842, w48843, w48844, w48845, w48846, w48847, w48848, w48849, w48850, w48851, w48852, w48853, w48854, w48855, w48856, w48857, w48858, w48859, w48860, w48861, w48862, w48863, w48864, w48865, w48866, w48867, w48868, w48869, w48870, w48871, w48872, w48873, w48874, w48875, w48876, w48877, w48878, w48879, w48880, w48881, w48882, w48883, w48884, w48885, w48886, w48887, w48888, w48889, w48890, w48891, w48892, w48893, w48894, w48895, w48896, w48897, w48898, w48899, w48900, w48901, w48902, w48903, w48904, w48905, w48906, w48907, w48908, w48909, w48910, w48911, w48912, w48913, w48914, w48915, w48916, w48917, w48918, w48919, w48920, w48921, w48922, w48923, w48924, w48925, w48926, w48927, w48928, w48929, w48930, w48931, w48932, w48933, w48934, w48935, w48936, w48937, w48938, w48939, w48940, w48941, w48942, w48943, w48944, w48945, w48946, w48947, w48948, w48949, w48950, w48951, w48952, w48953, w48954, w48955, w48956, w48957, w48958, w48959, w48960, w48961, w48962, w48963, w48964, w48965, w48966, w48967, w48968, w48969, w48970, w48971, w48972, w48973, w48974, w48975, w48976, w48977, w48978, w48979, w48980, w48981, w48982, w48983, w48984, w48985, w48986, w48987, w48988, w48989, w48990, w48991, w48992, w48993, w48994, w48995, w48996, w48997, w48998, w48999, w49000, w49001, w49002, w49003, w49004, w49005, w49006, w49007, w49008, w49009, w49010, w49011, w49012, w49013, w49014, w49015, w49016, w49017, w49018, w49019, w49020, w49021, w49022, w49023, w49024, w49025, w49026, w49027, w49028, w49029, w49030, w49031, w49032, w49033, w49034, w49035, w49036, w49037, w49038, w49039, w49040, w49041, w49042, w49043, w49044, w49045, w49046, w49047, w49048, w49049, w49050, w49051, w49052, w49053, w49054, w49055, w49056, w49057, w49058, w49059, w49060, w49061, w49062, w49063, w49064, w49065, w49066, w49067, w49068, w49069, w49070, w49071, w49072, w49073, w49074, w49075, w49076, w49077, w49078, w49079, w49080, w49081, w49082, w49083, w49084, w49085, w49086, w49087, w49088, w49089, w49090, w49091, w49092, w49093, w49094, w49095, w49096, w49097, w49098, w49099, w49100, w49101, w49102, w49103, w49104, w49105, w49106, w49107, w49108, w49109, w49110, w49111, w49112, w49113, w49114, w49115, w49116, w49117, w49118, w49119, w49120, w49121, w49122, w49123, w49124, w49125, w49126, w49127, w49128, w49129, w49130, w49131, w49132, w49133, w49134, w49135, w49136, w49137, w49138, w49139, w49140, w49141, w49142, w49143, w49144, w49145, w49146, w49147, w49148, w49149, w49150, w49151, w49152, w49153, w49154, w49155, w49156, w49157, w49158, w49159, w49160, w49161, w49162, w49163, w49164, w49165, w49166, w49167, w49168, w49169, w49170, w49171, w49172, w49173, w49174, w49175, w49176, w49177, w49178, w49179, w49180, w49181, w49182, w49183, w49184, w49185, w49186, w49187, w49188, w49189, w49190, w49191, w49192, w49193, w49194, w49195, w49196, w49197, w49198, w49199, w49200, w49201, w49202, w49203, w49204, w49205, w49206, w49207, w49208, w49209, w49210, w49211, w49212, w49213, w49214, w49215, w49216, w49217, w49218, w49219, w49220, w49221, w49222, w49223, w49224, w49225, w49226, w49227, w49228, w49229, w49230, w49231, w49232, w49233, w49234, w49235, w49236, w49237, w49238, w49239, w49240, w49241, w49242, w49243, w49244, w49245, w49246, w49247, w49248, w49249, w49250, w49251, w49252, w49253, w49254, w49255, w49256, w49257, w49258, w49259, w49260, w49261, w49262, w49263, w49264, w49265, w49266, w49267, w49268, w49269, w49270, w49271, w49272, w49273, w49274, w49275, w49276, w49277, w49278, w49279, w49280, w49281, w49282, w49283, w49284, w49285, w49286, w49287, w49288, w49289, w49290, w49291, w49292, w49293, w49294, w49295, w49296, w49297, w49298, w49299, w49300, w49301, w49302, w49303, w49304, w49305, w49306, w49307, w49308, w49309, w49310, w49311, w49312, w49313, w49314, w49315, w49316, w49317, w49318, w49319, w49320, w49321, w49322, w49323, w49324, w49325, w49326, w49327, w49328, w49329, w49330, w49331, w49332, w49333, w49334, w49335, w49336, w49337, w49338, w49339, w49340, w49341, w49342, w49343, w49344, w49345, w49346, w49347, w49348, w49349, w49350, w49351, w49352, w49353, w49354, w49355, w49356, w49357, w49358, w49359, w49360, w49361, w49362, w49363, w49364, w49365, w49366, w49367, w49368, w49369, w49370, w49371, w49372, w49373, w49374, w49375, w49376, w49377, w49378, w49379, w49380, w49381, w49382, w49383, w49384, w49385, w49386, w49387, w49388, w49389, w49390, w49391, w49392, w49393, w49394, w49395, w49396, w49397, w49398, w49399, w49400, w49401, w49402, w49403, w49404, w49405, w49406, w49407, w49408, w49409, w49410, w49411, w49412, w49413, w49414, w49415, w49416, w49417, w49418, w49419, w49420, w49421, w49422, w49423, w49424, w49425, w49426, w49427, w49428, w49429, w49430, w49431, w49432, w49433, w49434, w49435, w49436, w49437, w49438, w49439, w49440, w49441, w49442, w49443, w49444, w49445, w49446, w49447, w49448, w49449, w49450, w49451, w49452, w49453, w49454, w49455, w49456, w49457, w49458, w49459, w49460, w49461, w49462, w49463, w49464, w49465, w49466, w49467, w49468, w49469, w49470, w49471, w49472, w49473, w49474, w49475, w49476, w49477, w49478, w49479, w49480, w49481, w49482, w49483, w49484, w49485, w49486, w49487, w49488, w49489, w49490, w49491, w49492, w49493, w49494, w49495, w49496, w49497, w49498, w49499, w49500, w49501, w49502, w49503, w49504, w49505, w49506, w49507, w49508, w49509, w49510, w49511, w49512, w49513, w49514, w49515, w49516, w49517, w49518, w49519, w49520, w49521, w49522, w49523, w49524, w49525, w49526, w49527, w49528, w49529, w49530, w49531, w49532, w49533, w49534, w49535, w49536, w49537, w49538, w49539, w49540, w49541, w49542, w49543, w49544, w49545, w49546, w49547, w49548, w49549, w49550, w49551, w49552, w49553, w49554, w49555, w49556, w49557, w49558, w49559, w49560, w49561, w49562, w49563, w49564, w49565, w49566, w49567, w49568, w49569, w49570, w49571, w49572, w49573, w49574, w49575, w49576, w49577, w49578, w49579, w49580, w49581, w49582, w49583, w49584, w49585, w49586, w49587, w49588, w49589, w49590, w49591, w49592, w49593, w49594, w49595, w49596, w49597, w49598, w49599, w49600, w49601, w49602, w49603, w49604, w49605, w49606, w49607, w49608, w49609, w49610, w49611, w49612, w49613, w49614, w49615, w49616, w49617, w49618, w49619, w49620, w49621, w49622, w49623, w49624, w49625, w49626, w49627, w49628, w49629, w49630, w49631, w49632, w49633, w49634, w49635, w49636, w49637, w49638, w49639, w49640, w49641, w49642, w49643, w49644, w49645, w49646, w49647, w49648, w49649, w49650, w49651, w49652, w49653, w49654, w49655, w49656, w49657, w49658, w49659, w49660, w49661, w49662, w49663, w49664, w49665, w49666, w49667, w49668, w49669, w49670, w49671, w49672, w49673, w49674, w49675, w49676, w49677, w49678, w49679, w49680, w49681, w49682, w49683, w49684, w49685, w49686, w49687, w49688, w49689, w49690, w49691, w49692, w49693, w49694, w49695, w49696, w49697, w49698, w49699, w49700, w49701, w49702, w49703, w49704, w49705, w49706, w49707, w49708, w49709, w49710, w49711, w49712, w49713, w49714, w49715, w49716, w49717, w49718, w49719, w49720, w49721, w49722, w49723, w49724, w49725, w49726, w49727, w49728, w49729, w49730, w49731, w49732, w49733, w49734, w49735, w49736, w49737, w49738, w49739, w49740, w49741, w49742, w49743, w49744, w49745, w49746, w49747, w49748, w49749, w49750, w49751, w49752, w49753, w49754, w49755, w49756, w49757, w49758, w49759, w49760, w49761, w49762, w49763, w49764, w49765, w49766, w49767, w49768, w49769, w49770, w49771, w49772, w49773, w49774, w49775, w49776, w49777, w49778, w49779, w49780, w49781, w49782, w49783, w49784, w49785, w49786, w49787, w49788, w49789, w49790, w49791, w49792, w49793, w49794, w49795, w49796, w49797, w49798, w49799, w49800, w49801, w49802, w49803, w49804, w49805, w49806, w49807, w49808, w49809, w49810, w49811, w49812, w49813, w49814, w49815, w49816, w49817, w49818, w49819, w49820, w49821, w49822, w49823, w49824, w49825, w49826, w49827, w49828, w49829, w49830, w49831, w49832, w49833, w49834, w49835, w49836, w49837, w49838, w49839, w49840, w49841, w49842, w49843, w49844, w49845, w49846, w49847, w49848, w49849, w49850, w49851, w49852, w49853, w49854, w49855, w49856, w49857, w49858, w49859, w49860, w49861, w49862, w49863, w49864, w49865, w49866, w49867, w49868, w49869, w49870, w49871, w49872, w49873, w49874, w49875, w49876, w49877, w49878, w49879, w49880, w49881, w49882, w49883, w49884, w49885, w49886, w49887, w49888, w49889, w49890, w49891, w49892, w49893, w49894, w49895, w49896, w49897, w49898, w49899, w49900, w49901, w49902, w49903, w49904, w49905, w49906, w49907, w49908, w49909, w49910, w49911, w49912, w49913, w49914, w49915, w49916, w49917, w49918, w49919, w49920, w49921, w49922, w49923, w49924, w49925, w49926, w49927, w49928, w49929, w49930, w49931, w49932, w49933, w49934, w49935, w49936, w49937, w49938, w49939, w49940, w49941, w49942, w49943, w49944, w49945, w49946, w49947, w49948, w49949, w49950, w49951, w49952, w49953, w49954, w49955, w49956, w49957, w49958, w49959, w49960, w49961, w49962, w49963, w49964, w49965, w49966, w49967, w49968, w49969, w49970, w49971, w49972, w49973, w49974, w49975, w49976, w49977, w49978, w49979, w49980, w49981, w49982, w49983, w49984, w49985, w49986, w49987, w49988, w49989, w49990, w49991, w49992, w49993, w49994, w49995, w49996, w49997, w49998, w49999, w50000, w50001, w50002, w50003, w50004, w50005, w50006, w50007, w50008, w50009, w50010, w50011, w50012, w50013, w50014, w50015, w50016, w50017, w50018, w50019, w50020, w50021, w50022, w50023, w50024, w50025, w50026, w50027, w50028, w50029, w50030, w50031, w50032, w50033, w50034, w50035, w50036, w50037, w50038, w50039, w50040, w50041, w50042, w50043, w50044, w50045, w50046, w50047, w50048, w50049, w50050, w50051, w50052, w50053, w50054, w50055, w50056, w50057, w50058, w50059, w50060, w50061, w50062, w50063, w50064, w50065, w50066, w50067, w50068, w50069, w50070, w50071, w50072, w50073, w50074, w50075, w50076, w50077, w50078, w50079, w50080, w50081, w50082, w50083, w50084, w50085, w50086, w50087, w50088, w50089, w50090, w50091, w50092, w50093, w50094, w50095, w50096, w50097, w50098, w50099, w50100, w50101, w50102, w50103, w50104, w50105, w50106, w50107, w50108, w50109, w50110, w50111, w50112, w50113, w50114, w50115, w50116, w50117, w50118, w50119, w50120, w50121, w50122, w50123, w50124, w50125, w50126, w50127, w50128, w50129, w50130, w50131, w50132, w50133, w50134, w50135, w50136, w50137, w50138, w50139, w50140, w50141, w50142, w50143, w50144, w50145, w50146, w50147, w50148, w50149, w50150, w50151, w50152, w50153, w50154, w50155, w50156, w50157, w50158, w50159, w50160, w50161, w50162, w50163, w50164, w50165, w50166, w50167, w50168, w50169, w50170, w50171, w50172, w50173, w50174, w50175, w50176, w50177, w50178, w50179, w50180, w50181, w50182, w50183, w50184, w50185, w50186, w50187, w50188, w50189, w50190, w50191, w50192, w50193, w50194, w50195, w50196, w50197, w50198, w50199, w50200, w50201, w50202, w50203, w50204, w50205, w50206, w50207, w50208, w50209, w50210, w50211, w50212, w50213, w50214, w50215, w50216, w50217, w50218, w50219, w50220, w50221, w50222, w50223, w50224, w50225, w50226, w50227, w50228, w50229, w50230, w50231, w50232, w50233, w50234, w50235, w50236, w50237, w50238, w50239, w50240, w50241, w50242, w50243, w50244, w50245, w50246, w50247, w50248, w50249, w50250, w50251, w50252, w50253, w50254, w50255, w50256, w50257, w50258, w50259, w50260, w50261, w50262, w50263, w50264, w50265, w50266, w50267, w50268, w50269, w50270, w50271, w50272, w50273, w50274, w50275, w50276, w50277, w50278, w50279, w50280, w50281, w50282, w50283, w50284, w50285, w50286, w50287, w50288, w50289, w50290, w50291, w50292, w50293, w50294, w50295, w50296, w50297, w50298, w50299, w50300, w50301, w50302, w50303, w50304, w50305, w50306, w50307, w50308, w50309, w50310, w50311, w50312, w50313, w50314, w50315, w50316, w50317, w50318, w50319, w50320, w50321, w50322, w50323, w50324, w50325, w50326, w50327, w50328, w50329, w50330, w50331, w50332, w50333, w50334, w50335, w50336, w50337, w50338, w50339, w50340, w50341, w50342, w50343, w50344, w50345, w50346, w50347, w50348, w50349, w50350, w50351, w50352, w50353, w50354, w50355, w50356, w50357, w50358, w50359, w50360, w50361, w50362, w50363, w50364, w50365, w50366, w50367, w50368, w50369, w50370, w50371, w50372, w50373, w50374, w50375, w50376, w50377, w50378, w50379, w50380, w50381, w50382, w50383, w50384, w50385, w50386, w50387, w50388, w50389, w50390, w50391, w50392, w50393, w50394, w50395, w50396, w50397, w50398, w50399, w50400, w50401, w50402, w50403, w50404, w50405, w50406, w50407, w50408, w50409, w50410, w50411, w50412, w50413, w50414, w50415, w50416, w50417, w50418, w50419, w50420, w50421, w50422, w50423, w50424, w50425, w50426, w50427, w50428, w50429, w50430, w50431, w50432, w50433, w50434, w50435, w50436, w50437, w50438, w50439, w50440, w50441, w50442, w50443, w50444, w50445, w50446, w50447, w50448, w50449, w50450, w50451, w50452, w50453, w50454, w50455, w50456, w50457, w50458, w50459, w50460, w50461, w50462, w50463, w50464, w50465, w50466, w50467, w50468, w50469, w50470, w50471, w50472, w50473, w50474, w50475, w50476, w50477, w50478, w50479, w50480, w50481, w50482, w50483, w50484, w50485, w50486, w50487, w50488, w50489, w50490, w50491, w50492, w50493, w50494, w50495, w50496, w50497, w50498, w50499, w50500, w50501, w50502, w50503, w50504, w50505, w50506, w50507, w50508, w50509, w50510, w50511, w50512, w50513, w50514, w50515, w50516, w50517, w50518, w50519, w50520, w50521, w50522, w50523, w50524, w50525, w50526, w50527, w50528, w50529, w50530, w50531, w50532, w50533, w50534, w50535, w50536, w50537, w50538, w50539, w50540, w50541, w50542, w50543, w50544, w50545, w50546, w50547, w50548, w50549, w50550, w50551, w50552, w50553, w50554, w50555, w50556, w50557, w50558, w50559, w50560, w50561, w50562, w50563, w50564, w50565, w50566, w50567, w50568, w50569, w50570, w50571, w50572, w50573, w50574, w50575, w50576, w50577, w50578, w50579, w50580, w50581, w50582, w50583, w50584, w50585, w50586, w50587, w50588, w50589, w50590, w50591, w50592, w50593, w50594, w50595, w50596, w50597, w50598, w50599, w50600, w50601, w50602, w50603, w50604, w50605, w50606, w50607, w50608, w50609, w50610, w50611, w50612, w50613, w50614, w50615, w50616, w50617, w50618, w50619, w50620, w50621, w50622, w50623, w50624, w50625, w50626, w50627, w50628, w50629, w50630, w50631, w50632, w50633, w50634, w50635, w50636, w50637, w50638, w50639, w50640, w50641, w50642, w50643, w50644, w50645, w50646, w50647, w50648, w50649, w50650, w50651, w50652, w50653, w50654, w50655, w50656, w50657, w50658, w50659, w50660, w50661, w50662, w50663, w50664, w50665, w50666, w50667, w50668, w50669, w50670, w50671, w50672, w50673, w50674, w50675, w50676, w50677, w50678, w50679, w50680, w50681, w50682, w50683, w50684, w50685, w50686, w50687, w50688, w50689, w50690, w50691, w50692, w50693, w50694, w50695, w50696, w50697, w50698, w50699, w50700, w50701, w50702, w50703, w50704, w50705, w50706, w50707, w50708, w50709, w50710, w50711, w50712, w50713, w50714, w50715, w50716, w50717, w50718, w50719, w50720, w50721, w50722, w50723, w50724, w50725, w50726, w50727, w50728, w50729, w50730, w50731, w50732, w50733, w50734, w50735, w50736, w50737, w50738, w50739, w50740, w50741, w50742, w50743, w50744, w50745, w50746, w50747, w50748, w50749, w50750, w50751, w50752, w50753, w50754, w50755, w50756, w50757, w50758, w50759, w50760, w50761, w50762, w50763, w50764, w50765, w50766, w50767, w50768, w50769, w50770, w50771, w50772, w50773, w50774, w50775, w50776, w50777, w50778, w50779, w50780, w50781, w50782, w50783, w50784, w50785, w50786, w50787, w50788, w50789, w50790, w50791, w50792, w50793, w50794, w50795, w50796, w50797, w50798, w50799, w50800, w50801, w50802, w50803, w50804, w50805, w50806, w50807, w50808, w50809, w50810, w50811, w50812, w50813, w50814, w50815, w50816, w50817, w50818, w50819, w50820, w50821, w50822, w50823, w50824, w50825, w50826, w50827, w50828, w50829, w50830, w50831, w50832, w50833, w50834, w50835, w50836, w50837, w50838, w50839, w50840, w50841, w50842, w50843, w50844, w50845, w50846, w50847, w50848, w50849, w50850, w50851, w50852, w50853, w50854, w50855, w50856, w50857, w50858, w50859, w50860, w50861, w50862, w50863, w50864, w50865, w50866, w50867, w50868, w50869, w50870, w50871, w50872, w50873, w50874, w50875, w50876, w50877, w50878, w50879, w50880, w50881, w50882, w50883, w50884, w50885, w50886, w50887, w50888, w50889, w50890, w50891, w50892, w50893, w50894, w50895, w50896, w50897, w50898, w50899, w50900, w50901, w50902, w50903, w50904, w50905, w50906, w50907, w50908, w50909, w50910, w50911, w50912, w50913, w50914, w50915, w50916, w50917, w50918, w50919, w50920, w50921, w50922, w50923, w50924, w50925, w50926, w50927, w50928, w50929, w50930, w50931, w50932, w50933, w50934, w50935, w50936, w50937, w50938, w50939, w50940, w50941, w50942, w50943, w50944, w50945, w50946, w50947, w50948, w50949, w50950, w50951, w50952, w50953, w50954, w50955, w50956, w50957, w50958, w50959, w50960, w50961, w50962, w50963, w50964, w50965, w50966, w50967, w50968, w50969, w50970, w50971, w50972, w50973, w50974, w50975, w50976, w50977, w50978, w50979, w50980, w50981, w50982, w50983, w50984, w50985, w50986, w50987, w50988, w50989, w50990, w50991, w50992, w50993, w50994, w50995, w50996, w50997, w50998, w50999, w51000, w51001, w51002, w51003, w51004, w51005, w51006, w51007, w51008, w51009, w51010, w51011, w51012, w51013, w51014, w51015, w51016, w51017, w51018, w51019, w51020, w51021, w51022, w51023, w51024, w51025, w51026, w51027, w51028, w51029, w51030, w51031, w51032, w51033, w51034, w51035, w51036, w51037, w51038, w51039, w51040, w51041, w51042, w51043, w51044, w51045, w51046, w51047, w51048, w51049, w51050, w51051, w51052, w51053, w51054, w51055, w51056, w51057, w51058, w51059, w51060, w51061, w51062, w51063, w51064, w51065, w51066, w51067, w51068, w51069, w51070, w51071, w51072, w51073, w51074, w51075, w51076, w51077, w51078, w51079, w51080, w51081, w51082, w51083, w51084, w51085, w51086, w51087, w51088, w51089, w51090, w51091, w51092, w51093, w51094, w51095, w51096, w51097, w51098, w51099, w51100, w51101, w51102, w51103, w51104, w51105, w51106, w51107, w51108, w51109, w51110, w51111, w51112, w51113, w51114, w51115, w51116, w51117, w51118, w51119, w51120, w51121, w51122, w51123, w51124, w51125, w51126, w51127, w51128, w51129, w51130, w51131, w51132, w51133, w51134, w51135, w51136, w51137, w51138, w51139, w51140, w51141, w51142, w51143, w51144, w51145, w51146, w51147, w51148, w51149, w51150, w51151, w51152, w51153, w51154, w51155, w51156, w51157, w51158, w51159, w51160, w51161, w51162, w51163, w51164, w51165, w51166, w51167, w51168, w51169, w51170, w51171, w51172, w51173, w51174, w51175, w51176, w51177, w51178, w51179, w51180, w51181, w51182, w51183, w51184, w51185, w51186, w51187, w51188, w51189, w51190, w51191, w51192, w51193, w51194, w51195, w51196, w51197, w51198, w51199, w51200, w51201, w51202, w51203, w51204, w51205, w51206, w51207, w51208, w51209, w51210, w51211, w51212, w51213, w51214, w51215, w51216, w51217, w51218, w51219, w51220, w51221, w51222, w51223, w51224, w51225, w51226, w51227, w51228, w51229, w51230, w51231, w51232, w51233, w51234, w51235, w51236, w51237, w51238, w51239, w51240, w51241, w51242, w51243, w51244, w51245, w51246, w51247, w51248, w51249, w51250, w51251, w51252, w51253, w51254, w51255, w51256, w51257, w51258, w51259, w51260, w51261, w51262, w51263, w51264, w51265, w51266, w51267, w51268, w51269, w51270, w51271, w51272, w51273, w51274, w51275, w51276, w51277, w51278, w51279, w51280, w51281, w51282, w51283, w51284, w51285, w51286, w51287, w51288, w51289, w51290, w51291, w51292, w51293, w51294, w51295, w51296, w51297, w51298, w51299, w51300, w51301, w51302, w51303, w51304, w51305, w51306, w51307, w51308, w51309, w51310, w51311, w51312, w51313, w51314, w51315, w51316, w51317, w51318, w51319, w51320, w51321, w51322, w51323, w51324, w51325, w51326, w51327, w51328, w51329, w51330, w51331, w51332, w51333, w51334, w51335, w51336, w51337, w51338, w51339, w51340, w51341, w51342, w51343, w51344, w51345, w51346, w51347, w51348, w51349, w51350, w51351, w51352, w51353, w51354, w51355, w51356, w51357, w51358, w51359, w51360, w51361, w51362, w51363, w51364, w51365, w51366, w51367, w51368, w51369, w51370, w51371, w51372, w51373, w51374, w51375, w51376, w51377, w51378, w51379, w51380, w51381, w51382, w51383, w51384, w51385, w51386, w51387, w51388, w51389, w51390, w51391, w51392, w51393, w51394, w51395, w51396, w51397, w51398, w51399, w51400, w51401, w51402, w51403, w51404, w51405, w51406, w51407, w51408, w51409, w51410, w51411, w51412, w51413, w51414, w51415, w51416, w51417, w51418, w51419, w51420, w51421, w51422, w51423, w51424, w51425, w51426, w51427, w51428, w51429, w51430, w51431, w51432, w51433, w51434, w51435, w51436, w51437, w51438, w51439, w51440, w51441, w51442, w51443, w51444, w51445, w51446, w51447, w51448, w51449, w51450, w51451, w51452, w51453, w51454, w51455, w51456, w51457, w51458, w51459, w51460, w51461, w51462, w51463, w51464, w51465, w51466, w51467, w51468, w51469, w51470, w51471, w51472, w51473, w51474, w51475, w51476, w51477, w51478, w51479, w51480, w51481, w51482, w51483, w51484, w51485, w51486, w51487, w51488, w51489, w51490, w51491, w51492, w51493, w51494, w51495, w51496, w51497, w51498, w51499, w51500, w51501, w51502, w51503, w51504, w51505, w51506, w51507, w51508, w51509, w51510, w51511, w51512, w51513, w51514, w51515, w51516, w51517, w51518, w51519, w51520, w51521, w51522, w51523, w51524, w51525, w51526, w51527, w51528, w51529, w51530, w51531, w51532, w51533, w51534, w51535, w51536, w51537, w51538, w51539, w51540, w51541, w51542, w51543, w51544, w51545, w51546, w51547, w51548, w51549, w51550, w51551, w51552, w51553, w51554, w51555, w51556, w51557, w51558, w51559, w51560, w51561, w51562, w51563, w51564, w51565, w51566, w51567, w51568, w51569, w51570, w51571, w51572, w51573, w51574, w51575, w51576, w51577, w51578, w51579, w51580, w51581, w51582, w51583, w51584, w51585, w51586, w51587, w51588, w51589, w51590, w51591, w51592, w51593, w51594, w51595, w51596, w51597, w51598, w51599, w51600, w51601, w51602, w51603, w51604, w51605, w51606, w51607, w51608, w51609, w51610, w51611, w51612, w51613, w51614, w51615, w51616, w51617, w51618, w51619, w51620, w51621, w51622, w51623, w51624, w51625, w51626, w51627, w51628, w51629, w51630, w51631, w51632, w51633, w51634, w51635, w51636, w51637, w51638, w51639, w51640, w51641, w51642, w51643, w51644, w51645, w51646, w51647, w51648, w51649, w51650, w51651, w51652, w51653, w51654, w51655, w51656, w51657, w51658, w51659, w51660, w51661, w51662, w51663, w51664, w51665, w51666, w51667, w51668, w51669, w51670, w51671, w51672, w51673, w51674, w51675, w51676, w51677, w51678, w51679, w51680, w51681, w51682, w51683, w51684, w51685, w51686, w51687, w51688, w51689, w51690, w51691, w51692, w51693, w51694, w51695, w51696, w51697, w51698, w51699, w51700, w51701, w51702, w51703, w51704, w51705, w51706, w51707, w51708, w51709, w51710, w51711, w51712, w51713, w51714, w51715, w51716, w51717, w51718, w51719, w51720, w51721, w51722, w51723, w51724, w51725, w51726, w51727, w51728, w51729, w51730, w51731, w51732, w51733, w51734, w51735, w51736, w51737, w51738, w51739, w51740, w51741, w51742, w51743, w51744, w51745, w51746, w51747, w51748, w51749, w51750, w51751, w51752, w51753, w51754, w51755, w51756, w51757, w51758, w51759, w51760, w51761, w51762, w51763, w51764, w51765, w51766, w51767, w51768, w51769, w51770, w51771, w51772, w51773, w51774, w51775, w51776, w51777, w51778, w51779, w51780, w51781, w51782, w51783, w51784, w51785, w51786, w51787, w51788, w51789, w51790, w51791, w51792, w51793, w51794, w51795, w51796, w51797, w51798, w51799, w51800, w51801, w51802, w51803, w51804, w51805, w51806, w51807, w51808, w51809, w51810, w51811, w51812, w51813, w51814, w51815, w51816, w51817, w51818, w51819, w51820, w51821, w51822, w51823, w51824, w51825, w51826, w51827, w51828, w51829, w51830, w51831, w51832, w51833, w51834, w51835, w51836, w51837, w51838, w51839, w51840, w51841, w51842, w51843, w51844, w51845, w51846, w51847, w51848, w51849, w51850, w51851, w51852, w51853, w51854, w51855, w51856, w51857, w51858, w51859, w51860, w51861, w51862, w51863, w51864, w51865, w51866, w51867, w51868, w51869, w51870, w51871, w51872, w51873, w51874, w51875, w51876, w51877, w51878, w51879, w51880, w51881, w51882, w51883, w51884, w51885, w51886, w51887, w51888, w51889, w51890, w51891, w51892, w51893, w51894, w51895, w51896, w51897, w51898, w51899, w51900, w51901, w51902, w51903, w51904, w51905, w51906, w51907, w51908, w51909, w51910, w51911, w51912, w51913, w51914, w51915, w51916, w51917, w51918, w51919, w51920, w51921, w51922, w51923, w51924, w51925, w51926, w51927, w51928, w51929, w51930, w51931, w51932, w51933, w51934, w51935, w51936, w51937, w51938, w51939, w51940, w51941, w51942, w51943, w51944, w51945, w51946, w51947, w51948, w51949, w51950, w51951, w51952, w51953, w51954, w51955, w51956, w51957, w51958, w51959, w51960, w51961, w51962, w51963, w51964, w51965, w51966, w51967, w51968, w51969, w51970, w51971, w51972, w51973, w51974, w51975, w51976, w51977, w51978, w51979, w51980, w51981, w51982, w51983, w51984, w51985, w51986, w51987, w51988, w51989, w51990, w51991, w51992, w51993, w51994, w51995, w51996, w51997, w51998, w51999, w52000, w52001, w52002, w52003, w52004, w52005, w52006, w52007, w52008, w52009, w52010, w52011, w52012, w52013, w52014, w52015, w52016, w52017, w52018, w52019, w52020, w52021, w52022, w52023, w52024, w52025, w52026, w52027, w52028, w52029, w52030, w52031, w52032, w52033, w52034, w52035, w52036, w52037, w52038, w52039, w52040, w52041, w52042, w52043, w52044, w52045, w52046, w52047, w52048, w52049, w52050, w52051, w52052, w52053, w52054, w52055, w52056, w52057, w52058, w52059, w52060, w52061, w52062, w52063, w52064, w52065, w52066, w52067, w52068, w52069, w52070, w52071, w52072, w52073, w52074, w52075, w52076, w52077, w52078, w52079, w52080, w52081, w52082, w52083, w52084, w52085, w52086, w52087, w52088, w52089, w52090, w52091, w52092, w52093, w52094, w52095, w52096, w52097, w52098, w52099, w52100, w52101, w52102, w52103, w52104, w52105, w52106, w52107, w52108, w52109, w52110, w52111, w52112, w52113, w52114, w52115, w52116, w52117, w52118, w52119, w52120, w52121, w52122, w52123, w52124, w52125, w52126, w52127, w52128, w52129, w52130, w52131, w52132, w52133, w52134, w52135, w52136, w52137, w52138, w52139, w52140, w52141, w52142, w52143, w52144, w52145, w52146, w52147, w52148, w52149, w52150, w52151, w52152, w52153, w52154, w52155, w52156, w52157, w52158, w52159, w52160, w52161, w52162, w52163, w52164, w52165, w52166, w52167, w52168, w52169, w52170, w52171, w52172, w52173, w52174, w52175, w52176, w52177, w52178, w52179, w52180, w52181, w52182, w52183, w52184, w52185, w52186, w52187, w52188, w52189, w52190, w52191, w52192, w52193, w52194, w52195, w52196, w52197, w52198, w52199, w52200, w52201, w52202, w52203, w52204, w52205, w52206, w52207, w52208, w52209, w52210, w52211, w52212, w52213, w52214, w52215, w52216, w52217, w52218, w52219, w52220, w52221, w52222, w52223, w52224, w52225, w52226, w52227, w52228, w52229, w52230, w52231, w52232, w52233, w52234, w52235, w52236, w52237, w52238, w52239, w52240, w52241, w52242, w52243, w52244, w52245, w52246, w52247, w52248, w52249, w52250, w52251, w52252, w52253, w52254, w52255, w52256, w52257, w52258, w52259, w52260, w52261, w52262, w52263, w52264, w52265, w52266, w52267, w52268, w52269, w52270, w52271, w52272, w52273, w52274, w52275, w52276, w52277, w52278, w52279, w52280, w52281, w52282, w52283, w52284, w52285, w52286, w52287, w52288, w52289, w52290, w52291, w52292, w52293, w52294, w52295, w52296, w52297, w52298, w52299, w52300, w52301, w52302, w52303, w52304, w52305, w52306, w52307, w52308, w52309, w52310, w52311, w52312, w52313, w52314, w52315, w52316, w52317, w52318, w52319, w52320, w52321, w52322, w52323, w52324, w52325, w52326, w52327, w52328, w52329, w52330, w52331, w52332, w52333, w52334, w52335, w52336, w52337, w52338, w52339, w52340, w52341, w52342, w52343, w52344, w52345, w52346, w52347, w52348, w52349, w52350, w52351, w52352, w52353, w52354, w52355, w52356, w52357, w52358, w52359, w52360, w52361, w52362, w52363, w52364, w52365, w52366, w52367, w52368, w52369, w52370, w52371, w52372, w52373, w52374, w52375, w52376, w52377, w52378, w52379, w52380, w52381, w52382, w52383, w52384, w52385, w52386, w52387, w52388, w52389, w52390, w52391, w52392, w52393, w52394, w52395, w52396, w52397, w52398, w52399, w52400, w52401, w52402, w52403, w52404, w52405, w52406, w52407, w52408, w52409, w52410, w52411, w52412, w52413, w52414, w52415, w52416, w52417, w52418, w52419, w52420, w52421, w52422, w52423, w52424, w52425, w52426, w52427, w52428, w52429, w52430, w52431, w52432, w52433, w52434, w52435, w52436, w52437, w52438, w52439, w52440, w52441, w52442, w52443, w52444, w52445, w52446, w52447, w52448, w52449, w52450, w52451, w52452, w52453, w52454, w52455, w52456, w52457, w52458, w52459, w52460, w52461, w52462, w52463, w52464, w52465, w52466, w52467, w52468, w52469, w52470, w52471, w52472, w52473, w52474, w52475, w52476, w52477, w52478, w52479, w52480, w52481, w52482, w52483, w52484, w52485, w52486, w52487, w52488, w52489, w52490, w52491, w52492, w52493, w52494, w52495, w52496, w52497, w52498, w52499, w52500, w52501, w52502, w52503, w52504, w52505, w52506, w52507, w52508, w52509, w52510, w52511, w52512, w52513, w52514, w52515, w52516, w52517, w52518, w52519, w52520, w52521, w52522, w52523, w52524, w52525, w52526, w52527, w52528, w52529, w52530, w52531, w52532, w52533, w52534, w52535, w52536, w52537, w52538, w52539, w52540, w52541, w52542, w52543, w52544, w52545, w52546, w52547, w52548, w52549, w52550, w52551, w52552, w52553, w52554, w52555, w52556, w52557, w52558, w52559, w52560, w52561, w52562, w52563, w52564, w52565, w52566, w52567, w52568, w52569, w52570, w52571, w52572, w52573, w52574, w52575, w52576, w52577, w52578, w52579, w52580, w52581, w52582, w52583, w52584, w52585, w52586, w52587, w52588, w52589, w52590, w52591, w52592, w52593, w52594, w52595, w52596, w52597, w52598, w52599, w52600, w52601, w52602, w52603, w52604, w52605, w52606, w52607, w52608, w52609, w52610, w52611, w52612, w52613, w52614, w52615, w52616, w52617, w52618, w52619, w52620, w52621, w52622, w52623, w52624, w52625, w52626, w52627, w52628, w52629, w52630, w52631, w52632, w52633, w52634, w52635, w52636, w52637, w52638, w52639, w52640, w52641, w52642, w52643, w52644, w52645, w52646, w52647, w52648, w52649, w52650, w52651, w52652, w52653, w52654, w52655, w52656, w52657, w52658, w52659, w52660, w52661, w52662, w52663, w52664, w52665, w52666, w52667, w52668, w52669, w52670, w52671, w52672, w52673, w52674, w52675, w52676, w52677, w52678, w52679, w52680, w52681, w52682, w52683, w52684, w52685, w52686, w52687, w52688, w52689, w52690, w52691, w52692, w52693, w52694, w52695, w52696, w52697, w52698, w52699, w52700, w52701, w52702, w52703, w52704, w52705, w52706, w52707, w52708, w52709, w52710, w52711, w52712, w52713, w52714, w52715, w52716, w52717, w52718, w52719, w52720, w52721, w52722, w52723, w52724, w52725, w52726, w52727, w52728, w52729, w52730, w52731, w52732, w52733, w52734, w52735, w52736, w52737, w52738, w52739, w52740, w52741, w52742, w52743, w52744, w52745, w52746, w52747, w52748, w52749, w52750, w52751, w52752, w52753, w52754, w52755, w52756, w52757, w52758, w52759, w52760, w52761, w52762, w52763, w52764, w52765, w52766, w52767, w52768, w52769, w52770, w52771, w52772, w52773, w52774, w52775, w52776, w52777, w52778, w52779, w52780, w52781, w52782, w52783, w52784, w52785, w52786, w52787, w52788, w52789, w52790, w52791, w52792, w52793, w52794, w52795, w52796, w52797, w52798, w52799, w52800, w52801, w52802, w52803, w52804, w52805, w52806, w52807, w52808, w52809, w52810, w52811, w52812, w52813, w52814, w52815, w52816, w52817, w52818, w52819, w52820, w52821, w52822, w52823, w52824, w52825, w52826, w52827, w52828, w52829, w52830, w52831, w52832, w52833, w52834, w52835, w52836, w52837, w52838, w52839, w52840, w52841, w52842, w52843, w52844, w52845, w52846, w52847, w52848, w52849, w52850, w52851, w52852, w52853, w52854, w52855, w52856, w52857, w52858, w52859, w52860, w52861, w52862, w52863, w52864, w52865, w52866, w52867, w52868, w52869, w52870, w52871, w52872, w52873, w52874, w52875, w52876, w52877, w52878, w52879, w52880, w52881, w52882, w52883, w52884, w52885, w52886, w52887, w52888, w52889, w52890, w52891, w52892, w52893, w52894, w52895, w52896, w52897, w52898, w52899, w52900, w52901, w52902, w52903, w52904, w52905, w52906, w52907, w52908, w52909, w52910, w52911, w52912, w52913, w52914, w52915, w52916, w52917, w52918, w52919, w52920, w52921, w52922, w52923, w52924, w52925, w52926, w52927, w52928, w52929, w52930, w52931, w52932, w52933, w52934, w52935, w52936, w52937, w52938, w52939, w52940, w52941, w52942, w52943, w52944, w52945, w52946, w52947, w52948, w52949, w52950, w52951, w52952, w52953, w52954, w52955, w52956, w52957, w52958, w52959, w52960, w52961, w52962, w52963, w52964, w52965, w52966, w52967, w52968, w52969, w52970, w52971, w52972, w52973, w52974, w52975, w52976, w52977, w52978, w52979, w52980, w52981, w52982, w52983, w52984, w52985, w52986, w52987, w52988, w52989, w52990, w52991, w52992, w52993, w52994, w52995, w52996, w52997, w52998, w52999, w53000, w53001, w53002, w53003, w53004, w53005, w53006, w53007, w53008, w53009, w53010, w53011, w53012, w53013, w53014, w53015, w53016, w53017, w53018, w53019, w53020, w53021, w53022, w53023, w53024, w53025, w53026, w53027, w53028, w53029, w53030, w53031, w53032, w53033, w53034, w53035, w53036, w53037, w53038, w53039, w53040, w53041, w53042, w53043, w53044, w53045, w53046, w53047, w53048, w53049, w53050, w53051, w53052, w53053, w53054, w53055, w53056, w53057, w53058, w53059, w53060, w53061, w53062, w53063, w53064, w53065, w53066, w53067, w53068, w53069, w53070, w53071, w53072, w53073, w53074, w53075, w53076, w53077, w53078, w53079, w53080, w53081, w53082, w53083, w53084, w53085, w53086, w53087, w53088, w53089, w53090, w53091, w53092, w53093, w53094, w53095, w53096, w53097, w53098, w53099, w53100, w53101, w53102, w53103, w53104, w53105, w53106, w53107, w53108, w53109, w53110, w53111, w53112, w53113, w53114, w53115, w53116, w53117, w53118, w53119, w53120, w53121, w53122, w53123, w53124, w53125, w53126, w53127, w53128, w53129, w53130, w53131, w53132, w53133, w53134, w53135, w53136, w53137, w53138, w53139, w53140, w53141, w53142, w53143, w53144, w53145, w53146, w53147, w53148, w53149, w53150, w53151, w53152, w53153, w53154, w53155, w53156, w53157, w53158, w53159, w53160, w53161, w53162, w53163, w53164, w53165, w53166, w53167, w53168, w53169, w53170, w53171, w53172, w53173, w53174, w53175, w53176, w53177, w53178, w53179, w53180, w53181, w53182, w53183, w53184, w53185, w53186, w53187, w53188, w53189, w53190, w53191, w53192, w53193, w53194, w53195, w53196, w53197, w53198, w53199, w53200, w53201, w53202, w53203, w53204, w53205, w53206, w53207, w53208, w53209, w53210, w53211, w53212, w53213, w53214, w53215, w53216, w53217, w53218, w53219, w53220, w53221, w53222, w53223, w53224, w53225, w53226, w53227, w53228, w53229, w53230, w53231, w53232, w53233, w53234, w53235, w53236, w53237, w53238, w53239, w53240, w53241, w53242, w53243, w53244, w53245, w53246, w53247, w53248, w53249, w53250, w53251, w53252, w53253, w53254, w53255, w53256, w53257, w53258, w53259, w53260, w53261, w53262, w53263, w53264, w53265, w53266, w53267, w53268, w53269, w53270, w53271, w53272, w53273, w53274, w53275, w53276, w53277, w53278, w53279, w53280, w53281, w53282, w53283, w53284, w53285, w53286, w53287, w53288, w53289, w53290, w53291, w53292, w53293, w53294, w53295, w53296, w53297, w53298, w53299, w53300, w53301, w53302, w53303, w53304, w53305, w53306, w53307, w53308, w53309, w53310, w53311, w53312, w53313, w53314, w53315, w53316, w53317, w53318, w53319, w53320, w53321, w53322, w53323, w53324, w53325, w53326, w53327, w53328, w53329, w53330, w53331, w53332, w53333, w53334, w53335, w53336, w53337, w53338, w53339, w53340, w53341, w53342, w53343, w53344, w53345, w53346, w53347, w53348, w53349, w53350, w53351, w53352, w53353, w53354, w53355, w53356, w53357, w53358, w53359, w53360, w53361, w53362, w53363, w53364, w53365, w53366, w53367, w53368, w53369, w53370, w53371, w53372, w53373, w53374, w53375, w53376, w53377, w53378, w53379, w53380, w53381, w53382, w53383, w53384, w53385, w53386, w53387, w53388, w53389, w53390, w53391, w53392, w53393, w53394, w53395, w53396, w53397, w53398, w53399, w53400, w53401, w53402, w53403, w53404, w53405, w53406, w53407, w53408, w53409, w53410, w53411, w53412, w53413, w53414, w53415, w53416, w53417, w53418, w53419, w53420, w53421, w53422, w53423, w53424, w53425, w53426, w53427, w53428, w53429, w53430, w53431, w53432, w53433, w53434, w53435, w53436, w53437, w53438, w53439, w53440, w53441, w53442, w53443, w53444, w53445, w53446, w53447, w53448, w53449, w53450, w53451, w53452, w53453, w53454, w53455, w53456, w53457, w53458, w53459, w53460, w53461, w53462, w53463, w53464, w53465, w53466, w53467, w53468, w53469, w53470, w53471, w53472, w53473, w53474, w53475, w53476, w53477, w53478, w53479, w53480, w53481, w53482, w53483, w53484, w53485, w53486, w53487, w53488, w53489, w53490, w53491, w53492, w53493, w53494, w53495, w53496, w53497, w53498, w53499, w53500, w53501, w53502, w53503, w53504, w53505, w53506, w53507, w53508, w53509, w53510, w53511, w53512, w53513, w53514, w53515, w53516, w53517, w53518, w53519, w53520, w53521, w53522, w53523, w53524, w53525, w53526, w53527, w53528, w53529, w53530, w53531, w53532, w53533, w53534, w53535, w53536, w53537, w53538, w53539, w53540, w53541, w53542, w53543, w53544, w53545, w53546, w53547, w53548, w53549, w53550, w53551, w53552, w53553, w53554, w53555, w53556, w53557, w53558, w53559, w53560, w53561, w53562, w53563, w53564, w53565, w53566, w53567, w53568, w53569, w53570, w53571, w53572, w53573, w53574, w53575, w53576, w53577, w53578, w53579, w53580, w53581, w53582, w53583, w53584, w53585, w53586, w53587, w53588, w53589, w53590, w53591, w53592, w53593, w53594, w53595, w53596, w53597, w53598, w53599, w53600, w53601, w53602, w53603, w53604, w53605, w53606, w53607, w53608, w53609, w53610, w53611, w53612, w53613, w53614, w53615, w53616, w53617, w53618, w53619, w53620, w53621, w53622, w53623, w53624, w53625, w53626, w53627, w53628, w53629, w53630, w53631, w53632, w53633, w53634, w53635, w53636, w53637, w53638, w53639, w53640, w53641, w53642, w53643, w53644, w53645, w53646, w53647, w53648, w53649, w53650, w53651, w53652, w53653, w53654, w53655, w53656, w53657, w53658, w53659, w53660, w53661, w53662, w53663, w53664, w53665, w53666, w53667, w53668, w53669, w53670, w53671, w53672, w53673, w53674, w53675, w53676, w53677, w53678, w53679, w53680, w53681, w53682, w53683, w53684, w53685, w53686, w53687, w53688, w53689, w53690, w53691, w53692, w53693, w53694, w53695, w53696, w53697, w53698, w53699, w53700, w53701, w53702, w53703, w53704, w53705, w53706, w53707, w53708, w53709, w53710, w53711, w53712, w53713, w53714, w53715, w53716, w53717, w53718, w53719, w53720, w53721, w53722, w53723, w53724, w53725, w53726, w53727, w53728, w53729, w53730, w53731, w53732, w53733, w53734, w53735, w53736, w53737, w53738, w53739, w53740, w53741, w53742, w53743, w53744, w53745, w53746, w53747, w53748, w53749, w53750, w53751, w53752, w53753, w53754, w53755, w53756, w53757, w53758, w53759, w53760, w53761, w53762, w53763, w53764, w53765, w53766, w53767, w53768, w53769, w53770, w53771, w53772, w53773, w53774, w53775, w53776, w53777, w53778, w53779, w53780, w53781, w53782, w53783, w53784, w53785, w53786, w53787, w53788, w53789, w53790, w53791, w53792, w53793, w53794, w53795, w53796, w53797, w53798, w53799, w53800, w53801, w53802, w53803, w53804, w53805, w53806, w53807, w53808, w53809, w53810, w53811, w53812, w53813, w53814, w53815, w53816, w53817, w53818, w53819, w53820, w53821, w53822, w53823, w53824, w53825, w53826, w53827, w53828, w53829, w53830, w53831, w53832, w53833, w53834, w53835, w53836, w53837, w53838, w53839, w53840, w53841, w53842, w53843, w53844, w53845, w53846, w53847, w53848, w53849, w53850, w53851, w53852, w53853, w53854, w53855, w53856, w53857, w53858, w53859, w53860, w53861, w53862, w53863, w53864, w53865, w53866, w53867, w53868, w53869, w53870, w53871, w53872, w53873, w53874, w53875, w53876, w53877, w53878, w53879, w53880, w53881, w53882, w53883, w53884, w53885, w53886, w53887, w53888, w53889, w53890, w53891, w53892, w53893, w53894, w53895, w53896, w53897, w53898, w53899, w53900, w53901, w53902, w53903, w53904, w53905, w53906, w53907, w53908, w53909, w53910, w53911, w53912, w53913, w53914, w53915, w53916, w53917, w53918, w53919, w53920, w53921, w53922, w53923, w53924, w53925, w53926, w53927, w53928, w53929, w53930, w53931, w53932, w53933, w53934, w53935, w53936, w53937, w53938, w53939, w53940, w53941, w53942, w53943, w53944, w53945, w53946, w53947, w53948, w53949, w53950, w53951, w53952, w53953, w53954, w53955, w53956, w53957, w53958, w53959, w53960, w53961, w53962, w53963, w53964, w53965, w53966, w53967, w53968, w53969, w53970, w53971, w53972, w53973, w53974, w53975, w53976, w53977, w53978, w53979, w53980, w53981, w53982, w53983, w53984, w53985, w53986, w53987, w53988, w53989, w53990, w53991, w53992, w53993, w53994, w53995, w53996, w53997, w53998, w53999, w54000, w54001, w54002, w54003, w54004, w54005, w54006, w54007, w54008, w54009, w54010, w54011, w54012, w54013, w54014, w54015, w54016, w54017, w54018, w54019, w54020, w54021, w54022, w54023, w54024, w54025, w54026, w54027, w54028, w54029, w54030, w54031, w54032, w54033, w54034, w54035, w54036, w54037, w54038, w54039, w54040, w54041, w54042, w54043, w54044, w54045, w54046, w54047, w54048, w54049, w54050, w54051, w54052, w54053, w54054, w54055, w54056, w54057, w54058, w54059, w54060, w54061, w54062, w54063, w54064, w54065, w54066, w54067, w54068, w54069, w54070, w54071, w54072, w54073, w54074, w54075, w54076, w54077, w54078, w54079, w54080, w54081, w54082, w54083, w54084, w54085, w54086, w54087, w54088, w54089, w54090, w54091, w54092, w54093, w54094, w54095, w54096, w54097, w54098, w54099, w54100, w54101, w54102, w54103, w54104, w54105, w54106, w54107, w54108, w54109, w54110, w54111, w54112, w54113, w54114, w54115, w54116, w54117, w54118, w54119, w54120, w54121, w54122, w54123, w54124, w54125, w54126, w54127, w54128, w54129, w54130, w54131, w54132, w54133, w54134, w54135, w54136, w54137, w54138, w54139, w54140, w54141, w54142, w54143, w54144, w54145, w54146, w54147, w54148, w54149, w54150, w54151, w54152, w54153, w54154, w54155, w54156, w54157, w54158, w54159, w54160, w54161, w54162, w54163, w54164, w54165, w54166, w54167, w54168, w54169, w54170, w54171, w54172, w54173, w54174, w54175, w54176, w54177, w54178, w54179, w54180, w54181, w54182, w54183, w54184, w54185, w54186, w54187, w54188, w54189, w54190, w54191, w54192, w54193, w54194, w54195, w54196, w54197, w54198, w54199, w54200, w54201, w54202, w54203, w54204, w54205, w54206, w54207, w54208, w54209, w54210, w54211, w54212, w54213, w54214, w54215, w54216, w54217, w54218, w54219, w54220, w54221, w54222, w54223, w54224, w54225, w54226, w54227, w54228, w54229, w54230, w54231, w54232, w54233, w54234, w54235, w54236, w54237, w54238, w54239, w54240, w54241, w54242, w54243, w54244, w54245, w54246, w54247, w54248, w54249, w54250, w54251, w54252, w54253, w54254, w54255, w54256, w54257, w54258, w54259, w54260, w54261, w54262, w54263, w54264, w54265, w54266, w54267, w54268, w54269, w54270, w54271, w54272, w54273, w54274, w54275, w54276, w54277, w54278, w54279, w54280, w54281, w54282, w54283, w54284, w54285, w54286, w54287, w54288, w54289, w54290, w54291, w54292, w54293, w54294, w54295, w54296, w54297, w54298, w54299, w54300, w54301, w54302, w54303, w54304, w54305, w54306, w54307, w54308, w54309, w54310, w54311, w54312, w54313, w54314, w54315, w54316, w54317, w54318, w54319, w54320, w54321, w54322, w54323, w54324, w54325, w54326, w54327, w54328, w54329, w54330, w54331, w54332, w54333, w54334, w54335, w54336, w54337, w54338, w54339, w54340, w54341, w54342, w54343, w54344, w54345, w54346, w54347, w54348, w54349, w54350, w54351, w54352, w54353, w54354, w54355, w54356, w54357, w54358, w54359, w54360, w54361, w54362, w54363, w54364, w54365, w54366, w54367, w54368, w54369, w54370, w54371, w54372, w54373, w54374, w54375, w54376, w54377, w54378, w54379, w54380, w54381, w54382, w54383, w54384, w54385, w54386, w54387, w54388, w54389, w54390, w54391, w54392, w54393, w54394, w54395, w54396, w54397, w54398, w54399, w54400, w54401, w54402, w54403, w54404, w54405, w54406, w54407, w54408, w54409, w54410, w54411, w54412, w54413, w54414, w54415, w54416, w54417, w54418, w54419, w54420, w54421, w54422, w54423, w54424, w54425, w54426, w54427, w54428, w54429, w54430, w54431, w54432, w54433, w54434, w54435, w54436, w54437, w54438, w54439, w54440, w54441, w54442, w54443, w54444, w54445, w54446, w54447, w54448, w54449, w54450, w54451, w54452, w54453, w54454, w54455, w54456, w54457, w54458, w54459, w54460, w54461, w54462, w54463, w54464, w54465, w54466, w54467, w54468, w54469, w54470, w54471, w54472, w54473, w54474, w54475, w54476, w54477, w54478, w54479, w54480, w54481, w54482, w54483, w54484, w54485, w54486, w54487, w54488, w54489, w54490, w54491, w54492, w54493, w54494, w54495, w54496, w54497, w54498, w54499, w54500, w54501, w54502, w54503, w54504, w54505, w54506, w54507, w54508, w54509, w54510, w54511, w54512, w54513, w54514, w54515, w54516, w54517, w54518, w54519, w54520, w54521, w54522, w54523, w54524, w54525, w54526, w54527, w54528, w54529, w54530, w54531, w54532, w54533, w54534, w54535, w54536, w54537, w54538, w54539, w54540, w54541, w54542, w54543, w54544, w54545, w54546, w54547, w54548, w54549, w54550, w54551, w54552, w54553, w54554, w54555, w54556, w54557, w54558, w54559, w54560, w54561, w54562, w54563, w54564, w54565, w54566, w54567, w54568, w54569, w54570, w54571, w54572, w54573, w54574, w54575, w54576, w54577, w54578, w54579, w54580, w54581, w54582, w54583, w54584, w54585, w54586, w54587, w54588, w54589, w54590, w54591, w54592, w54593, w54594, w54595, w54596, w54597, w54598, w54599, w54600, w54601, w54602, w54603, w54604, w54605, w54606, w54607, w54608, w54609, w54610, w54611, w54612, w54613, w54614, w54615, w54616, w54617, w54618, w54619, w54620, w54621, w54622, w54623, w54624, w54625, w54626, w54627, w54628, w54629, w54630, w54631, w54632, w54633, w54634, w54635, w54636, w54637, w54638, w54639, w54640, w54641, w54642, w54643, w54644, w54645, w54646, w54647, w54648, w54649, w54650, w54651, w54652, w54653, w54654, w54655, w54656, w54657, w54658, w54659, w54660, w54661, w54662, w54663, w54664, w54665, w54666, w54667, w54668, w54669, w54670, w54671, w54672, w54673, w54674, w54675, w54676, w54677, w54678, w54679, w54680, w54681, w54682, w54683, w54684, w54685, w54686, w54687, w54688, w54689, w54690, w54691, w54692, w54693, w54694, w54695, w54696, w54697, w54698, w54699, w54700, w54701, w54702, w54703, w54704, w54705, w54706, w54707, w54708, w54709, w54710, w54711, w54712, w54713, w54714, w54715, w54716, w54717, w54718, w54719, w54720, w54721, w54722, w54723, w54724, w54725, w54726, w54727, w54728, w54729, w54730, w54731, w54732, w54733, w54734, w54735, w54736, w54737, w54738, w54739, w54740, w54741, w54742, w54743, w54744, w54745, w54746, w54747, w54748, w54749, w54750, w54751, w54752, w54753, w54754, w54755, w54756, w54757, w54758, w54759, w54760, w54761, w54762, w54763, w54764, w54765, w54766, w54767, w54768, w54769, w54770, w54771, w54772, w54773, w54774, w54775, w54776, w54777, w54778, w54779, w54780, w54781, w54782, w54783, w54784, w54785, w54786, w54787, w54788, w54789, w54790, w54791, w54792, w54793, w54794, w54795, w54796, w54797, w54798, w54799, w54800, w54801, w54802, w54803, w54804, w54805, w54806, w54807, w54808, w54809, w54810, w54811, w54812, w54813, w54814, w54815, w54816, w54817, w54818, w54819, w54820, w54821, w54822, w54823, w54824, w54825, w54826, w54827, w54828, w54829, w54830, w54831, w54832, w54833, w54834, w54835, w54836, w54837, w54838, w54839, w54840, w54841, w54842, w54843, w54844, w54845, w54846, w54847, w54848, w54849, w54850, w54851, w54852, w54853, w54854, w54855, w54856, w54857, w54858, w54859, w54860, w54861, w54862, w54863, w54864, w54865, w54866, w54867, w54868, w54869, w54870, w54871, w54872, w54873, w54874, w54875, w54876, w54877, w54878, w54879, w54880, w54881, w54882, w54883, w54884, w54885, w54886, w54887, w54888, w54889, w54890, w54891, w54892, w54893, w54894, w54895, w54896, w54897, w54898, w54899, w54900, w54901, w54902, w54903, w54904, w54905, w54906, w54907, w54908, w54909, w54910, w54911, w54912, w54913, w54914, w54915, w54916, w54917, w54918, w54919, w54920, w54921, w54922, w54923, w54924, w54925, w54926, w54927, w54928, w54929, w54930, w54931, w54932, w54933, w54934, w54935, w54936, w54937, w54938, w54939, w54940, w54941, w54942, w54943, w54944, w54945, w54946, w54947, w54948, w54949, w54950, w54951, w54952, w54953, w54954, w54955, w54956, w54957, w54958, w54959, w54960, w54961, w54962, w54963, w54964, w54965, w54966, w54967, w54968, w54969, w54970, w54971, w54972, w54973, w54974, w54975, w54976, w54977, w54978, w54979, w54980, w54981, w54982, w54983, w54984, w54985, w54986, w54987, w54988, w54989, w54990, w54991, w54992, w54993, w54994, w54995, w54996, w54997, w54998, w54999, w55000, w55001, w55002, w55003, w55004, w55005, w55006, w55007, w55008, w55009, w55010, w55011, w55012, w55013, w55014, w55015, w55016, w55017, w55018, w55019, w55020, w55021, w55022, w55023, w55024, w55025, w55026, w55027, w55028, w55029, w55030, w55031, w55032, w55033, w55034, w55035, w55036, w55037, w55038, w55039, w55040, w55041, w55042, w55043, w55044, w55045, w55046, w55047, w55048, w55049, w55050, w55051, w55052, w55053, w55054, w55055, w55056, w55057, w55058, w55059, w55060, w55061, w55062, w55063, w55064, w55065, w55066, w55067, w55068, w55069, w55070, w55071, w55072, w55073, w55074, w55075, w55076, w55077, w55078, w55079, w55080, w55081, w55082, w55083, w55084, w55085, w55086, w55087, w55088, w55089, w55090, w55091, w55092, w55093, w55094, w55095, w55096, w55097, w55098, w55099, w55100, w55101, w55102, w55103, w55104, w55105, w55106, w55107, w55108, w55109, w55110, w55111, w55112, w55113, w55114, w55115, w55116, w55117, w55118, w55119, w55120, w55121, w55122, w55123, w55124, w55125, w55126, w55127, w55128, w55129, w55130, w55131, w55132, w55133, w55134, w55135, w55136, w55137, w55138, w55139, w55140, w55141, w55142, w55143, w55144, w55145, w55146, w55147, w55148, w55149, w55150, w55151, w55152, w55153, w55154, w55155, w55156, w55157, w55158, w55159, w55160, w55161, w55162, w55163, w55164, w55165, w55166, w55167, w55168, w55169, w55170, w55171, w55172, w55173, w55174, w55175, w55176, w55177, w55178, w55179, w55180, w55181, w55182, w55183, w55184, w55185, w55186, w55187, w55188, w55189, w55190, w55191, w55192, w55193, w55194, w55195, w55196, w55197, w55198, w55199, w55200, w55201, w55202, w55203, w55204, w55205, w55206, w55207, w55208, w55209, w55210, w55211, w55212, w55213, w55214, w55215, w55216, w55217, w55218, w55219, w55220, w55221, w55222, w55223, w55224, w55225, w55226, w55227, w55228, w55229, w55230, w55231, w55232, w55233, w55234, w55235, w55236, w55237, w55238, w55239, w55240, w55241, w55242, w55243, w55244, w55245, w55246, w55247, w55248, w55249, w55250, w55251, w55252, w55253, w55254, w55255, w55256, w55257, w55258, w55259, w55260, w55261, w55262, w55263, w55264, w55265, w55266, w55267, w55268, w55269, w55270, w55271, w55272, w55273, w55274, w55275, w55276, w55277, w55278, w55279, w55280, w55281, w55282, w55283, w55284, w55285, w55286, w55287, w55288, w55289, w55290, w55291, w55292, w55293, w55294, w55295, w55296, w55297, w55298, w55299, w55300, w55301, w55302, w55303, w55304, w55305, w55306, w55307, w55308, w55309, w55310, w55311, w55312, w55313, w55314, w55315, w55316, w55317, w55318, w55319, w55320, w55321, w55322, w55323, w55324, w55325, w55326, w55327, w55328, w55329, w55330, w55331, w55332, w55333, w55334, w55335, w55336, w55337, w55338, w55339, w55340, w55341, w55342, w55343, w55344, w55345, w55346, w55347, w55348, w55349, w55350, w55351, w55352, w55353, w55354, w55355, w55356, w55357, w55358, w55359, w55360, w55361, w55362, w55363, w55364, w55365, w55366, w55367, w55368, w55369, w55370, w55371, w55372, w55373, w55374, w55375, w55376, w55377, w55378, w55379, w55380, w55381, w55382, w55383, w55384, w55385, w55386, w55387, w55388, w55389, w55390, w55391, w55392, w55393, w55394, w55395, w55396, w55397, w55398, w55399, w55400, w55401, w55402, w55403, w55404, w55405, w55406, w55407, w55408, w55409, w55410, w55411, w55412, w55413, w55414, w55415, w55416, w55417, w55418, w55419, w55420, w55421, w55422, w55423, w55424, w55425, w55426, w55427, w55428, w55429, w55430, w55431, w55432, w55433, w55434, w55435, w55436, w55437, w55438, w55439, w55440, w55441, w55442, w55443, w55444, w55445, w55446, w55447, w55448, w55449, w55450, w55451, w55452, w55453, w55454, w55455, w55456, w55457, w55458, w55459, w55460, w55461, w55462, w55463, w55464, w55465, w55466, w55467, w55468, w55469, w55470, w55471, w55472, w55473, w55474, w55475, w55476, w55477, w55478, w55479, w55480, w55481, w55482, w55483, w55484, w55485, w55486, w55487, w55488, w55489, w55490, w55491, w55492, w55493, w55494, w55495, w55496, w55497, w55498, w55499, w55500, w55501, w55502, w55503, w55504, w55505, w55506, w55507, w55508, w55509, w55510, w55511, w55512, w55513, w55514, w55515, w55516, w55517, w55518, w55519, w55520, w55521, w55522, w55523, w55524, w55525, w55526, w55527, w55528, w55529, w55530, w55531, w55532, w55533, w55534, w55535, w55536, w55537, w55538, w55539, w55540, w55541, w55542, w55543, w55544, w55545, w55546, w55547, w55548, w55549, w55550, w55551, w55552, w55553, w55554, w55555, w55556, w55557, w55558, w55559, w55560, w55561, w55562, w55563, w55564, w55565, w55566, w55567, w55568, w55569, w55570, w55571, w55572, w55573, w55574, w55575, w55576, w55577, w55578, w55579, w55580, w55581, w55582, w55583, w55584, w55585, w55586, w55587, w55588, w55589, w55590, w55591, w55592, w55593, w55594, w55595, w55596, w55597, w55598, w55599, w55600, w55601, w55602, w55603, w55604, w55605, w55606, w55607, w55608, w55609, w55610, w55611, w55612, w55613, w55614, w55615, w55616, w55617, w55618, w55619, w55620, w55621, w55622, w55623, w55624, w55625, w55626, w55627, w55628, w55629, w55630, w55631, w55632, w55633, w55634, w55635, w55636, w55637, w55638, w55639, w55640, w55641, w55642, w55643, w55644, w55645, w55646, w55647, w55648, w55649, w55650, w55651, w55652, w55653, w55654, w55655, w55656, w55657, w55658, w55659, w55660, w55661, w55662, w55663, w55664, w55665, w55666, w55667, w55668, w55669, w55670, w55671, w55672, w55673, w55674, w55675, w55676, w55677, w55678, w55679, w55680, w55681, w55682, w55683, w55684, w55685, w55686, w55687, w55688, w55689, w55690, w55691, w55692, w55693, w55694, w55695, w55696, w55697, w55698, w55699, w55700, w55701, w55702, w55703, w55704, w55705, w55706, w55707, w55708, w55709, w55710, w55711, w55712, w55713, w55714, w55715, w55716, w55717, w55718, w55719, w55720, w55721, w55722, w55723, w55724, w55725, w55726, w55727, w55728, w55729, w55730, w55731, w55732, w55733, w55734, w55735, w55736, w55737, w55738, w55739, w55740, w55741, w55742, w55743, w55744, w55745, w55746, w55747, w55748, w55749, w55750, w55751, w55752, w55753, w55754, w55755, w55756, w55757, w55758, w55759, w55760, w55761, w55762, w55763, w55764, w55765, w55766, w55767, w55768, w55769, w55770, w55771, w55772, w55773, w55774, w55775, w55776, w55777, w55778, w55779, w55780, w55781, w55782, w55783, w55784, w55785, w55786, w55787, w55788, w55789, w55790, w55791, w55792, w55793, w55794, w55795, w55796, w55797, w55798, w55799, w55800, w55801, w55802, w55803, w55804, w55805, w55806, w55807, w55808, w55809, w55810, w55811, w55812, w55813, w55814, w55815, w55816, w55817, w55818, w55819, w55820, w55821, w55822, w55823, w55824, w55825, w55826, w55827, w55828, w55829, w55830, w55831, w55832, w55833, w55834, w55835, w55836, w55837, w55838, w55839, w55840, w55841, w55842, w55843, w55844, w55845, w55846, w55847, w55848, w55849, w55850, w55851, w55852, w55853, w55854, w55855, w55856, w55857, w55858, w55859, w55860, w55861, w55862, w55863, w55864, w55865, w55866, w55867, w55868, w55869, w55870, w55871, w55872, w55873, w55874, w55875, w55876, w55877, w55878, w55879, w55880, w55881, w55882, w55883, w55884, w55885, w55886, w55887, w55888, w55889, w55890, w55891, w55892, w55893, w55894, w55895, w55896, w55897, w55898, w55899, w55900, w55901, w55902, w55903, w55904, w55905, w55906, w55907, w55908, w55909, w55910, w55911, w55912, w55913, w55914, w55915, w55916, w55917, w55918, w55919, w55920, w55921, w55922, w55923, w55924, w55925, w55926, w55927, w55928, w55929, w55930, w55931, w55932, w55933, w55934, w55935, w55936, w55937, w55938, w55939, w55940, w55941, w55942, w55943, w55944, w55945, w55946, w55947, w55948, w55949, w55950, w55951, w55952, w55953, w55954, w55955, w55956, w55957, w55958, w55959, w55960, w55961, w55962, w55963, w55964, w55965, w55966, w55967, w55968, w55969, w55970, w55971, w55972, w55973, w55974, w55975, w55976, w55977, w55978, w55979, w55980, w55981, w55982, w55983, w55984, w55985, w55986, w55987, w55988, w55989, w55990, w55991, w55992, w55993, w55994, w55995, w55996, w55997, w55998, w55999, w56000, w56001, w56002, w56003, w56004, w56005, w56006, w56007, w56008, w56009, w56010, w56011, w56012, w56013, w56014, w56015, w56016, w56017, w56018, w56019, w56020, w56021, w56022, w56023, w56024, w56025, w56026, w56027, w56028, w56029, w56030, w56031, w56032, w56033, w56034, w56035, w56036, w56037, w56038, w56039, w56040, w56041, w56042, w56043, w56044, w56045, w56046, w56047, w56048, w56049, w56050, w56051, w56052, w56053, w56054, w56055, w56056, w56057, w56058, w56059, w56060, w56061, w56062, w56063, w56064, w56065, w56066, w56067, w56068, w56069, w56070, w56071, w56072, w56073, w56074, w56075, w56076, w56077, w56078, w56079, w56080, w56081, w56082, w56083, w56084, w56085, w56086, w56087, w56088, w56089, w56090, w56091, w56092, w56093, w56094, w56095, w56096, w56097, w56098, w56099, w56100, w56101, w56102, w56103, w56104, w56105, w56106, w56107, w56108, w56109, w56110, w56111, w56112, w56113, w56114, w56115, w56116, w56117, w56118, w56119, w56120, w56121, w56122, w56123, w56124, w56125, w56126, w56127, w56128, w56129, w56130, w56131, w56132, w56133, w56134, w56135, w56136, w56137, w56138, w56139, w56140, w56141, w56142, w56143, w56144, w56145, w56146, w56147, w56148, w56149, w56150, w56151, w56152, w56153, w56154, w56155, w56156, w56157, w56158, w56159, w56160, w56161, w56162, w56163, w56164, w56165, w56166, w56167, w56168, w56169, w56170, w56171, w56172, w56173, w56174, w56175, w56176, w56177, w56178, w56179, w56180, w56181, w56182, w56183, w56184, w56185, w56186, w56187, w56188, w56189, w56190, w56191, w56192, w56193, w56194, w56195, w56196, w56197, w56198, w56199, w56200, w56201, w56202, w56203, w56204, w56205, w56206, w56207, w56208, w56209, w56210, w56211, w56212, w56213, w56214, w56215, w56216, w56217, w56218, w56219, w56220, w56221, w56222, w56223, w56224, w56225, w56226, w56227, w56228, w56229, w56230, w56231, w56232, w56233, w56234, w56235, w56236, w56237, w56238, w56239, w56240, w56241, w56242, w56243, w56244, w56245, w56246, w56247, w56248, w56249, w56250, w56251, w56252, w56253, w56254, w56255, w56256, w56257, w56258, w56259, w56260, w56261, w56262, w56263, w56264, w56265, w56266, w56267, w56268, w56269, w56270, w56271, w56272, w56273, w56274, w56275, w56276, w56277, w56278, w56279, w56280, w56281, w56282, w56283, w56284, w56285, w56286, w56287, w56288, w56289, w56290, w56291, w56292, w56293, w56294, w56295, w56296, w56297, w56298, w56299, w56300, w56301, w56302, w56303, w56304, w56305, w56306, w56307, w56308, w56309, w56310, w56311, w56312, w56313, w56314, w56315, w56316, w56317, w56318, w56319, w56320, w56321, w56322, w56323, w56324, w56325, w56326, w56327, w56328, w56329, w56330, w56331, w56332, w56333, w56334, w56335, w56336, w56337, w56338, w56339, w56340, w56341, w56342, w56343, w56344, w56345, w56346, w56347, w56348, w56349, w56350, w56351, w56352, w56353, w56354, w56355, w56356, w56357, w56358, w56359, w56360, w56361, w56362, w56363, w56364, w56365, w56366, w56367, w56368, w56369, w56370, w56371, w56372, w56373, w56374, w56375, w56376, w56377, w56378, w56379, w56380, w56381, w56382, w56383, w56384, w56385, w56386, w56387, w56388, w56389, w56390, w56391, w56392, w56393, w56394, w56395, w56396, w56397, w56398, w56399, w56400, w56401, w56402, w56403, w56404, w56405, w56406, w56407, w56408, w56409, w56410, w56411, w56412, w56413, w56414, w56415, w56416, w56417, w56418, w56419, w56420, w56421, w56422, w56423, w56424, w56425, w56426, w56427, w56428, w56429, w56430, w56431, w56432, w56433, w56434, w56435, w56436, w56437, w56438, w56439, w56440, w56441, w56442, w56443, w56444, w56445, w56446, w56447, w56448, w56449, w56450, w56451, w56452, w56453, w56454, w56455, w56456, w56457, w56458, w56459, w56460, w56461, w56462, w56463, w56464, w56465, w56466, w56467, w56468, w56469, w56470, w56471, w56472, w56473, w56474, w56475, w56476, w56477, w56478, w56479, w56480, w56481, w56482, w56483, w56484, w56485, w56486, w56487, w56488, w56489, w56490, w56491, w56492, w56493, w56494, w56495, w56496, w56497, w56498, w56499, w56500, w56501, w56502, w56503, w56504, w56505, w56506, w56507, w56508, w56509, w56510, w56511, w56512, w56513, w56514, w56515, w56516, w56517, w56518, w56519, w56520, w56521, w56522, w56523, w56524, w56525, w56526, w56527, w56528, w56529, w56530, w56531, w56532, w56533, w56534, w56535, w56536, w56537, w56538, w56539, w56540, w56541, w56542, w56543, w56544, w56545, w56546, w56547, w56548, w56549, w56550, w56551, w56552, w56553, w56554, w56555, w56556, w56557, w56558, w56559, w56560, w56561, w56562, w56563, w56564, w56565, w56566, w56567, w56568, w56569, w56570, w56571, w56572, w56573, w56574, w56575, w56576, w56577, w56578, w56579, w56580, w56581, w56582, w56583, w56584, w56585, w56586, w56587, w56588, w56589, w56590, w56591, w56592, w56593, w56594, w56595, w56596, w56597, w56598, w56599, w56600, w56601, w56602, w56603, w56604, w56605, w56606, w56607, w56608, w56609, w56610, w56611, w56612, w56613, w56614, w56615, w56616, w56617, w56618, w56619, w56620, w56621, w56622, w56623, w56624, w56625, w56626, w56627, w56628, w56629, w56630, w56631, w56632, w56633, w56634, w56635, w56636, w56637, w56638, w56639, w56640, w56641, w56642, w56643, w56644, w56645, w56646, w56647, w56648, w56649, w56650, w56651, w56652, w56653, w56654, w56655, w56656, w56657, w56658, w56659, w56660, w56661, w56662, w56663, w56664, w56665, w56666, w56667, w56668, w56669, w56670, w56671, w56672, w56673, w56674, w56675, w56676, w56677, w56678, w56679, w56680, w56681, w56682, w56683, w56684, w56685, w56686, w56687, w56688, w56689, w56690, w56691, w56692, w56693, w56694, w56695, w56696, w56697, w56698, w56699, w56700, w56701, w56702, w56703, w56704, w56705, w56706, w56707, w56708, w56709, w56710, w56711, w56712, w56713, w56714, w56715, w56716, w56717, w56718, w56719, w56720, w56721, w56722, w56723, w56724, w56725, w56726, w56727, w56728, w56729, w56730, w56731, w56732, w56733, w56734, w56735, w56736, w56737, w56738, w56739, w56740, w56741, w56742, w56743, w56744, w56745, w56746, w56747, w56748, w56749, w56750, w56751, w56752, w56753, w56754, w56755, w56756, w56757, w56758, w56759, w56760, w56761, w56762, w56763, w56764, w56765, w56766, w56767, w56768, w56769, w56770, w56771, w56772, w56773, w56774, w56775, w56776, w56777, w56778, w56779, w56780, w56781, w56782, w56783, w56784, w56785, w56786, w56787, w56788, w56789, w56790, w56791, w56792, w56793, w56794, w56795, w56796, w56797, w56798, w56799, w56800, w56801, w56802, w56803, w56804, w56805, w56806, w56807, w56808, w56809, w56810, w56811, w56812, w56813, w56814, w56815, w56816, w56817, w56818, w56819, w56820, w56821, w56822, w56823, w56824, w56825, w56826, w56827, w56828, w56829, w56830, w56831, w56832, w56833, w56834, w56835, w56836, w56837, w56838, w56839, w56840, w56841, w56842, w56843, w56844, w56845, w56846, w56847, w56848, w56849, w56850, w56851, w56852, w56853, w56854, w56855, w56856, w56857, w56858, w56859, w56860, w56861, w56862, w56863, w56864, w56865, w56866, w56867, w56868, w56869, w56870, w56871, w56872, w56873, w56874, w56875, w56876, w56877, w56878, w56879, w56880, w56881, w56882, w56883, w56884, w56885, w56886, w56887, w56888, w56889, w56890, w56891, w56892, w56893, w56894, w56895, w56896, w56897, w56898, w56899, w56900, w56901, w56902, w56903, w56904, w56905, w56906, w56907, w56908, w56909, w56910, w56911, w56912, w56913, w56914, w56915, w56916, w56917, w56918, w56919, w56920, w56921, w56922, w56923, w56924, w56925, w56926, w56927, w56928, w56929, w56930, w56931, w56932, w56933, w56934, w56935, w56936, w56937, w56938, w56939, w56940, w56941, w56942, w56943, w56944, w56945, w56946, w56947, w56948, w56949, w56950, w56951, w56952, w56953, w56954, w56955, w56956, w56957, w56958, w56959, w56960, w56961, w56962, w56963, w56964, w56965, w56966, w56967, w56968, w56969, w56970, w56971, w56972, w56973, w56974, w56975, w56976, w56977, w56978, w56979, w56980, w56981, w56982, w56983, w56984, w56985, w56986, w56987, w56988, w56989, w56990, w56991, w56992, w56993, w56994, w56995, w56996, w56997, w56998, w56999, w57000, w57001, w57002, w57003, w57004, w57005, w57006, w57007, w57008, w57009, w57010, w57011, w57012, w57013, w57014, w57015, w57016, w57017, w57018, w57019, w57020, w57021, w57022, w57023, w57024, w57025, w57026, w57027, w57028, w57029, w57030, w57031, w57032, w57033, w57034, w57035, w57036, w57037, w57038, w57039, w57040, w57041, w57042, w57043, w57044, w57045, w57046, w57047, w57048, w57049, w57050, w57051, w57052, w57053, w57054, w57055, w57056, w57057, w57058, w57059, w57060, w57061, w57062, w57063, w57064, w57065, w57066, w57067, w57068, w57069, w57070, w57071, w57072, w57073, w57074, w57075, w57076, w57077, w57078, w57079, w57080, w57081, w57082, w57083, w57084, w57085, w57086, w57087, w57088, w57089, w57090, w57091, w57092, w57093, w57094, w57095, w57096, w57097, w57098, w57099, w57100, w57101, w57102, w57103, w57104, w57105, w57106, w57107, w57108, w57109, w57110, w57111, w57112, w57113, w57114, w57115, w57116, w57117, w57118, w57119, w57120, w57121, w57122, w57123, w57124, w57125, w57126, w57127, w57128, w57129, w57130, w57131, w57132, w57133, w57134, w57135, w57136, w57137, w57138, w57139, w57140, w57141, w57142, w57143, w57144, w57145, w57146, w57147, w57148, w57149, w57150, w57151, w57152, w57153, w57154, w57155, w57156, w57157, w57158, w57159, w57160, w57161, w57162, w57163, w57164, w57165, w57166, w57167, w57168, w57169, w57170, w57171, w57172, w57173, w57174, w57175, w57176, w57177, w57178, w57179, w57180, w57181, w57182, w57183, w57184, w57185, w57186, w57187, w57188, w57189, w57190, w57191, w57192, w57193, w57194, w57195, w57196, w57197, w57198, w57199, w57200, w57201, w57202, w57203, w57204, w57205, w57206, w57207, w57208, w57209, w57210, w57211, w57212, w57213, w57214, w57215, w57216, w57217, w57218, w57219, w57220, w57221, w57222, w57223, w57224, w57225, w57226, w57227, w57228, w57229, w57230, w57231, w57232, w57233, w57234, w57235, w57236, w57237, w57238, w57239, w57240, w57241, w57242, w57243, w57244, w57245, w57246, w57247, w57248, w57249, w57250, w57251, w57252, w57253, w57254, w57255, w57256, w57257, w57258, w57259, w57260, w57261, w57262, w57263, w57264, w57265, w57266, w57267, w57268, w57269, w57270, w57271, w57272, w57273, w57274, w57275, w57276, w57277, w57278, w57279, w57280, w57281, w57282, w57283, w57284, w57285, w57286, w57287, w57288, w57289, w57290, w57291, w57292, w57293, w57294, w57295, w57296, w57297, w57298, w57299, w57300, w57301, w57302, w57303, w57304, w57305, w57306, w57307, w57308, w57309, w57310, w57311, w57312, w57313, w57314, w57315, w57316, w57317, w57318, w57319, w57320, w57321, w57322, w57323, w57324, w57325, w57326, w57327, w57328, w57329, w57330, w57331, w57332, w57333, w57334, w57335, w57336, w57337, w57338, w57339, w57340, w57341, w57342, w57343, w57344, w57345, w57346, w57347, w57348, w57349, w57350, w57351, w57352, w57353, w57354, w57355, w57356, w57357, w57358, w57359, w57360, w57361, w57362, w57363, w57364, w57365, w57366, w57367, w57368, w57369, w57370, w57371, w57372, w57373, w57374, w57375, w57376, w57377, w57378, w57379, w57380, w57381, w57382, w57383, w57384, w57385, w57386, w57387, w57388, w57389, w57390, w57391, w57392, w57393, w57394, w57395, w57396, w57397, w57398, w57399, w57400, w57401, w57402, w57403, w57404, w57405, w57406, w57407, w57408, w57409, w57410, w57411, w57412, w57413, w57414, w57415, w57416, w57417, w57418, w57419, w57420, w57421, w57422, w57423, w57424, w57425, w57426, w57427, w57428, w57429, w57430, w57431, w57432, w57433, w57434, w57435, w57436, w57437, w57438, w57439, w57440, w57441, w57442, w57443, w57444, w57445, w57446, w57447, w57448, w57449, w57450, w57451, w57452, w57453, w57454, w57455, w57456, w57457, w57458, w57459, w57460, w57461, w57462, w57463, w57464, w57465, w57466, w57467, w57468, w57469, w57470, w57471, w57472, w57473, w57474, w57475, w57476, w57477, w57478, w57479, w57480, w57481, w57482, w57483, w57484, w57485, w57486, w57487, w57488, w57489, w57490, w57491, w57492, w57493, w57494, w57495, w57496, w57497, w57498, w57499, w57500, w57501, w57502, w57503, w57504, w57505, w57506, w57507, w57508, w57509, w57510, w57511, w57512, w57513, w57514, w57515, w57516, w57517, w57518, w57519, w57520, w57521, w57522, w57523, w57524, w57525, w57526, w57527, w57528, w57529, w57530, w57531, w57532, w57533, w57534, w57535, w57536, w57537, w57538, w57539, w57540, w57541, w57542, w57543, w57544, w57545, w57546, w57547, w57548, w57549, w57550, w57551, w57552, w57553, w57554, w57555, w57556, w57557, w57558, w57559, w57560, w57561, w57562, w57563, w57564, w57565, w57566, w57567, w57568, w57569, w57570, w57571, w57572, w57573, w57574, w57575, w57576, w57577, w57578, w57579, w57580, w57581, w57582, w57583, w57584, w57585, w57586, w57587, w57588, w57589, w57590, w57591, w57592, w57593, w57594, w57595, w57596, w57597, w57598, w57599, w57600, w57601, w57602, w57603, w57604, w57605, w57606, w57607, w57608, w57609, w57610, w57611, w57612, w57613, w57614, w57615, w57616, w57617, w57618, w57619, w57620, w57621, w57622, w57623, w57624, w57625, w57626, w57627, w57628, w57629, w57630, w57631, w57632, w57633, w57634, w57635, w57636, w57637, w57638, w57639, w57640, w57641, w57642, w57643, w57644, w57645, w57646, w57647, w57648, w57649, w57650, w57651, w57652, w57653, w57654, w57655, w57656, w57657, w57658, w57659, w57660, w57661, w57662, w57663, w57664, w57665, w57666, w57667, w57668, w57669, w57670, w57671, w57672, w57673, w57674, w57675, w57676, w57677, w57678, w57679, w57680, w57681, w57682, w57683, w57684, w57685, w57686, w57687, w57688, w57689, w57690, w57691, w57692, w57693, w57694, w57695, w57696, w57697, w57698, w57699, w57700, w57701, w57702, w57703, w57704, w57705, w57706, w57707, w57708, w57709, w57710, w57711, w57712, w57713, w57714, w57715, w57716, w57717, w57718, w57719, w57720, w57721, w57722, w57723, w57724, w57725, w57726, w57727, w57728, w57729, w57730, w57731, w57732, w57733, w57734, w57735, w57736, w57737, w57738, w57739, w57740, w57741, w57742, w57743, w57744, w57745, w57746, w57747, w57748, w57749, w57750, w57751, w57752, w57753, w57754, w57755, w57756, w57757, w57758, w57759, w57760, w57761, w57762, w57763, w57764, w57765, w57766, w57767, w57768, w57769, w57770, w57771, w57772, w57773, w57774, w57775, w57776, w57777, w57778, w57779, w57780, w57781, w57782, w57783, w57784, w57785, w57786, w57787, w57788, w57789, w57790, w57791, w57792, w57793, w57794, w57795, w57796, w57797, w57798, w57799, w57800, w57801, w57802, w57803, w57804, w57805, w57806, w57807, w57808, w57809, w57810, w57811, w57812, w57813, w57814, w57815, w57816, w57817, w57818, w57819, w57820, w57821, w57822, w57823, w57824, w57825, w57826, w57827, w57828, w57829, w57830, w57831, w57832, w57833, w57834, w57835, w57836, w57837, w57838, w57839, w57840, w57841, w57842, w57843, w57844, w57845, w57846, w57847, w57848, w57849, w57850, w57851, w57852, w57853, w57854, w57855, w57856, w57857, w57858, w57859, w57860, w57861, w57862, w57863, w57864, w57865, w57866, w57867, w57868, w57869, w57870, w57871, w57872, w57873, w57874, w57875, w57876, w57877, w57878, w57879, w57880, w57881, w57882, w57883, w57884, w57885, w57886, w57887, w57888, w57889, w57890, w57891, w57892, w57893, w57894, w57895, w57896, w57897, w57898, w57899, w57900, w57901, w57902, w57903, w57904, w57905, w57906, w57907, w57908, w57909, w57910, w57911, w57912, w57913, w57914, w57915, w57916, w57917, w57918, w57919, w57920, w57921, w57922, w57923, w57924, w57925, w57926, w57927, w57928, w57929, w57930, w57931, w57932, w57933, w57934, w57935, w57936, w57937, w57938, w57939, w57940, w57941, w57942, w57943, w57944, w57945, w57946, w57947, w57948, w57949, w57950, w57951, w57952, w57953, w57954, w57955, w57956, w57957, w57958;
assign w0 = ~pi00965 & pi01260;
assign w1 = pi00855 & pi01258;
assign w2 = ~pi00966 & pi01254;
assign w3 = pi00853 & pi01259;
assign w4 = ~pi00964 & pi01255;
assign w5 = pi00856 & pi01257;
assign w6 = pi00854 & pi01256;
assign w7 = ~w0 & ~w1;
assign w8 = ~w2 & ~w3;
assign w9 = ~w4 & ~w5;
assign w10 = ~w6 & w9;
assign w11 = w7 & w8;
assign w12 = w10 & w11;
assign w13 = ~pi00000 & ~pi00250;
assign w14 = ~pi00234 & ~pi00235;
assign w15 = ~pi00236 & ~pi00237;
assign w16 = ~pi00238 & ~pi00239;
assign w17 = ~pi00242 & ~pi00243;
assign w18 = ~pi00244 & ~pi00245;
assign w19 = ~pi00246 & ~pi00247;
assign w20 = ~pi00248 & w19;
assign w21 = w17 & w18;
assign w22 = w15 & w16;
assign w23 = w14 & w22;
assign w24 = w20 & w21;
assign w25 = w23 & w24;
assign w26 = ~pi00233 & ~pi00240;
assign w27 = w25 & w54865;
assign w28 = pi00002 & pi00003;
assign w29 = ~pi00004 & pi00023;
assign w30 = pi00026 & pi00027;
assign w31 = pi00041 & pi00051;
assign w32 = pi00054 & pi00058;
assign w33 = pi00060 & pi00061;
assign w34 = pi00064 & pi00069;
assign w35 = pi00070 & pi00073;
assign w36 = pi00141 & pi00186;
assign w37 = pi00187 & ~pi00205;
assign w38 = pi00231 & pi00343;
assign w39 = pi00360 & pi00361;
assign w40 = pi00366 & pi00373;
assign w41 = pi00465 & pi00472;
assign w42 = pi00610 & pi00879;
assign w43 = pi01166 & pi01167;
assign w44 = w42 & w43;
assign w45 = w40 & w41;
assign w46 = w38 & w39;
assign w47 = w36 & w37;
assign w48 = w34 & w35;
assign w49 = w32 & w33;
assign w50 = w30 & w31;
assign w51 = w28 & w29;
assign w52 = w50 & w51;
assign w53 = w48 & w49;
assign w54 = w46 & w47;
assign w55 = w44 & w45;
assign w56 = w54 & w55;
assign w57 = w52 & w53;
assign w58 = w56 & w57;
assign w59 = ~w27 & ~w58;
assign w60 = pi00250 & ~w59;
assign w61 = ~pi00188 & ~w13;
assign w62 = ~w60 & w61;
assign w63 = ~pi00274 & ~pi10577;
assign w64 = ~pi00233 & pi00240;
assign w65 = pi00250 & w64;
assign w66 = w25 & w54866;
assign w67 = (w63 & ~w25) | (w63 & w54867) | (~w25 & w54867);
assign w68 = pi00001 & w67;
assign w69 = w25 & w54868;
assign w70 = ~pi00003 & w69;
assign w71 = ~w68 & ~w70;
assign w72 = ~pi09912 & ~pi09926;
assign w73 = (pi09819 & ~w72) | (pi09819 & w43508) | (~w72 & w43508);
assign w74 = w72 & w54745;
assign w75 = pi09969 & ~w74;
assign w76 = (~pi00188 & ~w75) | (~pi00188 & w54869) | (~w75 & w54869);
assign w77 = pi00003 & w76;
assign w78 = ~pi00249 & ~pi00250;
assign w79 = pi00241 & ~pi09800;
assign w80 = ~pi00246 & pi09888;
assign w81 = ~pi00243 & pi09882;
assign w82 = ~pi00244 & pi09883;
assign w83 = pi00239 & ~pi09980;
assign w84 = pi00242 & ~pi09881;
assign w85 = pi00244 & ~pi09883;
assign w86 = pi00233 & ~pi09877;
assign w87 = pi00240 & ~pi09879;
assign w88 = ~w86 & ~w87;
assign w89 = pi00247 & ~pi09948;
assign w90 = ~pi00247 & pi09948;
assign w91 = ~pi00242 & pi09881;
assign w92 = pi00246 & ~pi09888;
assign w93 = pi00243 & ~pi09882;
assign w94 = ~pi00248 & pi09971;
assign w95 = pi00248 & ~pi09971;
assign w96 = pi00238 & ~pi09979;
assign w97 = ~pi00234 & pi09972;
assign w98 = ~pi00241 & pi09800;
assign w99 = pi00235 & ~pi09974;
assign w100 = ~pi00237 & pi09944;
assign w101 = pi00234 & ~pi09972;
assign w102 = pi00237 & ~pi09944;
assign w103 = pi00236 & ~pi09978;
assign w104 = ~pi00235 & pi09974;
assign w105 = pi00245 & ~pi09799;
assign w106 = ~pi00238 & pi09979;
assign w107 = ~pi00236 & pi09978;
assign w108 = ~pi00233 & pi09877;
assign w109 = ~pi00239 & pi09980;
assign w110 = ~pi00245 & pi09799;
assign w111 = ~pi00240 & pi09879;
assign w112 = ~pi09949 & ~w79;
assign w113 = ~w80 & ~w81;
assign w114 = ~w82 & ~w83;
assign w115 = ~w84 & ~w85;
assign w116 = ~w89 & ~w90;
assign w117 = ~w91 & ~w92;
assign w118 = ~w93 & ~w94;
assign w119 = ~w95 & ~w96;
assign w120 = ~w97 & ~w98;
assign w121 = ~w99 & ~w100;
assign w122 = ~w101 & ~w102;
assign w123 = ~w103 & ~w104;
assign w124 = ~w105 & ~w106;
assign w125 = ~w107 & ~w108;
assign w126 = ~w109 & ~w110;
assign w127 = ~w111 & w126;
assign w128 = w124 & w125;
assign w129 = w122 & w123;
assign w130 = w120 & w121;
assign w131 = w118 & w119;
assign w132 = w116 & w117;
assign w133 = w114 & w115;
assign w134 = w112 & w113;
assign w135 = w88 & w134;
assign w136 = w132 & w133;
assign w137 = w130 & w131;
assign w138 = w128 & w129;
assign w139 = w127 & w138;
assign w140 = w136 & w137;
assign w141 = w135 & w140;
assign w142 = pi10444 & pi10585;
assign w143 = ~pi09872 & ~w142;
assign w144 = pi09872 & ~pi10447;
assign w145 = ~w143 & ~w144;
assign w146 = (w145 & ~w141) | (w145 & w54870) | (~w141 & w54870);
assign w147 = pi09872 & pi10370;
assign w148 = ~pi09872 & pi10670;
assign w149 = ~w147 & ~w148;
assign w150 = pi00205 & ~w149;
assign w151 = ~pi00205 & w149;
assign w152 = ~w150 & ~w151;
assign w153 = w146 & w54873;
assign w154 = (w146 & w54874) | (w146 & w54875) | (w54874 & w54875);
assign w155 = ~w153 & w154;
assign w156 = pi09872 & pi10372;
assign w157 = ~pi09872 & pi10669;
assign w158 = ~w156 & ~w157;
assign w159 = pi00026 & ~w158;
assign w160 = ~pi00026 & w158;
assign w161 = ~w159 & ~w160;
assign w162 = w146 & w54878;
assign w163 = (w146 & w54879) | (w146 & w54880) | (w54879 & w54880);
assign w164 = ~w162 & w163;
assign w165 = pi00005 & w67;
assign w166 = pi00041 & w69;
assign w167 = ~w165 & ~w166;
assign w168 = ~pi10235 & ~pi10237;
assign w169 = ~pi10026 & ~pi10027;
assign w170 = pi10234 & ~w169;
assign w171 = w168 & ~w170;
assign w172 = ~w170 & w54695;
assign w173 = ~pi10025 & w172;
assign w174 = w172 & w54700;
assign w175 = (~pi10235 & w169) | (~pi10235 & w54701) | (w169 & w54701);
assign w176 = pi10237 & ~w175;
assign w177 = (~pi00018 & w174) | (~pi00018 & w54721) | (w174 & w54721);
assign w178 = ~w169 & w54702;
assign w179 = ~w175 & ~w178;
assign w180 = (pi00017 & ~w172) | (pi00017 & w54722) | (~w172 & w54722);
assign w181 = ~w179 & ~w180;
assign w182 = ~pi10234 & w169;
assign w183 = ~w170 & ~w182;
assign w184 = pi10026 & pi10027;
assign w185 = ~w169 & ~w184;
assign w186 = pi00015 & w185;
assign w187 = ~pi00015 & ~w185;
assign w188 = pi00006 & pi00014;
assign w189 = ~pi00006 & ~pi00014;
assign w190 = pi10027 & ~w189;
assign w191 = ~w188 & ~w190;
assign w192 = ~w187 & ~w191;
assign w193 = (~w183 & w192) | (~w183 & w54723) | (w192 & w54723);
assign w194 = (pi00016 & w192) | (pi00016 & w54746) | (w192 & w54746);
assign w195 = ~w193 & ~w194;
assign w196 = ~w177 & ~w181;
assign w197 = ~w195 & w196;
assign w198 = pi00017 & pi00018;
assign w199 = w179 & w198;
assign w200 = (pi00020 & w172) | (pi00020 & w54724) | (w172 & w54724);
assign w201 = (pi10236 & w170) | (pi10236 & w54704) | (w170 & w54704);
assign w202 = ~w172 & ~w201;
assign w203 = pi00019 & w202;
assign w204 = (~w173 & w203) | (~w173 & w54725) | (w203 & w54725);
assign w205 = (~pi00018 & ~w179) | (~pi00018 & w54726) | (~w179 & w54726);
assign w206 = ~w171 & ~w176;
assign w207 = ~w205 & w206;
assign w208 = ~w199 & ~w207;
assign w209 = ~w204 & w208;
assign w210 = ~w197 & w209;
assign w211 = ~w172 & w54881;
assign w212 = ~w170 & w54882;
assign w213 = (~w212 & w202) | (~w212 & w54883) | (w202 & w54883);
assign w214 = ~w204 & ~w213;
assign w215 = w172 & w54727;
assign w216 = (pi10024 & ~w172) | (pi10024 & w54728) | (~w172 & w54728);
assign w217 = ~w215 & ~w216;
assign w218 = (~w211 & w217) | (~w211 & w54884) | (w217 & w54884);
assign w219 = ~w214 & w218;
assign w220 = pi00021 & w217;
assign w221 = (~w220 & w210) | (~w220 & w54729) | (w210 & w54729);
assign w222 = ~pi10023 & ~pi10024;
assign w223 = ~pi10025 & w222;
assign w224 = w172 & w223;
assign w225 = w172 & w54705;
assign w226 = (pi10239 & ~w172) | (pi10239 & w54747) | (~w172 & w54747);
assign w227 = ~w225 & ~w226;
assign w228 = ~pi00008 & ~w227;
assign w229 = w172 & w54730;
assign w230 = (pi10238 & ~w172) | (pi10238 & w54748) | (~w172 & w54748);
assign w231 = ~w229 & ~w230;
assign w232 = ~pi00009 & ~w231;
assign w233 = pi10021 & ~w229;
assign w234 = ~pi10021 & ~pi10234;
assign w235 = ~pi10236 & ~pi10238;
assign w236 = ~pi10239 & w235;
assign w237 = w168 & w234;
assign w238 = w236 & w237;
assign w239 = w223 & w238;
assign w240 = ~w233 & ~w239;
assign w241 = (~pi00010 & ~w240) | (~pi00010 & w54731) | (~w240 & w54731);
assign w242 = ~w232 & ~w241;
assign w243 = (pi10023 & ~w172) | (pi10023 & w54885) | (~w172 & w54885);
assign w244 = ~w224 & ~w243;
assign w245 = ~w228 & w244;
assign w246 = w242 & w245;
assign w247 = (pi00022 & w227) | (pi00022 & w54886) | (w227 & w54886);
assign w248 = ~w241 & w54887;
assign w249 = (~w54729 & w54888) | (~w54729 & w54889) | (w54888 & w54889);
assign w250 = pi00008 & w227;
assign w251 = ~w241 & w54890;
assign w252 = pi00009 & w231;
assign w253 = ~w233 & w54891;
assign w254 = ~w252 & ~w253;
assign w255 = w229 & w54749;
assign w256 = (w240 & w54892) | (w240 & w54893) | (w54892 & w54893);
assign w257 = ~w254 & w256;
assign w258 = ~w251 & ~w257;
assign w259 = ~w249 & w258;
assign w260 = (pi10241 & ~w229) | (pi10241 & w54894) | (~w229 & w54894);
assign w261 = w229 & w54750;
assign w262 = ~pi10240 & ~pi10241;
assign w263 = w238 & w54832;
assign w264 = (pi10240 & ~w229) | (pi10240 & w54833) | (~w229 & w54833);
assign w265 = ~w263 & ~w264;
assign w266 = (~pi00012 & w264) | (~pi00012 & w54895) | (w264 & w54895);
assign w267 = ~w260 & ~w261;
assign w268 = ~w266 & w267;
assign w269 = w229 & w54773;
assign w270 = (pi00011 & ~w229) | (pi00011 & w54897) | (~w229 & w54897);
assign w271 = ~w266 & w270;
assign w272 = ~w268 & ~w271;
assign w273 = (~w272 & ~w259) | (~w272 & w54733) | (~w259 & w54733);
assign w274 = (~pi10242 & w269) | (~pi10242 & w54834) | (w269 & w54834);
assign w275 = ~w269 & w54835;
assign w276 = ~w274 & ~w275;
assign w277 = pi00013 & w276;
assign w278 = pi00011 & w268;
assign w279 = (pi00012 & ~w229) | (pi00012 & w54898) | (~w229 & w54898);
assign w280 = w265 & w279;
assign w281 = ~w277 & ~w280;
assign w282 = ~w278 & w281;
assign w283 = ~pi00013 & ~w276;
assign w284 = ~pi10022 & ~w274;
assign w285 = pi10022 & w274;
assign w286 = ~w284 & ~w285;
assign w287 = ~w283 & ~w286;
assign w288 = ~pi09967 & pi10387;
assign w289 = pi09924 & ~pi10418;
assign w290 = pi10380 & pi10418;
assign w291 = ~w289 & ~w290;
assign w292 = pi09964 & ~w288;
assign w293 = ~w291 & w292;
assign w294 = ~pi00138 & ~pi09970;
assign w295 = w293 & w54899;
assign w296 = ~pi00137 & ~pi09950;
assign w297 = ~pi10535 & w296;
assign w298 = (~w297 & w293) | (~w297 & w54900) | (w293 & w54900);
assign w299 = (w273 & w54800) | (w273 & w54801) | (w54800 & w54801);
assign w300 = w293 & w297;
assign w301 = pi00015 & w188;
assign w302 = w188 & w54901;
assign w303 = ~pi00036 & ~pi09847;
assign w304 = pi00036 & pi09847;
assign w305 = ~pi00033 & ~pi09814;
assign w306 = pi00033 & pi09814;
assign w307 = pi00034 & ~pi09846;
assign w308 = ~pi00034 & pi09846;
assign w309 = ~w307 & ~w308;
assign w310 = ~pi00035 & ~pi09813;
assign w311 = pi00035 & pi09813;
assign w312 = ~w303 & ~w304;
assign w313 = ~w305 & ~w306;
assign w314 = ~w310 & ~w311;
assign w315 = w313 & w314;
assign w316 = ~w309 & w312;
assign w317 = w315 & w316;
assign w318 = pi10263 & ~w317;
assign w319 = (w302 & w317) | (w302 & w54902) | (w317 & w54902);
assign w320 = ~pi00024 & ~w288;
assign w321 = ~w288 & w54903;
assign w322 = ~w320 & ~w321;
assign w323 = pi00831 & ~pi09879;
assign w324 = ~pi00838 & ~pi09948;
assign w325 = pi00838 & pi09948;
assign w326 = ~w324 & ~w325;
assign w327 = ~pi00830 & pi09944;
assign w328 = pi00837 & ~pi09888;
assign w329 = ~pi00836 & pi09799;
assign w330 = ~pi00831 & pi09879;
assign w331 = pi00834 & ~pi09882;
assign w332 = pi00830 & ~pi09944;
assign w333 = ~pi00840 & pi09979;
assign w334 = ~pi00834 & pi09882;
assign w335 = pi00827 & ~pi09877;
assign w336 = pi00829 & ~pi09978;
assign w337 = ~pi00829 & pi09978;
assign w338 = ~pi00538 & pi09980;
assign w339 = pi00835 & pi09883;
assign w340 = ~pi00835 & ~pi09883;
assign w341 = ~w339 & ~w340;
assign w342 = ~pi00828 & pi09972;
assign w343 = ~pi00839 & pi09971;
assign w344 = ~pi00827 & pi09877;
assign w345 = pi00836 & ~pi09799;
assign w346 = pi00840 & ~pi09979;
assign w347 = ~pi00826 & pi09974;
assign w348 = pi00826 & ~pi09974;
assign w349 = pi00833 & ~pi09881;
assign w350 = pi00839 & ~pi09971;
assign w351 = pi00832 & ~pi09800;
assign w352 = pi00538 & ~pi09980;
assign w353 = pi00828 & ~pi09972;
assign w354 = ~pi00833 & pi09881;
assign w355 = ~pi00832 & pi09800;
assign w356 = ~pi00837 & pi09888;
assign w357 = ~pi09949 & ~w323;
assign w358 = ~w327 & ~w328;
assign w359 = ~w329 & ~w330;
assign w360 = ~w331 & ~w332;
assign w361 = ~w333 & ~w334;
assign w362 = ~w335 & ~w336;
assign w363 = ~w337 & ~w338;
assign w364 = ~w342 & ~w343;
assign w365 = ~w344 & ~w345;
assign w366 = ~w346 & ~w347;
assign w367 = ~w348 & ~w349;
assign w368 = ~w350 & ~w351;
assign w369 = ~w352 & ~w353;
assign w370 = ~w354 & ~w355;
assign w371 = ~w356 & w370;
assign w372 = w368 & w369;
assign w373 = w366 & w367;
assign w374 = w364 & w365;
assign w375 = w362 & w363;
assign w376 = w360 & w361;
assign w377 = w358 & w359;
assign w378 = ~w326 & w357;
assign w379 = ~w341 & w378;
assign w380 = w376 & w377;
assign w381 = w374 & w375;
assign w382 = w372 & w373;
assign w383 = w371 & w382;
assign w384 = w380 & w381;
assign w385 = w379 & w384;
assign w386 = w383 & w385;
assign w387 = w385 & w54836;
assign w388 = ~w319 & ~w387;
assign w389 = w301 & w320;
assign w390 = w293 & w54904;
assign w391 = ~w389 & ~w390;
assign w392 = ~pi00444 & ~pi00475;
assign w393 = ~pi00609 & ~pi00817;
assign w394 = ~pi00878 & ~pi01273;
assign w395 = ~pi09929 & ~pi10264;
assign w396 = ~pi10363 & ~pi10384;
assign w397 = w395 & w396;
assign w398 = w393 & w394;
assign w399 = w392 & w398;
assign w400 = (~pi09952 & ~w399) | (~pi09952 & w54905) | (~w399 & w54905);
assign w401 = w302 & ~w400;
assign w402 = pi00835 & ~pi01273;
assign w403 = w188 & w54837;
assign w404 = w198 & w403;
assign w405 = w403 & w54906;
assign w406 = ~pi00038 & w405;
assign w407 = ~pi00835 & pi01273;
assign w408 = ~pi00817 & pi00837;
assign w409 = ~pi00834 & pi09929;
assign w410 = pi00444 & ~pi00827;
assign w411 = ~pi00832 & pi10363;
assign w412 = ~pi00475 & pi00839;
assign w413 = pi00609 & pi00838;
assign w414 = ~pi00609 & ~pi00838;
assign w415 = ~w413 & ~w414;
assign w416 = ~pi00836 & pi00878;
assign w417 = ~pi00444 & pi00827;
assign w418 = pi00833 & ~pi10264;
assign w419 = ~pi00833 & pi10264;
assign w420 = pi00817 & ~pi00837;
assign w421 = pi00834 & ~pi09929;
assign w422 = pi00836 & ~pi00878;
assign w423 = pi00832 & ~pi10363;
assign w424 = pi00475 & ~pi00839;
assign w425 = pi00831 & ~pi10384;
assign w426 = ~pi00831 & pi10384;
assign w427 = ~w402 & ~w407;
assign w428 = ~w408 & ~w409;
assign w429 = ~w410 & ~w411;
assign w430 = ~w412 & ~w416;
assign w431 = ~w417 & ~w418;
assign w432 = ~w419 & ~w420;
assign w433 = ~w421 & ~w422;
assign w434 = ~w423 & ~w424;
assign w435 = ~w425 & ~w426;
assign w436 = w434 & w435;
assign w437 = w432 & w433;
assign w438 = w430 & w431;
assign w439 = w428 & w429;
assign w440 = ~w415 & w427;
assign w441 = w439 & w440;
assign w442 = w437 & w438;
assign w443 = w436 & w442;
assign w444 = w443 & w54907;
assign w445 = ~pi09967 & ~pi10452;
assign w446 = pi00019 & ~pi01269;
assign w447 = ~pi00019 & pi01461;
assign w448 = ~pi00017 & pi01460;
assign w449 = ~pi00018 & pi01278;
assign w450 = ~w448 & ~w449;
assign w451 = pi00006 & ~pi01456;
assign w452 = pi00015 & ~pi01458;
assign w453 = pi00014 & ~pi01457;
assign w454 = ~w452 & ~w453;
assign w455 = pi00019 & ~pi01461;
assign w456 = pi00018 & ~pi01278;
assign w457 = ~w455 & ~w456;
assign w458 = pi00016 & ~pi01459;
assign w459 = pi00017 & ~pi01460;
assign w460 = ~w458 & ~w459;
assign w461 = ~pi00014 & pi01457;
assign w462 = ~pi00016 & pi01459;
assign w463 = ~pi00015 & pi01458;
assign w464 = ~w462 & ~w463;
assign w465 = ~pi00006 & pi01456;
assign w466 = ~w461 & ~w465;
assign w467 = w464 & w466;
assign w468 = ~w447 & ~w451;
assign w469 = w450 & w468;
assign w470 = w454 & w457;
assign w471 = w460 & w470;
assign w472 = w467 & w469;
assign w473 = w471 & w472;
assign w474 = ~pi00019 & pi01269;
assign w475 = ~pi00018 & pi01268;
assign w476 = pi00018 & ~pi01268;
assign w477 = pi00017 & ~pi01267;
assign w478 = ~pi00016 & pi01266;
assign w479 = ~pi00017 & pi01267;
assign w480 = pi00016 & ~pi01266;
assign w481 = pi00015 & ~pi01265;
assign w482 = ~pi00015 & pi01265;
assign w483 = pi00014 & ~pi01264;
assign w484 = ~pi00014 & pi01264;
assign w485 = pi00006 & ~pi01263;
assign w486 = ~w484 & w485;
assign w487 = (~w482 & w486) | (~w482 & w54908) | (w486 & w54908);
assign w488 = ~w480 & ~w481;
assign w489 = ~w478 & ~w479;
assign w490 = (w489 & w487) | (w489 & w54909) | (w487 & w54909);
assign w491 = ~w476 & ~w477;
assign w492 = ~w474 & ~w475;
assign w493 = (w492 & w490) | (w492 & w54910) | (w490 & w54910);
assign w494 = ~pi00032 & ~pi10434;
assign w495 = w445 & w494;
assign w496 = ~w446 & w495;
assign w497 = ~w473 & w496;
assign w498 = ~w493 & w497;
assign w499 = ~w444 & w54911;
assign w500 = w388 & w499;
assign w501 = ~w288 & w54912;
assign w502 = pi00963 & w403;
assign w503 = ~pi09964 & ~pi10354;
assign w504 = pi00024 & w503;
assign w505 = w503 & w536;
assign w506 = (w288 & w502) | (w288 & w54913) | (w502 & w54913);
assign w507 = ~w501 & ~w506;
assign w508 = pi00008 & ~pi00009;
assign w509 = pi00010 & ~pi00011;
assign w510 = ~pi00016 & ~pi00019;
assign w511 = pi00020 & pi00021;
assign w512 = pi00022 & ~pi09968;
assign w513 = w511 & w512;
assign w514 = w509 & w510;
assign w515 = w198 & w508;
assign w516 = w514 & w515;
assign w517 = w301 & w513;
assign w518 = w516 & w517;
assign w519 = ~w518 & w54914;
assign w520 = pi10381 & pi10418;
assign w521 = pi00845 & ~pi01303;
assign w522 = ~pi10418 & w521;
assign w523 = ~w520 & ~w522;
assign w524 = w518 & w54915;
assign w525 = ~pi00038 & pi10476;
assign w526 = pi00007 & ~w525;
assign w527 = ~w302 & w526;
assign w528 = ~w502 & w527;
assign w529 = ~w519 & w528;
assign w530 = w529 & w54916;
assign w531 = w500 & w54838;
assign w532 = (~w273 & w54802) | (~w273 & w54803) | (w54802 & w54803);
assign w533 = ~w299 & w532;
assign w534 = ~w518 & w54751;
assign w535 = ~pi00963 & w503;
assign w536 = pi00024 & pi00031;
assign w537 = w535 & w536;
assign w538 = w535 & w54778;
assign w539 = pi00032 & pi00038;
assign w540 = w538 & w539;
assign w541 = (pi00006 & w534) | (pi00006 & w54917) | (w534 & w54917);
assign w542 = ~w534 & w54918;
assign w543 = ~w541 & ~w542;
assign w544 = w533 & w543;
assign w545 = ~pi00019 & pi01467;
assign w546 = pi00019 & ~pi01467;
assign w547 = ~pi00018 & pi01468;
assign w548 = pi00018 & ~pi01468;
assign w549 = ~pi00017 & pi01466;
assign w550 = pi00016 & ~pi01465;
assign w551 = pi00017 & ~pi01466;
assign w552 = ~pi00016 & pi01465;
assign w553 = ~pi00015 & pi01464;
assign w554 = pi00015 & ~pi01464;
assign w555 = ~pi00014 & pi01462;
assign w556 = ~pi00006 & pi01478;
assign w557 = ~w555 & ~w556;
assign w558 = pi00014 & ~pi01462;
assign w559 = ~w554 & ~w558;
assign w560 = ~w557 & w559;
assign w561 = ~w552 & ~w553;
assign w562 = ~w550 & ~w551;
assign w563 = (w562 & w560) | (w562 & w54919) | (w560 & w54919);
assign w564 = (~w548 & w563) | (~w548 & w54920) | (w563 & w54920);
assign w565 = pi10434 & ~w545;
assign w566 = (~w564 & w54922) | (~w564 & w54923) | (w54922 & w54923);
assign w567 = ~w454 & w464;
assign w568 = w460 & ~w467;
assign w569 = (w450 & ~w568) | (w450 & w54924) | (~w568 & w54924);
assign w570 = ~pi10434 & ~w447;
assign w571 = (w570 & w569) | (w570 & w54925) | (w569 & w54925);
assign w572 = ~w566 & ~w571;
assign w573 = (~pi00007 & w522) | (~pi00007 & w54926) | (w522 & w54926);
assign w574 = ~w445 & w573;
assign w575 = ~pi00007 & w445;
assign w576 = ~w525 & ~w575;
assign w577 = w500 & w54839;
assign w578 = (~w273 & w54804) | (~w273 & w54805) | (w54804 & w54805);
assign w579 = (~w572 & w54927) | (~w572 & w54928) | (w54927 & w54928);
assign w580 = w578 & w579;
assign w581 = (w405 & w534) | (w405 & w54929) | (w534 & w54929);
assign w582 = (w54779 & w534) | (w54779 & w54930) | (w534 & w54930);
assign w583 = (w54806 & w534) | (w54806 & w54840) | (w534 & w54840);
assign w584 = pi00022 & w583;
assign w585 = w583 & w54886;
assign w586 = (~pi00008 & ~w583) | (~pi00008 & w54931) | (~w583 & w54931);
assign w587 = ~w585 & ~w586;
assign w588 = w533 & w587;
assign w589 = (~pi00009 & ~w583) | (~pi00009 & w54932) | (~w583 & w54932);
assign w590 = w583 & w54933;
assign w591 = ~w589 & ~w590;
assign w592 = w533 & w591;
assign w593 = (~pi00010 & ~w583) | (~pi00010 & w54934) | (~w583 & w54934);
assign w594 = w583 & w54935;
assign w595 = ~w593 & ~w594;
assign w596 = w533 & w595;
assign w597 = w583 & w54936;
assign w598 = (~pi00011 & ~w583) | (~pi00011 & w54937) | (~w583 & w54937);
assign w599 = ~w597 & ~w598;
assign w600 = w533 & w599;
assign w601 = (~pi00012 & ~w583) | (~pi00012 & w54938) | (~w583 & w54938);
assign w602 = w583 & w54939;
assign w603 = ~w601 & ~w602;
assign w604 = w533 & w603;
assign w605 = (~pi00013 & ~w583) | (~pi00013 & w54940) | (~w583 & w54940);
assign w606 = w583 & w54941;
assign w607 = ~w605 & ~w606;
assign w608 = w533 & w607;
assign w609 = ~pi00014 & ~w541;
assign w610 = (w188 & w534) | (w188 & w54942) | (w534 & w54942);
assign w611 = ~w609 & ~w610;
assign w612 = w533 & w611;
assign w613 = ~pi00015 & ~w610;
assign w614 = (w301 & w534) | (w301 & w54943) | (w534 & w54943);
assign w615 = ~w613 & ~w614;
assign w616 = w533 & w615;
assign w617 = ~pi00016 & ~w614;
assign w618 = pi00016 & w614;
assign w619 = ~w617 & ~w618;
assign w620 = w533 & w619;
assign w621 = w614 & w54944;
assign w622 = (~pi00017 & ~w614) | (~pi00017 & w54945) | (~w614 & w54945);
assign w623 = ~w621 & ~w622;
assign w624 = w533 & w623;
assign w625 = (w404 & w534) | (w404 & w54946) | (w534 & w54946);
assign w626 = (~w625 & w621) | (~w625 & w54947) | (w621 & w54947);
assign w627 = w533 & w626;
assign w628 = ~pi00019 & ~w625;
assign w629 = ~w581 & ~w628;
assign w630 = w533 & w629;
assign w631 = ~pi00020 & ~w581;
assign w632 = ~w582 & ~w631;
assign w633 = w533 & w632;
assign w634 = ~pi00021 & ~w582;
assign w635 = ~w583 & ~w634;
assign w636 = w533 & w635;
assign w637 = ~pi00022 & ~w583;
assign w638 = ~w584 & ~w637;
assign w639 = w533 & w638;
assign w640 = pi00961 & pi09872;
assign w641 = ~pi09872 & pi10671;
assign w642 = ~w640 & ~w641;
assign w643 = pi00004 & ~w642;
assign w644 = ~pi00004 & w642;
assign w645 = ~w643 & ~w644;
assign w646 = w152 & w645;
assign w647 = ~w152 & ~w645;
assign w648 = ~w646 & ~w647;
assign w649 = w146 & w54948;
assign w650 = pi00051 & w649;
assign w651 = (w76 & w649) | (w76 & w54949) | (w649 & w54949);
assign w652 = ~w650 & w651;
assign w653 = (~w273 & w54841) | (~w273 & w54842) | (w54841 & w54842);
assign w654 = (~w273 & w54843) | (~w273 & w54844) | (w54843 & w54844);
assign w655 = ~w653 & w654;
assign w656 = ~w317 & w54950;
assign w657 = w400 & w656;
assign w658 = ~w506 & w54951;
assign w659 = ~w657 & ~w658;
assign w660 = w578 & w659;
assign w661 = ~pi00041 & w76;
assign w662 = w146 & w54952;
assign w663 = w146 & w54953;
assign w664 = ~w662 & ~w663;
assign w665 = ~pi00054 & w664;
assign w666 = (w76 & w664) | (w76 & w54954) | (w664 & w54954);
assign w667 = ~w665 & w666;
assign w668 = ~pi02656 & ~pi09822;
assign w669 = pi00007 & ~pi00963;
assign w670 = ~pi02666 & w669;
assign w671 = w668 & w670;
assign w672 = ~pi00040 & w671;
assign w673 = ~pi00039 & w671;
assign w674 = (~w273 & w54845) | (~w273 & w54846) | (w54845 & w54846);
assign w675 = ~w519 & ~w674;
assign w676 = (w273 & w54847) | (w273 & w54848) | (w54847 & w54848);
assign w677 = (~w273 & w54863) | (~w273 & w54864) | (w54863 & w54864);
assign w678 = ~w676 & w677;
assign w679 = (pi00032 & w518) | (pi00032 & w54955) | (w518 & w54955);
assign w680 = (~w679 & w572) | (~w679 & w54956) | (w572 & w54956);
assign w681 = w578 & w680;
assign w682 = (~pi00033 & w444) | (~pi00033 & w54957) | (w444 & w54957);
assign w683 = ~w444 & w54958;
assign w684 = (~w273 & w54809) | (~w273 & w54810) | (w54809 & w54810);
assign w685 = (~pi00929 & w522) | (~pi00929 & w54959) | (w522 & w54959);
assign w686 = w518 & w54960;
assign w687 = ~pi10476 & ~w686;
assign w688 = ~w387 & w54961;
assign w689 = (~w273 & w54849) | (~w273 & w54850) | (w54849 & w54850);
assign w690 = ~w682 & ~w683;
assign w691 = w689 & w690;
assign w692 = pi00034 & ~w682;
assign w693 = ~pi00033 & ~pi00034;
assign w694 = (w693 & w444) | (w693 & w54962) | (w444 & w54962);
assign w695 = ~w692 & ~w694;
assign w696 = w689 & w695;
assign w697 = pi00035 & ~w694;
assign w698 = ~pi00035 & w694;
assign w699 = ~w697 & ~w698;
assign w700 = w689 & w699;
assign w701 = (pi00036 & ~w694) | (pi00036 & w13020) | (~w694 & w13020);
assign w702 = w694 & w54963;
assign w703 = ~w701 & ~w702;
assign w704 = w689 & w703;
assign w705 = (pi00038 & ~w656) | (pi00038 & w54964) | (~w656 & w54964);
assign w706 = w578 & ~w705;
assign w707 = pi09964 & ~pi10354;
assign w708 = w707 & w54965;
assign w709 = pi10354 & ~pi10418;
assign w710 = pi00447 & w709;
assign w711 = pi10354 & pi10418;
assign w712 = pi00851 & w711;
assign w713 = w707 & w54966;
assign w714 = ~w710 & ~w712;
assign w715 = w714 & w54967;
assign w716 = ~pi00028 & ~w715;
assign w717 = pi00028 & w715;
assign w718 = ~w716 & ~w717;
assign w719 = w707 & w54968;
assign w720 = pi01449 & w711;
assign w721 = pi00450 & w709;
assign w722 = w707 & w54969;
assign w723 = ~w720 & ~w721;
assign w724 = w723 & w54970;
assign w725 = ~pi00043 & ~w724;
assign w726 = pi00043 & w724;
assign w727 = ~w725 & ~w726;
assign w728 = ~w718 & ~w727;
assign w729 = w718 & w727;
assign w730 = ~w728 & ~w729;
assign w731 = w730 & w54972;
assign w732 = (w730 & w54973) | (w730 & w54974) | (w54973 & w54974);
assign w733 = ~w731 & w732;
assign w734 = w707 & w54975;
assign w735 = pi00449 & w709;
assign w736 = pi09921 & w711;
assign w737 = w707 & w54976;
assign w738 = ~w735 & ~w736;
assign w739 = w738 & w54977;
assign w740 = ~pi00044 & ~w739;
assign w741 = pi00044 & w739;
assign w742 = ~w740 & ~w741;
assign w743 = pi00024 & ~w742;
assign w744 = ~w742 & w54979;
assign w745 = (~w742 & w54980) | (~w742 & w54981) | (w54980 & w54981);
assign w746 = ~w744 & w745;
assign w747 = pi09872 & pi09933;
assign w748 = ~pi09872 & pi10668;
assign w749 = ~w747 & ~w748;
assign w750 = pi00002 & ~w749;
assign w751 = ~pi00002 & w749;
assign w752 = ~w750 & ~w751;
assign w753 = w645 & w752;
assign w754 = ~w645 & ~w752;
assign w755 = ~w753 & ~w754;
assign w756 = w146 & w54982;
assign w757 = pi00060 & w756;
assign w758 = (w76 & w756) | (w76 & w54983) | (w756 & w54983);
assign w759 = ~w757 & w758;
assign w760 = ~w318 & ~w507;
assign w761 = ~w387 & ~w501;
assign w762 = ~w387 & w54984;
assign w763 = ~w686 & w762;
assign w764 = w684 & w763;
assign w765 = w707 & w54985;
assign w766 = pi09807 & w711;
assign w767 = pi00448 & w709;
assign w768 = w707 & w54986;
assign w769 = ~w766 & ~w767;
assign w770 = w769 & w54987;
assign w771 = ~pi00029 & ~w770;
assign w772 = pi00029 & w770;
assign w773 = ~w771 & ~w772;
assign w774 = ~w773 & w54989;
assign w775 = (~w773 & w54990) | (~w773 & w54991) | (w54990 & w54991);
assign w776 = ~w774 & w775;
assign w777 = ~w718 & w54993;
assign w778 = (~w718 & w54994) | (~w718 & w54995) | (w54994 & w54995);
assign w779 = ~w777 & w778;
assign w780 = pi10263 & w760;
assign w781 = ~pi10263 & w506;
assign w782 = w146 & w54998;
assign w783 = (w146 & w54999) | (w146 & w55000) | (w54999 & w55000);
assign w784 = ~w782 & w783;
assign w785 = pi01253 & pi10380;
assign w786 = (w273 & w54851) | (w273 & w54852) | (w54851 & w54852);
assign w787 = ~pi00052 & ~pi10465;
assign w788 = ~w786 & ~w787;
assign w789 = (pi00849 & w522) | (pi00849 & w55001) | (w522 & w55001);
assign w790 = (~w273 & w54853) | (~w273 & w54854) | (w54853 & w54854);
assign w791 = ~w789 & ~w790;
assign w792 = pi00058 & w76;
assign w793 = pi00024 & ~w727;
assign w794 = ~w727 & w55003;
assign w795 = (~w727 & w55004) | (~w727 & w55005) | (w55004 & w55005);
assign w796 = ~w794 & w795;
assign w797 = ~w742 & ~w773;
assign w798 = w742 & w773;
assign w799 = ~w797 & ~w798;
assign w800 = w799 & w55007;
assign w801 = (w799 & w55008) | (w799 & w55009) | (w55008 & w55009);
assign w802 = ~w800 & w801;
assign w803 = ~w727 & ~w742;
assign w804 = ~w743 & ~w793;
assign w805 = ~w803 & ~w804;
assign w806 = (pi00066 & w804) | (pi00066 & w55010) | (w804 & w55010);
assign w807 = ~w804 & w55011;
assign w808 = w671 & ~w806;
assign w809 = ~w807 & w808;
assign w810 = w146 & w55012;
assign w811 = w146 & w55014;
assign w812 = (w146 & w55015) | (w146 & w55016) | (w55015 & w55016);
assign w813 = ~w811 & w812;
assign w814 = ~w718 & ~w773;
assign w815 = w718 & w773;
assign w816 = ~w814 & ~w815;
assign w817 = w816 & w55018;
assign w818 = (w816 & w55019) | (w816 & w55020) | (w55019 & w55020);
assign w819 = ~w817 & w818;
assign w820 = w146 & w55022;
assign w821 = (w146 & w55023) | (w146 & w55024) | (w55023 & w55024);
assign w822 = ~w820 & w821;
assign w823 = w146 & w55026;
assign w824 = (w146 & w55027) | (w146 & w55028) | (w55027 & w55028);
assign w825 = ~w823 & w824;
assign w826 = pi09839 & pi10539;
assign w827 = pi09997 & w826;
assign w828 = pi10266 & ~pi10542;
assign w829 = pi10467 & pi10515;
assign w830 = ~w828 & ~w829;
assign w831 = ~pi01481 & pi10020;
assign w832 = w830 & ~w831;
assign w833 = (~pi00062 & ~w826) | (~pi00062 & w55029) | (~w826 & w55029);
assign w834 = w832 & w833;
assign w835 = ~pi00371 & ~pi00372;
assign w836 = pi00369 & ~w835;
assign w837 = ~pi00321 & ~pi00344;
assign w838 = ~pi00345 & ~pi00346;
assign w839 = ~pi00347 & ~pi00362;
assign w840 = ~pi00363 & ~pi00364;
assign w841 = ~pi00367 & ~pi00368;
assign w842 = ~pi00370 & ~pi10558;
assign w843 = ~pi10561 & w842;
assign w844 = w840 & w841;
assign w845 = w838 & w839;
assign w846 = w837 & w845;
assign w847 = w843 & w844;
assign w848 = ~w836 & w847;
assign w849 = w826 & w55030;
assign w850 = (w849 & ~w848) | (w849 & w55031) | (~w848 & w55031);
assign w851 = ~w834 & ~w850;
assign w852 = pi00376 & ~pi00814;
assign w853 = ~pi00310 & w852;
assign w854 = w852 & w55032;
assign w855 = (~pi10516 & ~w854) | (~pi10516 & w55033) | (~w854 & w55033);
assign w856 = ~pi00308 & ~pi00309;
assign w857 = ~pi10483 & ~pi10486;
assign w858 = pi10492 & pi10495;
assign w859 = pi10520 & w858;
assign w860 = pi10489 & pi10505;
assign w861 = w859 & w860;
assign w862 = w859 & w55034;
assign w863 = w857 & w862;
assign w864 = pi09895 & ~pi10483;
assign w865 = pi09891 & ~pi10492;
assign w866 = ~pi09891 & pi10492;
assign w867 = ~w865 & ~w866;
assign w868 = ~pi09874 & pi10511;
assign w869 = pi09876 & pi10489;
assign w870 = ~pi09895 & pi10483;
assign w871 = pi09874 & ~pi10511;
assign w872 = ~pi09878 & ~pi10520;
assign w873 = pi09878 & pi10520;
assign w874 = ~pi09801 & pi10495;
assign w875 = pi09801 & ~pi10495;
assign w876 = ~w874 & ~w875;
assign w877 = ~pi09880 & ~pi10486;
assign w878 = pi09880 & pi10486;
assign w879 = ~w877 & ~w878;
assign w880 = ~pi09876 & ~pi10489;
assign w881 = ~pi09894 & pi10505;
assign w882 = pi09894 & ~pi10505;
assign w883 = ~w881 & ~w882;
assign w884 = ~w864 & ~w868;
assign w885 = ~w869 & ~w870;
assign w886 = ~w871 & ~w872;
assign w887 = ~w873 & ~w880;
assign w888 = w886 & w887;
assign w889 = w884 & w885;
assign w890 = ~w867 & ~w876;
assign w891 = ~w879 & ~w883;
assign w892 = w890 & w891;
assign w893 = w888 & w889;
assign w894 = w892 & w893;
assign w895 = (w856 & w894) | (w856 & w55035) | (w894 & w55035);
assign w896 = pi00308 & ~pi00309;
assign w897 = pi10511 & w857;
assign w898 = w861 & w897;
assign w899 = ~pi02802 & ~pi10492;
assign w900 = ~pi02797 & ~pi10511;
assign w901 = pi02797 & pi10511;
assign w902 = ~w900 & ~w901;
assign w903 = pi02800 & ~pi10486;
assign w904 = pi02803 & pi10505;
assign w905 = ~pi02799 & ~pi10520;
assign w906 = pi02802 & pi10492;
assign w907 = ~pi02800 & pi10486;
assign w908 = pi02799 & pi10520;
assign w909 = ~pi02801 & pi10495;
assign w910 = pi02801 & ~pi10495;
assign w911 = ~w909 & ~w910;
assign w912 = pi02798 & ~pi10489;
assign w913 = ~pi02798 & pi10489;
assign w914 = ~w912 & ~w913;
assign w915 = ~pi02803 & ~pi10505;
assign w916 = pi02804 & pi10483;
assign w917 = ~pi02804 & ~pi10483;
assign w918 = ~w916 & ~w917;
assign w919 = ~w899 & ~w903;
assign w920 = ~w904 & ~w905;
assign w921 = ~w906 & ~w907;
assign w922 = ~w908 & ~w915;
assign w923 = w921 & w922;
assign w924 = w919 & w920;
assign w925 = ~w902 & ~w911;
assign w926 = ~w914 & ~w918;
assign w927 = w925 & w926;
assign w928 = w923 & w924;
assign w929 = w927 & w928;
assign w930 = (w896 & w929) | (w896 & w55036) | (w929 & w55036);
assign w931 = pi00295 & ~w895;
assign w932 = (w854 & ~w931) | (w854 & w55037) | (~w931 & w55037);
assign w933 = ~w855 & ~w932;
assign w934 = pi10483 & ~pi10486;
assign w935 = w862 & w934;
assign w936 = pi01472 & pi10495;
assign w937 = ~pi01472 & ~pi10495;
assign w938 = ~pi01476 & ~pi10492;
assign w939 = ~pi01474 & pi10483;
assign w940 = pi01471 & ~pi10486;
assign w941 = ~pi01471 & pi10486;
assign w942 = pi01475 & ~pi10511;
assign w943 = pi01476 & pi10492;
assign w944 = ~pi01475 & pi10511;
assign w945 = ~pi01473 & pi10505;
assign w946 = pi01473 & ~pi10505;
assign w947 = ~w945 & ~w946;
assign w948 = pi01470 & ~pi10520;
assign w949 = ~pi01470 & pi10520;
assign w950 = ~w948 & ~w949;
assign w951 = pi01474 & ~pi10483;
assign w952 = ~pi01469 & pi10489;
assign w953 = pi01469 & ~pi10489;
assign w954 = ~w952 & ~w953;
assign w955 = ~w936 & ~w937;
assign w956 = ~w938 & ~w939;
assign w957 = ~w940 & ~w941;
assign w958 = ~w942 & ~w943;
assign w959 = ~w944 & ~w951;
assign w960 = w958 & w959;
assign w961 = w956 & w957;
assign w962 = ~w947 & w955;
assign w963 = ~w950 & ~w954;
assign w964 = w962 & w963;
assign w965 = w960 & w961;
assign w966 = w964 & w965;
assign w967 = (w896 & w966) | (w896 & w55038) | (w966 & w55038);
assign w968 = ~pi00295 & ~pi00296;
assign w969 = w853 & w968;
assign w970 = pi09981 & ~pi10511;
assign w971 = ~pi09981 & pi10511;
assign w972 = ~pi09939 & ~pi10495;
assign w973 = ~pi09941 & pi10486;
assign w974 = ~pi09984 & ~pi10492;
assign w975 = pi09939 & pi10495;
assign w976 = ~pi09982 & ~pi10520;
assign w977 = pi09982 & pi10520;
assign w978 = pi09984 & pi10492;
assign w979 = ~pi09942 & pi10489;
assign w980 = pi09942 & ~pi10489;
assign w981 = ~w979 & ~w980;
assign w982 = ~pi09988 & ~pi10483;
assign w983 = pi09988 & pi10483;
assign w984 = ~w982 & ~w983;
assign w985 = ~pi09985 & pi10505;
assign w986 = pi09985 & ~pi10505;
assign w987 = ~w985 & ~w986;
assign w988 = pi09941 & ~pi10486;
assign w989 = ~w970 & ~w971;
assign w990 = ~w972 & ~w973;
assign w991 = ~w974 & ~w975;
assign w992 = ~w976 & ~w977;
assign w993 = ~w978 & ~w988;
assign w994 = w992 & w993;
assign w995 = w990 & w991;
assign w996 = ~w981 & w989;
assign w997 = ~w984 & ~w987;
assign w998 = w996 & w997;
assign w999 = w994 & w995;
assign w1000 = w998 & w999;
assign w1001 = ~pi10489 & ~pi10505;
assign w1002 = ~pi10511 & w1001;
assign w1003 = w934 & w1002;
assign w1004 = (~pi00308 & ~w1003) | (~pi00308 & w55039) | (~w1003 & w55039);
assign w1005 = ~pi09901 & ~pi10492;
assign w1006 = pi09903 & ~pi10483;
assign w1007 = pi09899 & ~pi10486;
assign w1008 = pi09901 & pi10492;
assign w1009 = ~pi09899 & pi10486;
assign w1010 = ~pi09896 & pi10511;
assign w1011 = pi09896 & ~pi10511;
assign w1012 = pi09897 & pi10489;
assign w1013 = ~pi09897 & ~pi10489;
assign w1014 = ~pi09900 & pi10495;
assign w1015 = pi09900 & ~pi10495;
assign w1016 = ~w1014 & ~w1015;
assign w1017 = pi09898 & ~pi10520;
assign w1018 = ~pi09898 & pi10520;
assign w1019 = ~w1017 & ~w1018;
assign w1020 = ~pi09902 & pi10505;
assign w1021 = pi09902 & ~pi10505;
assign w1022 = ~w1020 & ~w1021;
assign w1023 = ~pi09903 & pi10483;
assign w1024 = ~w1005 & ~w1006;
assign w1025 = ~w1007 & ~w1008;
assign w1026 = ~w1009 & ~w1010;
assign w1027 = ~w1011 & ~w1012;
assign w1028 = ~w1013 & ~w1023;
assign w1029 = w1027 & w1028;
assign w1030 = w1025 & w1026;
assign w1031 = ~w1016 & w1024;
assign w1032 = ~w1019 & ~w1022;
assign w1033 = w1031 & w1032;
assign w1034 = w1029 & w1030;
assign w1035 = w1033 & w1034;
assign w1036 = (pi00308 & ~w862) | (pi00308 & w55040) | (~w862 & w55040);
assign w1037 = ~w1035 & w1036;
assign w1038 = (pi00309 & w1000) | (pi00309 & w55041) | (w1000 & w55041);
assign w1039 = ~w1037 & w1038;
assign w1040 = ~w967 & w969;
assign w1041 = ~w1039 & w1040;
assign w1042 = pi00063 & ~w1041;
assign w1043 = ~w933 & w1042;
assign w1044 = ~pi02792 & pi10483;
assign w1045 = pi02790 & pi10492;
assign w1046 = pi02787 & ~pi10511;
assign w1047 = pi02789 & pi10495;
assign w1048 = pi02053 & ~pi10520;
assign w1049 = ~pi02053 & pi10520;
assign w1050 = ~w1048 & ~w1049;
assign w1051 = ~pi02788 & pi10489;
assign w1052 = pi02788 & ~pi10489;
assign w1053 = ~w1051 & ~w1052;
assign w1054 = ~pi02789 & ~pi10495;
assign w1055 = pi02791 & pi10486;
assign w1056 = ~pi02791 & ~pi10486;
assign w1057 = ~w1055 & ~w1056;
assign w1058 = pi02792 & ~pi10483;
assign w1059 = ~pi02050 & pi10505;
assign w1060 = pi02050 & ~pi10505;
assign w1061 = ~w1059 & ~w1060;
assign w1062 = ~pi02790 & ~pi10492;
assign w1063 = ~pi02787 & pi10511;
assign w1064 = ~w1044 & ~w1045;
assign w1065 = ~w1046 & ~w1047;
assign w1066 = ~w1054 & ~w1058;
assign w1067 = ~w1062 & ~w1063;
assign w1068 = w1066 & w1067;
assign w1069 = w1064 & w1065;
assign w1070 = ~w1050 & ~w1053;
assign w1071 = ~w1057 & ~w1061;
assign w1072 = w1070 & w1071;
assign w1073 = w1068 & w1069;
assign w1074 = w1072 & w1073;
assign w1075 = w853 & w55042;
assign w1076 = (w1075 & w1074) | (w1075 & w55043) | (w1074 & w55043);
assign w1077 = ~w1043 & ~w1076;
assign w1078 = ~w161 & w752;
assign w1079 = w161 & ~w752;
assign w1080 = ~w1078 & ~w1079;
assign w1081 = w146 & w55044;
assign w1082 = ~w152 & w1081;
assign w1083 = w146 & w55045;
assign w1084 = ~w1082 & ~w1083;
assign w1085 = (pi00141 & w1082) | (pi00141 & w55046) | (w1082 & w55046);
assign w1086 = ~w1082 & w55047;
assign w1087 = w76 & ~w1085;
assign w1088 = ~w1086 & w1087;
assign w1089 = (pi00184 & w773) | (pi00184 & w55048) | (w773 & w55048);
assign w1090 = ~w773 & w55049;
assign w1091 = w671 & ~w1089;
assign w1092 = ~w1090 & w1091;
assign w1093 = ~w718 & w55051;
assign w1094 = (~w718 & w55052) | (~w718 & w55053) | (w55052 & w55053);
assign w1095 = ~w1093 & w1094;
assign w1096 = ~pi00100 & w671;
assign w1097 = ~pi00101 & w671;
assign w1098 = ~w161 & w649;
assign w1099 = w146 & w55054;
assign w1100 = ~w1098 & ~w1099;
assign w1101 = (~pi00187 & w1098) | (~pi00187 & w55055) | (w1098 & w55055);
assign w1102 = ~w1098 & w55056;
assign w1103 = w76 & ~w1101;
assign w1104 = ~w1102 & w1103;
assign w1105 = (pi00186 & ~w146) | (pi00186 & w55057) | (~w146 & w55057);
assign w1106 = w146 & w55058;
assign w1107 = w76 & ~w1105;
assign w1108 = ~w1106 & w1107;
assign w1109 = pi00310 & w968;
assign w1110 = ~pi00814 & w856;
assign w1111 = w1109 & w1110;
assign w1112 = w861 & w55059;
assign w1113 = pi00295 & pi00296;
assign w1114 = w853 & w55060;
assign w1115 = (~pi00071 & w1112) | (~pi00071 & w55061) | (w1112 & w55061);
assign w1116 = ~pi00308 & pi00309;
assign w1117 = w853 & w55062;
assign w1118 = w863 & w1117;
assign w1119 = ~w1115 & ~w1118;
assign w1120 = ~w1111 & ~w1119;
assign w1121 = ~pi00814 & ~pi01272;
assign w1122 = pi10345 & w1121;
assign w1123 = w1121 & w55063;
assign w1124 = pi00089 & w1123;
assign w1125 = pi00203 & pi00230;
assign w1126 = pi00320 & pi00342;
assign w1127 = pi10345 & pi10435;
assign w1128 = ~pi00814 & w1127;
assign w1129 = w1127 & w55064;
assign w1130 = (w1125 & w1129) | (w1125 & w55065) | (w1129 & w55065);
assign w1131 = ~w1124 & ~w1130;
assign w1132 = pi00072 & w1131;
assign w1133 = ~pi00348 & ~pi00365;
assign w1134 = pi00342 & ~w1133;
assign w1135 = ~w1131 & ~w1134;
assign w1136 = pi00348 & ~w1131;
assign w1137 = ~w1131 & w55066;
assign w1138 = ~w1135 & ~w1137;
assign w1139 = pi00400 & ~w1138;
assign w1140 = ~w1132 & ~w1139;
assign w1141 = ~w152 & w756;
assign w1142 = w146 & w55067;
assign w1143 = (pi00231 & w1141) | (pi00231 & w55068) | (w1141 & w55068);
assign w1144 = ~w1141 & w55069;
assign w1145 = w76 & ~w1143;
assign w1146 = ~w1144 & w1145;
assign w1147 = pi00074 & w1131;
assign w1148 = pi00377 & ~w1138;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = pi00075 & w1131;
assign w1151 = pi00378 & ~w1138;
assign w1152 = ~w1150 & ~w1151;
assign w1153 = pi00076 & w1131;
assign w1154 = pi00380 & ~w1138;
assign w1155 = ~w1153 & ~w1154;
assign w1156 = pi00077 & w1131;
assign w1157 = pi00381 & ~w1138;
assign w1158 = ~w1156 & ~w1157;
assign w1159 = pi00078 & w1131;
assign w1160 = pi00382 & ~w1138;
assign w1161 = ~w1159 & ~w1160;
assign w1162 = pi00079 & w1131;
assign w1163 = ~w1131 & w55070;
assign w1164 = ~w1162 & ~w1163;
assign w1165 = pi00080 & w1131;
assign w1166 = pi00379 & ~w1138;
assign w1167 = ~w1165 & ~w1166;
assign w1168 = pi00081 & w1131;
assign w1169 = ~w1131 & w55071;
assign w1170 = ~w1168 & ~w1169;
assign w1171 = pi00082 & w1131;
assign w1172 = ~w1131 & w55072;
assign w1173 = ~w1171 & ~w1172;
assign w1174 = pi00083 & w1131;
assign w1175 = ~w1131 & w55073;
assign w1176 = ~w1174 & ~w1175;
assign w1177 = pi00084 & w1131;
assign w1178 = ~w1131 & w55074;
assign w1179 = ~w1177 & ~w1178;
assign w1180 = pi00085 & w1131;
assign w1181 = ~w1131 & w55075;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = pi00086 & w1131;
assign w1184 = pi00399 & ~w1138;
assign w1185 = ~w1183 & ~w1184;
assign w1186 = pi00087 & w1131;
assign w1187 = ~w1131 & w55076;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = pi00088 & w1131;
assign w1190 = ~w1131 & w55077;
assign w1191 = ~w1189 & ~w1190;
assign w1192 = pi00461 & pi10581;
assign w1193 = pi09966 & pi10480;
assign w1194 = pi10471 & w1193;
assign w1195 = (~pi00089 & ~w1193) | (~pi00089 & w55078) | (~w1193 & w55078);
assign w1196 = w1193 & w55079;
assign w1197 = ~w1192 & ~w1195;
assign w1198 = ~w1196 & w1197;
assign w1199 = pi09928 & w1193;
assign w1200 = w1193 & w55080;
assign w1201 = (pi00090 & ~w1193) | (pi00090 & w55081) | (~w1193 & w55081);
assign w1202 = ~pi10471 & ~w1200;
assign w1203 = ~w1201 & w1202;
assign w1204 = pi10579 & pi10580;
assign w1205 = ~pi10664 & ~pi10665;
assign w1206 = ~pi10666 & ~pi10667;
assign w1207 = w1205 & w1206;
assign w1208 = ~pi10663 & ~w1207;
assign w1209 = ~w1207 & w55082;
assign w1210 = ~pi10662 & w1209;
assign w1211 = w1209 & w55083;
assign w1212 = (~pi10575 & ~w1209) | (~pi10575 & w55084) | (~w1209 & w55084);
assign w1213 = pi10658 & ~pi10660;
assign w1214 = ~pi10659 & ~pi10661;
assign w1215 = w1214 & w55085;
assign w1216 = ~pi10654 & ~pi10656;
assign w1217 = w1215 & w55086;
assign w1218 = pi09878 & w1217;
assign w1219 = w1214 & w55087;
assign w1220 = ~pi10658 & ~pi10660;
assign w1221 = w1220 & w55088;
assign w1222 = w1219 & w1221;
assign w1223 = ~pi09834 & w1222;
assign w1224 = ~pi10654 & pi10656;
assign w1225 = w1220 & w1224;
assign w1226 = w1214 & w55089;
assign w1227 = w1225 & w1226;
assign w1228 = pi10410 & w1227;
assign w1229 = w1214 & w55090;
assign w1230 = w1225 & w1229;
assign w1231 = pi09972 & w1230;
assign w1232 = w1215 & w55091;
assign w1233 = pi09943 & w1232;
assign w1234 = w1216 & w1220;
assign w1235 = w1215 & w1234;
assign w1236 = pi09967 & w1235;
assign w1237 = w1219 & w1225;
assign w1238 = pi09858 & w1237;
assign w1239 = pi10654 & ~pi10656;
assign w1240 = w1215 & w55092;
assign w1241 = pi02053 & w1240;
assign w1242 = w1229 & w55092;
assign w1243 = pi09992 & w1242;
assign w1244 = w1229 & w55086;
assign w1245 = pi09986 & w1244;
assign w1246 = ~w1223 & ~w1228;
assign w1247 = ~w1231 & ~w1236;
assign w1248 = ~w1238 & w1247;
assign w1249 = w1211 & w1246;
assign w1250 = ~w1218 & ~w1233;
assign w1251 = ~w1241 & ~w1243;
assign w1252 = ~w1245 & w1251;
assign w1253 = w1249 & w1250;
assign w1254 = w1253 & w55093;
assign w1255 = ~w1212 & ~w1254;
assign w1256 = (~pi10568 & ~w1209) | (~pi10568 & w55094) | (~w1209 & w55094);
assign w1257 = pi09881 & w1230;
assign w1258 = w1220 & w1239;
assign w1259 = w1215 & w1258;
assign w1260 = pi00854 & w1259;
assign w1261 = pi09829 & w1222;
assign w1262 = pi09803 & w1235;
assign w1263 = pi10414 & w1227;
assign w1264 = w1229 & w1258;
assign w1265 = pi01465 & w1264;
assign w1266 = w1221 & w1229;
assign w1267 = pi09842 & w1266;
assign w1268 = w1215 & w1221;
assign w1269 = pi01459 & w1268;
assign w1270 = pi09907 & w1244;
assign w1271 = pi02800 & w1217;
assign w1272 = pi09916 & w1242;
assign w1273 = pi01471 & w1240;
assign w1274 = pi09887 & w1232;
assign w1275 = w1226 & w1234;
assign w1276 = pi09805 & w1275;
assign w1277 = w1219 & w1234;
assign w1278 = pi00478 & w1277;
assign w1279 = w1215 & w1225;
assign w1280 = pi01266 & w1279;
assign w1281 = w1229 & w1234;
assign w1282 = pi01256 & w1281;
assign w1283 = ~pi09852 & w1237;
assign w1284 = ~w1257 & ~w1260;
assign w1285 = ~w1261 & ~w1262;
assign w1286 = ~w1263 & ~w1265;
assign w1287 = ~w1267 & ~w1269;
assign w1288 = ~w1276 & ~w1278;
assign w1289 = ~w1280 & ~w1282;
assign w1290 = ~w1283 & w1289;
assign w1291 = w1287 & w1288;
assign w1292 = w1285 & w1286;
assign w1293 = w1211 & w1284;
assign w1294 = ~w1270 & ~w1271;
assign w1295 = ~w1272 & ~w1273;
assign w1296 = ~w1274 & w1295;
assign w1297 = w1293 & w1294;
assign w1298 = w1291 & w1292;
assign w1299 = w1290 & w1298;
assign w1300 = w1296 & w1297;
assign w1301 = w1299 & w1300;
assign w1302 = ~w1256 & ~w1301;
assign w1303 = (~pi10559 & ~w1209) | (~pi10559 & w55095) | (~w1209 & w55095);
assign w1304 = pi01255 & w1281;
assign w1305 = pi09915 & w1242;
assign w1306 = pi09906 & w1244;
assign w1307 = pi00482 & w1277;
assign w1308 = pi01464 & w1264;
assign w1309 = pi09886 & w1232;
assign w1310 = pi09851 & w1237;
assign w1311 = pi09860 & w1275;
assign w1312 = pi09828 & w1222;
assign w1313 = w1219 & w1258;
assign w1314 = pi01253 & w1313;
assign w1315 = pi01470 & w1240;
assign w1316 = pi02799 & w1217;
assign w1317 = ~pi00964 & w1259;
assign w1318 = pi09800 & w1230;
assign w1319 = pi01458 & w1268;
assign w1320 = w1226 & w1258;
assign w1321 = pi00843 & w1320;
assign w1322 = ~pi09841 & w1266;
assign w1323 = w1221 & w1226;
assign w1324 = pi10355 & w1323;
assign w1325 = ~pi09869 & w1235;
assign w1326 = pi10402 & w1227;
assign w1327 = pi01265 & w1279;
assign w1328 = ~w1304 & ~w1307;
assign w1329 = ~w1308 & ~w1310;
assign w1330 = ~w1311 & ~w1312;
assign w1331 = ~w1314 & ~w1317;
assign w1332 = ~w1318 & ~w1319;
assign w1333 = ~w1321 & ~w1322;
assign w1334 = ~w1324 & ~w1325;
assign w1335 = ~w1326 & ~w1327;
assign w1336 = w1334 & w1335;
assign w1337 = w1332 & w1333;
assign w1338 = w1330 & w1331;
assign w1339 = w1328 & w1329;
assign w1340 = w1211 & ~w1305;
assign w1341 = ~w1306 & ~w1309;
assign w1342 = ~w1315 & ~w1316;
assign w1343 = w1341 & w1342;
assign w1344 = w1339 & w1340;
assign w1345 = w1337 & w1338;
assign w1346 = w1336 & w1345;
assign w1347 = w1343 & w1344;
assign w1348 = w1346 & w1347;
assign w1349 = ~w1303 & ~w1348;
assign w1350 = pi00095 & w1192;
assign w1351 = w1192 & w54696;
assign w1352 = pi00119 & w1351;
assign w1353 = w1351 & w54706;
assign w1354 = pi00121 & pi00180;
assign w1355 = w1351 & w54734;
assign w1356 = (~pi00094 & ~w1355) | (~pi00094 & w55098) | (~w1355 & w55098);
assign w1357 = (~w1194 & ~w1355) | (~w1194 & w55099) | (~w1355 & w55099);
assign w1358 = ~w1356 & w1357;
assign w1359 = w1193 & w55100;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = ~pi00095 & ~w1192;
assign w1362 = ~w1194 & ~w1350;
assign w1363 = ~w1361 & w1362;
assign w1364 = w1193 & w55101;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = (~pi00096 & ~w1192) | (~pi00096 & w55102) | (~w1192 & w55102);
assign w1367 = ~w1194 & ~w1351;
assign w1368 = ~w1366 & w1367;
assign w1369 = w1193 & w55103;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = pi10432 & w826;
assign w1372 = w826 & w55104;
assign w1373 = ~pi00435 & ~pi10430;
assign w1374 = pi00098 & w1373;
assign w1375 = w1373 & w54697;
assign w1376 = pi00124 & w1375;
assign w1377 = w1375 & w54707;
assign w1378 = w1375 & w54735;
assign w1379 = w1378 & w54752;
assign w1380 = (~pi00097 & ~w1378) | (~pi00097 & w55106) | (~w1378 & w55106);
assign w1381 = pi00097 & pi00130;
assign w1382 = (~w1371 & ~w1378) | (~w1371 & w55108) | (~w1378 & w55108);
assign w1383 = ~w1380 & w1382;
assign w1384 = ~w1372 & ~w1383;
assign w1385 = ~pi00098 & ~w1373;
assign w1386 = ~w1371 & ~w1374;
assign w1387 = ~w1385 & w1386;
assign w1388 = w826 & w55109;
assign w1389 = ~w1387 & ~w1388;
assign w1390 = (~pi00099 & ~w1373) | (~pi00099 & w55110) | (~w1373 & w55110);
assign w1391 = ~w1371 & ~w1375;
assign w1392 = ~w1390 & w1391;
assign w1393 = w826 & w55111;
assign w1394 = ~w1392 & ~w1393;
assign w1395 = ~w727 & w55113;
assign w1396 = (~w727 & w55114) | (~w727 & w55115) | (w55114 & w55115);
assign w1397 = ~w1395 & w1396;
assign w1398 = ~w742 & w55117;
assign w1399 = (~w742 & w55118) | (~w742 & w55119) | (w55118 & w55119);
assign w1400 = ~w1398 & w1399;
assign w1401 = ~pi10449 & pi10509;
assign w1402 = ~pi00102 & ~w1401;
assign w1403 = pi00241 & pi09969;
assign w1404 = pi00242 & w1403;
assign w1405 = w1403 & w2598;
assign w1406 = pi00244 & w1405;
assign w1407 = w1405 & w54736;
assign w1408 = w1405 & w54753;
assign w1409 = ~pi00247 & ~w1408;
assign w1410 = pi00245 & pi00246;
assign w1411 = pi00247 & w1410;
assign w1412 = w1406 & w1411;
assign w1413 = ~w1409 & ~w1412;
assign w1414 = pi10023 & ~w1413;
assign w1415 = (~pi00248 & ~w1406) | (~pi00248 & w54754) | (~w1406 & w54754);
assign w1416 = w1406 & w1482;
assign w1417 = ~w1415 & ~w1416;
assign w1418 = pi10239 & ~w1417;
assign w1419 = ~pi10023 & w1413;
assign w1420 = (~pi00246 & ~w1405) | (~pi00246 & w54755) | (~w1405 & w54755);
assign w1421 = ~w1408 & ~w1420;
assign w1422 = ~pi10024 & w1421;
assign w1423 = (~pi00245 & ~w1405) | (~pi00245 & w18) | (~w1405 & w18);
assign w1424 = ~w1407 & ~w1423;
assign w1425 = pi10025 & ~w1424;
assign w1426 = pi10024 & ~w1421;
assign w1427 = ~pi10025 & w1424;
assign w1428 = ~pi00244 & ~w1405;
assign w1429 = ~w1406 & ~w1428;
assign w1430 = pi10236 & ~w1429;
assign w1431 = ~pi00241 & ~pi09969;
assign w1432 = ~w1403 & ~w1431;
assign w1433 = ~pi10234 & w1432;
assign w1434 = ~pi00242 & ~w1403;
assign w1435 = ~w1404 & ~w1434;
assign w1436 = ~pi10235 & w1435;
assign w1437 = pi10234 & ~w1432;
assign w1438 = ~pi00240 & pi10026;
assign w1439 = pi00240 & ~pi10026;
assign w1440 = ~pi00233 & pi10027;
assign w1441 = ~w1439 & w1440;
assign w1442 = ~w1438 & ~w1441;
assign w1443 = ~w1437 & w1442;
assign w1444 = ~w1433 & ~w1436;
assign w1445 = ~w1443 & w1444;
assign w1446 = pi10235 & ~w1435;
assign w1447 = (~pi00243 & ~w1403) | (~pi00243 & w17) | (~w1403 & w17);
assign w1448 = ~w1405 & ~w1447;
assign w1449 = pi10237 & ~w1448;
assign w1450 = ~w1446 & ~w1449;
assign w1451 = ~w1445 & w1450;
assign w1452 = ~pi10236 & w1429;
assign w1453 = ~pi10237 & w1448;
assign w1454 = ~w1452 & ~w1453;
assign w1455 = (~w1430 & w1451) | (~w1430 & w54708) | (w1451 & w54708);
assign w1456 = ~w1425 & ~w1426;
assign w1457 = ~w1419 & ~w1422;
assign w1458 = (~w1455 & w54756) | (~w1455 & w54757) | (w54756 & w54757);
assign w1459 = ~w1414 & ~w1418;
assign w1460 = (~pi00234 & ~w1406) | (~pi00234 & w54780) | (~w1406 & w54780);
assign w1461 = w1406 & w54781;
assign w1462 = ~w1460 & ~w1461;
assign w1463 = ~pi10238 & w1462;
assign w1464 = ~pi10239 & w1417;
assign w1465 = ~w1463 & ~w1464;
assign w1466 = pi10238 & ~w1462;
assign w1467 = ~pi00235 & ~w1461;
assign w1468 = pi00234 & pi00235;
assign w1469 = w1406 & w54783;
assign w1470 = (pi10021 & w1467) | (pi10021 & w54855) | (w1467 & w54855);
assign w1471 = ~w1466 & ~w1470;
assign w1472 = (~w1458 & w54811) | (~w1458 & w54812) | (w54811 & w54812);
assign w1473 = ~pi00236 & ~w1469;
assign w1474 = pi00236 & w1469;
assign w1475 = ~w1473 & ~w1474;
assign w1476 = ~pi10241 & w1475;
assign w1477 = ~w1467 & w55120;
assign w1478 = ~w1476 & ~w1477;
assign w1479 = pi10241 & ~w1475;
assign w1480 = (~pi00237 & ~w1469) | (~pi00237 & w15) | (~w1469 & w15);
assign w1481 = pi00236 & w1468;
assign w1482 = w1410 & w54758;
assign w1483 = w1468 & w54759;
assign w1484 = w1482 & w1483;
assign w1485 = w1406 & w1484;
assign w1486 = (pi10240 & w1480) | (pi10240 & w55121) | (w1480 & w55121);
assign w1487 = ~w1479 & ~w1486;
assign w1488 = pi00238 & w1485;
assign w1489 = (pi00239 & ~w1485) | (pi00239 & w54857) | (~w1485 & w54857);
assign w1490 = w1485 & w54858;
assign w1491 = ~w1489 & ~w1490;
assign w1492 = ~pi10022 & ~w1491;
assign w1493 = ~pi00238 & ~w1485;
assign w1494 = ~w1488 & ~w1493;
assign w1495 = ~pi10242 & w1494;
assign w1496 = ~w1480 & w55122;
assign w1497 = ~w1492 & ~w1495;
assign w1498 = ~w1496 & w1497;
assign w1499 = (~w1472 & w55123) | (~w1472 & w55124) | (w55123 & w55124);
assign w1500 = ~pi09980 & ~w1491;
assign w1501 = ~pi09972 & w1462;
assign w1502 = ~pi09971 & w1417;
assign w1503 = pi09948 & ~w1413;
assign w1504 = pi09971 & ~w1417;
assign w1505 = ~pi09888 & w1421;
assign w1506 = ~pi09948 & w1413;
assign w1507 = ~pi09882 & w1448;
assign w1508 = ~pi09881 & w1435;
assign w1509 = ~w88 & w54709;
assign w1510 = ~w1432 & ~w1509;
assign w1511 = pi09881 & ~w1435;
assign w1512 = (pi09800 & w88) | (pi09800 & w54710) | (w88 & w54710);
assign w1513 = ~w1511 & ~w1512;
assign w1514 = ~w1510 & w1513;
assign w1515 = ~w1507 & ~w1508;
assign w1516 = ~w1514 & w1515;
assign w1517 = pi09883 & ~w1429;
assign w1518 = pi09882 & ~w1448;
assign w1519 = ~w1517 & ~w1518;
assign w1520 = ~w1516 & w1519;
assign w1521 = ~pi09799 & w1424;
assign w1522 = ~pi09883 & w1429;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = pi09799 & ~w1424;
assign w1525 = pi09888 & ~w1421;
assign w1526 = ~w1524 & ~w1525;
assign w1527 = (w1526 & w1520) | (w1526 & w54738) | (w1520 & w54738);
assign w1528 = ~w1505 & ~w1506;
assign w1529 = ~w1503 & ~w1504;
assign w1530 = ~w1501 & ~w1502;
assign w1531 = (~w1527 & w54760) | (~w1527 & w54761) | (w54760 & w54761);
assign w1532 = (pi09974 & w1467) | (pi09974 & w55125) | (w1467 & w55125);
assign w1533 = pi09972 & ~w1462;
assign w1534 = ~w1532 & ~w1533;
assign w1535 = ~pi09978 & w1475;
assign w1536 = ~pi09979 & w1494;
assign w1537 = ~w1480 & w55126;
assign w1538 = ~w1536 & ~w1537;
assign w1539 = ~w1467 & w55127;
assign w1540 = ~w1535 & ~w1539;
assign w1541 = w1538 & w1540;
assign w1542 = (w1541 & w1531) | (w1541 & w54859) | (w1531 & w54859);
assign w1543 = pi09979 & ~w1494;
assign w1544 = (pi09944 & w1480) | (pi09944 & w55128) | (w1480 & w55128);
assign w1545 = pi09978 & ~w1475;
assign w1546 = ~w1544 & ~w1545;
assign w1547 = w1538 & ~w1546;
assign w1548 = pi09980 & w1491;
assign w1549 = ~w1543 & ~w1548;
assign w1550 = pi10022 & w1491;
assign w1551 = pi10242 & ~w1494;
assign w1552 = ~w1492 & w1551;
assign w1553 = ~w1550 & ~w1552;
assign w1554 = ~pi00000 & pi00338;
assign w1555 = pi01252 & pi10516;
assign w1556 = w1554 & w1555;
assign w1557 = ~w1552 & w55129;
assign w1558 = (w1542 & w54813) | (w1542 & w54814) | (w54813 & w54814);
assign w1559 = ~w1499 & w1558;
assign w1560 = ~w1402 & ~w1559;
assign w1561 = w1558 & w55130;
assign w1562 = ~pi00104 & ~pi00145;
assign w1563 = ~pi00103 & ~pi00147;
assign w1564 = ~pi00149 & ~pi00155;
assign w1565 = ~pi00151 & ~pi00154;
assign w1566 = ~pi00142 & ~pi00143;
assign w1567 = ~pi00144 & pi00146;
assign w1568 = ~pi00148 & ~pi00150;
assign w1569 = ~pi00152 & pi00153;
assign w1570 = w1568 & w1569;
assign w1571 = w1566 & w1567;
assign w1572 = w1562 & w1563;
assign w1573 = w1564 & w1565;
assign w1574 = w1572 & w1573;
assign w1575 = w1570 & w1571;
assign w1576 = w1574 & w1575;
assign w1577 = pi01252 & pi01303;
assign w1578 = pi10377 & w1577;
assign w1579 = w1577 & w54712;
assign w1580 = pi10386 & w1579;
assign w1581 = w1579 & w54713;
assign w1582 = w1579 & w54739;
assign w1583 = pi10361 & w1582;
assign w1584 = w1582 & w54762;
assign w1585 = w1562 & ~w1576;
assign w1586 = w1585 & w55131;
assign w1587 = pi00103 & ~w1586;
assign w1588 = w1585 & w54763;
assign w1589 = ~w1587 & ~w1588;
assign w1590 = (w1589 & ~w1558) | (w1589 & w55132) | (~w1558 & w55132);
assign w1591 = ~w1561 & ~w1590;
assign w1592 = w1558 & w55133;
assign w1593 = w1582 & w55134;
assign w1594 = (pi00104 & ~w1582) | (pi00104 & w55135) | (~w1582 & w55135);
assign w1595 = ~w1593 & ~w1594;
assign w1596 = ~w1576 & ~w1595;
assign w1597 = (w1596 & ~w1558) | (w1596 & w55136) | (~w1558 & w55136);
assign w1598 = ~w1592 & ~w1597;
assign w1599 = (~pi00105 & ~w1193) | (~pi00105 & w55137) | (~w1193 & w55137);
assign w1600 = w1193 & w55138;
assign w1601 = ~w1192 & ~w1599;
assign w1602 = ~w1600 & w1601;
assign w1603 = (~pi10571 & ~w1209) | (~pi10571 & w55139) | (~w1209 & w55139);
assign w1604 = pi09973 & w1232;
assign w1605 = pi10405 & w1227;
assign w1606 = pi09974 & w1230;
assign w1607 = pi09857 & w1237;
assign w1608 = pi02791 & w1240;
assign w1609 = ~pi09835 & w1222;
assign w1610 = pi09951 & w1235;
assign w1611 = pi09987 & w1244;
assign w1612 = pi09935 & w1242;
assign w1613 = pi09880 & w1217;
assign w1614 = ~w1605 & ~w1606;
assign w1615 = ~w1607 & ~w1609;
assign w1616 = ~w1610 & w1615;
assign w1617 = w1211 & w1614;
assign w1618 = ~w1604 & ~w1608;
assign w1619 = ~w1611 & ~w1612;
assign w1620 = ~w1613 & w1619;
assign w1621 = w1617 & w1618;
assign w1622 = w1621 & w55140;
assign w1623 = ~w1603 & ~w1622;
assign w1624 = (~pi10570 & ~w1209) | (~pi10570 & w55141) | (~w1209 & w55141);
assign w1625 = pi09936 & w1242;
assign w1626 = pi10396 & w1227;
assign w1627 = pi09971 & w1230;
assign w1628 = pi09968 & w1235;
assign w1629 = pi02788 & w1240;
assign w1630 = pi09811 & w1237;
assign w1631 = ~pi09833 & w1222;
assign w1632 = pi09946 & w1232;
assign w1633 = pi09940 & w1244;
assign w1634 = pi09876 & w1217;
assign w1635 = ~w1626 & ~w1627;
assign w1636 = ~w1628 & ~w1630;
assign w1637 = ~w1631 & w1636;
assign w1638 = w1211 & w1635;
assign w1639 = ~w1625 & ~w1629;
assign w1640 = ~w1632 & ~w1633;
assign w1641 = ~w1634 & w1640;
assign w1642 = w1638 & w1639;
assign w1643 = w1642 & w55142;
assign w1644 = ~w1624 & ~w1643;
assign w1645 = (~pi10564 & ~w1209) | (~pi10564 & w55143) | (~w1209 & w55143);
assign w1646 = pi10394 & w1227;
assign w1647 = pi09874 & w1217;
assign w1648 = pi09991 & w1242;
assign w1649 = pi09854 & w1237;
assign w1650 = pi02787 & w1240;
assign w1651 = pi09832 & w1222;
assign w1652 = pi09863 & w1275;
assign w1653 = pi09983 & w1244;
assign w1654 = pi09948 & w1230;
assign w1655 = pi09952 & w1235;
assign w1656 = pi09947 & w1232;
assign w1657 = ~w1646 & ~w1649;
assign w1658 = ~w1651 & ~w1652;
assign w1659 = ~w1654 & ~w1655;
assign w1660 = w1658 & w1659;
assign w1661 = w1211 & w1657;
assign w1662 = ~w1647 & ~w1648;
assign w1663 = ~w1650 & ~w1653;
assign w1664 = ~w1656 & w1663;
assign w1665 = w1661 & w1662;
assign w1666 = w1665 & w55144;
assign w1667 = ~w1645 & ~w1666;
assign w1668 = (~pi10562 & ~w1209) | (~pi10562 & w55145) | (~w1209 & w55145);
assign w1669 = pi09864 & w1275;
assign w1670 = pi09919 & w1242;
assign w1671 = pi02804 & w1217;
assign w1672 = pi09888 & w1230;
assign w1673 = pi09911 & w1244;
assign w1674 = pi00483 & w1277;
assign w1675 = pi09872 & w1235;
assign w1676 = pi01474 & w1240;
assign w1677 = pi09816 & w1222;
assign w1678 = pi10417 & w1227;
assign w1679 = pi09893 & w1232;
assign w1680 = ~w1669 & ~w1672;
assign w1681 = ~w1674 & ~w1675;
assign w1682 = ~w1677 & ~w1678;
assign w1683 = w1681 & w1682;
assign w1684 = w1211 & w1680;
assign w1685 = ~w1670 & ~w1671;
assign w1686 = ~w1673 & ~w1676;
assign w1687 = ~w1679 & w1686;
assign w1688 = w1684 & w1685;
assign w1689 = w1688 & w55146;
assign w1690 = ~w1668 & ~w1689;
assign w1691 = (~pi10567 & ~w1209) | (~pi10567 & w55147) | (~w1209 & w55147);
assign w1692 = pi01268 & w1279;
assign w1693 = pi09798 & w1242;
assign w1694 = pi01476 & w1240;
assign w1695 = pi09909 & w1244;
assign w1696 = pi02802 & w1217;
assign w1697 = pi10415 & w1227;
assign w1698 = pi00479 & w1277;
assign w1699 = pi00855 & w1259;
assign w1700 = pi01258 & w1281;
assign w1701 = pi01278 & w1268;
assign w1702 = pi09830 & w1222;
assign w1703 = pi09862 & w1275;
assign w1704 = pi09871 & w1235;
assign w1705 = pi01468 & w1264;
assign w1706 = pi09883 & w1230;
assign w1707 = pi09890 & w1232;
assign w1708 = ~pi09844 & w1266;
assign w1709 = ~w1692 & ~w1697;
assign w1710 = ~w1698 & ~w1699;
assign w1711 = ~w1700 & ~w1701;
assign w1712 = ~w1702 & ~w1703;
assign w1713 = ~w1704 & ~w1705;
assign w1714 = ~w1706 & ~w1708;
assign w1715 = w1713 & w1714;
assign w1716 = w1711 & w1712;
assign w1717 = w1709 & w1710;
assign w1718 = w1211 & ~w1693;
assign w1719 = ~w1694 & ~w1695;
assign w1720 = ~w1696 & ~w1707;
assign w1721 = w1719 & w1720;
assign w1722 = w1717 & w1718;
assign w1723 = w1715 & w1716;
assign w1724 = w1722 & w1723;
assign w1725 = w1721 & w1724;
assign w1726 = ~w1691 & ~w1725;
assign w1727 = (~pi10573 & ~w1209) | (~pi10573 & w55148) | (~w1209 & w55148);
assign w1728 = pi02789 & w1240;
assign w1729 = pi09810 & w1237;
assign w1730 = ~pi09815 & w1222;
assign w1731 = pi09969 & w1235;
assign w1732 = pi09938 & w1244;
assign w1733 = pi09978 & w1230;
assign w1734 = pi10411 & w1227;
assign w1735 = pi09801 & w1217;
assign w1736 = pi09975 & w1232;
assign w1737 = pi09993 & w1242;
assign w1738 = ~w1729 & ~w1730;
assign w1739 = ~w1731 & ~w1733;
assign w1740 = ~w1734 & w1739;
assign w1741 = w1211 & w1738;
assign w1742 = ~w1728 & ~w1732;
assign w1743 = ~w1735 & ~w1736;
assign w1744 = ~w1737 & w1743;
assign w1745 = w1741 & w1742;
assign w1746 = w1745 & w55149;
assign w1747 = ~w1727 & ~w1746;
assign w1748 = (~pi10560 & ~w1209) | (~pi10560 & w55150) | (~w1209 & w55150);
assign w1749 = pi09882 & w1230;
assign w1750 = pi00480 & w1277;
assign w1751 = pi00856 & w1259;
assign w1752 = pi09861 & w1275;
assign w1753 = pi01267 & w1279;
assign w1754 = ~pi09870 & w1235;
assign w1755 = ~pi09853 & w1237;
assign w1756 = pi01466 & w1264;
assign w1757 = pi02801 & w1217;
assign w1758 = pi09889 & w1232;
assign w1759 = pi09908 & w1244;
assign w1760 = pi01472 & w1240;
assign w1761 = pi09917 & w1242;
assign w1762 = pi01460 & w1268;
assign w1763 = ~pi09843 & w1266;
assign w1764 = pi01257 & w1281;
assign w1765 = pi09817 & w1222;
assign w1766 = pi10416 & w1227;
assign w1767 = ~w1749 & ~w1750;
assign w1768 = ~w1751 & ~w1752;
assign w1769 = ~w1753 & ~w1754;
assign w1770 = ~w1755 & ~w1756;
assign w1771 = ~w1762 & ~w1763;
assign w1772 = ~w1764 & ~w1765;
assign w1773 = ~w1766 & w1772;
assign w1774 = w1770 & w1771;
assign w1775 = w1768 & w1769;
assign w1776 = w1211 & w1767;
assign w1777 = ~w1757 & ~w1758;
assign w1778 = ~w1759 & ~w1760;
assign w1779 = ~w1761 & w1778;
assign w1780 = w1776 & w1777;
assign w1781 = w1774 & w1775;
assign w1782 = w1773 & w1781;
assign w1783 = w1779 & w1780;
assign w1784 = w1782 & w1783;
assign w1785 = ~w1748 & ~w1784;
assign w1786 = (~pi00113 & ~w826) | (~pi00113 & w55151) | (~w826 & w55151);
assign w1787 = w826 & w55152;
assign w1788 = ~w1786 & ~w1787;
assign w1789 = pi00460 & pi10581;
assign w1790 = ~w1371 & w55153;
assign w1791 = ~w1787 & ~w1790;
assign w1792 = (~pi00115 & ~w1355) | (~pi00115 & w55154) | (~w1355 & w55154);
assign w1793 = (~w1194 & ~w1355) | (~w1194 & w55155) | (~w1355 & w55155);
assign w1794 = ~w1792 & w1793;
assign w1795 = w1193 & w55156;
assign w1796 = ~w1794 & ~w1795;
assign w1797 = (~pi10566 & ~w1209) | (~pi10566 & w55157) | (~w1209 & w55157);
assign w1798 = ~pi09836 & w1222;
assign w1799 = pi09979 & w1230;
assign w1800 = pi10412 & w1227;
assign w1801 = pi09990 & w1244;
assign w1802 = pi09949 & w1235;
assign w1803 = pi09994 & w1242;
assign w1804 = pi09894 & w1217;
assign w1805 = pi02050 & w1240;
assign w1806 = pi09976 & w1232;
assign w1807 = ~w1798 & ~w1799;
assign w1808 = ~w1800 & ~w1802;
assign w1809 = w1807 & w1808;
assign w1810 = w1211 & ~w1801;
assign w1811 = ~w1803 & ~w1804;
assign w1812 = ~w1805 & ~w1806;
assign w1813 = w1811 & w1812;
assign w1814 = w1809 & w1810;
assign w1815 = w1813 & w1814;
assign w1816 = ~w1797 & ~w1815;
assign w1817 = w1355 & w55158;
assign w1818 = ~pi00117 & ~w1817;
assign w1819 = (~w1194 & ~w1817) | (~w1194 & w55159) | (~w1817 & w55159);
assign w1820 = ~w1818 & w1819;
assign w1821 = w1193 & w55160;
assign w1822 = ~w1820 & ~w1821;
assign w1823 = (~pi10569 & ~w1209) | (~pi10569 & w55161) | (~w1209 & w55161);
assign w1824 = pi09950 & w1235;
assign w1825 = ~pi09838 & w1222;
assign w1826 = pi09944 & w1230;
assign w1827 = pi09891 & w1217;
assign w1828 = pi10401 & w1227;
assign w1829 = pi09934 & w1242;
assign w1830 = pi09945 & w1232;
assign w1831 = pi09989 & w1244;
assign w1832 = pi02790 & w1240;
assign w1833 = ~w1824 & ~w1825;
assign w1834 = ~w1826 & ~w1828;
assign w1835 = w1833 & w1834;
assign w1836 = w1211 & ~w1827;
assign w1837 = ~w1829 & ~w1830;
assign w1838 = ~w1831 & ~w1832;
assign w1839 = w1837 & w1838;
assign w1840 = w1835 & w1836;
assign w1841 = w1839 & w1840;
assign w1842 = ~w1823 & ~w1841;
assign w1843 = ~pi00119 & ~w1351;
assign w1844 = ~w1194 & ~w1352;
assign w1845 = ~w1843 & w1844;
assign w1846 = w1193 & w55162;
assign w1847 = ~w1845 & ~w1846;
assign w1848 = (~pi00120 & ~w1351) | (~pi00120 & w55163) | (~w1351 & w55163);
assign w1849 = ~w1194 & ~w1353;
assign w1850 = ~w1848 & w1849;
assign w1851 = w1193 & w55164;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = w1193 & w55165;
assign w1854 = w1351 & w55166;
assign w1855 = ~pi00121 & ~w1854;
assign w1856 = ~w1194 & ~w1355;
assign w1857 = ~w1855 & w1856;
assign w1858 = ~w1853 & ~w1857;
assign w1859 = w1378 & w54785;
assign w1860 = pi00123 & w1859;
assign w1861 = (~pi00122 & ~w1859) | (~pi00122 & w55169) | (~w1859 & w55169);
assign w1862 = (~w1371 & ~w1859) | (~w1371 & w55170) | (~w1859 & w55170);
assign w1863 = ~w1861 & w1862;
assign w1864 = w826 & w55171;
assign w1865 = ~w1863 & ~w1864;
assign w1866 = ~pi00123 & ~w1859;
assign w1867 = (~w1371 & ~w1859) | (~w1371 & w55172) | (~w1859 & w55172);
assign w1868 = ~w1866 & w1867;
assign w1869 = w826 & w55173;
assign w1870 = ~w1868 & ~w1869;
assign w1871 = ~pi00124 & ~w1375;
assign w1872 = ~w1371 & ~w1376;
assign w1873 = ~w1871 & w1872;
assign w1874 = w826 & w55174;
assign w1875 = ~w1873 & ~w1874;
assign w1876 = pi00094 & pi00117;
assign w1877 = pi00128 & pi00129;
assign w1878 = w1876 & w1877;
assign w1879 = w1355 & w55175;
assign w1880 = ~pi00125 & ~w1879;
assign w1881 = (~w1194 & ~w1879) | (~w1194 & w55176) | (~w1879 & w55176);
assign w1882 = ~w1880 & w1881;
assign w1883 = w1193 & w55177;
assign w1884 = ~w1882 & ~w1883;
assign w1885 = (~pi00126 & ~w1375) | (~pi00126 & w55178) | (~w1375 & w55178);
assign w1886 = ~w1371 & ~w1377;
assign w1887 = ~w1885 & w1886;
assign w1888 = w826 & w55179;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = ~pi00127 & ~w1378;
assign w1891 = (~w1371 & ~w1378) | (~w1371 & w55180) | (~w1378 & w55180);
assign w1892 = ~w1890 & w1891;
assign w1893 = w826 & w55181;
assign w1894 = ~w1892 & ~w1893;
assign w1895 = (~pi00128 & ~w1355) | (~pi00128 & w55182) | (~w1355 & w55182);
assign w1896 = ~w1194 & ~w1817;
assign w1897 = ~w1895 & w1896;
assign w1898 = w1193 & w55183;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = w1193 & w55184;
assign w1901 = (~pi00129 & ~w1817) | (~pi00129 & w55185) | (~w1817 & w55185);
assign w1902 = ~w1194 & ~w1879;
assign w1903 = ~w1901 & w1902;
assign w1904 = ~w1900 & ~w1903;
assign w1905 = (~pi00130 & ~w1378) | (~pi00130 & w55186) | (~w1378 & w55186);
assign w1906 = (~w1371 & ~w1378) | (~w1371 & w55187) | (~w1378 & w55187);
assign w1907 = ~w1905 & w1906;
assign w1908 = w826 & w55188;
assign w1909 = ~w1907 & ~w1908;
assign w1910 = ~pi00131 & ~w1355;
assign w1911 = (~w1194 & ~w1355) | (~w1194 & w55189) | (~w1355 & w55189);
assign w1912 = ~w1910 & w1911;
assign w1913 = w1193 & w55190;
assign w1914 = ~w1912 & ~w1913;
assign w1915 = (pi00132 & ~w1193) | (pi00132 & w55191) | (~w1193 & w55191);
assign w1916 = w1193 & w55192;
assign w1917 = ~w1915 & ~w1916;
assign w1918 = (pi00133 & ~w1193) | (pi00133 & w55193) | (~w1193 & w55193);
assign w1919 = w1193 & w55194;
assign w1920 = ~w1918 & ~w1919;
assign w1921 = (~pi00134 & ~w1378) | (~pi00134 & w55195) | (~w1378 & w55195);
assign w1922 = ~w1371 & ~w1859;
assign w1923 = ~w1921 & w1922;
assign w1924 = w826 & w55196;
assign w1925 = ~w1923 & ~w1924;
assign w1926 = (~pi00135 & ~w1859) | (~pi00135 & w55197) | (~w1859 & w55197);
assign w1927 = (~w1371 & ~w1859) | (~w1371 & w55198) | (~w1859 & w55198);
assign w1928 = ~w1926 & w1927;
assign w1929 = w826 & w55199;
assign w1930 = ~w1928 & ~w1929;
assign w1931 = (~pi00136 & ~w1378) | (~pi00136 & w55200) | (~w1378 & w55200);
assign w1932 = ~w1371 & ~w1379;
assign w1933 = ~w1931 & w1932;
assign w1934 = w826 & w55201;
assign w1935 = ~w1933 & ~w1934;
assign w1936 = (pi00137 & ~w826) | (pi00137 & w55202) | (~w826 & w55202);
assign w1937 = w826 & w55203;
assign w1938 = ~w1936 & ~w1937;
assign w1939 = (pi00138 & ~w826) | (pi00138 & w55204) | (~w826 & w55204);
assign w1940 = w826 & w55205;
assign w1941 = ~w1939 & ~w1940;
assign w1942 = (pi00139 & ~w826) | (pi00139 & w55206) | (~w826 & w55206);
assign w1943 = w826 & w55207;
assign w1944 = ~w1942 & ~w1943;
assign w1945 = (pi00140 & ~w826) | (pi00140 & w55208) | (~w826 & w55208);
assign w1946 = w826 & w55209;
assign w1947 = ~w1945 & ~w1946;
assign w1948 = pi00343 & w664;
assign w1949 = (w76 & w664) | (w76 & w55210) | (w664 & w55210);
assign w1950 = ~w1948 & w1949;
assign w1951 = w1585 & w54786;
assign w1952 = w1585 & w54815;
assign w1953 = ~pi00148 & w1952;
assign w1954 = w1952 & w54860;
assign w1955 = (pi00142 & ~w1952) | (pi00142 & w55211) | (~w1952 & w55211);
assign w1956 = w1952 & w55212;
assign w1957 = ~w1955 & ~w1956;
assign w1958 = (w1957 & ~w1558) | (w1957 & w55213) | (~w1558 & w55213);
assign w1959 = w1558 & w55214;
assign w1960 = ~w1958 & ~w1959;
assign w1961 = (pi00143 & ~w1952) | (pi00143 & w55215) | (~w1952 & w55215);
assign w1962 = w1952 & w55216;
assign w1963 = ~w1961 & ~w1962;
assign w1964 = (w1963 & ~w1558) | (w1963 & w55217) | (~w1558 & w55217);
assign w1965 = w1558 & w55218;
assign w1966 = ~w1964 & ~w1965;
assign w1967 = w1952 & w55219;
assign w1968 = (pi00144 & ~w1952) | (pi00144 & w55220) | (~w1952 & w55220);
assign w1969 = w1952 & w55221;
assign w1970 = ~w1968 & ~w1969;
assign w1971 = (w1970 & ~w1558) | (w1970 & w55222) | (~w1558 & w55222);
assign w1972 = w1558 & w55223;
assign w1973 = ~w1971 & ~w1972;
assign w1974 = w1558 & w55224;
assign w1975 = (pi00145 & ~w1582) | (pi00145 & w55225) | (~w1582 & w55225);
assign w1976 = (~w1975 & ~w1585) | (~w1975 & w55226) | (~w1585 & w55226);
assign w1977 = (w1976 & ~w1558) | (w1976 & w55227) | (~w1558 & w55227);
assign w1978 = ~w1974 & ~w1977;
assign w1979 = w1558 & w55228;
assign w1980 = pi00153 & w1969;
assign w1981 = (w54715 & ~w1558) | (w54715 & w55229) | (~w1558 & w55229);
assign w1982 = ~w1979 & ~w1981;
assign w1983 = (pi00147 & ~w1585) | (pi00147 & w55230) | (~w1585 & w55230);
assign w1984 = ~w1586 & ~w1983;
assign w1985 = (w1984 & ~w1558) | (w1984 & w55231) | (~w1558 & w55231);
assign w1986 = w1558 & w55232;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = pi00148 & ~w1952;
assign w1989 = ~w1953 & ~w1988;
assign w1990 = (w1989 & ~w1558) | (w1989 & w55233) | (~w1558 & w55233);
assign w1991 = w1558 & w55234;
assign w1992 = ~w1990 & ~w1991;
assign w1993 = w1558 & w55235;
assign w1994 = w1952 & w55236;
assign w1995 = (pi00149 & ~w1952) | (pi00149 & w55237) | (~w1952 & w55237);
assign w1996 = ~w1954 & ~w1995;
assign w1997 = (w1996 & ~w1558) | (w1996 & w55238) | (~w1558 & w55238);
assign w1998 = ~w1993 & ~w1997;
assign w1999 = (pi00150 & ~w1585) | (pi00150 & w55239) | (~w1585 & w55239);
assign w2000 = ~w1951 & ~w1999;
assign w2001 = (w2000 & ~w1558) | (w2000 & w55240) | (~w1558 & w55240);
assign w2002 = w1558 & w55241;
assign w2003 = ~w2001 & ~w2002;
assign w2004 = (pi00151 & ~w1585) | (pi00151 & w55242) | (~w1585 & w55242);
assign w2005 = w1585 & w55243;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = (w2006 & ~w1558) | (w2006 & w55244) | (~w1558 & w55244);
assign w2008 = w1558 & w55245;
assign w2009 = ~w2007 & ~w2008;
assign w2010 = (pi00152 & ~w1952) | (pi00152 & w55246) | (~w1952 & w55246);
assign w2011 = ~w1967 & ~w2010;
assign w2012 = (w2011 & ~w1558) | (w2011 & w55247) | (~w1558 & w55247);
assign w2013 = w1558 & w55248;
assign w2014 = ~w2012 & ~w2013;
assign w2015 = ~pi00153 & ~w1969;
assign w2016 = (w54716 & ~w1558) | (w54716 & w55249) | (~w1558 & w55249);
assign w2017 = w1558 & w55250;
assign w2018 = ~w2016 & ~w2017;
assign w2019 = w1558 & w55251;
assign w2020 = pi00154 & ~w2005;
assign w2021 = ~w1952 & ~w2020;
assign w2022 = (w2021 & ~w1558) | (w2021 & w55252) | (~w1558 & w55252);
assign w2023 = ~w2019 & ~w2022;
assign w2024 = (pi00155 & ~w1952) | (pi00155 & w55253) | (~w1952 & w55253);
assign w2025 = ~w1994 & ~w2024;
assign w2026 = (w2025 & ~w1558) | (w2025 & w55254) | (~w1558 & w55254);
assign w2027 = w1558 & w55255;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = ~pi00209 & ~pi00267;
assign w2030 = ~pi00268 & w2029;
assign w2031 = ~pi00229 & ~pi00269;
assign w2032 = ~pi00270 & w2031;
assign w2033 = ~pi00189 & ~pi00190;
assign w2034 = ~pi00191 & ~pi00202;
assign w2035 = w2033 & w2034;
assign w2036 = w2032 & w2035;
assign w2037 = ~pi00156 & pi00201;
assign w2038 = ~pi00206 & ~pi00208;
assign w2039 = w2037 & w2038;
assign w2040 = w2036 & w2039;
assign w2041 = w2036 & w54764;
assign w2042 = ~w827 & ~w1789;
assign w2043 = (~w2042 & w2041) | (~w2042 & w55256) | (w2041 & w55256);
assign w2044 = ~w2041 & w54787;
assign w2045 = ~w2041 & w54816;
assign w2046 = w2045 & w55257;
assign w2047 = ~w2041 & w54817;
assign w2048 = pi00291 & pi00292;
assign w2049 = ~pi00291 & ~pi00292;
assign w2050 = ~w2048 & ~w2049;
assign w2051 = ~pi00114 & w2050;
assign w2052 = (~w2048 & ~w2050) | (~w2048 & w55258) | (~w2050 & w55258);
assign w2053 = (~w2042 & ~w2047) | (~w2042 & w54818) | (~w2047 & w54818);
assign w2054 = ~w2046 & w2053;
assign w2055 = w54819 & w55259;
assign w2056 = w2036 & w2055;
assign w2057 = pi00156 & ~w2043;
assign w2058 = w826 & w55261;
assign w2059 = w2055 & w55262;
assign w2060 = (w2055 & w55263) | (w2055 & w55264) | (w55263 & w55264);
assign w2061 = ~w2059 & w2060;
assign w2062 = pi00391 & ~w1131;
assign w2063 = pi00157 & w1131;
assign w2064 = ~w2062 & ~w2063;
assign w2065 = pi00392 & ~w1131;
assign w2066 = pi00158 & w1131;
assign w2067 = ~w2065 & ~w2066;
assign w2068 = pi00393 & ~w1131;
assign w2069 = pi00159 & w1131;
assign w2070 = ~w2068 & ~w2069;
assign w2071 = pi00394 & ~w1131;
assign w2072 = pi00160 & w1131;
assign w2073 = ~w2071 & ~w2072;
assign w2074 = pi00395 & ~w1131;
assign w2075 = pi00161 & w1131;
assign w2076 = ~w2074 & ~w2075;
assign w2077 = pi00396 & ~w1131;
assign w2078 = pi00162 & w1131;
assign w2079 = ~w2077 & ~w2078;
assign w2080 = pi00397 & ~w1131;
assign w2081 = pi00163 & w1131;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = pi00398 & ~w1131;
assign w2084 = pi00164 & w1131;
assign w2085 = ~w2083 & ~w2084;
assign w2086 = pi00165 & w1131;
assign w2087 = ~w1135 & ~w1136;
assign w2088 = pi00383 & ~w2087;
assign w2089 = ~w2086 & ~w2088;
assign w2090 = pi00166 & w1131;
assign w2091 = pi00384 & ~w2087;
assign w2092 = ~w2090 & ~w2091;
assign w2093 = pi00167 & w1131;
assign w2094 = pi00386 & ~w2087;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = pi00168 & w1131;
assign w2097 = pi00387 & ~w2087;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = pi00169 & w1131;
assign w2100 = pi00388 & ~w2087;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = pi00170 & w1131;
assign w2103 = pi00389 & ~w2087;
assign w2104 = ~w2102 & ~w2103;
assign w2105 = pi00171 & w1131;
assign w2106 = pi00390 & ~w2087;
assign w2107 = ~w2105 & ~w2106;
assign w2108 = pi00172 & w1131;
assign w2109 = pi00385 & ~w2087;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = pi10483 & w856;
assign w2112 = pi00173 & ~pi10483;
assign w2113 = w896 & w2112;
assign w2114 = ~w2111 & ~w2113;
assign w2115 = w853 & w55265;
assign w2116 = ~w2114 & w2115;
assign w2117 = w862 & w2116;
assign w2118 = w853 & w55266;
assign w2119 = pi00173 & ~pi10516;
assign w2120 = ~w2118 & w2119;
assign w2121 = ~w2117 & ~w2120;
assign w2122 = (~pi00174 & ~w826) | (~pi00174 & w55267) | (~w826 & w55267);
assign w2123 = ~w2058 & ~w2122;
assign w2124 = ~w1371 & w55268;
assign w2125 = pi10572 & w1371;
assign w2126 = ~w2124 & ~w2125;
assign w2127 = (~pi10565 & ~w1209) | (~pi10565 & w55269) | (~w1209 & w55269);
assign w2128 = pi09831 & w1222;
assign w2129 = pi00853 & w1259;
assign w2130 = pi02803 & w1217;
assign w2131 = pi01473 & w1240;
assign w2132 = pi10403 & w1227;
assign w2133 = pi01461 & w1268;
assign w2134 = pi09918 & w1242;
assign w2135 = pi09910 & w1244;
assign w2136 = pi09892 & w1232;
assign w2137 = pi09799 & w1230;
assign w2138 = pi09873 & w1235;
assign w2139 = pi09808 & w1275;
assign w2140 = pi01269 & w1279;
assign w2141 = pi00481 & w1277;
assign w2142 = pi01467 & w1264;
assign w2143 = pi01259 & w1281;
assign w2144 = ~w2128 & ~w2129;
assign w2145 = ~w2132 & ~w2133;
assign w2146 = ~w2137 & ~w2138;
assign w2147 = ~w2139 & ~w2140;
assign w2148 = ~w2141 & ~w2142;
assign w2149 = ~w2143 & w2148;
assign w2150 = w2146 & w2147;
assign w2151 = w2144 & w2145;
assign w2152 = w1211 & ~w2130;
assign w2153 = ~w2131 & ~w2134;
assign w2154 = ~w2135 & ~w2136;
assign w2155 = w2153 & w2154;
assign w2156 = w2151 & w2152;
assign w2157 = w2149 & w2150;
assign w2158 = w2156 & w2157;
assign w2159 = w2155 & w2158;
assign w2160 = ~w2127 & ~w2159;
assign w2161 = (~pi00177 & ~w826) | (~pi00177 & w55270) | (~w826 & w55270);
assign w2162 = ~w2125 & ~w2161;
assign w2163 = (~pi10574 & ~w1209) | (~pi10574 & w55271) | (~w1209 & w55271);
assign w2164 = ~pi09840 & w1266;
assign w2165 = pi09879 & w1230;
assign w2166 = pi01469 & w1240;
assign w2167 = pi09885 & w1232;
assign w2168 = pi02798 & w1217;
assign w2169 = w1220 & w55272;
assign w2170 = pi09809 & w1234;
assign w2171 = (w1226 & w2170) | (w1226 & w55273) | (w2170 & w55273);
assign w2172 = ~pi00966 & w1259;
assign w2173 = pi09827 & w1222;
assign w2174 = pi09905 & w1244;
assign w2175 = pi00477 & w1277;
assign w2176 = pi10413 & w1227;
assign w2177 = pi01457 & w1268;
assign w2178 = ~pi10357 & ~pi10439;
assign w2179 = ~pi00843 & ~pi00962;
assign w2180 = ~pi02658 & ~pi02660;
assign w2181 = ~pi10001 & ~pi10355;
assign w2182 = w2180 & w2181;
assign w2183 = w2178 & w2179;
assign w2184 = w2182 & w2183;
assign w2185 = w1323 & ~w2184;
assign w2186 = pi01252 & w1313;
assign w2187 = pi01462 & w1264;
assign w2188 = pi09850 & w1237;
assign w2189 = pi09804 & w1235;
assign w2190 = pi01254 & w1281;
assign w2191 = pi01264 & w1279;
assign w2192 = pi09914 & w1242;
assign w2193 = ~w2164 & ~w2165;
assign w2194 = ~w2171 & ~w2172;
assign w2195 = ~w2173 & ~w2175;
assign w2196 = ~w2176 & ~w2177;
assign w2197 = ~w2185 & ~w2186;
assign w2198 = ~w2187 & ~w2188;
assign w2199 = ~w2189 & ~w2190;
assign w2200 = ~w2191 & w2199;
assign w2201 = w2197 & w2198;
assign w2202 = w2195 & w2196;
assign w2203 = w2193 & w2194;
assign w2204 = w1211 & ~w2166;
assign w2205 = ~w2167 & ~w2168;
assign w2206 = ~w2174 & ~w2192;
assign w2207 = w2205 & w2206;
assign w2208 = w2203 & w2204;
assign w2209 = w2201 & w2202;
assign w2210 = w2200 & w2209;
assign w2211 = w2207 & w2208;
assign w2212 = w2210 & w2211;
assign w2213 = ~w2163 & ~w2212;
assign w2214 = (~pi10563 & ~w1209) | (~pi10563 & w55274) | (~w1209 & w55274);
assign w2215 = pi09970 & w1235;
assign w2216 = pi10395 & w1227;
assign w2217 = pi09980 & w1230;
assign w2218 = pi09977 & w1232;
assign w2219 = ~pi09837 & w1222;
assign w2220 = pi09937 & w1244;
assign w2221 = pi09895 & w1217;
assign w2222 = pi09995 & w1242;
assign w2223 = pi02792 & w1240;
assign w2224 = ~w2215 & ~w2216;
assign w2225 = ~w2217 & ~w2219;
assign w2226 = w2224 & w2225;
assign w2227 = w1211 & ~w2218;
assign w2228 = ~w2220 & ~w2221;
assign w2229 = ~w2222 & ~w2223;
assign w2230 = w2228 & w2229;
assign w2231 = w2226 & w2227;
assign w2232 = w2230 & w2231;
assign w2233 = ~w2214 & ~w2232;
assign w2234 = (~pi00180 & ~w1351) | (~pi00180 & w55275) | (~w1351 & w55275);
assign w2235 = ~w1194 & ~w1854;
assign w2236 = ~w2234 & w2235;
assign w2237 = w1193 & w55276;
assign w2238 = ~w2236 & ~w2237;
assign w2239 = (~pi00181 & ~w1375) | (~pi00181 & w55277) | (~w1375 & w55277);
assign w2240 = ~w1371 & ~w1378;
assign w2241 = ~w2239 & w2240;
assign w2242 = w826 & w55278;
assign w2243 = ~w2241 & ~w2242;
assign w2244 = w1193 & w55279;
assign w2245 = (~pi00182 & ~w1879) | (~pi00182 & w55280) | (~w1879 & w55280);
assign w2246 = pi00115 & pi00125;
assign w2247 = pi00131 & pi00182;
assign w2248 = w2246 & w2247;
assign w2249 = w1878 & w2248;
assign w2250 = w1355 & w2249;
assign w2251 = ~w1194 & ~w2250;
assign w2252 = ~w2245 & w2251;
assign w2253 = ~w2244 & ~w2252;
assign w2254 = (~pi00183 & ~w1859) | (~pi00183 & w55281) | (~w1859 & w55281);
assign w2255 = w1859 & w55282;
assign w2256 = ~w1371 & ~w2254;
assign w2257 = ~w2255 & w2256;
assign w2258 = w826 & w55283;
assign w2259 = ~w2257 & ~w2258;
assign w2260 = w816 & w55285;
assign w2261 = (w816 & w55286) | (w816 & w55287) | (w55286 & w55287);
assign w2262 = ~w2260 & w2261;
assign w2263 = (pi00359 & w718) | (pi00359 & w55288) | (w718 & w55288);
assign w2264 = ~w718 & w55289;
assign w2265 = w671 & ~w2263;
assign w2266 = ~w2264 & w2265;
assign w2267 = ~pi00361 & w1081;
assign w2268 = (w76 & w1081) | (w76 & w55290) | (w1081 & w55290);
assign w2269 = ~w2267 & w2268;
assign w2270 = (~pi00360 & w1141) | (~pi00360 & w55291) | (w1141 & w55291);
assign w2271 = ~w1141 & w55292;
assign w2272 = w76 & ~w2270;
assign w2273 = ~w2271 & w2272;
assign w2274 = ~pi00813 & ~pi09967;
assign w2275 = pi00274 & ~w2274;
assign w2276 = (~pi00271 & ~w145) | (~pi00271 & w55293) | (~w145 & w55293);
assign w2277 = ~w149 & w158;
assign w2278 = ~w749 & w2277;
assign w2279 = w2278 & w55294;
assign w2280 = ~w2276 & w2279;
assign w2281 = (pi00188 & ~w145) | (pi00188 & w55295) | (~w145 & w55295);
assign w2282 = ~w2280 & ~w2281;
assign w2283 = pi00188 & ~w642;
assign w2284 = w2278 & w55296;
assign w2285 = ~pi00249 & ~w2284;
assign w2286 = ~pi00188 & ~pi00271;
assign w2287 = ~pi00276 & w78;
assign w2288 = w2286 & w2287;
assign w2289 = ~w145 & ~w2288;
assign w2290 = pi00274 & w2274;
assign w2291 = ~pi00272 & pi00273;
assign w2292 = pi00275 & ~pi00277;
assign w2293 = ~pi00301 & w2292;
assign w2294 = (~pi09873 & ~w2293) | (~pi09873 & w55297) | (~w2293 & w55297);
assign w2295 = w141 & w54820;
assign w2296 = (~w2290 & ~w2284) | (~w2290 & w55298) | (~w2284 & w55298);
assign w2297 = (w145 & w2295) | (w145 & w55299) | (w2295 & w55299);
assign w2298 = ~w2289 & ~w2297;
assign w2299 = ~w2297 & w55300;
assign w2300 = ~w2282 & w2299;
assign w2301 = pi00189 & ~w2043;
assign w2302 = w826 & w55302;
assign w2303 = w2055 & w55303;
assign w2304 = (w2055 & w55304) | (w2055 & w55305) | (w55304 & w55305);
assign w2305 = ~w2303 & w2304;
assign w2306 = ~w2041 & w55307;
assign w2307 = w826 & w55309;
assign w2308 = w2055 & w55310;
assign w2309 = (w2055 & w55311) | (w2055 & w55312) | (w55311 & w55312);
assign w2310 = ~w2308 & w2309;
assign w2311 = pi00191 & ~w2043;
assign w2312 = (w2311 & ~w2055) | (w2311 & w55313) | (~w2055 & w55313);
assign w2313 = w826 & w55314;
assign w2314 = (~w2313 & ~w2055) | (~w2313 & w55315) | (~w2055 & w55315);
assign w2315 = ~w2312 & w2314;
assign w2316 = w1211 & w55316;
assign w2317 = w1211 & w1244;
assign w2318 = w1211 & w55317;
assign w2319 = (pi00321 & ~w1209) | (pi00321 & w55318) | (~w1209 & w55318);
assign w2320 = w1211 & w55319;
assign w2321 = w1211 & w1230;
assign w2322 = w1211 & w55320;
assign w2323 = ~w2316 & ~w2319;
assign w2324 = ~w2318 & ~w2320;
assign w2325 = ~w2322 & w2324;
assign w2326 = w2323 & w2325;
assign w2327 = (~pi00193 & ~w826) | (~pi00193 & w55321) | (~w826 & w55321);
assign w2328 = ~w2307 & ~w2327;
assign w2329 = (~pi00194 & ~w826) | (~pi00194 & w55322) | (~w826 & w55322);
assign w2330 = w826 & w55323;
assign w2331 = ~w2329 & ~w2330;
assign w2332 = (~pi00195 & ~w826) | (~pi00195 & w55324) | (~w826 & w55324);
assign w2333 = w826 & w55325;
assign w2334 = ~w2332 & ~w2333;
assign w2335 = (~pi00196 & ~w826) | (~pi00196 & w55326) | (~w826 & w55326);
assign w2336 = ~w2302 & ~w2335;
assign w2337 = (~pi00197 & ~w826) | (~pi00197 & w55327) | (~w826 & w55327);
assign w2338 = ~w2313 & ~w2337;
assign w2339 = (~pi10572 & ~w1209) | (~pi10572 & w55328) | (~w1209 & w55328);
assign w2340 = pi01456 & w1268;
assign w2341 = pi09904 & w1244;
assign w2342 = pi09884 & w1232;
assign w2343 = ~pi02724 & w1323;
assign w2344 = pi09877 & w1230;
assign w2345 = pi01475 & w1240;
assign w2346 = ~pi00965 & w1259;
assign w2347 = ~pi09859 & w1275;
assign w2348 = pi01478 & w1264;
assign w2349 = pi01251 & w1313;
assign w2350 = pi02797 & w1217;
assign w2351 = pi09913 & w1242;
assign w2352 = pi01263 & w1279;
assign w2353 = ~pi00872 & w1320;
assign w2354 = pi10404 & w1227;
assign w2355 = pi09849 & w1237;
assign w2356 = pi00484 & w1277;
assign w2357 = pi01260 & w1281;
assign w2358 = ~pi09845 & w1266;
assign w2359 = pi09826 & w1222;
assign w2360 = pi09868 & w1235;
assign w2361 = ~w2340 & ~w2343;
assign w2362 = ~w2344 & ~w2346;
assign w2363 = ~w2347 & ~w2348;
assign w2364 = ~w2349 & ~w2352;
assign w2365 = ~w2353 & ~w2354;
assign w2366 = ~w2355 & ~w2356;
assign w2367 = ~w2357 & ~w2358;
assign w2368 = ~w2359 & ~w2360;
assign w2369 = w2367 & w2368;
assign w2370 = w2365 & w2366;
assign w2371 = w2363 & w2364;
assign w2372 = w2361 & w2362;
assign w2373 = w1211 & ~w2341;
assign w2374 = ~w2342 & ~w2345;
assign w2375 = ~w2350 & ~w2351;
assign w2376 = w2374 & w2375;
assign w2377 = w2372 & w2373;
assign w2378 = w2370 & w2371;
assign w2379 = w2369 & w2378;
assign w2380 = w2376 & w2377;
assign w2381 = w2379 & w2380;
assign w2382 = ~w2339 & ~w2381;
assign w2383 = pi00304 & pi00305;
assign w2384 = w1355 & w54717;
assign w2385 = w54717 & w54740;
assign w2386 = w2385 & w54788;
assign w2387 = pi00219 & pi00262;
assign w2388 = w2385 & w55329;
assign w2389 = w2388 & w55330;
assign w2390 = (~pi00199 & ~w2388) | (~pi00199 & w55332) | (~w2388 & w55332);
assign w2391 = (~w1194 & ~w2388) | (~w1194 & w55333) | (~w2388 & w55333);
assign w2392 = ~w2390 & w2391;
assign w2393 = w1193 & w55334;
assign w2394 = ~w2392 & ~w2393;
assign w2395 = pi00183 & pi00306;
assign w2396 = pi00307 & w2395;
assign w2397 = pi00264 & pi00287;
assign w2398 = pi00289 & pi00293;
assign w2399 = w2397 & w2398;
assign w2400 = w1860 & w55335;
assign w2401 = pi00227 & pi00228;
assign w2402 = pi00265 & pi00288;
assign w2403 = w2401 & w2402;
assign w2404 = w2400 & w2403;
assign w2405 = pi00224 & pi00225;
assign w2406 = (~pi00200 & ~w2400) | (~pi00200 & w55338) | (~w2400 & w55338);
assign w2407 = (~w1371 & ~w2400) | (~w1371 & w55339) | (~w2400 & w55339);
assign w2408 = ~w2406 & w2407;
assign w2409 = w826 & w55340;
assign w2410 = ~w2408 & ~w2409;
assign w2411 = w2055 & w55342;
assign w2412 = ~pi00201 & ~w2043;
assign w2413 = (w2412 & ~w2055) | (w2412 & w55343) | (~w2055 & w55343);
assign w2414 = ~w2333 & ~w2413;
assign w2415 = pi00202 & ~w2043;
assign w2416 = (~w2055 & w55344) | (~w2055 & w55345) | (w55344 & w55345);
assign w2417 = ~w2056 & ~w2330;
assign w2418 = ~w2416 & w2417;
assign w2419 = pi00294 & ~pi10446;
assign w2420 = (~pi00320 & ~w1127) | (~pi00320 & w55346) | (~w1127 & w55346);
assign w2421 = pi00230 & ~w2420;
assign w2422 = (~pi00203 & w2420) | (~pi00203 & w55347) | (w2420 & w55347);
assign w2423 = ~w2420 & w1125;
assign w2424 = ~w1122 & ~w2422;
assign w2425 = pi00089 & ~pi00105;
assign w2426 = ~pi00089 & pi00105;
assign w2427 = ~w2425 & ~w2426;
assign w2428 = w1122 & ~w2427;
assign w2429 = (~w2428 & ~w2424) | (~w2428 & w55348) | (~w2424 & w55348);
assign w2430 = w2419 & ~w2429;
assign w2431 = (pi00249 & w143) | (pi00249 & w55349) | (w143 & w55349);
assign w2432 = pi00250 & ~w146;
assign w2433 = (~w2431 & w146) | (~w2431 & w55350) | (w146 & w55350);
assign w2434 = w1553 & ~w2433;
assign w2435 = ~w1499 & w2434;
assign w2436 = (~w146 & w55353) | (~w146 & w55354) | (w55353 & w55354);
assign w2437 = ~w2435 & w2436;
assign w2438 = (pi00366 & ~w146) | (pi00366 & w55355) | (~w146 & w55355);
assign w2439 = w146 & w55356;
assign w2440 = w76 & ~w2438;
assign w2441 = ~w2439 & w2440;
assign w2442 = pi00206 & ~w2043;
assign w2443 = (w2442 & ~w2055) | (w2442 & w55357) | (~w2055 & w55357);
assign w2444 = w826 & w55358;
assign w2445 = (~w2444 & ~w2055) | (~w2444 & w55359) | (~w2055 & w55359);
assign w2446 = ~w2443 & w2445;
assign w2447 = ~pi00207 & pi10462;
assign w2448 = pi00357 & ~pi01251;
assign w2449 = ~pi00204 & ~pi09875;
assign w2450 = ~pi00374 & ~pi00434;
assign w2451 = ~pi02811 & ~w2447;
assign w2452 = ~w2448 & ~w2449;
assign w2453 = ~w2450 & w2452;
assign w2454 = w2451 & w2453;
assign w2455 = w826 & w55360;
assign w2456 = ~w2041 & w55361;
assign w2457 = (w2456 & ~w2055) | (w2456 & w55362) | (~w2055 & w55362);
assign w2458 = ~w2411 & ~w2455;
assign w2459 = ~w2457 & w2458;
assign w2460 = w826 & w55363;
assign w2461 = ~w2041 & w55364;
assign w2462 = w2054 & w55365;
assign w2463 = w2054 & w55366;
assign w2464 = pi00209 & ~w2043;
assign w2465 = ~w2463 & w2464;
assign w2466 = ~w2055 & ~w2460;
assign w2467 = ~w2465 & w2466;
assign w2468 = w1211 & w55367;
assign w2469 = w1211 & w55368;
assign w2470 = (pi00347 & ~w1209) | (pi00347 & w55369) | (~w1209 & w55369);
assign w2471 = w1211 & w55370;
assign w2472 = w1211 & w55371;
assign w2473 = ~w2468 & ~w2470;
assign w2474 = ~w2469 & ~w2471;
assign w2475 = ~w2472 & w2474;
assign w2476 = w2473 & w2475;
assign w2477 = w1211 & w55372;
assign w2478 = w1211 & w55373;
assign w2479 = (pi10558 & ~w1209) | (pi10558 & w55374) | (~w1209 & w55374);
assign w2480 = w1211 & w55375;
assign w2481 = w1211 & w55376;
assign w2482 = ~w2477 & ~w2479;
assign w2483 = ~w2478 & ~w2480;
assign w2484 = ~w2481 & w2483;
assign w2485 = w2482 & w2484;
assign w2486 = w1211 & w55377;
assign w2487 = w1211 & w55378;
assign w2488 = (pi00344 & ~w1209) | (pi00344 & w55379) | (~w1209 & w55379);
assign w2489 = w1211 & w55380;
assign w2490 = w1211 & w55381;
assign w2491 = ~w2486 & ~w2488;
assign w2492 = ~w2487 & ~w2489;
assign w2493 = ~w2490 & w2492;
assign w2494 = w2491 & w2493;
assign w2495 = w1211 & w55382;
assign w2496 = w1211 & w55383;
assign w2497 = (pi00346 & ~w1209) | (pi00346 & w55384) | (~w1209 & w55384);
assign w2498 = w1211 & w55385;
assign w2499 = w1211 & w55386;
assign w2500 = ~w2495 & ~w2497;
assign w2501 = ~w2496 & ~w2498;
assign w2502 = ~w2499 & w2501;
assign w2503 = w2500 & w2502;
assign w2504 = w1211 & w55387;
assign w2505 = w1211 & w55388;
assign w2506 = (pi00345 & ~w1209) | (pi00345 & w55389) | (~w1209 & w55389);
assign w2507 = w1211 & w55390;
assign w2508 = w1211 & w55391;
assign w2509 = ~w2504 & ~w2506;
assign w2510 = ~w2505 & ~w2507;
assign w2511 = ~w2508 & w2510;
assign w2512 = w2509 & w2511;
assign w2513 = (~pi00215 & ~w826) | (~pi00215 & w55392) | (~w826 & w55392);
assign w2514 = ~w2444 & ~w2513;
assign w2515 = (~pi00216 & ~w826) | (~pi00216 & w55393) | (~w826 & w55393);
assign w2516 = ~w2455 & ~w2515;
assign w2517 = (~pi00217 & ~w826) | (~pi00217 & w55394) | (~w826 & w55394);
assign w2518 = ~w2460 & ~w2517;
assign w2519 = (~pi00218 & ~w826) | (~pi00218 & w55395) | (~w826 & w55395);
assign w2520 = w826 & w55396;
assign w2521 = ~w2519 & ~w2520;
assign w2522 = w1193 & w55397;
assign w2523 = (~pi00219 & ~w2385) | (~pi00219 & w55399) | (~w2385 & w55399);
assign w2524 = (~w1194 & ~w2385) | (~w1194 & w55400) | (~w2385 & w55400);
assign w2525 = ~w2523 & w2524;
assign w2526 = ~w2522 & ~w2525;
assign w2527 = (~pi00220 & ~w2385) | (~pi00220 & w55401) | (~w2385 & w55401);
assign w2528 = ~w1194 & ~w2388;
assign w2529 = ~w2527 & w2528;
assign w2530 = w1193 & w55402;
assign w2531 = ~w2529 & ~w2530;
assign w2532 = ~pi00221 & ~w2388;
assign w2533 = (~w1194 & ~w2388) | (~w1194 & w55403) | (~w2388 & w55403);
assign w2534 = ~w2532 & w2533;
assign w2535 = w1193 & w55404;
assign w2536 = ~w2534 & ~w2535;
assign w2537 = (~pi00222 & ~w2388) | (~pi00222 & w55405) | (~w2388 & w55405);
assign w2538 = ~w1194 & ~w2389;
assign w2539 = ~w2537 & w2538;
assign w2540 = w1193 & w55406;
assign w2541 = ~w2539 & ~w2540;
assign w2542 = pi00199 & pi00263;
assign w2543 = w2388 & w55407;
assign w2544 = (~pi00223 & ~w2388) | (~pi00223 & w55409) | (~w2388 & w55409);
assign w2545 = w2388 & w55410;
assign w2546 = ~w2544 & ~w2545;
assign w2547 = ~w1194 & ~w2546;
assign w2548 = w1193 & w55411;
assign w2549 = ~w2547 & ~w2548;
assign w2550 = w826 & w55412;
assign w2551 = (~pi00224 & ~w2400) | (~pi00224 & w55414) | (~w2400 & w55414);
assign w2552 = (~w1371 & ~w2400) | (~w1371 & w55415) | (~w2400 & w55415);
assign w2553 = ~w2551 & w2552;
assign w2554 = ~w2550 & ~w2553;
assign w2555 = (~pi00225 & ~w2400) | (~pi00225 & w55416) | (~w2400 & w55416);
assign w2556 = (~w1371 & ~w2400) | (~w1371 & w55417) | (~w2400 & w55417);
assign w2557 = ~w2555 & w2556;
assign w2558 = w826 & w55418;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = pi00200 & pi00266;
assign w2561 = w2400 & w55419;
assign w2562 = (~pi00226 & ~w2561) | (~pi00226 & w55420) | (~w2561 & w55420);
assign w2563 = w2561 & w55421;
assign w2564 = ~w2562 & ~w2563;
assign w2565 = ~w1371 & ~w2564;
assign w2566 = w826 & w55422;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = (~pi00227 & ~w2400) | (~pi00227 & w55424) | (~w2400 & w55424);
assign w2569 = (~w1371 & ~w2400) | (~w1371 & w55425) | (~w2400 & w55425);
assign w2570 = ~w2568 & w2569;
assign w2571 = w826 & w55426;
assign w2572 = ~w2570 & ~w2571;
assign w2573 = w826 & w55427;
assign w2574 = (~pi00228 & ~w2400) | (~pi00228 & w55428) | (~w2400 & w55428);
assign w2575 = ~w1371 & ~w2404;
assign w2576 = ~w2574 & w2575;
assign w2577 = ~w2573 & ~w2576;
assign w2578 = ~pi00269 & w2055;
assign w2579 = pi00229 & ~w2043;
assign w2580 = (w2579 & ~w2055) | (w2579 & w55430) | (~w2055 & w55430);
assign w2581 = (~w2520 & ~w2055) | (~w2520 & w55431) | (~w2055 & w55431);
assign w2582 = ~w2580 & w2581;
assign w2583 = ~pi00230 & w2420;
assign w2584 = ~w2421 & ~w2583;
assign w2585 = (~w1123 & w2584) | (~w1123 & w55432) | (w2584 & w55432);
assign w2586 = w2419 & w2585;
assign w2587 = ~w645 & w1081;
assign w2588 = w146 & w55433;
assign w2589 = (~pi00373 & w2587) | (~pi00373 & w55434) | (w2587 & w55434);
assign w2590 = ~w2587 & w55435;
assign w2591 = w76 & ~w2589;
assign w2592 = ~w2590 & w2591;
assign w2593 = (~w1542 & w54823) | (~w1542 & w54824) | (w54823 & w54824);
assign w2594 = ~w2433 & ~w2593;
assign w2595 = (~w146 & w55438) | (~w146 & w55439) | (w55438 & w55439);
assign w2596 = ~w2594 & w2595;
assign w2597 = ~w2275 & w2286;
assign w2598 = pi00242 & pi00243;
assign w2599 = pi00233 & pi00240;
assign w2600 = pi00241 & w2599;
assign w2601 = pi00238 & pi00239;
assign w2602 = pi00244 & w2601;
assign w2603 = w2598 & w2602;
assign w2604 = w2600 & w2603;
assign w2605 = w1484 & w2604;
assign w2606 = (pi00249 & w74) | (pi00249 & w54793) | (w74 & w54793);
assign w2607 = (~w2605 & w55440) | (~w2605 & w55441) | (w55440 & w55441);
assign w2608 = (~w2605 & w54794) | (~w2605 & w54795) | (w54794 & w54795);
assign w2609 = (w145 & w2295) | (w145 & w55442) | (w2295 & w55442);
assign w2610 = ~pi00233 & ~w2607;
assign w2611 = ~w2608 & ~w2610;
assign w2612 = ~w2609 & w2611;
assign w2613 = pi00240 & w2608;
assign w2614 = w2608 & w54825;
assign w2615 = w2608 & w55443;
assign w2616 = w2608 & w55444;
assign w2617 = w2608 & w55445;
assign w2618 = (~pi00234 & ~w2608) | (~pi00234 & w55446) | (~w2608 & w55446);
assign w2619 = w2608 & w55447;
assign w2620 = ~w2609 & ~w2618;
assign w2621 = ~w2619 & w2620;
assign w2622 = (~pi00235 & ~w2608) | (~pi00235 & w55448) | (~w2608 & w55448);
assign w2623 = w2608 & w55449;
assign w2624 = ~w2609 & ~w2622;
assign w2625 = ~w2623 & w2624;
assign w2626 = ~pi00236 & ~w2623;
assign w2627 = w2608 & w55450;
assign w2628 = ~w2609 & ~w2627;
assign w2629 = ~w2626 & w2628;
assign w2630 = ~w2609 & w55451;
assign w2631 = (~pi00237 & ~w2608) | (~pi00237 & w55452) | (~w2608 & w55452);
assign w2632 = ~w2609 & ~w2630;
assign w2633 = ~w2631 & w2632;
assign w2634 = (~w2609 & ~w2630) | (~w2609 & w55453) | (~w2630 & w55453);
assign w2635 = ~pi00238 & ~w2630;
assign w2636 = w2634 & ~w2635;
assign w2637 = (~pi00239 & ~w2630) | (~pi00239 & w16) | (~w2630 & w16);
assign w2638 = pi00239 & ~w2634;
assign w2639 = ~w2637 & ~w2638;
assign w2640 = ~pi00240 & ~w2608;
assign w2641 = ~w2609 & ~w2613;
assign w2642 = ~w2640 & w2641;
assign w2643 = (~pi00241 & ~w2608) | (~pi00241 & w55454) | (~w2608 & w55454);
assign w2644 = ~w2609 & ~w2614;
assign w2645 = ~w2643 & w2644;
assign w2646 = (~pi00242 & ~w2608) | (~pi00242 & w55455) | (~w2608 & w55455);
assign w2647 = w2608 & w55456;
assign w2648 = ~w2609 & ~w2646;
assign w2649 = ~w2647 & w2648;
assign w2650 = (~pi00243 & ~w2608) | (~pi00243 & w55457) | (~w2608 & w55457);
assign w2651 = ~w2609 & ~w2615;
assign w2652 = ~w2650 & w2651;
assign w2653 = (~pi00244 & ~w2608) | (~pi00244 & w55458) | (~w2608 & w55458);
assign w2654 = ~w2609 & ~w2616;
assign w2655 = ~w2653 & w2654;
assign w2656 = (~pi00245 & ~w2608) | (~pi00245 & w55459) | (~w2608 & w55459);
assign w2657 = w2608 & w55460;
assign w2658 = ~w2609 & ~w2656;
assign w2659 = ~w2657 & w2658;
assign w2660 = (~pi00246 & ~w2608) | (~pi00246 & w55461) | (~w2608 & w55461);
assign w2661 = ~w2609 & w55462;
assign w2662 = ~w2609 & ~w2661;
assign w2663 = ~w2660 & w2662;
assign w2664 = ~pi00247 & ~w2661;
assign w2665 = (pi00247 & w2661) | (pi00247 & w55463) | (w2661 & w55463);
assign w2666 = ~w2664 & ~w2665;
assign w2667 = ~w2609 & w55464;
assign w2668 = ~pi00248 & ~w2667;
assign w2669 = ~w2609 & ~w2617;
assign w2670 = ~w2668 & w2669;
assign w2671 = pi00250 & w2299;
assign w2672 = (~pi00250 & w2284) | (~pi00250 & w55465) | (w2284 & w55465);
assign w2673 = w2298 & w2672;
assign w2674 = (pi00251 & ~w2388) | (pi00251 & w55466) | (~w2388 & w55466);
assign w2675 = (~w1194 & ~w2388) | (~w1194 & w55467) | (~w2388 & w55467);
assign w2676 = ~w2674 & w2675;
assign w2677 = w1193 & w55468;
assign w2678 = ~w2676 & ~w2677;
assign w2679 = (pi00252 & ~w2400) | (pi00252 & w55469) | (~w2400 & w55469);
assign w2680 = (~w1371 & ~w2561) | (~w1371 & w55470) | (~w2561 & w55470);
assign w2681 = ~w2679 & w2680;
assign w2682 = w826 & w55471;
assign w2683 = ~w2681 & ~w2682;
assign w2684 = w1211 & w55472;
assign w2685 = w1211 & w55473;
assign w2686 = (pi00363 & ~w1209) | (pi00363 & w55474) | (~w1209 & w55474);
assign w2687 = w1211 & w55475;
assign w2688 = w1211 & w55476;
assign w2689 = ~w2684 & ~w2686;
assign w2690 = ~w2685 & ~w2687;
assign w2691 = ~w2688 & w2690;
assign w2692 = w2689 & w2691;
assign w2693 = w1211 & w55477;
assign w2694 = w1211 & w55478;
assign w2695 = (pi00362 & ~w1209) | (pi00362 & w55479) | (~w1209 & w55479);
assign w2696 = w1211 & w55480;
assign w2697 = w1211 & w55481;
assign w2698 = ~w2693 & ~w2695;
assign w2699 = ~w2694 & ~w2696;
assign w2700 = ~w2697 & w2699;
assign w2701 = w2698 & w2700;
assign w2702 = w1211 & w55482;
assign w2703 = w1211 & w55483;
assign w2704 = (pi00364 & ~w1209) | (pi00364 & w55484) | (~w1209 & w55484);
assign w2705 = w1211 & w55485;
assign w2706 = w1211 & w55486;
assign w2707 = ~w2702 & ~w2704;
assign w2708 = ~w2703 & ~w2705;
assign w2709 = ~w2706 & w2708;
assign w2710 = w2707 & w2709;
assign w2711 = w1211 & w55487;
assign w2712 = w1211 & w55488;
assign w2713 = (pi10561 & ~w1209) | (pi10561 & w55489) | (~w1209 & w55489);
assign w2714 = w1211 & w55490;
assign w2715 = w1211 & w55491;
assign w2716 = ~w2711 & ~w2713;
assign w2717 = ~w2712 & ~w2714;
assign w2718 = ~w2715 & w2717;
assign w2719 = w2716 & w2718;
assign w2720 = (~pi00257 & ~w826) | (~pi00257 & w55492) | (~w826 & w55492);
assign w2721 = w826 & w55493;
assign w2722 = ~w2720 & ~w2721;
assign w2723 = (~pi00258 & ~w826) | (~pi00258 & w55494) | (~w826 & w55494);
assign w2724 = w826 & w55495;
assign w2725 = ~w2723 & ~w2724;
assign w2726 = (~pi00259 & ~w826) | (~pi00259 & w55496) | (~w826 & w55496);
assign w2727 = w826 & w55497;
assign w2728 = ~w2726 & ~w2727;
assign w2729 = (~pi00260 & ~w826) | (~pi00260 & w55498) | (~w826 & w55498);
assign w2730 = w826 & w55499;
assign w2731 = ~w2729 & ~w2730;
assign w2732 = (~pi00261 & ~w2385) | (~pi00261 & w55500) | (~w2385 & w55500);
assign w2733 = (~w1194 & ~w2385) | (~w1194 & w55501) | (~w2385 & w55501);
assign w2734 = ~w2732 & w2733;
assign w2735 = w1193 & w55502;
assign w2736 = ~w2734 & ~w2735;
assign w2737 = (~pi00262 & ~w2385) | (~pi00262 & w55503) | (~w2385 & w55503);
assign w2738 = (~w1194 & ~w2385) | (~w1194 & w55504) | (~w2385 & w55504);
assign w2739 = ~w2737 & w2738;
assign w2740 = w1193 & w55505;
assign w2741 = ~w2739 & ~w2740;
assign w2742 = w1193 & w55506;
assign w2743 = (~pi00263 & ~w2388) | (~pi00263 & w55507) | (~w2388 & w55507);
assign w2744 = ~w1194 & ~w2543;
assign w2745 = ~w2743 & w2744;
assign w2746 = ~w2742 & ~w2745;
assign w2747 = w826 & w55508;
assign w2748 = w1860 & w55509;
assign w2749 = w2748 & w2397;
assign w2750 = (w2748 & w55511) | (w2748 & w55512) | (w55511 & w55512);
assign w2751 = ~w2749 & w2750;
assign w2752 = ~w2747 & ~w2751;
assign w2753 = (~pi00265 & ~w2400) | (~pi00265 & w55513) | (~w2400 & w55513);
assign w2754 = (~w1371 & ~w2400) | (~w1371 & w55514) | (~w2400 & w55514);
assign w2755 = ~w2753 & w2754;
assign w2756 = w826 & w55515;
assign w2757 = ~w2755 & ~w2756;
assign w2758 = w826 & w55516;
assign w2759 = (~pi00266 & ~w2400) | (~pi00266 & w55517) | (~w2400 & w55517);
assign w2760 = ~w1371 & ~w2561;
assign w2761 = ~w2759 & w2760;
assign w2762 = ~w2758 & ~w2761;
assign w2763 = (~w2721 & w2054) | (~w2721 & w55518) | (w2054 & w55518);
assign w2764 = ~w2462 & w2763;
assign w2765 = (pi00268 & ~w2054) | (pi00268 & w55519) | (~w2054 & w55519);
assign w2766 = ~w2724 & ~w2765;
assign w2767 = ~w2463 & w2766;
assign w2768 = (pi00269 & ~w826) | (pi00269 & w55520) | (~w826 & w55520);
assign w2769 = (w2768 & ~w54819) | (w2768 & w55521) | (~w54819 & w55521);
assign w2770 = ~w2730 & ~w2769;
assign w2771 = ~w2578 & w2770;
assign w2772 = ~w2041 & w55522;
assign w2773 = ~w2578 & w2772;
assign w2774 = (~w2727 & ~w2055) | (~w2727 & w55523) | (~w2055 & w55523);
assign w2775 = ~w2773 & w2774;
assign w2776 = ~w2276 & ~w2279;
assign w2777 = w2298 & w2776;
assign w2778 = ~pi00276 & ~w2284;
assign w2779 = ~pi00274 & w2286;
assign w2780 = w2294 & w55524;
assign w2781 = ~pi00272 & ~w2780;
assign w2782 = pi00272 & w2780;
assign w2783 = w2778 & ~w2781;
assign w2784 = ~w2782 & w2783;
assign w2785 = w2780 & w55525;
assign w2786 = w2780 & w55526;
assign w2787 = (~pi00273 & ~w2780) | (~pi00273 & w55527) | (~w2780 & w55527);
assign w2788 = w2780 & w55528;
assign w2789 = w2778 & ~w2787;
assign w2790 = ~w2788 & w2789;
assign w2791 = w2287 & w2779;
assign w2792 = ~w145 & ~w2791;
assign w2793 = (~pi00275 & ~w2780) | (~pi00275 & w55529) | (~w2780 & w55529);
assign w2794 = w2778 & ~w2786;
assign w2795 = ~w2793 & w2794;
assign w2796 = ~w2295 & w55530;
assign w2797 = w145 & ~w2796;
assign w2798 = (~pi00277 & ~w2780) | (~pi00277 & w55531) | (~w2780 & w55531);
assign w2799 = w2778 & ~w2785;
assign w2800 = ~w2798 & w2799;
assign w2801 = w1211 & w55532;
assign w2802 = w1211 & w55533;
assign w2803 = (pi00368 & ~w1209) | (pi00368 & w55534) | (~w1209 & w55534);
assign w2804 = w1211 & w55535;
assign w2805 = w1211 & w55536;
assign w2806 = ~w2801 & ~w2803;
assign w2807 = ~w2802 & ~w2804;
assign w2808 = ~w2805 & w2807;
assign w2809 = w2806 & w2808;
assign w2810 = w1211 & w55537;
assign w2811 = w1211 & w55538;
assign w2812 = (pi00367 & ~w1209) | (pi00367 & w55539) | (~w1209 & w55539);
assign w2813 = w1211 & w55540;
assign w2814 = w1211 & w55541;
assign w2815 = ~w2810 & ~w2812;
assign w2816 = ~w2811 & ~w2813;
assign w2817 = ~w2814 & w2816;
assign w2818 = w2815 & w2817;
assign w2819 = (~pi00280 & ~w826) | (~pi00280 & w55542) | (~w826 & w55542);
assign w2820 = w826 & w55543;
assign w2821 = ~w2819 & ~w2820;
assign w2822 = (~pi00281 & ~w826) | (~pi00281 & w55544) | (~w826 & w55544);
assign w2823 = w826 & w55545;
assign w2824 = ~w2822 & ~w2823;
assign w2825 = w1211 & w55546;
assign w2826 = w1211 & w55547;
assign w2827 = w1211 & w55548;
assign w2828 = (pi00369 & ~w1209) | (pi00369 & w55549) | (~w1209 & w55549);
assign w2829 = w1211 & w55550;
assign w2830 = w1211 & w55551;
assign w2831 = ~w2825 & ~w2828;
assign w2832 = ~w2826 & ~w2827;
assign w2833 = ~w2829 & ~w2830;
assign w2834 = w2832 & w2833;
assign w2835 = w2831 & w2834;
assign w2836 = w1211 & w55552;
assign w2837 = w1211 & w55553;
assign w2838 = w1211 & w55554;
assign w2839 = (pi00370 & ~w1209) | (pi00370 & w55555) | (~w1209 & w55555);
assign w2840 = w1211 & w55556;
assign w2841 = w1211 & w55557;
assign w2842 = ~w2836 & ~w2839;
assign w2843 = ~w2837 & ~w2838;
assign w2844 = ~w2840 & ~w2841;
assign w2845 = w2843 & w2844;
assign w2846 = w2842 & w2845;
assign w2847 = ~pi00284 & ~w2385;
assign w2848 = (~w1194 & ~w2385) | (~w1194 & w55558) | (~w2385 & w55558);
assign w2849 = ~w2847 & w2848;
assign w2850 = w1193 & w55559;
assign w2851 = ~w2849 & ~w2850;
assign w2852 = (~pi00285 & ~w2385) | (~pi00285 & w55560) | (~w2385 & w55560);
assign w2853 = ~w1194 & ~w2386;
assign w2854 = ~w2852 & w2853;
assign w2855 = w1193 & w55561;
assign w2856 = ~w2854 & ~w2855;
assign w2857 = (~pi00286 & ~w2385) | (~pi00286 & w55562) | (~w2385 & w55562);
assign w2858 = (~w1194 & ~w2385) | (~w1194 & w55563) | (~w2385 & w55563);
assign w2859 = ~w2857 & w2858;
assign w2860 = w1193 & w55564;
assign w2861 = ~w2859 & ~w2860;
assign w2862 = ~pi00287 & ~w2748;
assign w2863 = (~w1371 & ~w2748) | (~w1371 & w55565) | (~w2748 & w55565);
assign w2864 = ~w2862 & w2863;
assign w2865 = w826 & w55566;
assign w2866 = ~w2864 & ~w2865;
assign w2867 = ~pi00288 & ~w2400;
assign w2868 = (~w1371 & ~w2400) | (~w1371 & w55567) | (~w2400 & w55567);
assign w2869 = ~w2867 & w2868;
assign w2870 = w826 & w55568;
assign w2871 = ~w2869 & ~w2870;
assign w2872 = w826 & w55569;
assign w2873 = (~pi00289 & ~w2748) | (~pi00289 & w55570) | (~w2748 & w55570);
assign w2874 = ~w1371 & ~w2400;
assign w2875 = ~w2873 & w2874;
assign w2876 = ~w2872 & ~w2875;
assign w2877 = (~pi00290 & ~w54717) | (~pi00290 & w55571) | (~w54717 & w55571);
assign w2878 = ~w1194 & ~w2385;
assign w2879 = ~w2877 & w2878;
assign w2880 = w1193 & w55572;
assign w2881 = ~w2879 & ~w2880;
assign w2882 = ~w2042 & ~w2045;
assign w2883 = (pi00291 & w2045) | (pi00291 & w55573) | (w2045 & w55573);
assign w2884 = (~w2820 & ~w2047) | (~w2820 & w55574) | (~w2047 & w55574);
assign w2885 = ~w2883 & w2884;
assign w2886 = pi00114 & ~w2050;
assign w2887 = ~w2051 & ~w2886;
assign w2888 = (~pi00292 & ~w2045) | (~pi00292 & w55575) | (~w2045 & w55575);
assign w2889 = ~w2046 & ~w2882;
assign w2890 = ~w2888 & w2889;
assign w2891 = (~w2823 & ~w2047) | (~w2823 & w55576) | (~w2047 & w55576);
assign w2892 = ~w2890 & w2891;
assign w2893 = (~pi00293 & ~w1860) | (~pi00293 & w55577) | (~w1860 & w55577);
assign w2894 = ~w1371 & ~w2748;
assign w2895 = ~w2893 & w2894;
assign w2896 = w826 & w55578;
assign w2897 = ~w2895 & ~w2896;
assign w2898 = pi10426 & pi10458;
assign w2899 = ~pi00294 & ~w2898;
assign w2900 = ~pi00814 & pi00841;
assign w2901 = pi10435 & w1125;
assign w2902 = (~pi00320 & ~w2901) | (~pi00320 & w55579) | (~w2901 & w55579);
assign w2903 = (~w2899 & w1131) | (~w2899 & w55580) | (w1131 & w55580);
assign w2904 = ~pi10446 & ~w2903;
assign w2905 = ~pi00341 & pi09969;
assign w2906 = w852 & ~w2905;
assign w2907 = w2906 & w55581;
assign w2908 = (~pi00295 & ~w2906) | (~pi00295 & w55582) | (~w2906 & w55582);
assign w2909 = w2906 & w55583;
assign w2910 = ~pi00841 & ~w2908;
assign w2911 = ~w2909 & w2910;
assign w2912 = pi00296 & w2909;
assign w2913 = (~pi00841 & w2909) | (~pi00841 & w55584) | (w2909 & w55584);
assign w2914 = ~w2912 & w2913;
assign w2915 = (~w793 & ~w799) | (~w793 & w55585) | (~w799 & w55585);
assign w2916 = ~w727 & w799;
assign w2917 = ~w2915 & ~w2916;
assign w2918 = ~pi00402 & w2917;
assign w2919 = (w671 & w2917) | (w671 & w55586) | (w2917 & w55586);
assign w2920 = ~w2918 & w2919;
assign w2921 = w816 & w55587;
assign w2922 = w743 & ~w816;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = pi00401 & w2923;
assign w2925 = (w671 & w2923) | (w671 & w55588) | (w2923 & w55588);
assign w2926 = ~w2924 & w2925;
assign w2927 = ~pi00841 & ~pi02811;
assign w2928 = ~pi00299 & w2927;
assign w2929 = pi00233 & ~pi00240;
assign w2930 = pi00250 & w2929;
assign w2931 = (~w2928 & ~w25) | (~w2928 & w55590) | (~w25 & w55590);
assign w2932 = pi00812 & pi00886;
assign w2933 = pi10367 & pi10383;
assign w2934 = pi10427 & pi10429;
assign w2935 = pi10464 & pi10534;
assign w2936 = w2934 & w2935;
assign w2937 = w2932 & w2933;
assign w2938 = w2936 & w2937;
assign w2939 = (pi00250 & ~w2599) | (pi00250 & w55591) | (~w2599 & w55591);
assign w2940 = ~w2938 & w2939;
assign w2941 = w25 & w2940;
assign w2942 = ~w2931 & ~w2941;
assign w2943 = pi00240 & ~w78;
assign w2944 = w25 & w55592;
assign w2945 = ~pi00233 & w1074;
assign w2946 = pi00300 & w2599;
assign w2947 = w966 & w2946;
assign w2948 = ~w2945 & ~w2947;
assign w2949 = w2944 & ~w2948;
assign w2950 = w25 & w55593;
assign w2951 = w26 & w1000;
assign w2952 = w929 & w2599;
assign w2953 = w1035 & w2929;
assign w2954 = w64 & w894;
assign w2955 = ~w2952 & ~w2953;
assign w2956 = (~w2944 & ~w2955) | (~w2944 & w55594) | (~w2955 & w55594);
assign w2957 = w2927 & ~w2944;
assign w2958 = ~w2950 & w2957;
assign w2959 = (~w2956 & w55596) | (~w2956 & w55597) | (w55596 & w55597);
assign w2960 = pi00300 & ~w2959;
assign w2961 = ~w2949 & ~w2960;
assign w2962 = (~pi00301 & ~w2294) | (~pi00301 & w55598) | (~w2294 & w55598);
assign w2963 = ~w2780 & ~w2962;
assign w2964 = w2778 & w2963;
assign w2965 = pi01261 & w1232;
assign w2966 = pi09814 & w1266;
assign w2967 = pi09875 & w1235;
assign w2968 = pi10027 & w1230;
assign w2969 = pi10243 & w1244;
assign w2970 = pi09896 & w1217;
assign w2971 = pi10254 & w1242;
assign w2972 = ~w2966 & ~w2967;
assign w2973 = ~w2968 & w2972;
assign w2974 = ~w2965 & ~w2969;
assign w2975 = ~w2970 & ~w2971;
assign w2976 = w2974 & w2975;
assign w2977 = w2973 & w2976;
assign w2978 = w1211 & ~w2977;
assign w2979 = (pi00371 & ~w1209) | (pi00371 & w55599) | (~w1209 & w55599);
assign w2980 = ~w2978 & ~w2979;
assign w2981 = w1211 & w55600;
assign w2982 = pi10244 & w2317;
assign w2983 = w1211 & w55601;
assign w2984 = pi00372 & ~w1211;
assign w2985 = w1211 & w55602;
assign w2986 = pi10026 & w2321;
assign w2987 = ~w2981 & ~w2984;
assign w2988 = ~w2982 & ~w2983;
assign w2989 = ~w2985 & ~w2986;
assign w2990 = w2988 & w2989;
assign w2991 = w2987 & w2990;
assign w2992 = ~pi00304 & ~w2250;
assign w2993 = (~w1194 & ~w2250) | (~w1194 & w55603) | (~w2250 & w55603);
assign w2994 = ~w2992 & w2993;
assign w2995 = w1193 & w55604;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = w1193 & w55605;
assign w2998 = (~pi00305 & ~w2250) | (~pi00305 & w55606) | (~w2250 & w55606);
assign w2999 = ~w1194 & ~w2384;
assign w3000 = ~w2998 & w2999;
assign w3001 = ~w2997 & ~w3000;
assign w3002 = w1859 & w55607;
assign w3003 = (~pi00306 & ~w1859) | (~pi00306 & w55608) | (~w1859 & w55608);
assign w3004 = ~w1371 & ~w3002;
assign w3005 = ~w3003 & w3004;
assign w3006 = w826 & w55609;
assign w3007 = ~w3005 & ~w3006;
assign w3008 = w826 & w55610;
assign w3009 = ~pi00307 & ~w3002;
assign w3010 = (~w1371 & ~w1860) | (~w1371 & w55611) | (~w1860 & w55611);
assign w3011 = ~w3009 & w3010;
assign w3012 = ~w3008 & ~w3011;
assign w3013 = ~pi00308 & ~w2906;
assign w3014 = w1109 & w55612;
assign w3015 = (~pi00841 & ~w2906) | (~pi00841 & w55613) | (~w2906 & w55613);
assign w3016 = ~w3013 & w3015;
assign w3017 = ~w3014 & w3016;
assign w3018 = (~pi00309 & ~w2906) | (~pi00309 & w856) | (~w2906 & w856);
assign w3019 = ~pi00841 & ~w2907;
assign w3020 = ~w3018 & w3019;
assign w3021 = w2909 & w55614;
assign w3022 = (w2909 & w55615) | (w2909 & w55616) | (w55615 & w55616);
assign w3023 = ~w3021 & w3022;
assign w3024 = ~pi00311 & ~pi10468;
assign w3025 = w1131 & ~w3024;
assign w3026 = ~pi10446 & ~w3025;
assign w3027 = w1109 & w55617;
assign w3028 = ~w3027 & w55618;
assign w3029 = pi01272 & w3027;
assign w3030 = w3027 & w55619;
assign w3031 = ~w3028 & ~w3030;
assign w3032 = ~w3027 & w55620;
assign w3033 = w3027 & w55621;
assign w3034 = ~w3032 & ~w3033;
assign w3035 = ~w3027 & w55622;
assign w3036 = w3027 & w55623;
assign w3037 = ~w3035 & ~w3036;
assign w3038 = ~w3027 & w55624;
assign w3039 = w3027 & w55625;
assign w3040 = ~w3038 & ~w3039;
assign w3041 = ~w3027 & w55626;
assign w3042 = w3027 & w55627;
assign w3043 = ~w3041 & ~w3042;
assign w3044 = ~w3027 & w55628;
assign w3045 = w3027 & w55629;
assign w3046 = ~w3044 & ~w3045;
assign w3047 = ~w3027 & w55630;
assign w3048 = w3027 & w55631;
assign w3049 = ~w3047 & ~w3048;
assign w3050 = ~w3027 & w55632;
assign w3051 = ~pi10489 & w3029;
assign w3052 = ~w3050 & ~w3051;
assign w3053 = (pi00320 & ~w1125) | (pi00320 & w55633) | (~w1125 & w55633);
assign w3054 = ~w1125 & w1127;
assign w3055 = w2900 & w3054;
assign w3056 = ~w3053 & ~w3055;
assign w3057 = ~pi10446 & ~w3056;
assign w3058 = ~pi10549 & pi10551;
assign w3059 = ~pi10554 & pi10555;
assign w3060 = w3058 & w3059;
assign w3061 = pi10545 & ~pi10548;
assign w3062 = pi10544 & ~pi10557;
assign w3063 = w3061 & w3062;
assign w3064 = w3060 & w3063;
assign w3065 = pi03714 & w3064;
assign w3066 = pi10544 & pi10557;
assign w3067 = w3061 & w3066;
assign w3068 = pi10554 & ~pi10555;
assign w3069 = ~pi10549 & ~pi10551;
assign w3070 = w3068 & w3069;
assign w3071 = w3067 & w3070;
assign w3072 = pi03974 & w3071;
assign w3073 = pi10544 & pi10548;
assign w3074 = pi10545 & ~pi10557;
assign w3075 = w3073 & w3074;
assign w3076 = ~pi10554 & ~pi10555;
assign w3077 = w3069 & w3076;
assign w3078 = w3075 & w3077;
assign w3079 = pi06958 & w3078;
assign w3080 = ~pi10544 & pi10548;
assign w3081 = w3074 & w3080;
assign w3082 = w3070 & w3081;
assign w3083 = pi06897 & w3082;
assign w3084 = ~pi10545 & ~pi10557;
assign w3085 = w3080 & w3084;
assign w3086 = w3060 & w3085;
assign w3087 = pi04121 & w3086;
assign w3088 = pi10545 & pi10557;
assign w3089 = w3073 & w3088;
assign w3090 = pi10554 & pi10555;
assign w3091 = pi10549 & ~pi10551;
assign w3092 = w3090 & w3091;
assign w3093 = w3089 & w3092;
assign w3094 = pi07541 & w3093;
assign w3095 = w3073 & w3084;
assign w3096 = w3092 & w3095;
assign w3097 = pi09541 & w3096;
assign w3098 = ~pi10545 & ~pi10548;
assign w3099 = ~pi10544 & ~pi10557;
assign w3100 = w3098 & w3099;
assign w3101 = pi10549 & pi10551;
assign w3102 = w3090 & w3101;
assign w3103 = w3100 & w3102;
assign w3104 = pi03754 & w3103;
assign w3105 = w3058 & w3068;
assign w3106 = w3085 & w3105;
assign w3107 = pi07732 & w3106;
assign w3108 = w3058 & w3090;
assign w3109 = w3066 & w3098;
assign w3110 = w3108 & w3109;
assign w3111 = pi02085 & w3110;
assign w3112 = w3100 & w3105;
assign w3113 = pi09680 & w3112;
assign w3114 = w3059 & w3101;
assign w3115 = w3085 & w3114;
assign w3116 = pi04127 & w3115;
assign w3117 = w3068 & w3091;
assign w3118 = w3067 & w3117;
assign w3119 = pi03982 & w3118;
assign w3120 = ~pi10544 & pi10557;
assign w3121 = w3098 & w3120;
assign w3122 = w3108 & w3121;
assign w3123 = pi04231 & w3122;
assign w3124 = w3069 & w3090;
assign w3125 = w3089 & w3124;
assign w3126 = pi07535 & w3125;
assign w3127 = w3075 & w3108;
assign w3128 = pi07072 & w3127;
assign w3129 = w3063 & w3114;
assign w3130 = pi01671 & w3129;
assign w3131 = w3059 & w3069;
assign w3132 = w3067 & w3131;
assign w3133 = pi03956 & w3132;
assign w3134 = w3061 & w3120;
assign w3135 = w3070 & w3134;
assign w3136 = pi07157 & w3135;
assign w3137 = w3060 & w3081;
assign w3138 = pi03799 & w3137;
assign w3139 = w3075 & w3102;
assign w3140 = pi07079 & w3139;
assign w3141 = ~pi10545 & pi10557;
assign w3142 = w3080 & w3141;
assign w3143 = w3092 & w3142;
assign w3144 = pi02325 & w3143;
assign w3145 = w3059 & w3091;
assign w3146 = w3095 & w3145;
assign w3147 = pi04166 & w3146;
assign w3148 = w3121 & w3145;
assign w3149 = pi02303 & w3148;
assign w3150 = w3102 & w3109;
assign w3151 = pi08089 & w3150;
assign w3152 = w3076 & w3091;
assign w3153 = w3081 & w3152;
assign w3154 = pi09744 & w3153;
assign w3155 = w3068 & w3101;
assign w3156 = w3134 & w3155;
assign w3157 = pi09613 & w3156;
assign w3158 = w3070 & w3121;
assign w3159 = pi07962 & w3158;
assign w3160 = w3109 & w3131;
assign w3161 = pi08031 & w3160;
assign w3162 = w3109 & w3152;
assign w3163 = pi04242 & w3162;
assign w3164 = w3080 & w3088;
assign w3165 = w3145 & w3164;
assign w3166 = pi07336 & w3165;
assign w3167 = w3067 & w3102;
assign w3168 = pi07314 & w3167;
assign w3169 = w3117 & w3121;
assign w3170 = pi04212 & w3169;
assign w3171 = w3155 & w3164;
assign w3172 = pi07412 & w3171;
assign w3173 = w3085 & w3117;
assign w3174 = pi07708 & w3173;
assign w3175 = w3100 & w3131;
assign w3176 = pi07607 & w3175;
assign w3177 = w3109 & w3117;
assign w3178 = pi02468 & w3177;
assign w3179 = w3102 & w3121;
assign w3180 = pi08006 & w3179;
assign w3181 = w3070 & w3164;
assign w3182 = pi04039 & w3181;
assign w3183 = w3076 & w3101;
assign w3184 = w3109 & w3183;
assign w3185 = pi04262 & w3184;
assign w3186 = w3081 & w3155;
assign w3187 = pi06936 & w3186;
assign w3188 = w3095 & w3155;
assign w3189 = pi07851 & w3188;
assign w3190 = w3085 & w3092;
assign w3191 = pi04134 & w3190;
assign w3192 = w3089 & w3152;
assign w3193 = pi07447 & w3192;
assign w3194 = w3124 & w3164;
assign w3195 = pi07382 & w3194;
assign w3196 = w3073 & w3141;
assign w3197 = w3152 & w3196;
assign w3198 = pi03559 & w3197;
assign w3199 = w3063 & w3070;
assign w3200 = pi06818 & w3199;
assign w3201 = w3164 & w3183;
assign w3202 = pi07351 & w3201;
assign w3203 = w3100 & w3108;
assign w3204 = pi06805 & w3203;
assign w3205 = w3108 & w3134;
assign w3206 = pi07183 & w3205;
assign w3207 = w3089 & w3183;
assign w3208 = pi07485 & w3207;
assign w3209 = w3134 & w3183;
assign w3210 = pi03897 & w3209;
assign w3211 = w3105 & w3109;
assign w3212 = pi02392 & w3211;
assign w3213 = w3062 & w3098;
assign w3214 = w3108 & w3213;
assign w3215 = pi04107 & w3214;
assign w3216 = w3061 & w3099;
assign w3217 = w3152 & w3216;
assign w3218 = pi06662 & w3217;
assign w3219 = w3092 & w3100;
assign w3220 = pi06608 & w3219;
assign w3221 = w3067 & w3145;
assign w3222 = pi07224 & w3221;
assign w3223 = w3102 & w3213;
assign w3224 = pi07619 & w3223;
assign w3225 = w3067 & w3077;
assign w3226 = pi03113 & w3225;
assign w3227 = w3063 & w3155;
assign w3228 = pi06844 & w3227;
assign w3229 = w3077 & w3121;
assign w3230 = pi07880 & w3229;
assign w3231 = w3058 & w3076;
assign w3232 = w3142 & w3231;
assign w3233 = pi06484 & w3232;
assign w3234 = w3075 & w3155;
assign w3235 = pi07056 & w3234;
assign w3236 = w3063 & w3077;
assign w3237 = pi06766 & w3236;
assign w3238 = w3089 & w3105;
assign w3239 = pi07550 & w3238;
assign w3240 = w3114 & w3142;
assign w3241 = pi06491 & w3240;
assign w3242 = w3100 & w3117;
assign w3243 = pi01570 & w3242;
assign w3244 = w3075 & w3152;
assign w3245 = pi03838 & w3244;
assign w3246 = w3070 & w3100;
assign w3247 = pi08063 & w3246;
assign w3248 = w3108 & w3142;
assign w3249 = pi06539 & w3248;
assign w3250 = w3063 & w3183;
assign w3251 = pi03702 & w3250;
assign w3252 = w3114 & w3196;
assign w3253 = pi06600 & w3252;
assign w3254 = w3102 & w3134;
assign w3255 = pi07189 & w3254;
assign w3256 = w3075 & w3145;
assign w3257 = pi06975 & w3256;
assign w3258 = w3121 & w3155;
assign w3259 = pi04225 & w3258;
assign w3260 = w3081 & w3124;
assign w3261 = pi03819 & w3260;
assign w3262 = w3081 & w3114;
assign w3263 = pi03806 & w3262;
assign w3264 = w3095 & w3131;
assign w3265 = pi07773 & w3264;
assign w3266 = w3070 & w3142;
assign w3267 = pi02417 & w3266;
assign w3268 = w3117 & w3196;
assign w3269 = pi03599 & w3268;
assign w3270 = w3060 & w3089;
assign w3271 = pi07496 & w3270;
assign w3272 = w3060 & w3067;
assign w3273 = pi07246 & w3272;
assign w3274 = w3081 & w3131;
assign w3275 = pi03767 & w3274;
assign w3276 = w3067 & w3105;
assign w3277 = pi01716 & w3276;
assign w3278 = w3077 & w3213;
assign w3279 = pi06910 & w3278;
assign w3280 = w3070 & w3095;
assign w3281 = pi09564 & w3280;
assign w3282 = w3100 & w3231;
assign w3283 = pi01939 & w3282;
assign w3284 = w3081 & w3102;
assign w3285 = pi06949 & w3284;
assign w3286 = w3134 & w3231;
assign w3287 = pi02103 & w3286;
assign w3288 = w3102 & w3196;
assign w3289 = pi06648 & w3288;
assign w3290 = w3117 & w3213;
assign w3291 = pi04081 & w3290;
assign w3292 = w3081 & w3117;
assign w3293 = pi03812 & w3292;
assign w3294 = w3121 & w3231;
assign w3295 = pi07919 & w3294;
assign w3296 = w3081 & w3183;
assign w3297 = pi03791 & w3296;
assign w3298 = w3063 & w3152;
assign w3299 = pi01877 & w3298;
assign w3300 = w3075 & w3092;
assign w3301 = pi07040 & w3300;
assign w3302 = w3092 & w3121;
assign w3303 = pi04218 & w3302;
assign w3304 = w3063 & w3108;
assign w3305 = pi09788 & w3304;
assign w3306 = w3060 & w3142;
assign w3307 = pi03518 & w3306;
assign w3308 = w3142 & w3155;
assign w3309 = pi06520 & w3308;
assign w3310 = w3081 & w3108;
assign w3311 = pi03832 & w3310;
assign w3312 = w3077 & w3164;
assign w3313 = pi07321 & w3312;
assign w3314 = w3100 & w3155;
assign w3315 = pi06739 & w3314;
assign w3316 = w3121 & w3183;
assign w3317 = pi01917 & w3316;
assign w3318 = w3100 & w3183;
assign w3319 = pi04111 & w3318;
assign w3320 = w3077 & w3095;
assign w3321 = pi02284 & w3320;
assign w3322 = w3063 & w3105;
assign w3323 = pi03741 & w3322;
assign w3324 = w3060 & w3100;
assign w3325 = pi07941 & w3324;
assign w3326 = w3092 & w3213;
assign w3327 = pi04087 & w3326;
assign w3328 = w3085 & w3155;
assign w3329 = pi04140 & w3328;
assign w3330 = w3108 & w3216;
assign w3331 = pi03682 & w3330;
assign w3332 = w3060 & w3121;
assign w3333 = pi07949 & w3332;
assign w3334 = w3155 & w3213;
assign w3335 = pi04095 & w3334;
assign w3336 = w3131 & w3196;
assign w3337 = pi03568 & w3336;
assign w3338 = w3060 & w3134;
assign w3339 = pi03904 & w3338;
assign w3340 = w3131 & w3134;
assign w3341 = pi07101 & w3340;
assign w3342 = w3121 & w3131;
assign w3343 = pi07900 & w3342;
assign w3344 = w3145 & w3196;
assign w3345 = pi06569 & w3344;
assign w3346 = w3124 & w3142;
assign w3347 = pi03539 & w3346;
assign w3348 = w3117 & w3134;
assign w3349 = pi03916 & w3348;
assign w3350 = w3070 & w3075;
assign w3351 = pi03864 & w3350;
assign w3352 = w3089 & w3117;
assign w3353 = pi07522 & w3352;
assign w3354 = w3063 & w3131;
assign w3355 = pi06782 & w3354;
assign w3356 = w3145 & w3216;
assign w3357 = pi09737 & w3356;
assign w3358 = w3067 & w3124;
assign w3359 = pi07266 & w3358;
assign w3360 = w3089 & w3131;
assign w3361 = pi07457 & w3360;
assign w3362 = w3092 & w3216;
assign w3363 = pi03663 & w3362;
assign w3364 = w3092 & w3134;
assign w3365 = pi07163 & w3364;
assign w3366 = w3085 & w3183;
assign w3367 = pi07671 & w3366;
assign w3368 = w3077 & w3109;
assign w3369 = pi08023 & w3368;
assign w3370 = w3060 & w3095;
assign w3371 = pi04180 & w3370;
assign w3372 = w3060 & w3213;
assign w3373 = pi07359 & w3372;
assign w3374 = w3114 & w3164;
assign w3375 = pi07366 & w3374;
assign w3376 = w3067 & w3114;
assign w3377 = pi07254 & w3376;
assign w3378 = w3131 & w3216;
assign w3379 = pi06675 & w3378;
assign w3380 = w3117 & w3142;
assign w3381 = pi03532 & w3380;
assign w3382 = w3070 & w3089;
assign w3383 = pi07514 & w3382;
assign w3384 = w3075 & w3114;
assign w3385 = pi07011 & w3384;
assign w3386 = w3089 & w3114;
assign w3387 = pi07504 & w3386;
assign w3388 = w3070 & w3109;
assign w3389 = pi04279 & w3388;
assign w3390 = w3089 & w3145;
assign w3391 = pi07466 & w3390;
assign w3392 = w3063 & w3231;
assign w3393 = pi06795 & w3392;
assign w3394 = w3067 & w3231;
assign w3395 = pi03963 & w3394;
assign w3396 = w3092 & w3109;
assign w3397 = pi04305 & w3396;
assign w3398 = w3075 & w3105;
assign w3399 = pi07046 & w3398;
assign w3400 = w3063 & w3124;
assign w3401 = pi03734 & w3400;
assign w3402 = w3095 & w3108;
assign w3403 = pi07861 & w3402;
assign w3404 = w3155 & w3216;
assign w3405 = pi03676 & w3404;
assign w3406 = w3077 & w3134;
assign w3407 = pi07085 & w3406;
assign w3408 = w3142 & w3152;
assign w3409 = pi08109 & w3408;
assign w3410 = w3145 & w3213;
assign w3411 = pi01657 & w3410;
assign w3412 = w3095 & w3105;
assign w3413 = pi04199 & w3412;
assign w3414 = w3070 & w3216;
assign w3415 = pi06713 & w3414;
assign w3416 = w3060 & w3216;
assign w3417 = pi03643 & w3416;
assign w3418 = w3109 & w3114;
assign w3419 = pi08053 & w3418;
assign w3420 = w3100 & w3152;
assign w3421 = pi01492 & w3420;
assign w3422 = w3063 & w3092;
assign w3423 = pi06833 & w3422;
assign w3424 = w3081 & w3231;
assign w3425 = pi03781 & w3424;
assign w3426 = w3089 & w3155;
assign w3427 = pi07560 & w3426;
assign w3428 = w3164 & w3231;
assign w3429 = pi04015 & w3428;
assign w3430 = w3105 & w3164;
assign w3431 = pi07402 & w3430;
assign w3432 = w3075 & w3117;
assign w3433 = pi07024 & w3432;
assign w3434 = w3067 & w3155;
assign w3435 = pi07298 & w3434;
assign w3436 = w3100 & w3124;
assign w3437 = pi06529 & w3436;
assign w3438 = w3100 & w3114;
assign w3439 = pi08014 & w3438;
assign w3440 = w3085 & w3145;
assign w3441 = pi07652 & w3440;
assign w3442 = w3075 & w3183;
assign w3443 = pi01755 & w3442;
assign w3444 = w3085 & w3102;
assign w3445 = pi07746 & w3444;
assign w3446 = w3085 & w3152;
assign w3447 = pi07633 & w3446;
assign w3448 = w3067 & w3092;
assign w3449 = pi07275 & w3448;
assign w3450 = w3102 & w3216;
assign w3451 = pi06759 & w3450;
assign w3452 = w3092 & w3196;
assign w3453 = pi06621 & w3452;
assign w3454 = w3077 & w3089;
assign w3455 = pi04055 & w3454;
assign w3456 = w3124 & w3134;
assign w3457 = pi03926 & w3456;
assign w3458 = w3102 & w3164;
assign w3459 = pi07431 & w3458;
assign w3460 = w3216 & w3231;
assign w3461 = pi06694 & w3460;
assign w3462 = w3063 & w3102;
assign w3463 = pi06859 & w3462;
assign w3464 = w3089 & w3231;
assign w3465 = pi07476 & w3464;
assign w3466 = w3131 & w3213;
assign w3467 = pi07066 & w3466;
assign w3468 = w3070 & w3085;
assign w3469 = pi07699 & w3468;
assign w3470 = w3114 & w3216;
assign w3471 = pi03650 & w3470;
assign w3472 = w3213 & w3231;
assign w3473 = pi02652 & w3472;
assign w3474 = w3089 & w3102;
assign w3475 = pi07575 & w3474;
assign w3476 = w3108 & w3164;
assign w3477 = pi07421 & w3476;
assign w3478 = w3095 & w3152;
assign w3479 = pi02221 & w3478;
assign w3480 = w3077 & w3216;
assign w3481 = pi09758 & w3480;
assign w3482 = w3124 & w3216;
assign w3483 = pi06727 & w3482;
assign w3484 = w3085 & w3108;
assign w3485 = pi04147 & w3484;
assign w3486 = w3077 & w3100;
assign w3487 = pi02612 & w3486;
assign w3488 = w3142 & w3145;
assign w3489 = pi04330 & w3488;
assign w3490 = w3075 & w3231;
assign w3491 = pi03851 & w3490;
assign w3492 = w3183 & w3196;
assign w3493 = pi06580 & w3492;
assign w3494 = w3131 & w3164;
assign w3495 = pi04008 & w3494;
assign w3496 = w3077 & w3081;
assign w3497 = pi06870 & w3496;
assign w3498 = w3067 & w3152;
assign w3499 = pi03950 & w3498;
assign w3500 = w3070 & w3196;
assign w3501 = pi02029 & w3500;
assign w3502 = w3114 & w3213;
assign w3503 = pi04048 & w3502;
assign w3504 = w3109 & w3145;
assign w3505 = pi04251 & w3504;
assign w3506 = w3075 & w3124;
assign w3507 = pi07033 & w3506;
assign w3508 = w3067 & w3108;
assign w3509 = pi07307 & w3508;
assign w3510 = w3131 & w3142;
assign w3511 = pi01610 & w3510;
assign w3512 = w3095 & w3124;
assign w3513 = pi04192 & w3512;
assign w3514 = w3081 & w3092;
assign w3515 = pi06923 & w3514;
assign w3516 = w3089 & w3108;
assign w3517 = pi07567 & w3516;
assign w3518 = w3152 & w3213;
assign w3519 = pi06984 & w3518;
assign w3520 = w3105 & w3142;
assign w3521 = pi03551 & w3520;
assign w3522 = w3060 & w3164;
assign w3523 = pi09635 & w3522;
assign w3524 = w3109 & w3231;
assign w3525 = pi08042 & w3524;
assign w3526 = w3060 & w3075;
assign w3527 = pi03858 & w3526;
assign w3528 = w3105 & w3196;
assign w3529 = pi01665 & w3528;
assign w3530 = w3063 & w3145;
assign w3531 = pi03695 & w3530;
assign w3532 = w3124 & w3213;
assign w3533 = pi07585 & w3532;
assign w3534 = w3063 & w3117;
assign w3535 = pi03728 & w3534;
assign w3536 = w3081 & w3145;
assign w3537 = pi03773 & w3536;
assign w3538 = w3105 & w3216;
assign w3539 = pi02084 & w3538;
assign w3540 = w3117 & w3216;
assign w3541 = pi02324 & w3540;
assign w3542 = w3095 & w3114;
assign w3543 = pi07802 & w3542;
assign w3544 = w3196 & w3231;
assign w3545 = pi03578 & w3544;
assign w3546 = w3095 & w3231;
assign w3547 = pi01673 & w3546;
assign w3548 = w3075 & w3131;
assign w3549 = pi03845 & w3548;
assign w3550 = w3155 & w3196;
assign w3551 = pi06635 & w3550;
assign w3552 = w3114 & w3134;
assign w3553 = pi07130 & w3552;
assign w3554 = w3124 & w3196;
assign w3555 = pi01680 & w3554;
assign w3556 = w3060 & w3109;
assign w3557 = pi04271 & w3556;
assign w3558 = w3077 & w3142;
assign w3559 = pi01710 & w3558;
assign w3560 = w3121 & w3152;
assign w3561 = pi07890 & w3560;
assign w3562 = w3114 & w3121;
assign w3563 = pi04205 & w3562;
assign w3564 = w3095 & w3183;
assign w3565 = pi04173 & w3564;
assign w3566 = w3183 & w3213;
assign w3567 = pi07281 & w3566;
assign w3568 = w3108 & w3196;
assign w3569 = pi01499 & w3568;
assign w3570 = w3085 & w3131;
assign w3571 = pi09573 & w3570;
assign w3572 = w3134 & w3152;
assign w3573 = pi07092 & w3572;
assign w3574 = w3152 & w3164;
assign w3575 = pi04002 & w3574;
assign w3576 = w3134 & w3145;
assign w3577 = pi03890 & w3576;
assign w3578 = w3105 & w3121;
assign w3579 = pi07988 & w3578;
assign w3580 = w3095 & w3102;
assign w3581 = pi07870 & w3580;
assign w3582 = w3109 & w3155;
assign w3583 = pi04324 & w3582;
assign w3584 = w3085 & w3124;
assign w3585 = pi07719 & w3584;
assign w3586 = w3183 & w3216;
assign w3587 = pi06701 & w3586;
assign w3588 = w3109 & w3124;
assign w3589 = pi04297 & w3588;
assign w3590 = w3092 & w3164;
assign w3591 = pi07393 & w3590;
assign w3592 = w3105 & w3134;
assign w3593 = pi03937 & w3592;
assign w3594 = w3100 & w3145;
assign w3595 = pi07688 & w3594;
assign w3596 = w3070 & w3213;
assign w3597 = pi07528 & w3596;
assign w3598 = w3102 & w3142;
assign w3599 = pi06548 & w3598;
assign w3600 = w3117 & w3164;
assign w3601 = pi07373 & w3600;
assign w3602 = w3121 & w3124;
assign w3603 = pi07975 & w3602;
assign w3604 = w3077 & w3196;
assign w3605 = pi06559 & w3604;
assign w3606 = w3077 & w3085;
assign w3607 = pi07627 & w3606;
assign w3608 = w3085 & w3231;
assign w3609 = pi07661 & w3608;
assign w3610 = w3081 & w3105;
assign w3611 = pi03825 & w3610;
assign w3612 = w3060 & w3196;
assign w3613 = pi06590 & w3612;
assign w3614 = w3142 & w3183;
assign w3615 = pi03509 & w3614;
assign w3616 = w3105 & w3213;
assign w3617 = pi07600 & w3616;
assign w3618 = w3095 & w3117;
assign w3619 = pi04186 & w3618;
assign w3620 = w3067 & w3183;
assign w3621 = pi07237 & w3620;
assign w3622 = ~w3065 & ~w3072;
assign w3623 = ~w3079 & ~w3083;
assign w3624 = ~w3087 & ~w3094;
assign w3625 = ~w3097 & ~w3104;
assign w3626 = ~w3107 & ~w3111;
assign w3627 = ~w3113 & ~w3116;
assign w3628 = ~w3119 & ~w3123;
assign w3629 = ~w3126 & ~w3128;
assign w3630 = ~w3130 & ~w3133;
assign w3631 = ~w3136 & ~w3138;
assign w3632 = ~w3140 & ~w3144;
assign w3633 = ~w3147 & ~w3149;
assign w3634 = ~w3151 & ~w3154;
assign w3635 = ~w3157 & ~w3159;
assign w3636 = ~w3161 & ~w3163;
assign w3637 = ~w3166 & ~w3168;
assign w3638 = ~w3170 & ~w3172;
assign w3639 = ~w3174 & ~w3176;
assign w3640 = ~w3178 & ~w3180;
assign w3641 = ~w3182 & ~w3185;
assign w3642 = ~w3187 & ~w3189;
assign w3643 = ~w3191 & ~w3193;
assign w3644 = ~w3195 & ~w3198;
assign w3645 = ~w3200 & ~w3202;
assign w3646 = ~w3204 & ~w3206;
assign w3647 = ~w3208 & ~w3210;
assign w3648 = ~w3212 & ~w3215;
assign w3649 = ~w3218 & ~w3220;
assign w3650 = ~w3222 & ~w3224;
assign w3651 = ~w3226 & ~w3228;
assign w3652 = ~w3230 & ~w3233;
assign w3653 = ~w3235 & ~w3237;
assign w3654 = ~w3239 & ~w3241;
assign w3655 = ~w3243 & ~w3245;
assign w3656 = ~w3247 & ~w3249;
assign w3657 = ~w3251 & ~w3253;
assign w3658 = ~w3255 & ~w3257;
assign w3659 = ~w3259 & ~w3261;
assign w3660 = ~w3263 & ~w3265;
assign w3661 = ~w3267 & ~w3269;
assign w3662 = ~w3271 & ~w3273;
assign w3663 = ~w3275 & ~w3277;
assign w3664 = ~w3279 & ~w3281;
assign w3665 = ~w3283 & ~w3285;
assign w3666 = ~w3287 & ~w3289;
assign w3667 = ~w3291 & ~w3293;
assign w3668 = ~w3295 & ~w3297;
assign w3669 = ~w3299 & ~w3301;
assign w3670 = ~w3303 & ~w3305;
assign w3671 = ~w3307 & ~w3309;
assign w3672 = ~w3311 & ~w3313;
assign w3673 = ~w3315 & ~w3317;
assign w3674 = ~w3319 & ~w3321;
assign w3675 = ~w3323 & ~w3325;
assign w3676 = ~w3327 & ~w3329;
assign w3677 = ~w3331 & ~w3333;
assign w3678 = ~w3335 & ~w3337;
assign w3679 = ~w3339 & ~w3341;
assign w3680 = ~w3343 & ~w3345;
assign w3681 = ~w3347 & ~w3349;
assign w3682 = ~w3351 & ~w3353;
assign w3683 = ~w3355 & ~w3357;
assign w3684 = ~w3359 & ~w3361;
assign w3685 = ~w3363 & ~w3365;
assign w3686 = ~w3367 & ~w3369;
assign w3687 = ~w3371 & ~w3373;
assign w3688 = ~w3375 & ~w3377;
assign w3689 = ~w3379 & ~w3381;
assign w3690 = ~w3383 & ~w3385;
assign w3691 = ~w3387 & ~w3389;
assign w3692 = ~w3391 & ~w3393;
assign w3693 = ~w3395 & ~w3397;
assign w3694 = ~w3399 & ~w3401;
assign w3695 = ~w3403 & ~w3405;
assign w3696 = ~w3407 & ~w3409;
assign w3697 = ~w3411 & ~w3413;
assign w3698 = ~w3415 & ~w3417;
assign w3699 = ~w3419 & ~w3421;
assign w3700 = ~w3423 & ~w3425;
assign w3701 = ~w3427 & ~w3429;
assign w3702 = ~w3431 & ~w3433;
assign w3703 = ~w3435 & ~w3437;
assign w3704 = ~w3439 & ~w3441;
assign w3705 = ~w3443 & ~w3445;
assign w3706 = ~w3447 & ~w3449;
assign w3707 = ~w3451 & ~w3453;
assign w3708 = ~w3455 & ~w3457;
assign w3709 = ~w3459 & ~w3461;
assign w3710 = ~w3463 & ~w3465;
assign w3711 = ~w3467 & ~w3469;
assign w3712 = ~w3471 & ~w3473;
assign w3713 = ~w3475 & ~w3477;
assign w3714 = ~w3479 & ~w3481;
assign w3715 = ~w3483 & ~w3485;
assign w3716 = ~w3487 & ~w3489;
assign w3717 = ~w3491 & ~w3493;
assign w3718 = ~w3495 & ~w3497;
assign w3719 = ~w3499 & ~w3501;
assign w3720 = ~w3503 & ~w3505;
assign w3721 = ~w3507 & ~w3509;
assign w3722 = ~w3511 & ~w3513;
assign w3723 = ~w3515 & ~w3517;
assign w3724 = ~w3519 & ~w3521;
assign w3725 = ~w3523 & ~w3525;
assign w3726 = ~w3527 & ~w3529;
assign w3727 = ~w3531 & ~w3533;
assign w3728 = ~w3535 & ~w3537;
assign w3729 = ~w3539 & ~w3541;
assign w3730 = ~w3543 & ~w3545;
assign w3731 = ~w3547 & ~w3549;
assign w3732 = ~w3551 & ~w3553;
assign w3733 = ~w3555 & ~w3557;
assign w3734 = ~w3559 & ~w3561;
assign w3735 = ~w3563 & ~w3565;
assign w3736 = ~w3567 & ~w3569;
assign w3737 = ~w3571 & ~w3573;
assign w3738 = ~w3575 & ~w3577;
assign w3739 = ~w3579 & ~w3581;
assign w3740 = ~w3583 & ~w3585;
assign w3741 = ~w3587 & ~w3589;
assign w3742 = ~w3591 & ~w3593;
assign w3743 = ~w3595 & ~w3597;
assign w3744 = ~w3599 & ~w3601;
assign w3745 = ~w3603 & ~w3605;
assign w3746 = ~w3607 & ~w3609;
assign w3747 = ~w3611 & ~w3613;
assign w3748 = ~w3615 & ~w3617;
assign w3749 = ~w3619 & ~w3621;
assign w3750 = w3748 & w3749;
assign w3751 = w3746 & w3747;
assign w3752 = w3744 & w3745;
assign w3753 = w3742 & w3743;
assign w3754 = w3740 & w3741;
assign w3755 = w3738 & w3739;
assign w3756 = w3736 & w3737;
assign w3757 = w3734 & w3735;
assign w3758 = w3732 & w3733;
assign w3759 = w3730 & w3731;
assign w3760 = w3728 & w3729;
assign w3761 = w3726 & w3727;
assign w3762 = w3724 & w3725;
assign w3763 = w3722 & w3723;
assign w3764 = w3720 & w3721;
assign w3765 = w3718 & w3719;
assign w3766 = w3716 & w3717;
assign w3767 = w3714 & w3715;
assign w3768 = w3712 & w3713;
assign w3769 = w3710 & w3711;
assign w3770 = w3708 & w3709;
assign w3771 = w3706 & w3707;
assign w3772 = w3704 & w3705;
assign w3773 = w3702 & w3703;
assign w3774 = w3700 & w3701;
assign w3775 = w3698 & w3699;
assign w3776 = w3696 & w3697;
assign w3777 = w3694 & w3695;
assign w3778 = w3692 & w3693;
assign w3779 = w3690 & w3691;
assign w3780 = w3688 & w3689;
assign w3781 = w3686 & w3687;
assign w3782 = w3684 & w3685;
assign w3783 = w3682 & w3683;
assign w3784 = w3680 & w3681;
assign w3785 = w3678 & w3679;
assign w3786 = w3676 & w3677;
assign w3787 = w3674 & w3675;
assign w3788 = w3672 & w3673;
assign w3789 = w3670 & w3671;
assign w3790 = w3668 & w3669;
assign w3791 = w3666 & w3667;
assign w3792 = w3664 & w3665;
assign w3793 = w3662 & w3663;
assign w3794 = w3660 & w3661;
assign w3795 = w3658 & w3659;
assign w3796 = w3656 & w3657;
assign w3797 = w3654 & w3655;
assign w3798 = w3652 & w3653;
assign w3799 = w3650 & w3651;
assign w3800 = w3648 & w3649;
assign w3801 = w3646 & w3647;
assign w3802 = w3644 & w3645;
assign w3803 = w3642 & w3643;
assign w3804 = w3640 & w3641;
assign w3805 = w3638 & w3639;
assign w3806 = w3636 & w3637;
assign w3807 = w3634 & w3635;
assign w3808 = w3632 & w3633;
assign w3809 = w3630 & w3631;
assign w3810 = w3628 & w3629;
assign w3811 = w3626 & w3627;
assign w3812 = w3624 & w3625;
assign w3813 = w3622 & w3623;
assign w3814 = w3812 & w3813;
assign w3815 = w3810 & w3811;
assign w3816 = w3808 & w3809;
assign w3817 = w3806 & w3807;
assign w3818 = w3804 & w3805;
assign w3819 = w3802 & w3803;
assign w3820 = w3800 & w3801;
assign w3821 = w3798 & w3799;
assign w3822 = w3796 & w3797;
assign w3823 = w3794 & w3795;
assign w3824 = w3792 & w3793;
assign w3825 = w3790 & w3791;
assign w3826 = w3788 & w3789;
assign w3827 = w3786 & w3787;
assign w3828 = w3784 & w3785;
assign w3829 = w3782 & w3783;
assign w3830 = w3780 & w3781;
assign w3831 = w3778 & w3779;
assign w3832 = w3776 & w3777;
assign w3833 = w3774 & w3775;
assign w3834 = w3772 & w3773;
assign w3835 = w3770 & w3771;
assign w3836 = w3768 & w3769;
assign w3837 = w3766 & w3767;
assign w3838 = w3764 & w3765;
assign w3839 = w3762 & w3763;
assign w3840 = w3760 & w3761;
assign w3841 = w3758 & w3759;
assign w3842 = w3756 & w3757;
assign w3843 = w3754 & w3755;
assign w3844 = w3752 & w3753;
assign w3845 = w3750 & w3751;
assign w3846 = w3844 & w3845;
assign w3847 = w3842 & w3843;
assign w3848 = w3840 & w3841;
assign w3849 = w3838 & w3839;
assign w3850 = w3836 & w3837;
assign w3851 = w3834 & w3835;
assign w3852 = w3832 & w3833;
assign w3853 = w3830 & w3831;
assign w3854 = w3828 & w3829;
assign w3855 = w3826 & w3827;
assign w3856 = w3824 & w3825;
assign w3857 = w3822 & w3823;
assign w3858 = w3820 & w3821;
assign w3859 = w3818 & w3819;
assign w3860 = w3816 & w3817;
assign w3861 = w3814 & w3815;
assign w3862 = w3860 & w3861;
assign w3863 = w3858 & w3859;
assign w3864 = w3856 & w3857;
assign w3865 = w3854 & w3855;
assign w3866 = w3852 & w3853;
assign w3867 = w3850 & w3851;
assign w3868 = w3848 & w3849;
assign w3869 = w3846 & w3847;
assign w3870 = w3868 & w3869;
assign w3871 = w3866 & w3867;
assign w3872 = w3864 & w3865;
assign w3873 = w3862 & w3863;
assign w3874 = w3872 & w3873;
assign w3875 = w3870 & w3871;
assign w3876 = w3874 & w3875;
assign w3877 = ~pi10577 & ~w3876;
assign w3878 = pi09953 & pi10540;
assign w3879 = pi09823 & w3878;
assign w3880 = ~w827 & ~w1194;
assign w3881 = ~w1199 & ~w1371;
assign w3882 = ~w3879 & w3881;
assign w3883 = w3880 & w3882;
assign w3884 = w3014 & w55634;
assign w3885 = (~pi10516 & ~w3014) | (~pi10516 & w55635) | (~w3014 & w55635);
assign w3886 = (~w3014 & w55636) | (~w3014 & w55637) | (w55636 & w55637);
assign w3887 = ~w3884 & ~w3886;
assign w3888 = w3014 & w55638;
assign w3889 = (~w3014 & w55639) | (~w3014 & w55640) | (w55639 & w55640);
assign w3890 = ~w3888 & ~w3889;
assign w3891 = w3014 & w55641;
assign w3892 = (~w3014 & w55642) | (~w3014 & w55643) | (w55642 & w55643);
assign w3893 = ~w3891 & ~w3892;
assign w3894 = w3014 & w55644;
assign w3895 = (~w3014 & w55645) | (~w3014 & w55646) | (w55645 & w55646);
assign w3896 = ~w3894 & ~w3895;
assign w3897 = w3014 & w55647;
assign w3898 = (~w3014 & w55648) | (~w3014 & w55649) | (w55648 & w55649);
assign w3899 = ~w3897 & ~w3898;
assign w3900 = w3014 & w55650;
assign w3901 = (~w3014 & w55651) | (~w3014 & w55652) | (w55651 & w55652);
assign w3902 = ~w3900 & ~w3901;
assign w3903 = w3014 & w55653;
assign w3904 = (~w3014 & w55654) | (~w3014 & w55655) | (w55654 & w55655);
assign w3905 = ~w3903 & ~w3904;
assign w3906 = w3014 & w55656;
assign w3907 = (~w3014 & w55657) | (~w3014 & w55658) | (w55657 & w55658);
assign w3908 = ~w3906 & ~w3907;
assign w3909 = w3014 & w55659;
assign w3910 = (~w3014 & w55660) | (~w3014 & w55661) | (w55660 & w55661);
assign w3911 = ~w3909 & ~w3910;
assign w3912 = w3014 & w55662;
assign w3913 = (~w3014 & w55663) | (~w3014 & w55664) | (w55663 & w55664);
assign w3914 = ~w3912 & ~w3913;
assign w3915 = w3014 & w55665;
assign w3916 = (~w3014 & w55666) | (~w3014 & w55667) | (w55666 & w55667);
assign w3917 = ~w3915 & ~w3916;
assign w3918 = w3014 & w55668;
assign w3919 = (~w3014 & w55669) | (~w3014 & w55670) | (w55669 & w55670);
assign w3920 = ~w3918 & ~w3919;
assign w3921 = w3014 & w55671;
assign w3922 = (~w3014 & w55672) | (~w3014 & w55673) | (w55672 & w55673);
assign w3923 = ~w3921 & ~w3922;
assign w3924 = w3014 & w55674;
assign w3925 = (~w3014 & w55675) | (~w3014 & w55676) | (w55675 & w55676);
assign w3926 = ~w3924 & ~w3925;
assign w3927 = w3014 & w55677;
assign w3928 = (~w3014 & w55678) | (~w3014 & w55679) | (w55678 & w55679);
assign w3929 = ~w3927 & ~w3928;
assign w3930 = w3014 & w55680;
assign w3931 = ~pi00337 & w3885;
assign w3932 = ~w3930 & ~w3931;
assign w3933 = ~pi00071 & pi00173;
assign w3934 = (~pi00338 & ~w1111) | (~pi00338 & w55682) | (~w1111 & w55682);
assign w3935 = ~pi10516 & ~w3934;
assign w3936 = ~pi00341 & ~pi00814;
assign w3937 = ~pi00339 & ~w3936;
assign w3938 = pi00339 & ~pi00841;
assign w3939 = w3936 & w3938;
assign w3940 = ~w2900 & ~w3939;
assign w3941 = ~w3937 & w3940;
assign w3942 = ~pi00340 & ~w3939;
assign w3943 = (pi00340 & w3939) | (pi00340 & w55683) | (w3939 & w55683);
assign w3944 = ~w3942 & ~w3943;
assign w3945 = (~pi00341 & ~w3939) | (~pi00341 & w55684) | (~w3939 & w55684);
assign w3946 = ~w2900 & ~w3945;
assign w3947 = ~pi00342 & w2902;
assign w3948 = w2419 & ~w3947;
assign w3949 = (~pi00879 & w1141) | (~pi00879 & w55685) | (w1141 & w55685);
assign w3950 = ~w1141 & w55686;
assign w3951 = w76 & ~w3949;
assign w3952 = ~w3950 & w3951;
assign w3953 = pi06534 & w3248;
assign w3954 = pi06604 & w3219;
assign w3955 = pi04248 & w3504;
assign w3956 = pi01658 & w3199;
assign w3957 = pi03725 & w3534;
assign w3958 = pi07563 & w3516;
assign w3959 = pi03679 & w3330;
assign w3960 = pi01895 & w3236;
assign w3961 = pi07915 & w3294;
assign w3962 = pi06918 & w3514;
assign w3963 = pi07293 & w3434;
assign w3964 = pi06709 & w3414;
assign w3965 = pi07726 & w3106;
assign w3966 = pi06776 & w3354;
assign w3967 = pi07241 & w3272;
assign w3968 = pi06755 & w3450;
assign w3969 = pi04209 & w3169;
assign w3970 = pi06789 & w3392;
assign w3971 = pi07109 & w3286;
assign w3972 = pi02469 & w3584;
assign w3973 = pi07742 & w3444;
assign w3974 = pi06514 & w3308;
assign w3975 = pi03960 & w3394;
assign w3976 = pi06954 & w3078;
assign w3977 = pi04163 & w3146;
assign w3978 = pi03855 & w3526;
assign w3979 = pi01625 & w3384;
assign w3980 = pi04328 & w3488;
assign w3981 = pi04202 & w3562;
assign w3982 = pi04170 & w3564;
assign w3983 = pi02066 & w3614;
assign w3984 = pi04283 & w3177;
assign w3985 = pi03647 & w3470;
assign w3986 = pi03822 & w3610;
assign w3987 = pi03861 & w3350;
assign w3988 = pi09761 & w3496;
assign w3989 = pi06980 & w3518;
assign w3990 = pi07075 & w3139;
assign w3991 = pi07657 & w3608;
assign w3992 = pi03660 & w3362;
assign w3993 = pi03529 & w3380;
assign w3994 = pi03584 & w3500;
assign w3995 = pi03692 & w3530;
assign w3996 = pi07856 & w3402;
assign w3997 = pi09752 & w3378;
assign w3998 = pi07525 & w3596;
assign w3999 = pi04034 & w3181;
assign w4000 = pi06905 & w3278;
assign w4001 = pi03887 & w3576;
assign w4002 = pi07630 & w3446;
assign w4003 = pi07667 & w3366;
assign w4004 = pi08010 & w3438;
assign w4005 = pi04012 & w3428;
assign w4006 = pi04183 & w3618;
assign w4007 = pi03638 & w3416;
assign w4008 = pi03999 & w3574;
assign w4009 = pi01491 & w3422;
assign w4010 = pi02313 & w3143;
assign w4011 = pi04084 & w3326;
assign w4012 = pi07362 & w3374;
assign w4013 = pi01864 & w3298;
assign w4014 = pi01697 & w3129;
assign w4015 = pi07781 & w3546;
assign w4016 = pi04222 & w3258;
assign w4017 = pi03894 & w3209;
assign w4018 = pi06469 & w3486;
assign w4019 = pi07904 & w3148;
assign w4020 = pi07019 & w3432;
assign w4021 = pi07218 & w3221;
assign w4022 = pi04078 & w3290;
assign w4023 = pi01677 & w3452;
assign w4024 = pi01486 & w3344;
assign w4025 = pi03513 & w3306;
assign w4026 = pi03546 & w3520;
assign w4027 = pi07531 & w3125;
assign w4028 = pi03709 & w3064;
assign w4029 = pi07377 & w3194;
assign w4030 = pi04118 & w3086;
assign w4031 = pi03829 & w3310;
assign w4032 = pi01795 & w3492;
assign w4033 = pi09528 & w3201;
assign w4034 = pi04228 & w3122;
assign w4035 = pi02466 & w3240;
assign w4036 = pi07875 & w3229;
assign w4037 = pi04124 & w3115;
assign w4038 = pi06892 & w3082;
assign w4039 = pi07923 & w3316;
assign w4040 = pi07846 & w3188;
assign w4041 = pi03556 & w3197;
assign w4042 = pi04144 & w3484;
assign w4043 = pi03777 & w3424;
assign w4044 = pi03671 & w3404;
assign w4045 = pi03953 & w3132;
assign w4046 = pi04052 & w3454;
assign w4047 = pi08144 & w3270;
assign w4048 = pi07595 & w3616;
assign w4049 = pi07097 & w3340;
assign w4050 = pi02312 & w3436;
assign w4051 = pi07703 & w3173;
assign w4052 = pi04104 & w3214;
assign w4053 = pi03764 & w3274;
assign w4054 = pi01667 & w3528;
assign w4055 = pi09768 & w3112;
assign w4056 = pi07332 & w3165;
assign w4057 = pi02503 & w3468;
assign w4058 = pi07769 & w3264;
assign w4059 = pi04189 & w3512;
assign w4060 = pi07051 & w3234;
assign w4061 = pi07153 & w3135;
assign w4062 = pi04137 & w3328;
assign w4063 = pi04257 & w3184;
assign w4064 = pi07461 & w3390;
assign w4065 = pi02655 & w3386;
assign w4066 = pi07310 & w3167;
assign w4067 = pi04019 & w3522;
assign w4068 = pi01507 & w3348;
assign w4069 = pi01577 & w3568;
assign w4070 = pi02260 & w3538;
assign w4071 = pi07582 & w3532;
assign w4072 = pi08113 & w3510;
assign w4073 = pi07571 & w3474;
assign w4074 = pi07369 & w3600;
assign w4075 = pi04215 & w3302;
assign w4076 = pi04320 & w3582;
assign w4077 = pi01861 & w3590;
assign w4078 = pi06969 & w3256;
assign w4079 = pi07636 & w3570;
assign w4080 = pi07756 & w3478;
assign w4081 = pi07088 & w3572;
assign w4082 = pi07270 & w3448;
assign w4083 = pi09791 & w3217;
assign w4084 = pi07958 & w3158;
assign w4085 = pi06993 & w3442;
assign w4086 = pi03562 & w3336;
assign w4087 = pi02096 & w3171;
assign w4088 = pi07069 & w3127;
assign w4089 = pi07179 & w3205;
assign w4090 = pi06681 & w3356;
assign w4091 = pi03816 & w3260;
assign w4092 = pi04176 & w3370;
assign w4093 = pi07934 & w3324;
assign w4094 = pi01771 & w3612;
assign w4095 = pi07555 & w3426;
assign w4096 = pi07832 & w3318;
assign w4097 = pi07082 & w3406;
assign w4098 = pi03835 & w3244;
assign w4099 = pi07160 & w3364;
assign w4100 = pi09750 & w3153;
assign w4101 = pi06944 & w3284;
assign w4102 = pi01644 & w3360;
assign w4103 = pi06479 & w3232;
assign w4104 = pi01729 & w3458;
assign w4105 = pi04196 & w3412;
assign w4106 = pi04238 & w3162;
assign w4107 = pi07036 & w3300;
assign w4108 = pi04045 & w3502;
assign w4109 = pi03795 & w3137;
assign w4110 = pi07615 & w3223;
assign w4111 = pi07303 & w3508;
assign w4112 = pi07518 & w3352;
assign w4113 = pi08049 & w3418;
assign w4114 = pi07043 & w3398;
assign w4115 = pi09763 & w3304;
assign w4116 = pi01504 & w3288;
assign w4117 = pi07170 & w3156;
assign w4118 = pi07806 & w3280;
assign w4119 = pi07317 & w3312;
assign w4120 = pi04309 & w3211;
assign w4121 = pi09764 & w3462;
assign w4122 = pi02565 & w3586;
assign w4123 = pi08020 & w3368;
assign w4124 = pi03595 & w3268;
assign w4125 = pi08126 & w3242;
assign w4126 = pi03535 & w3346;
assign w4127 = pi02314 & w3482;
assign w4128 = pi07284 & w3276;
assign w4129 = pi02198 & w3430;
assign w4130 = pi02152 & w3376;
assign w4131 = pi07231 & w3620;
assign w4132 = pi03803 & w3262;
assign w4133 = pi01891 & w3604;
assign w4134 = pi06543 & w3598;
assign w4135 = pi03575 & w3544;
assign w4136 = pi01748 & w3203;
assign w4137 = pi09615 & w3464;
assign w4138 = pi01918 & w3282;
assign w4139 = pi04294 & w3588;
assign w4140 = pi07145 & w3420;
assign w4141 = pi03979 & w3118;
assign w4142 = pi07193 & w3225;
assign w4143 = pi07545 & w3238;
assign w4144 = pi07895 & w3342;
assign w4145 = pi07125 & w3552;
assign w4146 = pi03738 & w3322;
assign w4147 = pi07480 & w3207;
assign w4148 = pi08084 & w3150;
assign w4149 = pi07983 & w3578;
assign w4150 = pi03848 & w3490;
assign w4151 = pi07797 & w3542;
assign w4152 = pi02280 & w3320;
assign w4153 = pi03900 & w3338;
assign w4154 = pi03842 & w3548;
assign w4155 = pi07538 & w3093;
assign w4156 = pi07061 & w3466;
assign w4157 = pi04275 & w3388;
assign w4158 = pi06594 & w3252;
assign w4159 = pi07441 & w3192;
assign w4160 = pi06735 & w3314;
assign w4161 = pi02580 & w3179;
assign w4162 = pi07205 & w3472;
assign w4163 = pi04131 & w3190;
assign w4164 = pi08026 & w3160;
assign w4165 = pi03770 & w3536;
assign w4166 = pi07945 & w3332;
assign w4167 = pi07278 & w3566;
assign w4168 = pi04267 & w3556;
assign w4169 = pi07355 & w3372;
assign w4170 = pi08094 & w3558;
assign w4171 = pi04005 & w3494;
assign w4172 = pi02556 & w3382;
assign w4173 = pi06931 & w3186;
assign w4174 = pi03968 & w3071;
assign w4175 = pi07865 & w3580;
assign w4176 = pi07884 & w3560;
assign w4177 = pi08039 & w3524;
assign w4178 = pi01483 & w3227;
assign w4179 = pi08074 & w3110;
assign w4180 = pi02317 & w3540;
assign w4181 = pi08104 & w3408;
assign w4182 = pi04092 & w3334;
assign w4183 = pi07971 & w3602;
assign w4184 = pi07186 & w3254;
assign w4185 = pi07823 & w3096;
assign w4186 = pi03751 & w3103;
assign w4187 = pi06690 & w3460;
assign w4188 = pi03947 & w3498;
assign w4189 = pi03699 & w3250;
assign w4190 = pi02363 & w3266;
assign w4191 = pi07029 & w3506;
assign w4192 = pi04301 & w3396;
assign w4193 = pi07416 & w3476;
assign w4194 = pi01619 & w3550;
assign w4195 = pi01495 & w3480;
assign w4196 = pi07623 & w3606;
assign w4197 = pi03809 & w3292;
assign w4198 = pi07646 & w3440;
assign w4199 = pi09789 & w3456;
assign w4200 = pi07684 & w3594;
assign w4201 = pi03786 & w3296;
assign w4202 = pi07135 & w3410;
assign w4203 = pi03934 & w3592;
assign w4204 = pi07260 & w3358;
assign w4205 = pi03731 & w3400;
assign w4206 = pi07604 & w3175;
assign w4207 = pi01675 & w3554;
assign w4208 = pi08059 & w3246;
assign w4209 = ~w3953 & ~w3954;
assign w4210 = ~w3955 & ~w3956;
assign w4211 = ~w3957 & ~w3958;
assign w4212 = ~w3959 & ~w3960;
assign w4213 = ~w3961 & ~w3962;
assign w4214 = ~w3963 & ~w3964;
assign w4215 = ~w3965 & ~w3966;
assign w4216 = ~w3967 & ~w3968;
assign w4217 = ~w3969 & ~w3970;
assign w4218 = ~w3971 & ~w3972;
assign w4219 = ~w3973 & ~w3974;
assign w4220 = ~w3975 & ~w3976;
assign w4221 = ~w3977 & ~w3978;
assign w4222 = ~w3979 & ~w3980;
assign w4223 = ~w3981 & ~w3982;
assign w4224 = ~w3983 & ~w3984;
assign w4225 = ~w3985 & ~w3986;
assign w4226 = ~w3987 & ~w3988;
assign w4227 = ~w3989 & ~w3990;
assign w4228 = ~w3991 & ~w3992;
assign w4229 = ~w3993 & ~w3994;
assign w4230 = ~w3995 & ~w3996;
assign w4231 = ~w3997 & ~w3998;
assign w4232 = ~w3999 & ~w4000;
assign w4233 = ~w4001 & ~w4002;
assign w4234 = ~w4003 & ~w4004;
assign w4235 = ~w4005 & ~w4006;
assign w4236 = ~w4007 & ~w4008;
assign w4237 = ~w4009 & ~w4010;
assign w4238 = ~w4011 & ~w4012;
assign w4239 = ~w4013 & ~w4014;
assign w4240 = ~w4015 & ~w4016;
assign w4241 = ~w4017 & ~w4018;
assign w4242 = ~w4019 & ~w4020;
assign w4243 = ~w4021 & ~w4022;
assign w4244 = ~w4023 & ~w4024;
assign w4245 = ~w4025 & ~w4026;
assign w4246 = ~w4027 & ~w4028;
assign w4247 = ~w4029 & ~w4030;
assign w4248 = ~w4031 & ~w4032;
assign w4249 = ~w4033 & ~w4034;
assign w4250 = ~w4035 & ~w4036;
assign w4251 = ~w4037 & ~w4038;
assign w4252 = ~w4039 & ~w4040;
assign w4253 = ~w4041 & ~w4042;
assign w4254 = ~w4043 & ~w4044;
assign w4255 = ~w4045 & ~w4046;
assign w4256 = ~w4047 & ~w4048;
assign w4257 = ~w4049 & ~w4050;
assign w4258 = ~w4051 & ~w4052;
assign w4259 = ~w4053 & ~w4054;
assign w4260 = ~w4055 & ~w4056;
assign w4261 = ~w4057 & ~w4058;
assign w4262 = ~w4059 & ~w4060;
assign w4263 = ~w4061 & ~w4062;
assign w4264 = ~w4063 & ~w4064;
assign w4265 = ~w4065 & ~w4066;
assign w4266 = ~w4067 & ~w4068;
assign w4267 = ~w4069 & ~w4070;
assign w4268 = ~w4071 & ~w4072;
assign w4269 = ~w4073 & ~w4074;
assign w4270 = ~w4075 & ~w4076;
assign w4271 = ~w4077 & ~w4078;
assign w4272 = ~w4079 & ~w4080;
assign w4273 = ~w4081 & ~w4082;
assign w4274 = ~w4083 & ~w4084;
assign w4275 = ~w4085 & ~w4086;
assign w4276 = ~w4087 & ~w4088;
assign w4277 = ~w4089 & ~w4090;
assign w4278 = ~w4091 & ~w4092;
assign w4279 = ~w4093 & ~w4094;
assign w4280 = ~w4095 & ~w4096;
assign w4281 = ~w4097 & ~w4098;
assign w4282 = ~w4099 & ~w4100;
assign w4283 = ~w4101 & ~w4102;
assign w4284 = ~w4103 & ~w4104;
assign w4285 = ~w4105 & ~w4106;
assign w4286 = ~w4107 & ~w4108;
assign w4287 = ~w4109 & ~w4110;
assign w4288 = ~w4111 & ~w4112;
assign w4289 = ~w4113 & ~w4114;
assign w4290 = ~w4115 & ~w4116;
assign w4291 = ~w4117 & ~w4118;
assign w4292 = ~w4119 & ~w4120;
assign w4293 = ~w4121 & ~w4122;
assign w4294 = ~w4123 & ~w4124;
assign w4295 = ~w4125 & ~w4126;
assign w4296 = ~w4127 & ~w4128;
assign w4297 = ~w4129 & ~w4130;
assign w4298 = ~w4131 & ~w4132;
assign w4299 = ~w4133 & ~w4134;
assign w4300 = ~w4135 & ~w4136;
assign w4301 = ~w4137 & ~w4138;
assign w4302 = ~w4139 & ~w4140;
assign w4303 = ~w4141 & ~w4142;
assign w4304 = ~w4143 & ~w4144;
assign w4305 = ~w4145 & ~w4146;
assign w4306 = ~w4147 & ~w4148;
assign w4307 = ~w4149 & ~w4150;
assign w4308 = ~w4151 & ~w4152;
assign w4309 = ~w4153 & ~w4154;
assign w4310 = ~w4155 & ~w4156;
assign w4311 = ~w4157 & ~w4158;
assign w4312 = ~w4159 & ~w4160;
assign w4313 = ~w4161 & ~w4162;
assign w4314 = ~w4163 & ~w4164;
assign w4315 = ~w4165 & ~w4166;
assign w4316 = ~w4167 & ~w4168;
assign w4317 = ~w4169 & ~w4170;
assign w4318 = ~w4171 & ~w4172;
assign w4319 = ~w4173 & ~w4174;
assign w4320 = ~w4175 & ~w4176;
assign w4321 = ~w4177 & ~w4178;
assign w4322 = ~w4179 & ~w4180;
assign w4323 = ~w4181 & ~w4182;
assign w4324 = ~w4183 & ~w4184;
assign w4325 = ~w4185 & ~w4186;
assign w4326 = ~w4187 & ~w4188;
assign w4327 = ~w4189 & ~w4190;
assign w4328 = ~w4191 & ~w4192;
assign w4329 = ~w4193 & ~w4194;
assign w4330 = ~w4195 & ~w4196;
assign w4331 = ~w4197 & ~w4198;
assign w4332 = ~w4199 & ~w4200;
assign w4333 = ~w4201 & ~w4202;
assign w4334 = ~w4203 & ~w4204;
assign w4335 = ~w4205 & ~w4206;
assign w4336 = ~w4207 & ~w4208;
assign w4337 = w4335 & w4336;
assign w4338 = w4333 & w4334;
assign w4339 = w4331 & w4332;
assign w4340 = w4329 & w4330;
assign w4341 = w4327 & w4328;
assign w4342 = w4325 & w4326;
assign w4343 = w4323 & w4324;
assign w4344 = w4321 & w4322;
assign w4345 = w4319 & w4320;
assign w4346 = w4317 & w4318;
assign w4347 = w4315 & w4316;
assign w4348 = w4313 & w4314;
assign w4349 = w4311 & w4312;
assign w4350 = w4309 & w4310;
assign w4351 = w4307 & w4308;
assign w4352 = w4305 & w4306;
assign w4353 = w4303 & w4304;
assign w4354 = w4301 & w4302;
assign w4355 = w4299 & w4300;
assign w4356 = w4297 & w4298;
assign w4357 = w4295 & w4296;
assign w4358 = w4293 & w4294;
assign w4359 = w4291 & w4292;
assign w4360 = w4289 & w4290;
assign w4361 = w4287 & w4288;
assign w4362 = w4285 & w4286;
assign w4363 = w4283 & w4284;
assign w4364 = w4281 & w4282;
assign w4365 = w4279 & w4280;
assign w4366 = w4277 & w4278;
assign w4367 = w4275 & w4276;
assign w4368 = w4273 & w4274;
assign w4369 = w4271 & w4272;
assign w4370 = w4269 & w4270;
assign w4371 = w4267 & w4268;
assign w4372 = w4265 & w4266;
assign w4373 = w4263 & w4264;
assign w4374 = w4261 & w4262;
assign w4375 = w4259 & w4260;
assign w4376 = w4257 & w4258;
assign w4377 = w4255 & w4256;
assign w4378 = w4253 & w4254;
assign w4379 = w4251 & w4252;
assign w4380 = w4249 & w4250;
assign w4381 = w4247 & w4248;
assign w4382 = w4245 & w4246;
assign w4383 = w4243 & w4244;
assign w4384 = w4241 & w4242;
assign w4385 = w4239 & w4240;
assign w4386 = w4237 & w4238;
assign w4387 = w4235 & w4236;
assign w4388 = w4233 & w4234;
assign w4389 = w4231 & w4232;
assign w4390 = w4229 & w4230;
assign w4391 = w4227 & w4228;
assign w4392 = w4225 & w4226;
assign w4393 = w4223 & w4224;
assign w4394 = w4221 & w4222;
assign w4395 = w4219 & w4220;
assign w4396 = w4217 & w4218;
assign w4397 = w4215 & w4216;
assign w4398 = w4213 & w4214;
assign w4399 = w4211 & w4212;
assign w4400 = w4209 & w4210;
assign w4401 = w4399 & w4400;
assign w4402 = w4397 & w4398;
assign w4403 = w4395 & w4396;
assign w4404 = w4393 & w4394;
assign w4405 = w4391 & w4392;
assign w4406 = w4389 & w4390;
assign w4407 = w4387 & w4388;
assign w4408 = w4385 & w4386;
assign w4409 = w4383 & w4384;
assign w4410 = w4381 & w4382;
assign w4411 = w4379 & w4380;
assign w4412 = w4377 & w4378;
assign w4413 = w4375 & w4376;
assign w4414 = w4373 & w4374;
assign w4415 = w4371 & w4372;
assign w4416 = w4369 & w4370;
assign w4417 = w4367 & w4368;
assign w4418 = w4365 & w4366;
assign w4419 = w4363 & w4364;
assign w4420 = w4361 & w4362;
assign w4421 = w4359 & w4360;
assign w4422 = w4357 & w4358;
assign w4423 = w4355 & w4356;
assign w4424 = w4353 & w4354;
assign w4425 = w4351 & w4352;
assign w4426 = w4349 & w4350;
assign w4427 = w4347 & w4348;
assign w4428 = w4345 & w4346;
assign w4429 = w4343 & w4344;
assign w4430 = w4341 & w4342;
assign w4431 = w4339 & w4340;
assign w4432 = w4337 & w4338;
assign w4433 = w4431 & w4432;
assign w4434 = w4429 & w4430;
assign w4435 = w4427 & w4428;
assign w4436 = w4425 & w4426;
assign w4437 = w4423 & w4424;
assign w4438 = w4421 & w4422;
assign w4439 = w4419 & w4420;
assign w4440 = w4417 & w4418;
assign w4441 = w4415 & w4416;
assign w4442 = w4413 & w4414;
assign w4443 = w4411 & w4412;
assign w4444 = w4409 & w4410;
assign w4445 = w4407 & w4408;
assign w4446 = w4405 & w4406;
assign w4447 = w4403 & w4404;
assign w4448 = w4401 & w4402;
assign w4449 = w4447 & w4448;
assign w4450 = w4445 & w4446;
assign w4451 = w4443 & w4444;
assign w4452 = w4441 & w4442;
assign w4453 = w4439 & w4440;
assign w4454 = w4437 & w4438;
assign w4455 = w4435 & w4436;
assign w4456 = w4433 & w4434;
assign w4457 = w4455 & w4456;
assign w4458 = w4453 & w4454;
assign w4459 = w4451 & w4452;
assign w4460 = w4449 & w4450;
assign w4461 = w4459 & w4460;
assign w4462 = w4457 & w4458;
assign w4463 = w4461 & w4462;
assign w4464 = ~pi10577 & ~w4463;
assign w4465 = pi02003 & w3470;
assign w4466 = pi07624 & w3606;
assign w4467 = pi07311 & w3167;
assign w4468 = pi09523 & w3086;
assign w4469 = pi06672 & w3378;
assign w4470 = pi02346 & w3342;
assign w4471 = pi09745 & w3356;
assign w4472 = pi09649 & w3574;
assign w4473 = pi06618 & w3452;
assign w4474 = pi06666 & w3112;
assign w4475 = pi01805 & w3292;
assign w4476 = pi06724 & w3482;
assign w4477 = pi06770 & w3298;
assign w4478 = pi06855 & w3462;
assign w4479 = pi07089 & w3572;
assign w4480 = pi02764 & w3302;
assign w4481 = pi02761 & w3562;
assign w4482 = pi02615 & w3388;
assign w4483 = pi07647 & w3440;
assign w4484 = pi06906 & w3278;
assign w4485 = pi09609 & w3454;
assign w4486 = pi01964 & w3400;
assign w4487 = pi02057 & w3380;
assign w4488 = pi07356 & w3372;
assign w4489 = pi07714 & w3584;
assign w4490 = pi07695 & w3468;
assign w4491 = pi02640 & w3368;
assign w4492 = pi07318 & w3312;
assign w4493 = pi07172 & w3156;
assign w4494 = pi02771 & w3618;
assign w4495 = pi01595 & w3242;
assign w4496 = pi07426 & w3458;
assign w4497 = pi07380 & w3194;
assign w4498 = pi02768 & w3412;
assign w4499 = pi09577 & w3326;
assign w4500 = pi07206 & w3472;
assign w4501 = pi07136 & w3410;
assign w4502 = pi01811 & w3260;
assign w4503 = pi07044 & w3398;
assign w4504 = pi02319 & w3340;
assign w4505 = pi06586 & w3612;
assign w4506 = pi02777 & w3146;
assign w4507 = pi07052 & w3234;
assign w4508 = pi09608 & w3502;
assign w4509 = pi08011 & w3438;
assign w4510 = pi07154 & w3135;
assign w4511 = pi06554 & w3604;
assign w4512 = pi09544 & w3214;
assign w4513 = pi07037 & w3300;
assign w4514 = pi06566 & w3344;
assign w4515 = pi01933 & w3536;
assign w4516 = pi01760 & w3244;
assign w4517 = pi08050 & w3418;
assign w4518 = pi04259 & w3184;
assign w4519 = pi02060 & w3286;
assign w4520 = pi04239 & w3162;
assign w4521 = pi02489 & w3229;
assign w4522 = pi02294 & w3426;
assign w4523 = pi06652 & w3480;
assign w4524 = pi07972 & w3602;
assign w4525 = pi04093 & w3334;
assign w4526 = pi07251 & w3376;
assign w4527 = pi07194 & w3225;
assign w4528 = pi02393 & w3488;
assign w4529 = pi02521 & w3580;
assign w4530 = pi06736 & w3314;
assign w4531 = pi09706 & w3132;
assign w4532 = pi03913 & w3348;
assign w4533 = pi02758 & w3122;
assign w4534 = pi02333 & w3148;
assign w4535 = pi01791 & w3610;
assign w4536 = pi06470 & w3486;
assign w4537 = pi07180 & w3205;
assign w4538 = pi07834 & w3318;
assign w4539 = pi06525 & w3436;
assign w4540 = pi07959 & w3158;
assign w4541 = pi07030 & w3506;
assign w4542 = pi09682 & w3118;
assign w4543 = pi07388 & w3590;
assign w4544 = pi09584 & w3290;
assign w4545 = pi01800 & w3532;
assign w4546 = pi02781 & w3484;
assign w4547 = pi01746 & w3526;
assign w4548 = pi07482 & w3207;
assign w4549 = pi06515 & w3308;
assign w4550 = pi06639 & w3568;
assign w4551 = pi06488 & w3240;
assign w4552 = pi03787 & w3296;
assign w4553 = pi07808 & w3280;
assign w4554 = pi09647 & w3428;
assign w4555 = pi07547 & w3238;
assign w4556 = pi03922 & w3456;
assign w4557 = pi02365 & w3402;
assign w4558 = pi02784 & w3190;
assign w4559 = pi01613 & w3324;
assign w4560 = pi02505 & w3396;
assign w4561 = pi02473 & w3160;
assign w4562 = pi07304 & w3508;
assign w4563 = pi06763 & w3236;
assign w4564 = pi07161 & w3364;
assign w4565 = pi06508 & w3143;
assign w4566 = pi07418 & w3476;
assign w4567 = pi02042 & w3336;
assign w4568 = pi01736 & w3350;
assign w4569 = pi02056 & w3346;
assign w4570 = pi06659 & w3217;
assign w4571 = pi06802 & w3203;
assign w4572 = pi07824 & w3096;
assign w4573 = pi01740 & w3490;
assign w4574 = pi07279 & w3566;
assign w4575 = pi01961 & w3322;
assign w4576 = pi07285 & w3276;
assign w4577 = pi02076 & w3256;
assign w4578 = pi01831 & w3442;
assign w4579 = pi07334 & w3165;
assign w4580 = pi01521 & w3338;
assign w4581 = pi07219 & w3221;
assign w4582 = pi06867 & w3496;
assign w4583 = pi01645 & w3432;
assign w4584 = pi06718 & w3540;
assign w4585 = pi06481 & w3232;
assign w4586 = pi09644 & w3494;
assign w4587 = pi07658 & w3608;
assign w4588 = pi07511 & w3382;
assign w4589 = pi06710 & w3414;
assign w4590 = pi06612 & w3554;
assign w4591 = pi07631 & w3446;
assign w4592 = pi07472 & w3464;
assign w4593 = pi07370 & w3600;
assign w4594 = pi04035 & w3181;
assign w4595 = pi03504 & w3614;
assign w4596 = pi06829 & w3422;
assign w4597 = pi07501 & w3386;
assign w4598 = pi06495 & w3266;
assign w4599 = pi01589 & w3576;
assign w4600 = pi02400 & w3582;
assign w4601 = pi01662 & w3408;
assign w4602 = pi06815 & w3199;
assign w4603 = pi04311 & w3211;
assign w4604 = pi03515 & w3306;
assign w4605 = pi06535 & w3248;
assign w4606 = pi02620 & w3556;
assign w4607 = pi06596 & w3252;
assign w4608 = pi06791 & w3392;
assign w4609 = pi02035 & w3500;
assign w4610 = pi06756 & w3450;
assign w4611 = pi06605 & w3219;
assign w4612 = pi02038 & w3544;
assign w4613 = pi02033 & w3268;
assign w4614 = pi07444 & w3192;
assign w4615 = pi03547 & w3520;
assign w4616 = pi07848 & w3188;
assign w4617 = pi07605 & w3175;
assign w4618 = pi02775 & w3564;
assign w4619 = pi07526 & w3596;
assign w4620 = pi07685 & w3594;
assign w4621 = pi02786 & w3115;
assign w4622 = pi02782 & w3328;
assign w4623 = pi07705 & w3173;
assign w4624 = pi02288 & w3294;
assign w4625 = pi07232 & w3620;
assign w4626 = pi01835 & w3137;
assign w4627 = pi01936 & w3274;
assign w4628 = pi06625 & w3528;
assign w4629 = pi06545 & w3598;
assign w4630 = pi02282 & w3246;
assign w4631 = pi01946 & w3103;
assign w4632 = pi03672 & w3404;
assign w4633 = pi02769 & w3512;
assign w4634 = pi02757 & w3504;
assign w4635 = pi06848 & w3304;
assign w4636 = pi07146 & w3420;
assign w4637 = pi07886 & w3560;
assign w4638 = pi08095 & w3558;
assign w4639 = pi06698 & w3586;
assign w4640 = pi07782 & w3546;
assign w4641 = pi07572 & w3474;
assign w4642 = pi07407 & w3171;
assign w4643 = pi07532 & w3125;
assign w4644 = pi03778 & w3424;
assign w4645 = pi02766 & w3169;
assign w4646 = pi07985 & w3578;
assign w4647 = pi07243 & w3272;
assign w4648 = pi06874 & w3153;
assign w4649 = pi01752 & w3548;
assign w4650 = pi06744 & w3538;
assign w4651 = pi03325 & w3366;
assign w4652 = pi07295 & w3434;
assign w4653 = pi07565 & w3516;
assign w4654 = pi07076 & w3139;
assign w4655 = pi03971 & w3071;
assign w4656 = pi07750 & w3320;
assign w4657 = pi03710 & w3064;
assign w4658 = pi06841 & w3227;
assign w4659 = pi02524 & w3588;
assign w4660 = pi07262 & w3358;
assign w4661 = pi07363 & w3374;
assign w4662 = pi08001 & w3179;
assign w4663 = pi07770 & w3264;
assign w4664 = pi07925 & w3316;
assign w4665 = pi07083 & w3406;
assign w4666 = pi01637 & w3542;
assign w4667 = pi07007 & w3384;
assign w4668 = pi02414 & w3524;
assign w4669 = pi03639 & w3416;
assign w4670 = pi02763 & w3258;
assign w4671 = pi01848 & w3262;
assign w4672 = pi02044 & w3197;
assign w4673 = pi09718 & w3498;
assign w4674 = pi07763 & w3282;
assign w4675 = pi02329 & w3186;
assign w4676 = pi01929 & w3150;
assign w4677 = pi07519 & w3352;
assign w4678 = pi06577 & w3492;
assign w4679 = pi09700 & w3394;
assign w4680 = pi07491 & w3270;
assign w4681 = pi02773 & w3370;
assign w4682 = pi01884 & w3518;
assign w4683 = pi06778 & w3354;
assign w4684 = pi09729 & w3592;
assign w4685 = pi07743 & w3444;
assign w4686 = pi07539 & w3093;
assign w4687 = pi06691 & w3460;
assign w4688 = pi07187 & w3254;
assign w4689 = pi07757 & w3478;
assign w4690 = pi02090 & w3110;
assign w4691 = pi01497 & w3209;
assign w4692 = pi01987 & w3250;
assign w4693 = pi07346 & w3201;
assign w4694 = pi01988 & w3530;
assign w4695 = pi02220 & w3078;
assign w4696 = pi07638 & w3570;
assign w4697 = pi07062 & w3466;
assign w4698 = pi07398 & w3430;
assign w4699 = pi06893 & w3082;
assign w4700 = pi06809 & w3129;
assign w4701 = pi06919 & w3514;
assign w4702 = pi04285 & w3177;
assign w4703 = pi04021 & w3522;
assign w4704 = pi07452 & w3360;
assign w4705 = pi01779 & w3552;
assign w4706 = pi02001 & w3362;
assign w4707 = pi07272 & w3448;
assign w4708 = pi06645 & w3288;
assign w4709 = pi01995 & w3330;
assign w4710 = pi01968 & w3534;
assign w4711 = pi07462 & w3390;
assign w4712 = pi01701 & w3616;
assign w4713 = pi01618 & w3510;
assign w4714 = pi07070 & w3127;
assign w4715 = pi01767 & w3310;
assign w4716 = pi06632 & w3550;
assign w4717 = pi06945 & w3284;
assign w4718 = pi01616 & w3332;
assign w4719 = pi01630 & w3223;
assign w4720 = pi02433 & w3106;
assign w4721 = ~w4465 & ~w4466;
assign w4722 = ~w4467 & ~w4468;
assign w4723 = ~w4469 & ~w4470;
assign w4724 = ~w4471 & ~w4472;
assign w4725 = ~w4473 & ~w4474;
assign w4726 = ~w4475 & ~w4476;
assign w4727 = ~w4477 & ~w4478;
assign w4728 = ~w4479 & ~w4480;
assign w4729 = ~w4481 & ~w4482;
assign w4730 = ~w4483 & ~w4484;
assign w4731 = ~w4485 & ~w4486;
assign w4732 = ~w4487 & ~w4488;
assign w4733 = ~w4489 & ~w4490;
assign w4734 = ~w4491 & ~w4492;
assign w4735 = ~w4493 & ~w4494;
assign w4736 = ~w4495 & ~w4496;
assign w4737 = ~w4497 & ~w4498;
assign w4738 = ~w4499 & ~w4500;
assign w4739 = ~w4501 & ~w4502;
assign w4740 = ~w4503 & ~w4504;
assign w4741 = ~w4505 & ~w4506;
assign w4742 = ~w4507 & ~w4508;
assign w4743 = ~w4509 & ~w4510;
assign w4744 = ~w4511 & ~w4512;
assign w4745 = ~w4513 & ~w4514;
assign w4746 = ~w4515 & ~w4516;
assign w4747 = ~w4517 & ~w4518;
assign w4748 = ~w4519 & ~w4520;
assign w4749 = ~w4521 & ~w4522;
assign w4750 = ~w4523 & ~w4524;
assign w4751 = ~w4525 & ~w4526;
assign w4752 = ~w4527 & ~w4528;
assign w4753 = ~w4529 & ~w4530;
assign w4754 = ~w4531 & ~w4532;
assign w4755 = ~w4533 & ~w4534;
assign w4756 = ~w4535 & ~w4536;
assign w4757 = ~w4537 & ~w4538;
assign w4758 = ~w4539 & ~w4540;
assign w4759 = ~w4541 & ~w4542;
assign w4760 = ~w4543 & ~w4544;
assign w4761 = ~w4545 & ~w4546;
assign w4762 = ~w4547 & ~w4548;
assign w4763 = ~w4549 & ~w4550;
assign w4764 = ~w4551 & ~w4552;
assign w4765 = ~w4553 & ~w4554;
assign w4766 = ~w4555 & ~w4556;
assign w4767 = ~w4557 & ~w4558;
assign w4768 = ~w4559 & ~w4560;
assign w4769 = ~w4561 & ~w4562;
assign w4770 = ~w4563 & ~w4564;
assign w4771 = ~w4565 & ~w4566;
assign w4772 = ~w4567 & ~w4568;
assign w4773 = ~w4569 & ~w4570;
assign w4774 = ~w4571 & ~w4572;
assign w4775 = ~w4573 & ~w4574;
assign w4776 = ~w4575 & ~w4576;
assign w4777 = ~w4577 & ~w4578;
assign w4778 = ~w4579 & ~w4580;
assign w4779 = ~w4581 & ~w4582;
assign w4780 = ~w4583 & ~w4584;
assign w4781 = ~w4585 & ~w4586;
assign w4782 = ~w4587 & ~w4588;
assign w4783 = ~w4589 & ~w4590;
assign w4784 = ~w4591 & ~w4592;
assign w4785 = ~w4593 & ~w4594;
assign w4786 = ~w4595 & ~w4596;
assign w4787 = ~w4597 & ~w4598;
assign w4788 = ~w4599 & ~w4600;
assign w4789 = ~w4601 & ~w4602;
assign w4790 = ~w4603 & ~w4604;
assign w4791 = ~w4605 & ~w4606;
assign w4792 = ~w4607 & ~w4608;
assign w4793 = ~w4609 & ~w4610;
assign w4794 = ~w4611 & ~w4612;
assign w4795 = ~w4613 & ~w4614;
assign w4796 = ~w4615 & ~w4616;
assign w4797 = ~w4617 & ~w4618;
assign w4798 = ~w4619 & ~w4620;
assign w4799 = ~w4621 & ~w4622;
assign w4800 = ~w4623 & ~w4624;
assign w4801 = ~w4625 & ~w4626;
assign w4802 = ~w4627 & ~w4628;
assign w4803 = ~w4629 & ~w4630;
assign w4804 = ~w4631 & ~w4632;
assign w4805 = ~w4633 & ~w4634;
assign w4806 = ~w4635 & ~w4636;
assign w4807 = ~w4637 & ~w4638;
assign w4808 = ~w4639 & ~w4640;
assign w4809 = ~w4641 & ~w4642;
assign w4810 = ~w4643 & ~w4644;
assign w4811 = ~w4645 & ~w4646;
assign w4812 = ~w4647 & ~w4648;
assign w4813 = ~w4649 & ~w4650;
assign w4814 = ~w4651 & ~w4652;
assign w4815 = ~w4653 & ~w4654;
assign w4816 = ~w4655 & ~w4656;
assign w4817 = ~w4657 & ~w4658;
assign w4818 = ~w4659 & ~w4660;
assign w4819 = ~w4661 & ~w4662;
assign w4820 = ~w4663 & ~w4664;
assign w4821 = ~w4665 & ~w4666;
assign w4822 = ~w4667 & ~w4668;
assign w4823 = ~w4669 & ~w4670;
assign w4824 = ~w4671 & ~w4672;
assign w4825 = ~w4673 & ~w4674;
assign w4826 = ~w4675 & ~w4676;
assign w4827 = ~w4677 & ~w4678;
assign w4828 = ~w4679 & ~w4680;
assign w4829 = ~w4681 & ~w4682;
assign w4830 = ~w4683 & ~w4684;
assign w4831 = ~w4685 & ~w4686;
assign w4832 = ~w4687 & ~w4688;
assign w4833 = ~w4689 & ~w4690;
assign w4834 = ~w4691 & ~w4692;
assign w4835 = ~w4693 & ~w4694;
assign w4836 = ~w4695 & ~w4696;
assign w4837 = ~w4697 & ~w4698;
assign w4838 = ~w4699 & ~w4700;
assign w4839 = ~w4701 & ~w4702;
assign w4840 = ~w4703 & ~w4704;
assign w4841 = ~w4705 & ~w4706;
assign w4842 = ~w4707 & ~w4708;
assign w4843 = ~w4709 & ~w4710;
assign w4844 = ~w4711 & ~w4712;
assign w4845 = ~w4713 & ~w4714;
assign w4846 = ~w4715 & ~w4716;
assign w4847 = ~w4717 & ~w4718;
assign w4848 = ~w4719 & ~w4720;
assign w4849 = w4847 & w4848;
assign w4850 = w4845 & w4846;
assign w4851 = w4843 & w4844;
assign w4852 = w4841 & w4842;
assign w4853 = w4839 & w4840;
assign w4854 = w4837 & w4838;
assign w4855 = w4835 & w4836;
assign w4856 = w4833 & w4834;
assign w4857 = w4831 & w4832;
assign w4858 = w4829 & w4830;
assign w4859 = w4827 & w4828;
assign w4860 = w4825 & w4826;
assign w4861 = w4823 & w4824;
assign w4862 = w4821 & w4822;
assign w4863 = w4819 & w4820;
assign w4864 = w4817 & w4818;
assign w4865 = w4815 & w4816;
assign w4866 = w4813 & w4814;
assign w4867 = w4811 & w4812;
assign w4868 = w4809 & w4810;
assign w4869 = w4807 & w4808;
assign w4870 = w4805 & w4806;
assign w4871 = w4803 & w4804;
assign w4872 = w4801 & w4802;
assign w4873 = w4799 & w4800;
assign w4874 = w4797 & w4798;
assign w4875 = w4795 & w4796;
assign w4876 = w4793 & w4794;
assign w4877 = w4791 & w4792;
assign w4878 = w4789 & w4790;
assign w4879 = w4787 & w4788;
assign w4880 = w4785 & w4786;
assign w4881 = w4783 & w4784;
assign w4882 = w4781 & w4782;
assign w4883 = w4779 & w4780;
assign w4884 = w4777 & w4778;
assign w4885 = w4775 & w4776;
assign w4886 = w4773 & w4774;
assign w4887 = w4771 & w4772;
assign w4888 = w4769 & w4770;
assign w4889 = w4767 & w4768;
assign w4890 = w4765 & w4766;
assign w4891 = w4763 & w4764;
assign w4892 = w4761 & w4762;
assign w4893 = w4759 & w4760;
assign w4894 = w4757 & w4758;
assign w4895 = w4755 & w4756;
assign w4896 = w4753 & w4754;
assign w4897 = w4751 & w4752;
assign w4898 = w4749 & w4750;
assign w4899 = w4747 & w4748;
assign w4900 = w4745 & w4746;
assign w4901 = w4743 & w4744;
assign w4902 = w4741 & w4742;
assign w4903 = w4739 & w4740;
assign w4904 = w4737 & w4738;
assign w4905 = w4735 & w4736;
assign w4906 = w4733 & w4734;
assign w4907 = w4731 & w4732;
assign w4908 = w4729 & w4730;
assign w4909 = w4727 & w4728;
assign w4910 = w4725 & w4726;
assign w4911 = w4723 & w4724;
assign w4912 = w4721 & w4722;
assign w4913 = w4911 & w4912;
assign w4914 = w4909 & w4910;
assign w4915 = w4907 & w4908;
assign w4916 = w4905 & w4906;
assign w4917 = w4903 & w4904;
assign w4918 = w4901 & w4902;
assign w4919 = w4899 & w4900;
assign w4920 = w4897 & w4898;
assign w4921 = w4895 & w4896;
assign w4922 = w4893 & w4894;
assign w4923 = w4891 & w4892;
assign w4924 = w4889 & w4890;
assign w4925 = w4887 & w4888;
assign w4926 = w4885 & w4886;
assign w4927 = w4883 & w4884;
assign w4928 = w4881 & w4882;
assign w4929 = w4879 & w4880;
assign w4930 = w4877 & w4878;
assign w4931 = w4875 & w4876;
assign w4932 = w4873 & w4874;
assign w4933 = w4871 & w4872;
assign w4934 = w4869 & w4870;
assign w4935 = w4867 & w4868;
assign w4936 = w4865 & w4866;
assign w4937 = w4863 & w4864;
assign w4938 = w4861 & w4862;
assign w4939 = w4859 & w4860;
assign w4940 = w4857 & w4858;
assign w4941 = w4855 & w4856;
assign w4942 = w4853 & w4854;
assign w4943 = w4851 & w4852;
assign w4944 = w4849 & w4850;
assign w4945 = w4943 & w4944;
assign w4946 = w4941 & w4942;
assign w4947 = w4939 & w4940;
assign w4948 = w4937 & w4938;
assign w4949 = w4935 & w4936;
assign w4950 = w4933 & w4934;
assign w4951 = w4931 & w4932;
assign w4952 = w4929 & w4930;
assign w4953 = w4927 & w4928;
assign w4954 = w4925 & w4926;
assign w4955 = w4923 & w4924;
assign w4956 = w4921 & w4922;
assign w4957 = w4919 & w4920;
assign w4958 = w4917 & w4918;
assign w4959 = w4915 & w4916;
assign w4960 = w4913 & w4914;
assign w4961 = w4959 & w4960;
assign w4962 = w4957 & w4958;
assign w4963 = w4955 & w4956;
assign w4964 = w4953 & w4954;
assign w4965 = w4951 & w4952;
assign w4966 = w4949 & w4950;
assign w4967 = w4947 & w4948;
assign w4968 = w4945 & w4946;
assign w4969 = w4967 & w4968;
assign w4970 = w4965 & w4966;
assign w4971 = w4963 & w4964;
assign w4972 = w4961 & w4962;
assign w4973 = w4971 & w4972;
assign w4974 = w4969 & w4970;
assign w4975 = w4973 & w4974;
assign w4976 = ~pi10577 & ~w4975;
assign w4977 = pi07045 & w3398;
assign w4978 = pi03797 & w3137;
assign w4979 = pi06725 & w3482;
assign w4980 = pi04006 & w3494;
assign w4981 = pi06803 & w3203;
assign w4982 = pi07758 & w3478;
assign w4983 = pi08096 & w3558;
assign w4984 = pi06526 & w3436;
assign w4985 = pi03700 & w3250;
assign w4986 = pi07399 & w3430;
assign w4987 = pi07639 & w3570;
assign w4988 = pi04046 & w3502;
assign w4989 = pi03586 & w3500;
assign w4990 = pi07878 & w3229;
assign w4991 = pi03856 & w3526;
assign w4992 = pi07835 & w3318;
assign w4993 = pi07937 & w3324;
assign w4994 = pi06745 & w3538;
assign w4995 = pi06660 & w3217;
assign w4996 = pi03789 & w3296;
assign w4997 = pi03849 & w3490;
assign w4998 = pi07445 & w3192;
assign w4999 = pi07783 & w3546;
assign w5000 = pi07288 & w3276;
assign w5001 = pi07031 & w3506;
assign w5002 = pi02499 & w3468;
assign w5003 = pi03914 & w3348;
assign w5004 = pi07849 & w3188;
assign w5005 = pi08012 & w3438;
assign w5006 = pi06792 & w3392;
assign w5007 = pi04085 & w3326;
assign w5008 = pi07419 & w3476;
assign w5009 = pi03902 & w3338;
assign w5010 = pi06606 & w3219;
assign w5011 = pi06868 & w3496;
assign w5012 = pi08076 & w3110;
assign w5013 = pi07906 & w3148;
assign w5014 = pi06653 & w3480;
assign w5015 = pi06673 & w3378;
assign w5016 = pi07502 & w3386;
assign w5017 = pi07533 & w3125;
assign w5018 = pi04269 & w3556;
assign w5019 = pi07428 & w3458;
assign w5020 = pi03516 & w3306;
assign w5021 = pi06619 & w3452;
assign w5022 = pi04164 & w3146;
assign w5023 = pi03961 & w3394;
assign w5024 = pi07409 & w3171;
assign w5025 = pi04178 & w3370;
assign w5026 = pi03530 & w3380;
assign w5027 = pi04132 & w3190;
assign w5028 = pi04119 & w3086;
assign w5029 = pi06613 & w3554;
assign w5030 = pi07022 & w3432;
assign w5031 = pi03549 & w3520;
assign w5032 = pi06946 & w3284;
assign w5033 = pi07744 & w3444;
assign w5034 = pi06849 & w3304;
assign w5035 = pi06667 & w3112;
assign w5036 = pi04053 & w3454;
assign w5037 = pi04210 & w3169;
assign w5038 = pi03680 & w3330;
assign w5039 = pi04240 & w3162;
assign w5040 = pi03732 & w3400;
assign w5041 = pi03576 & w3544;
assign w5042 = pi06633 & w3550;
assign w5043 = pi04138 & w3328;
assign w5044 = pi07887 & w3560;
assign w5045 = pi04022 & w3522;
assign w5046 = pi06810 & w3129;
assign w5047 = pi04277 & w3388;
assign w5048 = pi03506 & w3614;
assign w5049 = pi03752 & w3103;
assign w5050 = pi06598 & w3252;
assign w5051 = pi03935 & w3592;
assign w5052 = pi04322 & w3582;
assign w5053 = pi03810 & w3292;
assign w5054 = pi06588 & w3612;
assign w5055 = pi07868 & w3580;
assign w5056 = pi06842 & w3227;
assign w5057 = pi07617 & w3223;
assign w5058 = pi07926 & w3316;
assign w5059 = pi07054 & w3234;
assign w5060 = pi04295 & w3588;
assign w5061 = pi06995 & w3442;
assign w5062 = pi06489 & w3240;
assign w5063 = pi02449 & w3093;
assign w5064 = pi04260 & w3184;
assign w5065 = pi06907 & w3278;
assign w5066 = pi03661 & w3362;
assign w5067 = pi06771 & w3298;
assign w5068 = pi09556 & w3165;
assign w5069 = pi07112 & w3286;
assign w5070 = pi02307 & w3314;
assign w5071 = pi07917 & w3294;
assign w5072 = pi03726 & w3534;
assign w5073 = pi06972 & w3256;
assign w5074 = pi04249 & w3504;
assign w5075 = pi06856 & w3462;
assign w5076 = pi07162 & w3364;
assign w5077 = pi07800 & w3542;
assign w5078 = pi07483 & w3207;
assign w5079 = pi03765 & w3274;
assign w5080 = pi07764 & w3282;
assign w5081 = pi03924 & w3456;
assign w5082 = pi07127 & w3552;
assign w5083 = pi04145 & w3484;
assign w5084 = pi06779 & w3354;
assign w5085 = pi03739 & w3322;
assign w5086 = pi03771 & w3536;
assign w5087 = pi09558 & w3312;
assign w5088 = pi06757 & w3450;
assign w5089 = pi06816 & w3199;
assign w5090 = pi07273 & w3448;
assign w5091 = pi06982 & w3518;
assign w5092 = pi04333 & w3488;
assign w5093 = pi07391 & w3590;
assign w5094 = pi03804 & w3262;
assign w5095 = pi03888 & w3576;
assign w5096 = pi07090 & w3572;
assign w5097 = pi04287 & w3177;
assign w5098 = pi06682 & w3356;
assign w5099 = pi07686 & w3594;
assign w5100 = pi06764 & w3236;
assign w5101 = pi02041 & w3248;
assign w5102 = pi04190 & w3512;
assign w5103 = pi08115 & w3510;
assign w5104 = pi03537 & w3346;
assign w5105 = pi02472 & w3232;
assign w5106 = pi08087 & w3150;
assign w5107 = pi01682 & w3508;
assign w5108 = pi03648 & w3470;
assign w5109 = pi04312 & w3211;
assign w5110 = pi04171 & w3564;
assign w5111 = pi07960 & w3158;
assign w5112 = pi07155 & w3135;
assign w5113 = pi07137 & w3410;
assign w5114 = pi08105 & w3408;
assign w5115 = pi07188 & w3254;
assign w5116 = pi07063 & w3466;
assign w5117 = pi06933 & w3186;
assign w5118 = pi07253 & w3376;
assign w5119 = pi02649 & w3446;
assign w5120 = pi07706 & w3173;
assign w5121 = pi04036 & w3181;
assign w5122 = pi07771 & w3264;
assign w5123 = pi06920 & w3514;
assign w5124 = pi07625 & w3606;
assign w5125 = pi06711 & w3414;
assign w5126 = pi04184 & w3618;
assign w5127 = pi06626 & w3528;
assign w5128 = pi02644 & w3486;
assign w5129 = pi07084 & w3406;
assign w5130 = pi08040 & w3524;
assign w5131 = pi03836 & w3244;
assign w5132 = pi07038 & w3300;
assign w5133 = pi07947 & w3332;
assign w5134 = pi03895 & w3209;
assign w5135 = pi03712 & w3064;
assign w5136 = pi07263 & w3358;
assign w5137 = pi07825 & w3096;
assign w5138 = pi04079 & w3290;
assign w5139 = pi08021 & w3368;
assign w5140 = pi01775 & w3566;
assign w5141 = pi07597 & w3616;
assign w5142 = pi07659 & w3608;
assign w5143 = pi07751 & w3320;
assign w5144 = pi08051 & w3418;
assign w5145 = pi08003 & w3179;
assign w5146 = pi03843 & w3548;
assign w5147 = pi06875 & w3153;
assign w5148 = pi01660 & w3175;
assign w5149 = pi06509 & w3143;
assign w5150 = pi04125 & w3115;
assign w5151 = pi07548 & w3238;
assign w5152 = pi02793 & w3372;
assign w5153 = pi07009 & w3384;
assign w5154 = pi08061 & w3246;
assign w5155 = pi06517 & w3308;
assign w5156 = pi03564 & w3336;
assign w5157 = pi07077 & w3139;
assign w5158 = pi06546 & w3598;
assign w5159 = pi03948 & w3498;
assign w5160 = pi07235 & w3620;
assign w5161 = pi07147 & w3420;
assign w5162 = pi06699 & w3586;
assign w5163 = pi02495 & w3596;
assign w5164 = pi03597 & w3268;
assign w5165 = pi04105 & w3214;
assign w5166 = pi07809 & w3280;
assign w5167 = pi07716 & w3584;
assign w5168 = pi03862 & w3350;
assign w5169 = pi07573 & w3474;
assign w5170 = pi06567 & w3344;
assign w5171 = pi06956 & w3078;
assign w5172 = pi07195 & w3225;
assign w5173 = pi02287 & w3516;
assign w5174 = pi07859 & w3402;
assign w5175 = pi07221 & w3221;
assign w5176 = pi07312 & w3167;
assign w5177 = pi04197 & w3412;
assign w5178 = pi04000 & w3574;
assign w5179 = pi07583 & w3532;
assign w5180 = pi03693 & w3530;
assign w5181 = pi02447 & w3194;
assign w5182 = pi06640 & w3568;
assign w5183 = pi04303 & w3396;
assign w5184 = pi07557 & w3426;
assign w5185 = pi06556 & w3604;
assign w5186 = pi03674 & w3404;
assign w5187 = pi08562 & w3201;
assign w5188 = pi07520 & w3352;
assign w5189 = pi03830 & w3310;
assign w5190 = pi07474 & w3464;
assign w5191 = pi06830 & w3422;
assign w5192 = pi03779 & w3424;
assign w5193 = pi07364 & w3374;
assign w5194 = pi06719 & w3540;
assign w5195 = pi07463 & w3390;
assign w5196 = pi07513 & w3382;
assign w5197 = pi04229 & w3122;
assign w5198 = pi08028 & w3160;
assign w5199 = pi07973 & w3602;
assign w5200 = pi07729 & w3106;
assign w5201 = pi03823 & w3610;
assign w5202 = pi07208 & w3472;
assign w5203 = pi08128 & w3242;
assign w5204 = pi07071 & w3127;
assign w5205 = pi03972 & w3071;
assign w5206 = pi09675 & w3156;
assign w5207 = pi03817 & w3260;
assign w5208 = pi02291 & w3272;
assign w5209 = pi02514 & w3600;
assign w5210 = pi01643 & w3434;
assign w5211 = pi03641 & w3416;
assign w5212 = pi07669 & w3366;
assign w5213 = pi07493 & w3270;
assign w5214 = pi04203 & w3562;
assign w5215 = pi07648 & w3440;
assign w5216 = pi04013 & w3428;
assign w5217 = pi07897 & w3342;
assign w5218 = pi03954 & w3132;
assign w5219 = pi07454 & w3360;
assign w5220 = pi07181 & w3205;
assign w5221 = pi07986 & w3578;
assign w5222 = pi03557 & w3197;
assign w5223 = pi04094 & w3334;
assign w5224 = pi06692 & w3460;
assign w5225 = pi06496 & w3266;
assign w5226 = pi04216 & w3302;
assign w5227 = pi07098 & w3340;
assign w5228 = pi04223 & w3258;
assign w5229 = pi06646 & w3288;
assign w5230 = pi03980 & w3118;
assign w5231 = pi06894 & w3082;
assign w5232 = pi06578 & w3492;
assign w5233 = ~w4977 & ~w4978;
assign w5234 = ~w4979 & ~w4980;
assign w5235 = ~w4981 & ~w4982;
assign w5236 = ~w4983 & ~w4984;
assign w5237 = ~w4985 & ~w4986;
assign w5238 = ~w4987 & ~w4988;
assign w5239 = ~w4989 & ~w4990;
assign w5240 = ~w4991 & ~w4992;
assign w5241 = ~w4993 & ~w4994;
assign w5242 = ~w4995 & ~w4996;
assign w5243 = ~w4997 & ~w4998;
assign w5244 = ~w4999 & ~w5000;
assign w5245 = ~w5001 & ~w5002;
assign w5246 = ~w5003 & ~w5004;
assign w5247 = ~w5005 & ~w5006;
assign w5248 = ~w5007 & ~w5008;
assign w5249 = ~w5009 & ~w5010;
assign w5250 = ~w5011 & ~w5012;
assign w5251 = ~w5013 & ~w5014;
assign w5252 = ~w5015 & ~w5016;
assign w5253 = ~w5017 & ~w5018;
assign w5254 = ~w5019 & ~w5020;
assign w5255 = ~w5021 & ~w5022;
assign w5256 = ~w5023 & ~w5024;
assign w5257 = ~w5025 & ~w5026;
assign w5258 = ~w5027 & ~w5028;
assign w5259 = ~w5029 & ~w5030;
assign w5260 = ~w5031 & ~w5032;
assign w5261 = ~w5033 & ~w5034;
assign w5262 = ~w5035 & ~w5036;
assign w5263 = ~w5037 & ~w5038;
assign w5264 = ~w5039 & ~w5040;
assign w5265 = ~w5041 & ~w5042;
assign w5266 = ~w5043 & ~w5044;
assign w5267 = ~w5045 & ~w5046;
assign w5268 = ~w5047 & ~w5048;
assign w5269 = ~w5049 & ~w5050;
assign w5270 = ~w5051 & ~w5052;
assign w5271 = ~w5053 & ~w5054;
assign w5272 = ~w5055 & ~w5056;
assign w5273 = ~w5057 & ~w5058;
assign w5274 = ~w5059 & ~w5060;
assign w5275 = ~w5061 & ~w5062;
assign w5276 = ~w5063 & ~w5064;
assign w5277 = ~w5065 & ~w5066;
assign w5278 = ~w5067 & ~w5068;
assign w5279 = ~w5069 & ~w5070;
assign w5280 = ~w5071 & ~w5072;
assign w5281 = ~w5073 & ~w5074;
assign w5282 = ~w5075 & ~w5076;
assign w5283 = ~w5077 & ~w5078;
assign w5284 = ~w5079 & ~w5080;
assign w5285 = ~w5081 & ~w5082;
assign w5286 = ~w5083 & ~w5084;
assign w5287 = ~w5085 & ~w5086;
assign w5288 = ~w5087 & ~w5088;
assign w5289 = ~w5089 & ~w5090;
assign w5290 = ~w5091 & ~w5092;
assign w5291 = ~w5093 & ~w5094;
assign w5292 = ~w5095 & ~w5096;
assign w5293 = ~w5097 & ~w5098;
assign w5294 = ~w5099 & ~w5100;
assign w5295 = ~w5101 & ~w5102;
assign w5296 = ~w5103 & ~w5104;
assign w5297 = ~w5105 & ~w5106;
assign w5298 = ~w5107 & ~w5108;
assign w5299 = ~w5109 & ~w5110;
assign w5300 = ~w5111 & ~w5112;
assign w5301 = ~w5113 & ~w5114;
assign w5302 = ~w5115 & ~w5116;
assign w5303 = ~w5117 & ~w5118;
assign w5304 = ~w5119 & ~w5120;
assign w5305 = ~w5121 & ~w5122;
assign w5306 = ~w5123 & ~w5124;
assign w5307 = ~w5125 & ~w5126;
assign w5308 = ~w5127 & ~w5128;
assign w5309 = ~w5129 & ~w5130;
assign w5310 = ~w5131 & ~w5132;
assign w5311 = ~w5133 & ~w5134;
assign w5312 = ~w5135 & ~w5136;
assign w5313 = ~w5137 & ~w5138;
assign w5314 = ~w5139 & ~w5140;
assign w5315 = ~w5141 & ~w5142;
assign w5316 = ~w5143 & ~w5144;
assign w5317 = ~w5145 & ~w5146;
assign w5318 = ~w5147 & ~w5148;
assign w5319 = ~w5149 & ~w5150;
assign w5320 = ~w5151 & ~w5152;
assign w5321 = ~w5153 & ~w5154;
assign w5322 = ~w5155 & ~w5156;
assign w5323 = ~w5157 & ~w5158;
assign w5324 = ~w5159 & ~w5160;
assign w5325 = ~w5161 & ~w5162;
assign w5326 = ~w5163 & ~w5164;
assign w5327 = ~w5165 & ~w5166;
assign w5328 = ~w5167 & ~w5168;
assign w5329 = ~w5169 & ~w5170;
assign w5330 = ~w5171 & ~w5172;
assign w5331 = ~w5173 & ~w5174;
assign w5332 = ~w5175 & ~w5176;
assign w5333 = ~w5177 & ~w5178;
assign w5334 = ~w5179 & ~w5180;
assign w5335 = ~w5181 & ~w5182;
assign w5336 = ~w5183 & ~w5184;
assign w5337 = ~w5185 & ~w5186;
assign w5338 = ~w5187 & ~w5188;
assign w5339 = ~w5189 & ~w5190;
assign w5340 = ~w5191 & ~w5192;
assign w5341 = ~w5193 & ~w5194;
assign w5342 = ~w5195 & ~w5196;
assign w5343 = ~w5197 & ~w5198;
assign w5344 = ~w5199 & ~w5200;
assign w5345 = ~w5201 & ~w5202;
assign w5346 = ~w5203 & ~w5204;
assign w5347 = ~w5205 & ~w5206;
assign w5348 = ~w5207 & ~w5208;
assign w5349 = ~w5209 & ~w5210;
assign w5350 = ~w5211 & ~w5212;
assign w5351 = ~w5213 & ~w5214;
assign w5352 = ~w5215 & ~w5216;
assign w5353 = ~w5217 & ~w5218;
assign w5354 = ~w5219 & ~w5220;
assign w5355 = ~w5221 & ~w5222;
assign w5356 = ~w5223 & ~w5224;
assign w5357 = ~w5225 & ~w5226;
assign w5358 = ~w5227 & ~w5228;
assign w5359 = ~w5229 & ~w5230;
assign w5360 = ~w5231 & ~w5232;
assign w5361 = w5359 & w5360;
assign w5362 = w5357 & w5358;
assign w5363 = w5355 & w5356;
assign w5364 = w5353 & w5354;
assign w5365 = w5351 & w5352;
assign w5366 = w5349 & w5350;
assign w5367 = w5347 & w5348;
assign w5368 = w5345 & w5346;
assign w5369 = w5343 & w5344;
assign w5370 = w5341 & w5342;
assign w5371 = w5339 & w5340;
assign w5372 = w5337 & w5338;
assign w5373 = w5335 & w5336;
assign w5374 = w5333 & w5334;
assign w5375 = w5331 & w5332;
assign w5376 = w5329 & w5330;
assign w5377 = w5327 & w5328;
assign w5378 = w5325 & w5326;
assign w5379 = w5323 & w5324;
assign w5380 = w5321 & w5322;
assign w5381 = w5319 & w5320;
assign w5382 = w5317 & w5318;
assign w5383 = w5315 & w5316;
assign w5384 = w5313 & w5314;
assign w5385 = w5311 & w5312;
assign w5386 = w5309 & w5310;
assign w5387 = w5307 & w5308;
assign w5388 = w5305 & w5306;
assign w5389 = w5303 & w5304;
assign w5390 = w5301 & w5302;
assign w5391 = w5299 & w5300;
assign w5392 = w5297 & w5298;
assign w5393 = w5295 & w5296;
assign w5394 = w5293 & w5294;
assign w5395 = w5291 & w5292;
assign w5396 = w5289 & w5290;
assign w5397 = w5287 & w5288;
assign w5398 = w5285 & w5286;
assign w5399 = w5283 & w5284;
assign w5400 = w5281 & w5282;
assign w5401 = w5279 & w5280;
assign w5402 = w5277 & w5278;
assign w5403 = w5275 & w5276;
assign w5404 = w5273 & w5274;
assign w5405 = w5271 & w5272;
assign w5406 = w5269 & w5270;
assign w5407 = w5267 & w5268;
assign w5408 = w5265 & w5266;
assign w5409 = w5263 & w5264;
assign w5410 = w5261 & w5262;
assign w5411 = w5259 & w5260;
assign w5412 = w5257 & w5258;
assign w5413 = w5255 & w5256;
assign w5414 = w5253 & w5254;
assign w5415 = w5251 & w5252;
assign w5416 = w5249 & w5250;
assign w5417 = w5247 & w5248;
assign w5418 = w5245 & w5246;
assign w5419 = w5243 & w5244;
assign w5420 = w5241 & w5242;
assign w5421 = w5239 & w5240;
assign w5422 = w5237 & w5238;
assign w5423 = w5235 & w5236;
assign w5424 = w5233 & w5234;
assign w5425 = w5423 & w5424;
assign w5426 = w5421 & w5422;
assign w5427 = w5419 & w5420;
assign w5428 = w5417 & w5418;
assign w5429 = w5415 & w5416;
assign w5430 = w5413 & w5414;
assign w5431 = w5411 & w5412;
assign w5432 = w5409 & w5410;
assign w5433 = w5407 & w5408;
assign w5434 = w5405 & w5406;
assign w5435 = w5403 & w5404;
assign w5436 = w5401 & w5402;
assign w5437 = w5399 & w5400;
assign w5438 = w5397 & w5398;
assign w5439 = w5395 & w5396;
assign w5440 = w5393 & w5394;
assign w5441 = w5391 & w5392;
assign w5442 = w5389 & w5390;
assign w5443 = w5387 & w5388;
assign w5444 = w5385 & w5386;
assign w5445 = w5383 & w5384;
assign w5446 = w5381 & w5382;
assign w5447 = w5379 & w5380;
assign w5448 = w5377 & w5378;
assign w5449 = w5375 & w5376;
assign w5450 = w5373 & w5374;
assign w5451 = w5371 & w5372;
assign w5452 = w5369 & w5370;
assign w5453 = w5367 & w5368;
assign w5454 = w5365 & w5366;
assign w5455 = w5363 & w5364;
assign w5456 = w5361 & w5362;
assign w5457 = w5455 & w5456;
assign w5458 = w5453 & w5454;
assign w5459 = w5451 & w5452;
assign w5460 = w5449 & w5450;
assign w5461 = w5447 & w5448;
assign w5462 = w5445 & w5446;
assign w5463 = w5443 & w5444;
assign w5464 = w5441 & w5442;
assign w5465 = w5439 & w5440;
assign w5466 = w5437 & w5438;
assign w5467 = w5435 & w5436;
assign w5468 = w5433 & w5434;
assign w5469 = w5431 & w5432;
assign w5470 = w5429 & w5430;
assign w5471 = w5427 & w5428;
assign w5472 = w5425 & w5426;
assign w5473 = w5471 & w5472;
assign w5474 = w5469 & w5470;
assign w5475 = w5467 & w5468;
assign w5476 = w5465 & w5466;
assign w5477 = w5463 & w5464;
assign w5478 = w5461 & w5462;
assign w5479 = w5459 & w5460;
assign w5480 = w5457 & w5458;
assign w5481 = w5479 & w5480;
assign w5482 = w5477 & w5478;
assign w5483 = w5475 & w5476;
assign w5484 = w5473 & w5474;
assign w5485 = w5483 & w5484;
assign w5486 = w5481 & w5482;
assign w5487 = w5485 & w5486;
assign w5488 = ~pi10577 & ~w5487;
assign w5489 = pi02106 & w3376;
assign w5490 = pi03907 & w3338;
assign w5491 = pi06603 & w3252;
assign w5492 = pi04175 & w3564;
assign w5493 = pi08112 & w3408;
assign w5494 = pi03921 & w3348;
assign w5495 = pi02327 & w3406;
assign w5496 = pi07014 & w3384;
assign w5497 = pi07776 & w3264;
assign w5498 = pi07666 & w3608;
assign w5499 = pi07517 & w3382;
assign w5500 = pi03698 & w3530;
assign w5501 = pi08135 & w3242;
assign w5502 = pi03808 & w3262;
assign w5503 = pi09773 & w3300;
assign w5504 = pi06798 & w3392;
assign w5505 = pi06487 & w3232;
assign w5506 = pi09760 & w3506;
assign w5507 = pi04195 & w3512;
assign w5508 = pi06562 & w3604;
assign w5509 = pi06697 & w3460;
assign w5510 = pi04130 & w3115;
assign w5511 = pi03939 & w3592;
assign w5512 = pi04319 & w3211;
assign w5513 = pi08103 & w3558;
assign w5514 = pi03666 & w3362;
assign w5515 = pi07694 & w3594;
assign w5516 = pi07376 & w3600;
assign w5517 = pi07192 & w3254;
assign w5518 = pi03959 & w3132;
assign w5519 = pi03769 & w3274;
assign w5520 = pi04201 & w3412;
assign w5521 = pi07713 & w3173;
assign w5522 = pi07096 & w3572;
assign w5523 = pi06552 & w3598;
assign w5524 = pi08025 & w3368;
assign w5525 = pi06853 & w3304;
assign w5526 = pi07060 & w3234;
assign w5527 = pi07368 & w3374;
assign w5528 = pi03571 & w3336;
assign w5529 = pi07610 & w3175;
assign w5530 = pi03602 & w3268;
assign w5531 = pi08034 & w3160;
assign w5532 = pi04004 & w3574;
assign w5533 = pi04169 & w3146;
assign w5534 = pi06611 & w3219;
assign w5535 = pi06927 & w3514;
assign w5536 = pi07789 & w3546;
assign w5537 = pi07415 & w3171;
assign w5538 = pi06671 & w3112;
assign w5539 = pi02625 & w3420;
assign w5540 = pi04051 & w3502;
assign w5541 = pi04136 & w3190;
assign w5542 = pi04083 & w3290;
assign w5543 = pi02626 & w3466;
assign w5544 = pi07361 & w3372;
assign w5545 = pi07425 & w3476;
assign w5546 = pi03893 & w3576;
assign w5547 = pi08045 & w3524;
assign w5548 = pi06808 & w3203;
assign w5549 = pi04227 & w3258;
assign w5550 = pi07049 & w3398;
assign w5551 = pi06940 & w3186;
assign w5552 = pi07250 & w3272;
assign w5553 = pi03867 & w3350;
assign w5554 = pi07434 & w3458;
assign w5555 = pi07903 & w3342;
assign w5556 = pi08019 & w3438;
assign w5557 = pi03678 & w3404;
assign w5558 = pi06785 & w3354;
assign w5559 = pi07460 & w3360;
assign w5560 = pi04208 & w3562;
assign w5561 = pi07028 & w3432;
assign w5562 = pi07944 & w3324;
assign w5563 = pi01714 & w3276;
assign w5564 = pi02249 & w3436;
assign w5565 = pi06762 & w3450;
assign w5566 = pi06680 & w3378;
assign w5567 = pi06862 & w3462;
assign w5568 = pi03834 & w3310;
assign w5569 = pi06988 & w3518;
assign w5570 = pi08121 & w3510;
assign w5571 = pi02320 & w3482;
assign w5572 = pi04300 & w3588;
assign w5573 = pi07386 & w3194;
assign w5574 = pi03828 & w3610;
assign w5575 = pi03776 & w3536;
assign w5576 = pi07544 & w3093;
assign w5577 = pi07831 & w3096;
assign w5578 = pi06478 & w3486;
assign w5579 = pi06617 & w3554;
assign w5580 = pi03685 & w3330;
assign w5581 = pi09780 & w3135;
assign w5582 = pi07471 & w3390;
assign w5583 = pi04266 & w3184;
assign w5584 = pi06638 & w3550;
assign w5585 = pi03756 & w3103;
assign w5586 = pi04057 & w3454;
assign w5587 = pi07537 & w3125;
assign w5588 = pi07735 & w3106;
assign w5589 = pi06821 & w3199;
assign w5590 = pi07768 & w3282;
assign w5591 = pi02395 & w3266;
assign w5592 = pi07406 & w3430;
assign w5593 = pi07001 & w3442;
assign w5594 = pi04221 & w3302;
assign w5595 = pi06689 & w3356;
assign w5596 = pi03717 & w3064;
assign w5597 = pi07967 & w3158;
assign w5598 = pi06913 & w3278;
assign w5599 = pi06523 & w3308;
assign w5600 = pi07118 & w3286;
assign w5601 = pi01490 & w3298;
assign w5602 = pi07166 & w3364;
assign w5603 = pi04234 & w3122;
assign w5604 = pi04253 & w3504;
assign w5605 = pi08058 & w3418;
assign w5606 = pi03730 & w3534;
assign w5607 = pi03737 & w3400;
assign w5608 = pi07656 & w3440;
assign w5609 = pi02277 & w3426;
assign w5610 = pi04017 & w3428;
assign w5611 = pi04090 & w3326;
assign w5612 = pi01502 & w3422;
assign w5613 = pi06657 & w3480;
assign w5614 = pi07702 & w3468;
assign w5615 = pi07589 & w3532;
assign w5616 = pi07277 & w3448;
assign w5617 = pi08009 & w3179;
assign w5618 = pi08066 & w3246;
assign w5619 = pi08093 & w3150;
assign w5620 = pi09618 & w3156;
assign w5621 = pi02577 & w3225;
assign w5622 = pi06814 & w3129;
assign w5623 = pi06979 & w3256;
assign w5624 = pi07309 & w3508;
assign w5625 = pi03978 & w3071;
assign w5626 = pi07396 & w3590;
assign w5627 = pi07922 & w3294;
assign w5628 = pi04282 & w3388;
assign w5629 = pi07622 & w3223;
assign w5630 = pi06749 & w3538;
assign w5631 = pi03847 & w3548;
assign w5632 = pi03561 & w3197;
assign w5633 = pi07805 & w3542;
assign w5634 = pi07530 & w3596;
assign w5635 = pi06873 & w3496;
assign w5636 = pi07755 & w3320;
assign w5637 = pi06651 & w3288;
assign w5638 = pi02523 & w3127;
assign w5639 = pi03815 & w3292;
assign w5640 = pi04109 & w3214;
assign w5641 = pi06585 & w3492;
assign w5642 = pi07815 & w3280;
assign w5643 = pi04182 & w3370;
assign w5644 = pi04188 & w3618;
assign w5645 = pi07602 & w3616;
assign w5646 = pi07105 & w3340;
assign w5647 = pi07283 & w3566;
assign w5648 = pi03534 & w3380;
assign w5649 = pi02651 & w3472;
assign w5650 = pi06630 & w3528;
assign w5651 = pi03794 & w3296;
assign w5652 = pi04044 & w3181;
assign w5653 = pi02350 & w3139;
assign w5654 = pi07554 & w3238;
assign w5655 = pi07953 & w3332;
assign w5656 = pi07980 & w3602;
assign w5657 = pi07570 & w3516;
assign w5658 = pi07933 & w3316;
assign w5659 = pi03985 & w3118;
assign w5660 = pi07722 & w3584;
assign w5661 = pi06513 & w3143;
assign w5662 = pi07749 & w3444;
assign w5663 = pi03743 & w3322;
assign w5664 = pi06962 & w3078;
assign w5665 = pi03705 & w3250;
assign w5666 = pi04143 & w3328;
assign w5667 = pi07134 & w3552;
assign w5668 = pi03512 & w3614;
assign w5669 = pi06572 & w3344;
assign w5670 = pi07675 & w3366;
assign w5671 = pi07325 & w3312;
assign w5672 = pi07841 & w3318;
assign w5673 = pi07894 & w3560;
assign w5674 = pi04247 & w3162;
assign w5675 = pi07490 & w3207;
assign w5676 = pi09587 & w3205;
assign w5677 = pi03841 & w3244;
assign w5678 = pi07914 & w3148;
assign w5679 = pi03594 & w3500;
assign w5680 = pi06542 & w3248;
assign w5681 = pi07992 & w3578;
assign w5682 = pi08083 & w3110;
assign w5683 = pi06665 & w3217;
assign w5684 = pi07500 & w3270;
assign w5685 = pi03543 & w3346;
assign w5686 = pi07341 & w3165;
assign w5687 = pi03646 & w3416;
assign w5688 = pi07144 & w3410;
assign w5689 = pi06723 & w3540;
assign w5690 = pi03952 & w3498;
assign w5691 = pi07635 & w3446;
assign w5692 = pi04029 & w3522;
assign w5693 = pi06743 & w3314;
assign w5694 = pi04332 & w3488;
assign w5695 = pi01692 & w3434;
assign w5696 = pi03785 & w3424;
assign w5697 = pi03555 & w3520;
assign w5698 = pi06624 & w3452;
assign w5699 = pi07874 & w3580;
assign w5700 = pi06847 & w3227;
assign w5701 = pi04149 & w3484;
assign w5702 = pi03522 & w3306;
assign w5703 = pi03965 & w3394;
assign w5704 = pi03860 & w3526;
assign w5705 = pi07855 & w3188;
assign w5706 = pi06902 & w3082;
assign w5707 = pi07479 & w3464;
assign w5708 = pi07577 & w3474;
assign w5709 = pi07524 & w3352;
assign w5710 = pi06593 & w3612;
assign w5711 = pi06644 & w3568;
assign w5712 = pi04100 & w3334;
assign w5713 = pi03854 & w3490;
assign w5714 = pi04011 & w3494;
assign w5715 = pi07762 & w3478;
assign w5716 = pi04214 & w3169;
assign w5717 = pi04327 & w3582;
assign w5718 = pi07629 & w3606;
assign w5719 = pi07451 & w3192;
assign w5720 = pi03581 & w3544;
assign w5721 = pi03899 & w3209;
assign w5722 = pi06494 & w3240;
assign w5723 = pi03929 & w3456;
assign w5724 = pi06704 & w3586;
assign w5725 = pi06953 & w3284;
assign w5726 = pi04587 & w3201;
assign w5727 = pi06717 & w3414;
assign w5728 = pi04274 & w3556;
assign w5729 = pi04293 & w3177;
assign w5730 = pi07316 & w3167;
assign w5731 = pi07864 & w3402;
assign w5732 = pi07883 & w3229;
assign w5733 = pi03802 & w3137;
assign w5734 = pi03821 & w3260;
assign w5735 = pi07645 & w3570;
assign w5736 = pi06769 & w3236;
assign w5737 = pi03652 & w3470;
assign w5738 = pi07510 & w3386;
assign w5739 = pi06879 & w3153;
assign w5740 = pi04308 & w3396;
assign w5741 = pi02121 & w3620;
assign w5742 = pi01832 & w3358;
assign w5743 = pi04123 & w3086;
assign w5744 = pi07227 & w3221;
assign w5745 = ~w5489 & ~w5490;
assign w5746 = ~w5491 & ~w5492;
assign w5747 = ~w5493 & ~w5494;
assign w5748 = ~w5495 & ~w5496;
assign w5749 = ~w5497 & ~w5498;
assign w5750 = ~w5499 & ~w5500;
assign w5751 = ~w5501 & ~w5502;
assign w5752 = ~w5503 & ~w5504;
assign w5753 = ~w5505 & ~w5506;
assign w5754 = ~w5507 & ~w5508;
assign w5755 = ~w5509 & ~w5510;
assign w5756 = ~w5511 & ~w5512;
assign w5757 = ~w5513 & ~w5514;
assign w5758 = ~w5515 & ~w5516;
assign w5759 = ~w5517 & ~w5518;
assign w5760 = ~w5519 & ~w5520;
assign w5761 = ~w5521 & ~w5522;
assign w5762 = ~w5523 & ~w5524;
assign w5763 = ~w5525 & ~w5526;
assign w5764 = ~w5527 & ~w5528;
assign w5765 = ~w5529 & ~w5530;
assign w5766 = ~w5531 & ~w5532;
assign w5767 = ~w5533 & ~w5534;
assign w5768 = ~w5535 & ~w5536;
assign w5769 = ~w5537 & ~w5538;
assign w5770 = ~w5539 & ~w5540;
assign w5771 = ~w5541 & ~w5542;
assign w5772 = ~w5543 & ~w5544;
assign w5773 = ~w5545 & ~w5546;
assign w5774 = ~w5547 & ~w5548;
assign w5775 = ~w5549 & ~w5550;
assign w5776 = ~w5551 & ~w5552;
assign w5777 = ~w5553 & ~w5554;
assign w5778 = ~w5555 & ~w5556;
assign w5779 = ~w5557 & ~w5558;
assign w5780 = ~w5559 & ~w5560;
assign w5781 = ~w5561 & ~w5562;
assign w5782 = ~w5563 & ~w5564;
assign w5783 = ~w5565 & ~w5566;
assign w5784 = ~w5567 & ~w5568;
assign w5785 = ~w5569 & ~w5570;
assign w5786 = ~w5571 & ~w5572;
assign w5787 = ~w5573 & ~w5574;
assign w5788 = ~w5575 & ~w5576;
assign w5789 = ~w5577 & ~w5578;
assign w5790 = ~w5579 & ~w5580;
assign w5791 = ~w5581 & ~w5582;
assign w5792 = ~w5583 & ~w5584;
assign w5793 = ~w5585 & ~w5586;
assign w5794 = ~w5587 & ~w5588;
assign w5795 = ~w5589 & ~w5590;
assign w5796 = ~w5591 & ~w5592;
assign w5797 = ~w5593 & ~w5594;
assign w5798 = ~w5595 & ~w5596;
assign w5799 = ~w5597 & ~w5598;
assign w5800 = ~w5599 & ~w5600;
assign w5801 = ~w5601 & ~w5602;
assign w5802 = ~w5603 & ~w5604;
assign w5803 = ~w5605 & ~w5606;
assign w5804 = ~w5607 & ~w5608;
assign w5805 = ~w5609 & ~w5610;
assign w5806 = ~w5611 & ~w5612;
assign w5807 = ~w5613 & ~w5614;
assign w5808 = ~w5615 & ~w5616;
assign w5809 = ~w5617 & ~w5618;
assign w5810 = ~w5619 & ~w5620;
assign w5811 = ~w5621 & ~w5622;
assign w5812 = ~w5623 & ~w5624;
assign w5813 = ~w5625 & ~w5626;
assign w5814 = ~w5627 & ~w5628;
assign w5815 = ~w5629 & ~w5630;
assign w5816 = ~w5631 & ~w5632;
assign w5817 = ~w5633 & ~w5634;
assign w5818 = ~w5635 & ~w5636;
assign w5819 = ~w5637 & ~w5638;
assign w5820 = ~w5639 & ~w5640;
assign w5821 = ~w5641 & ~w5642;
assign w5822 = ~w5643 & ~w5644;
assign w5823 = ~w5645 & ~w5646;
assign w5824 = ~w5647 & ~w5648;
assign w5825 = ~w5649 & ~w5650;
assign w5826 = ~w5651 & ~w5652;
assign w5827 = ~w5653 & ~w5654;
assign w5828 = ~w5655 & ~w5656;
assign w5829 = ~w5657 & ~w5658;
assign w5830 = ~w5659 & ~w5660;
assign w5831 = ~w5661 & ~w5662;
assign w5832 = ~w5663 & ~w5664;
assign w5833 = ~w5665 & ~w5666;
assign w5834 = ~w5667 & ~w5668;
assign w5835 = ~w5669 & ~w5670;
assign w5836 = ~w5671 & ~w5672;
assign w5837 = ~w5673 & ~w5674;
assign w5838 = ~w5675 & ~w5676;
assign w5839 = ~w5677 & ~w5678;
assign w5840 = ~w5679 & ~w5680;
assign w5841 = ~w5681 & ~w5682;
assign w5842 = ~w5683 & ~w5684;
assign w5843 = ~w5685 & ~w5686;
assign w5844 = ~w5687 & ~w5688;
assign w5845 = ~w5689 & ~w5690;
assign w5846 = ~w5691 & ~w5692;
assign w5847 = ~w5693 & ~w5694;
assign w5848 = ~w5695 & ~w5696;
assign w5849 = ~w5697 & ~w5698;
assign w5850 = ~w5699 & ~w5700;
assign w5851 = ~w5701 & ~w5702;
assign w5852 = ~w5703 & ~w5704;
assign w5853 = ~w5705 & ~w5706;
assign w5854 = ~w5707 & ~w5708;
assign w5855 = ~w5709 & ~w5710;
assign w5856 = ~w5711 & ~w5712;
assign w5857 = ~w5713 & ~w5714;
assign w5858 = ~w5715 & ~w5716;
assign w5859 = ~w5717 & ~w5718;
assign w5860 = ~w5719 & ~w5720;
assign w5861 = ~w5721 & ~w5722;
assign w5862 = ~w5723 & ~w5724;
assign w5863 = ~w5725 & ~w5726;
assign w5864 = ~w5727 & ~w5728;
assign w5865 = ~w5729 & ~w5730;
assign w5866 = ~w5731 & ~w5732;
assign w5867 = ~w5733 & ~w5734;
assign w5868 = ~w5735 & ~w5736;
assign w5869 = ~w5737 & ~w5738;
assign w5870 = ~w5739 & ~w5740;
assign w5871 = ~w5741 & ~w5742;
assign w5872 = ~w5743 & ~w5744;
assign w5873 = w5871 & w5872;
assign w5874 = w5869 & w5870;
assign w5875 = w5867 & w5868;
assign w5876 = w5865 & w5866;
assign w5877 = w5863 & w5864;
assign w5878 = w5861 & w5862;
assign w5879 = w5859 & w5860;
assign w5880 = w5857 & w5858;
assign w5881 = w5855 & w5856;
assign w5882 = w5853 & w5854;
assign w5883 = w5851 & w5852;
assign w5884 = w5849 & w5850;
assign w5885 = w5847 & w5848;
assign w5886 = w5845 & w5846;
assign w5887 = w5843 & w5844;
assign w5888 = w5841 & w5842;
assign w5889 = w5839 & w5840;
assign w5890 = w5837 & w5838;
assign w5891 = w5835 & w5836;
assign w5892 = w5833 & w5834;
assign w5893 = w5831 & w5832;
assign w5894 = w5829 & w5830;
assign w5895 = w5827 & w5828;
assign w5896 = w5825 & w5826;
assign w5897 = w5823 & w5824;
assign w5898 = w5821 & w5822;
assign w5899 = w5819 & w5820;
assign w5900 = w5817 & w5818;
assign w5901 = w5815 & w5816;
assign w5902 = w5813 & w5814;
assign w5903 = w5811 & w5812;
assign w5904 = w5809 & w5810;
assign w5905 = w5807 & w5808;
assign w5906 = w5805 & w5806;
assign w5907 = w5803 & w5804;
assign w5908 = w5801 & w5802;
assign w5909 = w5799 & w5800;
assign w5910 = w5797 & w5798;
assign w5911 = w5795 & w5796;
assign w5912 = w5793 & w5794;
assign w5913 = w5791 & w5792;
assign w5914 = w5789 & w5790;
assign w5915 = w5787 & w5788;
assign w5916 = w5785 & w5786;
assign w5917 = w5783 & w5784;
assign w5918 = w5781 & w5782;
assign w5919 = w5779 & w5780;
assign w5920 = w5777 & w5778;
assign w5921 = w5775 & w5776;
assign w5922 = w5773 & w5774;
assign w5923 = w5771 & w5772;
assign w5924 = w5769 & w5770;
assign w5925 = w5767 & w5768;
assign w5926 = w5765 & w5766;
assign w5927 = w5763 & w5764;
assign w5928 = w5761 & w5762;
assign w5929 = w5759 & w5760;
assign w5930 = w5757 & w5758;
assign w5931 = w5755 & w5756;
assign w5932 = w5753 & w5754;
assign w5933 = w5751 & w5752;
assign w5934 = w5749 & w5750;
assign w5935 = w5747 & w5748;
assign w5936 = w5745 & w5746;
assign w5937 = w5935 & w5936;
assign w5938 = w5933 & w5934;
assign w5939 = w5931 & w5932;
assign w5940 = w5929 & w5930;
assign w5941 = w5927 & w5928;
assign w5942 = w5925 & w5926;
assign w5943 = w5923 & w5924;
assign w5944 = w5921 & w5922;
assign w5945 = w5919 & w5920;
assign w5946 = w5917 & w5918;
assign w5947 = w5915 & w5916;
assign w5948 = w5913 & w5914;
assign w5949 = w5911 & w5912;
assign w5950 = w5909 & w5910;
assign w5951 = w5907 & w5908;
assign w5952 = w5905 & w5906;
assign w5953 = w5903 & w5904;
assign w5954 = w5901 & w5902;
assign w5955 = w5899 & w5900;
assign w5956 = w5897 & w5898;
assign w5957 = w5895 & w5896;
assign w5958 = w5893 & w5894;
assign w5959 = w5891 & w5892;
assign w5960 = w5889 & w5890;
assign w5961 = w5887 & w5888;
assign w5962 = w5885 & w5886;
assign w5963 = w5883 & w5884;
assign w5964 = w5881 & w5882;
assign w5965 = w5879 & w5880;
assign w5966 = w5877 & w5878;
assign w5967 = w5875 & w5876;
assign w5968 = w5873 & w5874;
assign w5969 = w5967 & w5968;
assign w5970 = w5965 & w5966;
assign w5971 = w5963 & w5964;
assign w5972 = w5961 & w5962;
assign w5973 = w5959 & w5960;
assign w5974 = w5957 & w5958;
assign w5975 = w5955 & w5956;
assign w5976 = w5953 & w5954;
assign w5977 = w5951 & w5952;
assign w5978 = w5949 & w5950;
assign w5979 = w5947 & w5948;
assign w5980 = w5945 & w5946;
assign w5981 = w5943 & w5944;
assign w5982 = w5941 & w5942;
assign w5983 = w5939 & w5940;
assign w5984 = w5937 & w5938;
assign w5985 = w5983 & w5984;
assign w5986 = w5981 & w5982;
assign w5987 = w5979 & w5980;
assign w5988 = w5977 & w5978;
assign w5989 = w5975 & w5976;
assign w5990 = w5973 & w5974;
assign w5991 = w5971 & w5972;
assign w5992 = w5969 & w5970;
assign w5993 = w5991 & w5992;
assign w5994 = w5989 & w5990;
assign w5995 = w5987 & w5988;
assign w5996 = w5985 & w5986;
assign w5997 = w5995 & w5996;
assign w5998 = w5993 & w5994;
assign w5999 = w5997 & w5998;
assign w6000 = ~pi10577 & ~w5999;
assign w6001 = w1121 & ~w2427;
assign w6002 = ~pi00320 & ~pi00814;
assign w6003 = pi01272 & pi10435;
assign w6004 = w6002 & w6003;
assign w6005 = (~w1121 & ~w6004) | (~w1121 & w55687) | (~w6004 & w55687);
assign w6006 = pi00348 & w6005;
assign w6007 = w6004 & w55688;
assign w6008 = ~w6001 & ~w6007;
assign w6009 = ~w6006 & w6008;
assign w6010 = w1109 & w55689;
assign w6011 = ~w6010 & w55690;
assign w6012 = pi01272 & w6010;
assign w6013 = w6010 & w55631;
assign w6014 = ~w6011 & ~w6013;
assign w6015 = ~w6010 & w55691;
assign w6016 = w6010 & w55621;
assign w6017 = ~w6015 & ~w6016;
assign w6018 = ~w6010 & w55692;
assign w6019 = w6010 & w55625;
assign w6020 = ~w6018 & ~w6019;
assign w6021 = ~w6010 & w55693;
assign w6022 = w6010 & w55619;
assign w6023 = ~w6021 & ~w6022;
assign w6024 = ~w6010 & w55694;
assign w6025 = w6010 & w55627;
assign w6026 = ~w6024 & ~w6025;
assign w6027 = ~w6010 & w55695;
assign w6028 = w6010 & w55623;
assign w6029 = ~w6027 & ~w6028;
assign w6030 = ~w6010 & w55696;
assign w6031 = w6010 & w55697;
assign w6032 = ~w6030 & ~w6031;
assign w6033 = ~w6010 & w55698;
assign w6034 = pi10483 & w6012;
assign w6035 = ~w6033 & ~w6034;
assign w6036 = pi01251 & pi10466;
assign w6037 = (~pi00357 & ~w1111) | (~pi00357 & w55699) | (~w1111 & w55699);
assign w6038 = ~w2448 & ~w6036;
assign w6039 = ~w6037 & w6038;
assign w6040 = ~w727 & w816;
assign w6041 = (~w793 & ~w816) | (~w793 & w55585) | (~w816 & w55585);
assign w6042 = ~w6040 & ~w6041;
assign w6043 = ~pi00463 & w6042;
assign w6044 = (w671 & w6042) | (w671 & w55700) | (w6042 & w55700);
assign w6045 = ~w6043 & w6044;
assign w6046 = (~w743 & ~w730) | (~w743 & w55701) | (~w730 & w55701);
assign w6047 = w730 & ~w742;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = ~pi00464 & w6048;
assign w6050 = (w671 & w6048) | (w671 & w55702) | (w6048 & w55702);
assign w6051 = ~w6049 & w6050;
assign w6052 = (~pi01166 & w2587) | (~pi01166 & w55703) | (w2587 & w55703);
assign w6053 = ~w2587 & w55704;
assign w6054 = w76 & ~w6052;
assign w6055 = ~w6053 & w6054;
assign w6056 = (~pi00472 & w2587) | (~pi00472 & w55705) | (w2587 & w55705);
assign w6057 = ~w2587 & w55706;
assign w6058 = w76 & ~w6056;
assign w6059 = ~w6057 & w6058;
assign w6060 = pi09726 & w3518;
assign w6061 = pi03468 & w3396;
assign w6062 = pi02636 & w3292;
assign w6063 = pi05298 & w3538;
assign w6064 = pi02807 & w3610;
assign w6065 = pi01954 & w3298;
assign w6066 = pi03026 & w3310;
assign w6067 = pi05483 & w3300;
assign w6068 = pi03375 & w3169;
assign w6069 = pi06223 & w3402;
assign w6070 = pi06136 & w3264;
assign w6071 = pi06309 & w3158;
assign w6072 = pi05180 & w3219;
assign w6073 = pi02874 & w3500;
assign w6074 = pi03132 & w3118;
assign w6075 = pi05950 & w3616;
assign w6076 = pi03146 & w3494;
assign w6077 = pi05763 & w3430;
assign w6078 = pi05509 & w3127;
assign w6079 = pi06317 & w3602;
assign w6080 = pi05359 & w3422;
assign w6081 = pi05886 & w3596;
assign w6082 = pi05515 & w3139;
assign w6083 = pi06288 & w3324;
assign w6084 = pi03331 & w3618;
assign w6085 = pi02906 & w3404;
assign w6086 = pi03251 & w3334;
assign w6087 = pi06342 & w3179;
assign w6088 = pi03110 & w3132;
assign w6089 = pi06454 & w3510;
assign w6090 = pi05606 & w3472;
assign w6091 = pi06174 & w3280;
assign w6092 = pi09732 & w3382;
assign w6093 = pi03058 & w3350;
assign w6094 = pi05743 & w3600;
assign w6095 = pi02927 & w3250;
assign w6096 = pi05462 & w3384;
assign w6097 = pi03071 & w3209;
assign w6098 = pi05548 & w3552;
assign w6099 = pi05838 & w3207;
assign w6100 = pi03158 & w3428;
assign w6101 = pi01797 & w3304;
assign w6102 = pi05213 & w3568;
assign w6103 = pi06447 & w3408;
assign w6104 = pi06269 & w3294;
assign w6105 = pi05770 & w3171;
assign w6106 = pi06213 & w3188;
assign w6107 = pi06027 & w3366;
assign w6108 = pi05278 & w3540;
assign w6109 = pi05987 & w3606;
assign w6110 = pi05931 & w3474;
assign w6111 = pi03091 & w3456;
assign w6112 = pi03398 & w3122;
assign w6113 = pi05166 & w3612;
assign w6114 = pi02638 & w3242;
assign w6115 = pi03429 & w3184;
assign w6116 = pi05400 & w3082;
assign w6117 = pi05639 & w3358;
assign w6118 = pi05271 & w3414;
assign w6119 = pi03436 & w3556;
assign w6120 = pi05574 & w3364;
assign w6121 = pi05206 & w3550;
assign w6122 = pi03383 & w3302;
assign w6123 = pi05284 & w3482;
assign w6124 = pi05718 & w3372;
assign w6125 = pi02385 & w3167;
assign w6126 = pi02946 & w3400;
assign w6127 = pi05528 & w3572;
assign w6128 = pi03476 & w3211;
assign w6129 = pi05146 & w3604;
assign w6130 = pi05808 & w3360;
assign w6131 = pi06278 & w3316;
assign w6132 = pi05710 & w3201;
assign w6133 = pi03257 & w3214;
assign w6134 = pi06395 & w3418;
assign w6135 = pi05120 & w3308;
assign w6136 = pi03462 & w3588;
assign w6137 = pi05126 & w3436;
assign w6138 = pi05908 & w3238;
assign w6139 = pi03039 & w3548;
assign w6140 = pi03012 & w3260;
assign w6141 = pi06165 & w3542;
assign w6142 = pi05193 & w3452;
assign w6143 = pi06379 & w3524;
assign w6144 = pi06117 & w3478;
assign w6145 = pi05153 & w3344;
assign w6146 = pi01817 & w3227;
assign w6147 = pi02900 & w3362;
assign w6148 = pi06039 & w3594;
assign w6149 = pi05750 & w3194;
assign w6150 = pi02835 & w3380;
assign w6151 = pi05258 & w3460;
assign w6152 = pi06149 & w3546;
assign w6153 = pi03052 & w3526;
assign w6154 = pi06297 & w3332;
assign w6155 = pi02087 & w3177;
assign w6156 = pi09572 & w3516;
assign w6157 = pi03344 & w3412;
assign w6158 = pi05535 & w3340;
assign w6159 = pi06407 & w3246;
assign w6160 = pi05692 & w3312;
assign w6161 = pi02848 & w3520;
assign w6162 = pi05942 & w3532;
assign w6163 = pi03423 & w3504;
assign w6164 = pi06330 & w3578;
assign w6165 = pi02940 & w3534;
assign w6166 = pi05757 & w3590;
assign w6167 = pi05658 & w3276;
assign w6168 = pi06048 & w3468;
assign w6169 = pi05113 & w3143;
assign w6170 = pi05600 & w3225;
assign w6171 = pi06349 & w3438;
assign w6172 = pi02828 & w3306;
assign w6173 = pi01830 & w3458;
assign w6174 = pi05311 & w3236;
assign w6175 = pi06355 & w3368;
assign w6176 = pi03309 & w3146;
assign w6177 = pi02406 & w3508;
assign w6178 = pi05139 & w3598;
assign w6179 = pi03171 & w3522;
assign w6180 = pi05093 & w3232;
assign w6181 = pi05496 & w3234;
assign w6182 = pi03208 & w3454;
assign w6183 = pi03389 & w3258;
assign w6184 = pi03337 & w3512;
assign w6185 = pi01764 & w3282;
assign w6186 = pi06014 & w3440;
assign w6187 = pi03045 & w3490;
assign w6188 = pi05580 & w3156;
assign w6189 = pi03290 & w3190;
assign w6190 = pi01759 & w3462;
assign w6191 = pi05265 & w3586;
assign w6192 = pi06060 & w3173;
assign w6193 = pi05613 & w3221;
assign w6194 = pi05593 & w3254;
assign w6195 = pi02822 & w3614;
assign w6196 = pi05645 & w3448;
assign w6197 = pi05964 & w3175;
assign w6198 = pi03316 & w3564;
assign w6199 = pi03283 & w3115;
assign w6200 = pi05704 & w3165;
assign w6201 = pi02973 & w3536;
assign w6202 = pi06230 & w3580;
assign w6203 = pi06259 & w3148;
assign w6204 = pi05106 & w3266;
assign w6205 = pi05848 & w3270;
assign w6206 = pi05902 & w3093;
assign w6207 = pi05799 & w3192;
assign w6208 = pi05435 & w3078;
assign w6209 = pi05413 & w3514;
assign w6210 = pi05187 & w3554;
assign w6211 = pi05086 & w3486;
assign w6212 = pi01751 & w3153;
assign w6213 = pi05828 & w3464;
assign w6214 = pi03032 & w3244;
assign w6215 = pi05339 & w3203;
assign w6216 = pi05541 & w3286;
assign w6217 = pi05632 & w3376;
assign w6218 = pi03442 & w3388;
assign w6219 = pi05456 & w3442;
assign w6220 = pi09568 & w3137;
assign w6221 = pi05665 & w3434;
assign w6222 = pi05407 & w3278;
assign w6223 = pi05353 & w3199;
assign w6224 = pi05226 & w3480;
assign w6225 = pi03416 & w3162;
assign w6226 = pi02880 & w3268;
assign w6227 = pi05426 & w3284;
assign w6228 = pi01768 & w3496;
assign w6229 = pi01879 & w3584;
assign w6230 = pi05778 & w3476;
assign w6231 = pi05239 & w3112;
assign w6232 = pi02854 & w3197;
assign w6233 = pi03364 & w3562;
assign w6234 = pi03097 & w3592;
assign w6235 = pi03138 & w3574;
assign w6236 = pi06441 & w3558;
assign w6237 = pi02861 & w3336;
assign w6238 = pi05977 & w3223;
assign w6239 = pi05245 & w3378;
assign w6240 = pi02841 & w3346;
assign w6241 = pi02999 & w3262;
assign w6242 = pi03502 & w3488;
assign w6243 = pi03296 & w3328;
assign w6244 = pi06243 & w3560;
assign w6245 = pi09793 & w3150;
assign w6246 = pi05522 & w3406;
assign w6247 = pi05219 & w3288;
assign w6248 = pi01926 & w3450;
assign w6249 = pi03177 & w3181;
assign w6250 = pi02887 & w3416;
assign w6251 = pi02920 & w3530;
assign w6252 = pi05619 & w3620;
assign w6253 = pi05915 & w3426;
assign w6254 = pi05652 & w3566;
assign w6255 = pi06249 & w3342;
assign w6256 = pi03243 & w3326;
assign w6257 = pi03276 & w3086;
assign w6258 = pi05554 & w3410;
assign w6259 = pi09580 & w3424;
assign w6260 = pi06107 & w3320;
assign w6261 = pi05099 & w3240;
assign w6262 = pi05160 & w3492;
assign w6263 = pi02867 & w3544;
assign w6264 = pi05252 & w3356;
assign w6265 = pi05200 & w3528;
assign w6266 = pi05325 & w3354;
assign w6267 = pi05232 & w3217;
assign w6268 = pi05561 & w3420;
assign w6269 = pi05476 & w3506;
assign w6270 = pi06236 & w3229;
assign w6271 = pi06098 & w3444;
assign w6272 = pi05587 & w3205;
assign w6273 = pi03078 & w3338;
assign w6274 = pi03303 & w3484;
assign w6275 = pi02959 & w3103;
assign w6276 = pi09589 & w3274;
assign w6277 = pi03486 & w3582;
assign w6278 = pi06199 & w3318;
assign w6279 = pi02893 & w3470;
assign w6280 = pi06191 & w3096;
assign w6281 = pi05857 & w3386;
assign w6282 = pi06007 & w3570;
assign w6283 = pi06021 & w3608;
assign w6284 = pi02211 & w3502;
assign w6285 = pi05818 & w3390;
assign w6286 = pi05567 & w3135;
assign w6287 = pi05895 & w3125;
assign w6288 = pi05345 & w3129;
assign w6289 = pi09719 & w3352;
assign w6290 = pi01615 & w3160;
assign w6291 = pi02986 & w3296;
assign w6292 = pi05442 & w3256;
assign w6293 = pi05291 & w3314;
assign w6294 = pi05420 & w3186;
assign w6295 = pi05731 & w3374;
assign w6296 = pi03119 & w3394;
assign w6297 = pi03230 & w3290;
assign w6298 = pi05626 & w3272;
assign w6299 = pi03065 & w3576;
assign w6300 = pi06081 & w3106;
assign w6301 = pi05489 & w3398;
assign w6302 = pi05502 & w3466;
assign w6303 = pi03125 & w3071;
assign w6304 = pi01484 & w3110;
assign w6305 = pi03322 & w3370;
assign w6306 = pi05133 & w3248;
assign w6307 = pi03104 & w3498;
assign w6308 = pi03084 & w3348;
assign w6309 = pi05173 & w3252;
assign w6310 = pi02914 & w3330;
assign w6311 = pi05996 & w3446;
assign w6312 = pi05332 & w3392;
assign w6313 = pi02933 & w3064;
assign w6314 = pi05469 & w3432;
assign w6315 = pi02953 & w3322;
assign w6316 = ~w6060 & ~w6061;
assign w6317 = ~w6062 & ~w6063;
assign w6318 = ~w6064 & ~w6065;
assign w6319 = ~w6066 & ~w6067;
assign w6320 = ~w6068 & ~w6069;
assign w6321 = ~w6070 & ~w6071;
assign w6322 = ~w6072 & ~w6073;
assign w6323 = ~w6074 & ~w6075;
assign w6324 = ~w6076 & ~w6077;
assign w6325 = ~w6078 & ~w6079;
assign w6326 = ~w6080 & ~w6081;
assign w6327 = ~w6082 & ~w6083;
assign w6328 = ~w6084 & ~w6085;
assign w6329 = ~w6086 & ~w6087;
assign w6330 = ~w6088 & ~w6089;
assign w6331 = ~w6090 & ~w6091;
assign w6332 = ~w6092 & ~w6093;
assign w6333 = ~w6094 & ~w6095;
assign w6334 = ~w6096 & ~w6097;
assign w6335 = ~w6098 & ~w6099;
assign w6336 = ~w6100 & ~w6101;
assign w6337 = ~w6102 & ~w6103;
assign w6338 = ~w6104 & ~w6105;
assign w6339 = ~w6106 & ~w6107;
assign w6340 = ~w6108 & ~w6109;
assign w6341 = ~w6110 & ~w6111;
assign w6342 = ~w6112 & ~w6113;
assign w6343 = ~w6114 & ~w6115;
assign w6344 = ~w6116 & ~w6117;
assign w6345 = ~w6118 & ~w6119;
assign w6346 = ~w6120 & ~w6121;
assign w6347 = ~w6122 & ~w6123;
assign w6348 = ~w6124 & ~w6125;
assign w6349 = ~w6126 & ~w6127;
assign w6350 = ~w6128 & ~w6129;
assign w6351 = ~w6130 & ~w6131;
assign w6352 = ~w6132 & ~w6133;
assign w6353 = ~w6134 & ~w6135;
assign w6354 = ~w6136 & ~w6137;
assign w6355 = ~w6138 & ~w6139;
assign w6356 = ~w6140 & ~w6141;
assign w6357 = ~w6142 & ~w6143;
assign w6358 = ~w6144 & ~w6145;
assign w6359 = ~w6146 & ~w6147;
assign w6360 = ~w6148 & ~w6149;
assign w6361 = ~w6150 & ~w6151;
assign w6362 = ~w6152 & ~w6153;
assign w6363 = ~w6154 & ~w6155;
assign w6364 = ~w6156 & ~w6157;
assign w6365 = ~w6158 & ~w6159;
assign w6366 = ~w6160 & ~w6161;
assign w6367 = ~w6162 & ~w6163;
assign w6368 = ~w6164 & ~w6165;
assign w6369 = ~w6166 & ~w6167;
assign w6370 = ~w6168 & ~w6169;
assign w6371 = ~w6170 & ~w6171;
assign w6372 = ~w6172 & ~w6173;
assign w6373 = ~w6174 & ~w6175;
assign w6374 = ~w6176 & ~w6177;
assign w6375 = ~w6178 & ~w6179;
assign w6376 = ~w6180 & ~w6181;
assign w6377 = ~w6182 & ~w6183;
assign w6378 = ~w6184 & ~w6185;
assign w6379 = ~w6186 & ~w6187;
assign w6380 = ~w6188 & ~w6189;
assign w6381 = ~w6190 & ~w6191;
assign w6382 = ~w6192 & ~w6193;
assign w6383 = ~w6194 & ~w6195;
assign w6384 = ~w6196 & ~w6197;
assign w6385 = ~w6198 & ~w6199;
assign w6386 = ~w6200 & ~w6201;
assign w6387 = ~w6202 & ~w6203;
assign w6388 = ~w6204 & ~w6205;
assign w6389 = ~w6206 & ~w6207;
assign w6390 = ~w6208 & ~w6209;
assign w6391 = ~w6210 & ~w6211;
assign w6392 = ~w6212 & ~w6213;
assign w6393 = ~w6214 & ~w6215;
assign w6394 = ~w6216 & ~w6217;
assign w6395 = ~w6218 & ~w6219;
assign w6396 = ~w6220 & ~w6221;
assign w6397 = ~w6222 & ~w6223;
assign w6398 = ~w6224 & ~w6225;
assign w6399 = ~w6226 & ~w6227;
assign w6400 = ~w6228 & ~w6229;
assign w6401 = ~w6230 & ~w6231;
assign w6402 = ~w6232 & ~w6233;
assign w6403 = ~w6234 & ~w6235;
assign w6404 = ~w6236 & ~w6237;
assign w6405 = ~w6238 & ~w6239;
assign w6406 = ~w6240 & ~w6241;
assign w6407 = ~w6242 & ~w6243;
assign w6408 = ~w6244 & ~w6245;
assign w6409 = ~w6246 & ~w6247;
assign w6410 = ~w6248 & ~w6249;
assign w6411 = ~w6250 & ~w6251;
assign w6412 = ~w6252 & ~w6253;
assign w6413 = ~w6254 & ~w6255;
assign w6414 = ~w6256 & ~w6257;
assign w6415 = ~w6258 & ~w6259;
assign w6416 = ~w6260 & ~w6261;
assign w6417 = ~w6262 & ~w6263;
assign w6418 = ~w6264 & ~w6265;
assign w6419 = ~w6266 & ~w6267;
assign w6420 = ~w6268 & ~w6269;
assign w6421 = ~w6270 & ~w6271;
assign w6422 = ~w6272 & ~w6273;
assign w6423 = ~w6274 & ~w6275;
assign w6424 = ~w6276 & ~w6277;
assign w6425 = ~w6278 & ~w6279;
assign w6426 = ~w6280 & ~w6281;
assign w6427 = ~w6282 & ~w6283;
assign w6428 = ~w6284 & ~w6285;
assign w6429 = ~w6286 & ~w6287;
assign w6430 = ~w6288 & ~w6289;
assign w6431 = ~w6290 & ~w6291;
assign w6432 = ~w6292 & ~w6293;
assign w6433 = ~w6294 & ~w6295;
assign w6434 = ~w6296 & ~w6297;
assign w6435 = ~w6298 & ~w6299;
assign w6436 = ~w6300 & ~w6301;
assign w6437 = ~w6302 & ~w6303;
assign w6438 = ~w6304 & ~w6305;
assign w6439 = ~w6306 & ~w6307;
assign w6440 = ~w6308 & ~w6309;
assign w6441 = ~w6310 & ~w6311;
assign w6442 = ~w6312 & ~w6313;
assign w6443 = ~w6314 & ~w6315;
assign w6444 = w6442 & w6443;
assign w6445 = w6440 & w6441;
assign w6446 = w6438 & w6439;
assign w6447 = w6436 & w6437;
assign w6448 = w6434 & w6435;
assign w6449 = w6432 & w6433;
assign w6450 = w6430 & w6431;
assign w6451 = w6428 & w6429;
assign w6452 = w6426 & w6427;
assign w6453 = w6424 & w6425;
assign w6454 = w6422 & w6423;
assign w6455 = w6420 & w6421;
assign w6456 = w6418 & w6419;
assign w6457 = w6416 & w6417;
assign w6458 = w6414 & w6415;
assign w6459 = w6412 & w6413;
assign w6460 = w6410 & w6411;
assign w6461 = w6408 & w6409;
assign w6462 = w6406 & w6407;
assign w6463 = w6404 & w6405;
assign w6464 = w6402 & w6403;
assign w6465 = w6400 & w6401;
assign w6466 = w6398 & w6399;
assign w6467 = w6396 & w6397;
assign w6468 = w6394 & w6395;
assign w6469 = w6392 & w6393;
assign w6470 = w6390 & w6391;
assign w6471 = w6388 & w6389;
assign w6472 = w6386 & w6387;
assign w6473 = w6384 & w6385;
assign w6474 = w6382 & w6383;
assign w6475 = w6380 & w6381;
assign w6476 = w6378 & w6379;
assign w6477 = w6376 & w6377;
assign w6478 = w6374 & w6375;
assign w6479 = w6372 & w6373;
assign w6480 = w6370 & w6371;
assign w6481 = w6368 & w6369;
assign w6482 = w6366 & w6367;
assign w6483 = w6364 & w6365;
assign w6484 = w6362 & w6363;
assign w6485 = w6360 & w6361;
assign w6486 = w6358 & w6359;
assign w6487 = w6356 & w6357;
assign w6488 = w6354 & w6355;
assign w6489 = w6352 & w6353;
assign w6490 = w6350 & w6351;
assign w6491 = w6348 & w6349;
assign w6492 = w6346 & w6347;
assign w6493 = w6344 & w6345;
assign w6494 = w6342 & w6343;
assign w6495 = w6340 & w6341;
assign w6496 = w6338 & w6339;
assign w6497 = w6336 & w6337;
assign w6498 = w6334 & w6335;
assign w6499 = w6332 & w6333;
assign w6500 = w6330 & w6331;
assign w6501 = w6328 & w6329;
assign w6502 = w6326 & w6327;
assign w6503 = w6324 & w6325;
assign w6504 = w6322 & w6323;
assign w6505 = w6320 & w6321;
assign w6506 = w6318 & w6319;
assign w6507 = w6316 & w6317;
assign w6508 = w6506 & w6507;
assign w6509 = w6504 & w6505;
assign w6510 = w6502 & w6503;
assign w6511 = w6500 & w6501;
assign w6512 = w6498 & w6499;
assign w6513 = w6496 & w6497;
assign w6514 = w6494 & w6495;
assign w6515 = w6492 & w6493;
assign w6516 = w6490 & w6491;
assign w6517 = w6488 & w6489;
assign w6518 = w6486 & w6487;
assign w6519 = w6484 & w6485;
assign w6520 = w6482 & w6483;
assign w6521 = w6480 & w6481;
assign w6522 = w6478 & w6479;
assign w6523 = w6476 & w6477;
assign w6524 = w6474 & w6475;
assign w6525 = w6472 & w6473;
assign w6526 = w6470 & w6471;
assign w6527 = w6468 & w6469;
assign w6528 = w6466 & w6467;
assign w6529 = w6464 & w6465;
assign w6530 = w6462 & w6463;
assign w6531 = w6460 & w6461;
assign w6532 = w6458 & w6459;
assign w6533 = w6456 & w6457;
assign w6534 = w6454 & w6455;
assign w6535 = w6452 & w6453;
assign w6536 = w6450 & w6451;
assign w6537 = w6448 & w6449;
assign w6538 = w6446 & w6447;
assign w6539 = w6444 & w6445;
assign w6540 = w6538 & w6539;
assign w6541 = w6536 & w6537;
assign w6542 = w6534 & w6535;
assign w6543 = w6532 & w6533;
assign w6544 = w6530 & w6531;
assign w6545 = w6528 & w6529;
assign w6546 = w6526 & w6527;
assign w6547 = w6524 & w6525;
assign w6548 = w6522 & w6523;
assign w6549 = w6520 & w6521;
assign w6550 = w6518 & w6519;
assign w6551 = w6516 & w6517;
assign w6552 = w6514 & w6515;
assign w6553 = w6512 & w6513;
assign w6554 = w6510 & w6511;
assign w6555 = w6508 & w6509;
assign w6556 = w6554 & w6555;
assign w6557 = w6552 & w6553;
assign w6558 = w6550 & w6551;
assign w6559 = w6548 & w6549;
assign w6560 = w6546 & w6547;
assign w6561 = w6544 & w6545;
assign w6562 = w6542 & w6543;
assign w6563 = w6540 & w6541;
assign w6564 = w6562 & w6563;
assign w6565 = w6560 & w6561;
assign w6566 = w6558 & w6559;
assign w6567 = w6556 & w6557;
assign w6568 = w6566 & w6567;
assign w6569 = w6564 & w6565;
assign w6570 = w6568 & w6569;
assign w6571 = ~pi10577 & ~w6570;
assign w6572 = pi03951 & w3498;
assign w6573 = pi07701 & w3468;
assign w6574 = pi03898 & w3209;
assign w6575 = pi02443 & w3229;
assign w6576 = pi04299 & w3588;
assign w6577 = pi02281 & w3516;
assign w6578 = pi07292 & w3276;
assign w6579 = pi06583 & w3492;
assign w6580 = pi07931 & w3316;
assign w6581 = pi07414 & w3171;
assign w6582 = pi03820 & w3260;
assign w6583 = pi04252 & w3504;
assign w6584 = pi03827 & w3610;
assign w6585 = pi03560 & w3197;
assign w6586 = pi01659 & w3508;
assign w6587 = pi03906 & w3338;
assign w6588 = pi07767 & w3282;
assign w6589 = pi07692 & w3594;
assign w6590 = pi04226 & w3258;
assign w6591 = pi06687 & w3356;
assign w6592 = pi06560 & w3604;
assign w6593 = pi07143 & w3410;
assign w6594 = pi07059 & w3234;
assign w6595 = pi07747 & w3444;
assign w6596 = pi02272 & w3284;
assign w6597 = pi06571 & w3344;
assign w6598 = pi07081 & w3139;
assign w6599 = pi07200 & w3225;
assign w6600 = pi07911 & w3148;
assign w6601 = pi04273 & w3556;
assign w6602 = pi04245 & w3162;
assign w6603 = pi07469 & w3390;
assign w6604 = pi09565 & w3446;
assign w6605 = pi07248 & w3272;
assign w6606 = pi06742 & w3314;
assign w6607 = pi07433 & w3458;
assign w6608 = pi01732 & w3324;
assign w6609 = pi06852 & w3304;
assign w6610 = pi08024 & w3368;
assign w6611 = pi01641 & w3546;
assign w6612 = pi07159 & w3135;
assign w6613 = pi03801 & w3137;
assign w6614 = pi03729 & w3534;
assign w6615 = pi06477 & w3486;
assign w6616 = pi08101 & w3558;
assign w6617 = pi07840 & w3318;
assign w6618 = pi06664 & w3217;
assign w6619 = pi09633 & w3522;
assign w6620 = pi06629 & w3528;
assign w6621 = pi06900 & w3082;
assign w6622 = pi04220 & w3302;
assign w6623 = pi02389 & w3488;
assign w6624 = pi04213 & w3169;
assign w6625 = pi03859 & w3526;
assign w6626 = pi01882 & w3424;
assign w6627 = pi09769 & w3462;
assign w6628 = pi06493 & w3240;
assign w6629 = pi06592 & w3612;
assign w6630 = pi03775 & w3536;
assign w6631 = pi07268 & w3358;
assign w6632 = pi02491 & w3173;
assign w6633 = pi06679 & w3378;
assign w6634 = pi04108 & w3214;
assign w6635 = pi07488 & w3207;
assign w6636 = pi06643 & w3568;
assign w6637 = pi04050 & w3502;
assign w6638 = pi03768 & w3274;
assign w6639 = pi06729 & w3482;
assign w6640 = pi04089 & w3326;
assign w6641 = pi06872 & w3496;
assign w6642 = pi07395 & w3590;
assign w6643 = pi02321 & w3572;
assign w6644 = pi07965 & w3158;
assign w6645 = pi03664 & w3362;
assign w6646 = pi07562 & w3426;
assign w6647 = pi07814 & w3280;
assign w6648 = pi06637 & w3550;
assign w6649 = pi06761 & w3450;
assign w6650 = pi03592 & w3500;
assign w6651 = pi08119 & w3510;
assign w6652 = pi06999 & w3442;
assign w6653 = pi07384 & w3194;
assign w6654 = pi07013 & w3384;
assign w6655 = pi08008 & w3179;
assign w6656 = pi08056 & w3418;
assign w6657 = pi07035 & w3506;
assign w6658 = pi04181 & w3370;
assign w6659 = pi03570 & w3336;
assign w6660 = pi02412 & w3211;
assign w6661 = pi07133 & w3552;
assign w6662 = pi07375 & w3600;
assign w6663 = pi06512 & w3143;
assign w6664 = pi04082 & w3290;
assign w6665 = pi02545 & w3177;
assign w6666 = pi06623 & w3452;
assign w6667 = pi06960 & w3078;
assign w6668 = pi06485 & w3232;
assign w6669 = pi01560 & w3542;
assign w6670 = pi07761 & w3478;
assign w6671 = pi06878 & w3153;
assign w6672 = pi04056 & w3454;
assign w6673 = pi04010 & w3494;
assign w6674 = pi01549 & w3188;
assign w6675 = pi01913 & w3342;
assign w6676 = pi07951 & w3332;
assign w6677 = pi06836 & w3422;
assign w6678 = pi06499 & w3266;
assign w6679 = pi06846 & w3227;
assign w6680 = pi06715 & w3414;
assign w6681 = pi08017 & w3438;
assign w6682 = pi01742 & w3566;
assign w6683 = pi04174 & w3564;
assign w6684 = pi03697 & w3530;
assign w6685 = pi07104 & w3340;
assign w6686 = pi01638 & w3167;
assign w6687 = pi02451 & w3160;
assign w6688 = pi03716 & w3064;
assign w6689 = pi08092 & w3150;
assign w6690 = pi07323 & w3312;
assign w6691 = pi03541 & w3346;
assign w6692 = pi06768 & w3236;
assign w6693 = pi04016 & w3428;
assign w6694 = pi07165 & w3364;
assign w6695 = pi03846 & w3548;
assign w6696 = pi07068 & w3466;
assign w6697 = pi02616 & w3388;
assign w6698 = pi08081 & w3110;
assign w6699 = pi01782 & w3448;
assign w6700 = pi06616 & w3554;
assign w6701 = pi04207 & w3562;
assign w6702 = pi02283 & w3294;
assign w6703 = pi07404 & w3430;
assign w6704 = pi07893 & w3560;
assign w6705 = pi07499 & w3270;
assign w6706 = pi06522 & w3308;
assign w6707 = pi08065 & w3246;
assign w6708 = pi06656 & w3480;
assign w6709 = pi06696 & w3460;
assign w6710 = pi07754 & w3320;
assign w6711 = pi07116 & w3286;
assign w6712 = pi06421 & w3096;
assign w6713 = pi07543 & w3093;
assign w6714 = pi03520 & w3306;
assign w6715 = pi03938 & w3592;
assign w6716 = pi02588 & w3372;
assign w6717 = pi04168 & w3146;
assign w6718 = pi07873 & w3580;
assign w6719 = pi04003 & w3574;
assign w6720 = pi01605 & w3296;
assign w6721 = pi01695 & w3408;
assign w6722 = pi07256 & w3376;
assign w6723 = pi01921 & w3474;
assign w6724 = pi04194 & w3512;
assign w6725 = pi07734 & w3106;
assign w6726 = pi07664 & w3608;
assign w6727 = pi03840 & w3244;
assign w6728 = pi06703 & w3586;
assign w6729 = pi07609 & w3175;
assign w6730 = pi03580 & w3544;
assign w6731 = pi06775 & w3298;
assign w6732 = pi09347 & w3440;
assign w6733 = pi07300 & w3434;
assign w6734 = pi07178 & w3156;
assign w6735 = pi06813 & w3129;
assign w6736 = pi07449 & w3192;
assign w6737 = pi03892 & w3576;
assign w6738 = pi03866 & w3350;
assign w6739 = pi03853 & w3490;
assign w6740 = pi04326 & w3582;
assign w6741 = pi03807 & w3262;
assign w6742 = pi03964 & w3394;
assign w6743 = pi03645 & w3416;
assign w6744 = pi03958 & w3132;
assign w6745 = pi03511 & w3614;
assign w6746 = pi07588 & w3532;
assign w6747 = pi04129 & w3115;
assign w6748 = pi04187 & w3618;
assign w6749 = pi04135 & w3190;
assign w6750 = pi06610 & w3219;
assign w6751 = pi02496 & w3352;
assign w6752 = pi08132 & w3242;
assign w6753 = pi01856 & w3514;
assign w6754 = pi02471 & w3396;
assign w6755 = pi07074 & w3127;
assign w6756 = pi07553 & w3238;
assign w6757 = pi03928 & w3456;
assign w6758 = pi07601 & w3616;
assign w6759 = pi07507 & w3386;
assign w6760 = pi06602 & w3252;
assign w6761 = pi07027 & w3432;
assign w6762 = pi07226 & w3221;
assign w6763 = pi02629 & w3278;
assign w6764 = pi06541 & w3248;
assign w6765 = pi03684 & w3330;
assign w6766 = pi06807 & w3203;
assign w6767 = pi01860 & w3256;
assign w6768 = pi06748 & w3538;
assign w6769 = pi03833 & w3310;
assign w6770 = pi03736 & w3400;
assign w6771 = pi02440 & w3125;
assign w6772 = pi03601 & w3268;
assign w6773 = pi02538 & w3402;
assign w6774 = pi01585 & w3223;
assign w6775 = pi03984 & w3118;
assign w6776 = pi03554 & w3520;
assign w6777 = pi08044 & w3524;
assign w6778 = pi07213 & w3472;
assign w6779 = pi06551 & w3598;
assign w6780 = pi04042 & w3181;
assign w6781 = pi02530 & w3374;
assign w6782 = pi04098 & w3334;
assign w6783 = pi03677 & w3404;
assign w6784 = pi02624 & w3184;
assign w6785 = pi03755 & w3103;
assign w6786 = pi07459 & w3360;
assign w6787 = pi06650 & w3288;
assign w6788 = pi06986 & w3518;
assign w6789 = pi06722 & w3540;
assign w6790 = pi07478 & w3464;
assign w6791 = pi07087 & w3406;
assign w6792 = pi03742 & w3322;
assign w6793 = pi07423 & w3476;
assign w6794 = pi03533 & w3380;
assign w6795 = pi06670 & w3112;
assign w6796 = pi07152 & w3420;
assign w6797 = pi07990 & w3578;
assign w6798 = pi07240 & w3620;
assign w6799 = pi09681 & w3071;
assign w6800 = pi01554 & w3606;
assign w6801 = pi07185 & w3205;
assign w6802 = pi09762 & w3398;
assign w6803 = pi06784 & w3354;
assign w6804 = pi06532 & w3436;
assign w6805 = pi06820 & w3199;
assign w6806 = pi02548 & w3366;
assign w6807 = pi03651 & w3470;
assign w6808 = pi02531 & w3382;
assign w6809 = pi07644 & w3570;
assign w6810 = pi04233 & w3122;
assign w6811 = pi03703 & w3250;
assign w6812 = pi03814 & w3292;
assign w6813 = pi04200 & w3412;
assign w6814 = pi07775 & w3264;
assign w6815 = pi07191 & w3254;
assign w6816 = pi03919 & w3348;
assign w6817 = pi04122 & w3086;
assign w6818 = pi07338 & w3165;
assign w6819 = pi07042 & w3300;
assign w6820 = pi04148 & w3484;
assign w6821 = pi04142 & w3328;
assign w6822 = pi02481 & w3596;
assign w6823 = pi07353 & w3201;
assign w6824 = pi07978 & w3602;
assign w6825 = pi06797 & w3392;
assign w6826 = pi02315 & w3186;
assign w6827 = pi07721 & w3584;
assign w6828 = ~w6572 & ~w6573;
assign w6829 = ~w6574 & ~w6575;
assign w6830 = ~w6576 & ~w6577;
assign w6831 = ~w6578 & ~w6579;
assign w6832 = ~w6580 & ~w6581;
assign w6833 = ~w6582 & ~w6583;
assign w6834 = ~w6584 & ~w6585;
assign w6835 = ~w6586 & ~w6587;
assign w6836 = ~w6588 & ~w6589;
assign w6837 = ~w6590 & ~w6591;
assign w6838 = ~w6592 & ~w6593;
assign w6839 = ~w6594 & ~w6595;
assign w6840 = ~w6596 & ~w6597;
assign w6841 = ~w6598 & ~w6599;
assign w6842 = ~w6600 & ~w6601;
assign w6843 = ~w6602 & ~w6603;
assign w6844 = ~w6604 & ~w6605;
assign w6845 = ~w6606 & ~w6607;
assign w6846 = ~w6608 & ~w6609;
assign w6847 = ~w6610 & ~w6611;
assign w6848 = ~w6612 & ~w6613;
assign w6849 = ~w6614 & ~w6615;
assign w6850 = ~w6616 & ~w6617;
assign w6851 = ~w6618 & ~w6619;
assign w6852 = ~w6620 & ~w6621;
assign w6853 = ~w6622 & ~w6623;
assign w6854 = ~w6624 & ~w6625;
assign w6855 = ~w6626 & ~w6627;
assign w6856 = ~w6628 & ~w6629;
assign w6857 = ~w6630 & ~w6631;
assign w6858 = ~w6632 & ~w6633;
assign w6859 = ~w6634 & ~w6635;
assign w6860 = ~w6636 & ~w6637;
assign w6861 = ~w6638 & ~w6639;
assign w6862 = ~w6640 & ~w6641;
assign w6863 = ~w6642 & ~w6643;
assign w6864 = ~w6644 & ~w6645;
assign w6865 = ~w6646 & ~w6647;
assign w6866 = ~w6648 & ~w6649;
assign w6867 = ~w6650 & ~w6651;
assign w6868 = ~w6652 & ~w6653;
assign w6869 = ~w6654 & ~w6655;
assign w6870 = ~w6656 & ~w6657;
assign w6871 = ~w6658 & ~w6659;
assign w6872 = ~w6660 & ~w6661;
assign w6873 = ~w6662 & ~w6663;
assign w6874 = ~w6664 & ~w6665;
assign w6875 = ~w6666 & ~w6667;
assign w6876 = ~w6668 & ~w6669;
assign w6877 = ~w6670 & ~w6671;
assign w6878 = ~w6672 & ~w6673;
assign w6879 = ~w6674 & ~w6675;
assign w6880 = ~w6676 & ~w6677;
assign w6881 = ~w6678 & ~w6679;
assign w6882 = ~w6680 & ~w6681;
assign w6883 = ~w6682 & ~w6683;
assign w6884 = ~w6684 & ~w6685;
assign w6885 = ~w6686 & ~w6687;
assign w6886 = ~w6688 & ~w6689;
assign w6887 = ~w6690 & ~w6691;
assign w6888 = ~w6692 & ~w6693;
assign w6889 = ~w6694 & ~w6695;
assign w6890 = ~w6696 & ~w6697;
assign w6891 = ~w6698 & ~w6699;
assign w6892 = ~w6700 & ~w6701;
assign w6893 = ~w6702 & ~w6703;
assign w6894 = ~w6704 & ~w6705;
assign w6895 = ~w6706 & ~w6707;
assign w6896 = ~w6708 & ~w6709;
assign w6897 = ~w6710 & ~w6711;
assign w6898 = ~w6712 & ~w6713;
assign w6899 = ~w6714 & ~w6715;
assign w6900 = ~w6716 & ~w6717;
assign w6901 = ~w6718 & ~w6719;
assign w6902 = ~w6720 & ~w6721;
assign w6903 = ~w6722 & ~w6723;
assign w6904 = ~w6724 & ~w6725;
assign w6905 = ~w6726 & ~w6727;
assign w6906 = ~w6728 & ~w6729;
assign w6907 = ~w6730 & ~w6731;
assign w6908 = ~w6732 & ~w6733;
assign w6909 = ~w6734 & ~w6735;
assign w6910 = ~w6736 & ~w6737;
assign w6911 = ~w6738 & ~w6739;
assign w6912 = ~w6740 & ~w6741;
assign w6913 = ~w6742 & ~w6743;
assign w6914 = ~w6744 & ~w6745;
assign w6915 = ~w6746 & ~w6747;
assign w6916 = ~w6748 & ~w6749;
assign w6917 = ~w6750 & ~w6751;
assign w6918 = ~w6752 & ~w6753;
assign w6919 = ~w6754 & ~w6755;
assign w6920 = ~w6756 & ~w6757;
assign w6921 = ~w6758 & ~w6759;
assign w6922 = ~w6760 & ~w6761;
assign w6923 = ~w6762 & ~w6763;
assign w6924 = ~w6764 & ~w6765;
assign w6925 = ~w6766 & ~w6767;
assign w6926 = ~w6768 & ~w6769;
assign w6927 = ~w6770 & ~w6771;
assign w6928 = ~w6772 & ~w6773;
assign w6929 = ~w6774 & ~w6775;
assign w6930 = ~w6776 & ~w6777;
assign w6931 = ~w6778 & ~w6779;
assign w6932 = ~w6780 & ~w6781;
assign w6933 = ~w6782 & ~w6783;
assign w6934 = ~w6784 & ~w6785;
assign w6935 = ~w6786 & ~w6787;
assign w6936 = ~w6788 & ~w6789;
assign w6937 = ~w6790 & ~w6791;
assign w6938 = ~w6792 & ~w6793;
assign w6939 = ~w6794 & ~w6795;
assign w6940 = ~w6796 & ~w6797;
assign w6941 = ~w6798 & ~w6799;
assign w6942 = ~w6800 & ~w6801;
assign w6943 = ~w6802 & ~w6803;
assign w6944 = ~w6804 & ~w6805;
assign w6945 = ~w6806 & ~w6807;
assign w6946 = ~w6808 & ~w6809;
assign w6947 = ~w6810 & ~w6811;
assign w6948 = ~w6812 & ~w6813;
assign w6949 = ~w6814 & ~w6815;
assign w6950 = ~w6816 & ~w6817;
assign w6951 = ~w6818 & ~w6819;
assign w6952 = ~w6820 & ~w6821;
assign w6953 = ~w6822 & ~w6823;
assign w6954 = ~w6824 & ~w6825;
assign w6955 = ~w6826 & ~w6827;
assign w6956 = w6954 & w6955;
assign w6957 = w6952 & w6953;
assign w6958 = w6950 & w6951;
assign w6959 = w6948 & w6949;
assign w6960 = w6946 & w6947;
assign w6961 = w6944 & w6945;
assign w6962 = w6942 & w6943;
assign w6963 = w6940 & w6941;
assign w6964 = w6938 & w6939;
assign w6965 = w6936 & w6937;
assign w6966 = w6934 & w6935;
assign w6967 = w6932 & w6933;
assign w6968 = w6930 & w6931;
assign w6969 = w6928 & w6929;
assign w6970 = w6926 & w6927;
assign w6971 = w6924 & w6925;
assign w6972 = w6922 & w6923;
assign w6973 = w6920 & w6921;
assign w6974 = w6918 & w6919;
assign w6975 = w6916 & w6917;
assign w6976 = w6914 & w6915;
assign w6977 = w6912 & w6913;
assign w6978 = w6910 & w6911;
assign w6979 = w6908 & w6909;
assign w6980 = w6906 & w6907;
assign w6981 = w6904 & w6905;
assign w6982 = w6902 & w6903;
assign w6983 = w6900 & w6901;
assign w6984 = w6898 & w6899;
assign w6985 = w6896 & w6897;
assign w6986 = w6894 & w6895;
assign w6987 = w6892 & w6893;
assign w6988 = w6890 & w6891;
assign w6989 = w6888 & w6889;
assign w6990 = w6886 & w6887;
assign w6991 = w6884 & w6885;
assign w6992 = w6882 & w6883;
assign w6993 = w6880 & w6881;
assign w6994 = w6878 & w6879;
assign w6995 = w6876 & w6877;
assign w6996 = w6874 & w6875;
assign w6997 = w6872 & w6873;
assign w6998 = w6870 & w6871;
assign w6999 = w6868 & w6869;
assign w7000 = w6866 & w6867;
assign w7001 = w6864 & w6865;
assign w7002 = w6862 & w6863;
assign w7003 = w6860 & w6861;
assign w7004 = w6858 & w6859;
assign w7005 = w6856 & w6857;
assign w7006 = w6854 & w6855;
assign w7007 = w6852 & w6853;
assign w7008 = w6850 & w6851;
assign w7009 = w6848 & w6849;
assign w7010 = w6846 & w6847;
assign w7011 = w6844 & w6845;
assign w7012 = w6842 & w6843;
assign w7013 = w6840 & w6841;
assign w7014 = w6838 & w6839;
assign w7015 = w6836 & w6837;
assign w7016 = w6834 & w6835;
assign w7017 = w6832 & w6833;
assign w7018 = w6830 & w6831;
assign w7019 = w6828 & w6829;
assign w7020 = w7018 & w7019;
assign w7021 = w7016 & w7017;
assign w7022 = w7014 & w7015;
assign w7023 = w7012 & w7013;
assign w7024 = w7010 & w7011;
assign w7025 = w7008 & w7009;
assign w7026 = w7006 & w7007;
assign w7027 = w7004 & w7005;
assign w7028 = w7002 & w7003;
assign w7029 = w7000 & w7001;
assign w7030 = w6998 & w6999;
assign w7031 = w6996 & w6997;
assign w7032 = w6994 & w6995;
assign w7033 = w6992 & w6993;
assign w7034 = w6990 & w6991;
assign w7035 = w6988 & w6989;
assign w7036 = w6986 & w6987;
assign w7037 = w6984 & w6985;
assign w7038 = w6982 & w6983;
assign w7039 = w6980 & w6981;
assign w7040 = w6978 & w6979;
assign w7041 = w6976 & w6977;
assign w7042 = w6974 & w6975;
assign w7043 = w6972 & w6973;
assign w7044 = w6970 & w6971;
assign w7045 = w6968 & w6969;
assign w7046 = w6966 & w6967;
assign w7047 = w6964 & w6965;
assign w7048 = w6962 & w6963;
assign w7049 = w6960 & w6961;
assign w7050 = w6958 & w6959;
assign w7051 = w6956 & w6957;
assign w7052 = w7050 & w7051;
assign w7053 = w7048 & w7049;
assign w7054 = w7046 & w7047;
assign w7055 = w7044 & w7045;
assign w7056 = w7042 & w7043;
assign w7057 = w7040 & w7041;
assign w7058 = w7038 & w7039;
assign w7059 = w7036 & w7037;
assign w7060 = w7034 & w7035;
assign w7061 = w7032 & w7033;
assign w7062 = w7030 & w7031;
assign w7063 = w7028 & w7029;
assign w7064 = w7026 & w7027;
assign w7065 = w7024 & w7025;
assign w7066 = w7022 & w7023;
assign w7067 = w7020 & w7021;
assign w7068 = w7066 & w7067;
assign w7069 = w7064 & w7065;
assign w7070 = w7062 & w7063;
assign w7071 = w7060 & w7061;
assign w7072 = w7058 & w7059;
assign w7073 = w7056 & w7057;
assign w7074 = w7054 & w7055;
assign w7075 = w7052 & w7053;
assign w7076 = w7074 & w7075;
assign w7077 = w7072 & w7073;
assign w7078 = w7070 & w7071;
assign w7079 = w7068 & w7069;
assign w7080 = w7078 & w7079;
assign w7081 = w7076 & w7077;
assign w7082 = w7080 & w7081;
assign w7083 = ~pi10577 & ~w7082;
assign w7084 = pi03241 & w3326;
assign w7085 = pi05104 & w3266;
assign w7086 = pi06392 & w3418;
assign w7087 = pi05308 & w3236;
assign w7088 = pi02197 & w3112;
assign w7089 = pi05623 & w3272;
assign w7090 = pi01833 & w3179;
assign w7091 = pi05384 & w3496;
assign w7092 = pi05748 & w3194;
assign w7093 = pi05835 & w3207;
assign w7094 = pi03395 & w3122;
assign w7095 = pi01862 & w3528;
assign w7096 = pi09742 & w3382;
assign w7097 = pi03129 & w3118;
assign w7098 = pi05480 & w3300;
assign w7099 = pi05091 & w3232;
assign w7100 = pi05767 & w3171;
assign w7101 = pi02149 & w3356;
assign w7102 = pi03414 & w3162;
assign w7103 = pi05739 & w3600;
assign w7104 = pi03003 & w3292;
assign w7105 = pi09743 & w3544;
assign w7106 = pi06210 & w3188;
assign w7107 = pi09676 & w3336;
assign w7108 = pi05474 & w3506;
assign w7109 = pi05688 & w3312;
assign w7110 = pi02354 & w3554;
assign w7111 = pi05526 & w3572;
assign w7112 = pi05343 & w3129;
assign w7113 = pi05124 & w3436;
assign w7114 = pi05591 & w3254;
assign w7115 = pi01520 & w3520;
assign w7116 = pi05929 & w3474;
assign w7117 = pi05532 & w3340;
assign w7118 = pi03168 & w3522;
assign w7119 = pi05636 & w3358;
assign w7120 = pi09599 & w3530;
assign w7121 = pi05453 & w3442;
assign w7122 = pi03447 & w3177;
assign w7123 = pi05715 & w3372;
assign w7124 = pi05558 & w3420;
assign w7125 = pi05761 & w3430;
assign w7126 = pi05727 & w3374;
assign w7127 = pi02175 & w3217;
assign w7128 = pi05825 & w3464;
assign w7129 = pi02015 & w3314;
assign w7130 = pi03320 & w3370;
assign w7131 = pi05604 & w3472;
assign w7132 = pi01666 & w3546;
assign w7133 = pi09712 & w3268;
assign w7134 = pi05338 & w3203;
assign w7135 = pi09669 & w3125;
assign w7136 = pi09607 & w3064;
assign w7137 = pi03387 & w3258;
assign w7138 = pi09652 & w3362;
assign w7139 = pi01786 & w3390;
assign w7140 = pi02116 & w3586;
assign w7141 = pi02404 & w3508;
assign w7142 = pi05610 & w3221;
assign w7143 = pi01640 & w3514;
assign w7144 = pi05899 & w3093;
assign w7145 = pi03228 & w3290;
assign w7146 = pi02398 & w3342;
assign w7147 = pi05643 & w3448;
assign w7148 = pi06036 & w3594;
assign w7149 = pi01804 & w3360;
assign w7150 = pi01747 & w3264;
assign w7151 = pi06328 & w3578;
assign w7152 = pi02970 & w3536;
assign w7153 = pi01649 & w3246;
assign w7154 = pi02349 & w3452;
assign w7155 = pi09785 & w3078;
assign w7156 = pi05701 & w3165;
assign w7157 = pi05571 & w3364;
assign w7158 = pi06227 & w3580;
assign w7159 = pi05302 & w3450;
assign w7160 = pi03499 & w3488;
assign w7161 = pi05552 & w3410;
assign w7162 = pi03281 & w3115;
assign w7163 = pi05584 & w3205;
assign w7164 = pi03300 & w3484;
assign w7165 = pi03372 & w3169;
assign w7166 = pi03248 & w3334;
assign w7167 = pi05630 & w3376;
assign w7168 = pi05961 & w3175;
assign w7169 = pi05350 & w3199;
assign w7170 = pi03116 & w3394;
assign w7171 = pi05137 & w3598;
assign w7172 = pi05519 & w3406;
assign w7173 = pi09634 & w3404;
assign w7174 = pi03154 & w3428;
assign w7175 = pi05708 & w3201;
assign w7176 = pi05295 & w3538;
assign w7177 = pi05795 & w3192;
assign w7178 = pi05545 & w3552;
assign w7179 = pi05171 & w3252;
assign w7180 = pi06123 & w3282;
assign w7181 = pi01824 & w3422;
assign w7182 = pi06346 & w3438;
assign w7183 = pi06114 & w3478;
assign w7184 = pi05974 & w3223;
assign w7185 = pi03287 & w3190;
assign w7186 = pi05649 & w3566;
assign w7187 = pi03043 & w3490;
assign w7188 = pi05993 & w3446;
assign w7189 = pi05118 & w3308;
assign w7190 = pi02964 & w3274;
assign w7191 = pi05158 & w3492;
assign w7192 = pi06065 & w3584;
assign w7193 = pi02264 & w3288;
assign w7194 = pi01523 & w3346;
assign w7195 = pi02370 & w3167;
assign w7196 = pi03380 & w3302;
assign w7197 = pi03082 & w3348;
assign w7198 = pi03088 & w3456;
assign w7199 = pi03056 & w3350;
assign w7200 = pi05565 & w3135;
assign w7201 = pi03142 & w3494;
assign w7202 = pi05500 & w3466;
assign w7203 = pi02983 & w3296;
assign w7204 = pi06376 & w3524;
assign w7205 = pi01634 & w3270;
assign w7206 = pi05493 & w3234;
assign w7207 = pi09754 & w3408;
assign w7208 = pi02356 & w3219;
assign w7209 = pi06285 & w3324;
assign w7210 = pi09643 & w3238;
assign w7211 = pi09603 & w3322;
assign w7212 = pi03294 & w3328;
assign w7213 = pi06275 & w3316;
assign w7214 = pi05912 & w3426;
assign w7215 = pi05578 & w3156;
assign w7216 = pi03341 & w3412;
assign w7217 = pi02351 & w3440;
assign w7218 = pi06171 & w3280;
assign w7219 = pi03433 & w3556;
assign w7220 = pi06256 & w3148;
assign w7221 = pi02339 & w3550;
assign w7222 = pi01551 & w3306;
assign w7223 = pi05418 & w3186;
assign w7224 = pi05487 & w3398;
assign w7225 = pi05131 & w3248;
assign w7226 = pi03255 & w3214;
assign w7227 = pi03335 & w3512;
assign w7228 = pi03196 & w3502;
assign w7229 = pi06094 & w3444;
assign w7230 = pi03069 & w3209;
assign w7231 = pi06464 & w3242;
assign w7232 = pi05363 & w3227;
assign w7233 = pi03307 & w3146;
assign w7234 = pi06078 & w3106;
assign w7235 = pi06438 & w3558;
assign w7236 = pi05460 & w3384;
assign w7237 = pi03420 & w3504;
assign w7238 = pi03030 & w3244;
assign w7239 = pi02996 & w3262;
assign w7240 = pi05321 & w3354;
assign w7241 = pi03175 & w3181;
assign w7242 = pi03136 & w3574;
assign w7243 = pi05539 & w3286;
assign w7244 = pi03095 & w3592;
assign w7245 = pi09781 & w3197;
assign w7246 = pi09598 & w3103;
assign w7247 = pi05446 & w3518;
assign w7248 = pi05854 & w3386;
assign w7249 = pi05656 & w3276;
assign w7250 = pi02990 & w3137;
assign w7251 = pi06162 & w3542;
assign w7252 = pi05754 & w3590;
assign w7253 = pi05110 & w3143;
assign w7254 = pi03427 & w3184;
assign w7255 = pi02448 & w3229;
assign w7256 = pi06306 & w3158;
assign w7257 = pi02297 & w3366;
assign w7258 = pi05164 & w3612;
assign w7259 = pi06187 & w3096;
assign w7260 = pi06451 & w3510;
assign w7261 = pi09605 & w3400;
assign w7262 = pi03075 & w3338;
assign w7263 = pi05506 & w3127;
assign w7264 = pi06313 & w3602;
assign w7265 = pi02210 & w3480;
assign w7266 = pi06363 & w3160;
assign w7267 = pi03440 & w3388;
assign w7268 = pi06265 & w3294;
assign w7269 = pi02135 & w3460;
assign w7270 = pi03313 & w3564;
assign w7271 = pi06045 & w3468;
assign w7272 = pi01538 & w3380;
assign w7273 = pi03009 & w3260;
assign w7274 = pi09610 & w3534;
assign w7275 = pi03049 & w3526;
assign w7276 = pi05775 & w3476;
assign w7277 = pi05084 & w3486;
assign w7278 = pi06295 & w3332;
assign w7279 = pi06240 & w3560;
assign w7280 = pi05662 & w3434;
assign w7281 = pi02977 & w3424;
assign w7282 = pi02271 & w3568;
assign w7283 = pi01780 & w3368;
assign w7284 = pi05984 & w3606;
assign w7285 = pi05617 & w3620;
assign w7286 = pi05424 & w3284;
assign w7287 = pi05513 & w3139;
assign w7288 = pi09551 & w3516;
assign w7289 = pi03016 & w3610;
assign w7290 = pi05439 & w3256;
assign w7291 = pi02165 & w3086;
assign w7292 = pi06056 & w3173;
assign w7293 = pi02143 & w3378;
assign w7294 = pi05597 & w3225;
assign w7295 = pi05873 & w3352;
assign w7296 = pi05370 & w3304;
assign w7297 = pi03108 & w3132;
assign w7298 = pi03101 & w3498;
assign w7299 = pi05939 & w3532;
assign w7300 = pi03123 & w3071;
assign w7301 = pi06004 & w3570;
assign w7302 = pi03062 & w3576;
assign w7303 = pi05883 & w3596;
assign w7304 = pi05151 & w3344;
assign w7305 = pi06220 & w3402;
assign w7306 = pi02034 & w3482;
assign w7307 = pi05405 & w3278;
assign w7308 = pi05097 & w3240;
assign w7309 = pi09625 & w3250;
assign w7310 = pi05315 & w3298;
assign w7311 = pi06018 & w3608;
assign w7312 = pi06197 & w3318;
assign w7313 = pi02054 & w3414;
assign w7314 = pi03482 & w3582;
assign w7315 = pi05391 & w3153;
assign w7316 = pi03036 & w3548;
assign w7317 = pi09728 & w3500;
assign w7318 = pi01574 & w3614;
assign w7319 = pi05144 & w3604;
assign w7320 = pi03473 & w3211;
assign w7321 = pi03328 & w3618;
assign w7322 = pi06104 & w3320;
assign w7323 = pi03361 & w3562;
assign w7324 = pi02911 & w3330;
assign w7325 = pi05398 & w3082;
assign w7326 = pi03466 & w3396;
assign w7327 = pi03023 & w3310;
assign w7328 = pi05330 & w3392;
assign w7329 = pi03205 & w3454;
assign w7330 = pi05466 & w3432;
assign w7331 = pi03459 & w3588;
assign w7332 = pi01979 & w3540;
assign w7333 = pi06428 & w3150;
assign w7334 = pi01508 & w3110;
assign w7335 = pi09702 & w3416;
assign w7336 = pi09630 & w3470;
assign w7337 = pi01843 & w3458;
assign w7338 = pi05948 & w3616;
assign w7339 = pi05378 & w3462;
assign w7340 = ~w7084 & ~w7085;
assign w7341 = ~w7086 & ~w7087;
assign w7342 = ~w7088 & ~w7089;
assign w7343 = ~w7090 & ~w7091;
assign w7344 = ~w7092 & ~w7093;
assign w7345 = ~w7094 & ~w7095;
assign w7346 = ~w7096 & ~w7097;
assign w7347 = ~w7098 & ~w7099;
assign w7348 = ~w7100 & ~w7101;
assign w7349 = ~w7102 & ~w7103;
assign w7350 = ~w7104 & ~w7105;
assign w7351 = ~w7106 & ~w7107;
assign w7352 = ~w7108 & ~w7109;
assign w7353 = ~w7110 & ~w7111;
assign w7354 = ~w7112 & ~w7113;
assign w7355 = ~w7114 & ~w7115;
assign w7356 = ~w7116 & ~w7117;
assign w7357 = ~w7118 & ~w7119;
assign w7358 = ~w7120 & ~w7121;
assign w7359 = ~w7122 & ~w7123;
assign w7360 = ~w7124 & ~w7125;
assign w7361 = ~w7126 & ~w7127;
assign w7362 = ~w7128 & ~w7129;
assign w7363 = ~w7130 & ~w7131;
assign w7364 = ~w7132 & ~w7133;
assign w7365 = ~w7134 & ~w7135;
assign w7366 = ~w7136 & ~w7137;
assign w7367 = ~w7138 & ~w7139;
assign w7368 = ~w7140 & ~w7141;
assign w7369 = ~w7142 & ~w7143;
assign w7370 = ~w7144 & ~w7145;
assign w7371 = ~w7146 & ~w7147;
assign w7372 = ~w7148 & ~w7149;
assign w7373 = ~w7150 & ~w7151;
assign w7374 = ~w7152 & ~w7153;
assign w7375 = ~w7154 & ~w7155;
assign w7376 = ~w7156 & ~w7157;
assign w7377 = ~w7158 & ~w7159;
assign w7378 = ~w7160 & ~w7161;
assign w7379 = ~w7162 & ~w7163;
assign w7380 = ~w7164 & ~w7165;
assign w7381 = ~w7166 & ~w7167;
assign w7382 = ~w7168 & ~w7169;
assign w7383 = ~w7170 & ~w7171;
assign w7384 = ~w7172 & ~w7173;
assign w7385 = ~w7174 & ~w7175;
assign w7386 = ~w7176 & ~w7177;
assign w7387 = ~w7178 & ~w7179;
assign w7388 = ~w7180 & ~w7181;
assign w7389 = ~w7182 & ~w7183;
assign w7390 = ~w7184 & ~w7185;
assign w7391 = ~w7186 & ~w7187;
assign w7392 = ~w7188 & ~w7189;
assign w7393 = ~w7190 & ~w7191;
assign w7394 = ~w7192 & ~w7193;
assign w7395 = ~w7194 & ~w7195;
assign w7396 = ~w7196 & ~w7197;
assign w7397 = ~w7198 & ~w7199;
assign w7398 = ~w7200 & ~w7201;
assign w7399 = ~w7202 & ~w7203;
assign w7400 = ~w7204 & ~w7205;
assign w7401 = ~w7206 & ~w7207;
assign w7402 = ~w7208 & ~w7209;
assign w7403 = ~w7210 & ~w7211;
assign w7404 = ~w7212 & ~w7213;
assign w7405 = ~w7214 & ~w7215;
assign w7406 = ~w7216 & ~w7217;
assign w7407 = ~w7218 & ~w7219;
assign w7408 = ~w7220 & ~w7221;
assign w7409 = ~w7222 & ~w7223;
assign w7410 = ~w7224 & ~w7225;
assign w7411 = ~w7226 & ~w7227;
assign w7412 = ~w7228 & ~w7229;
assign w7413 = ~w7230 & ~w7231;
assign w7414 = ~w7232 & ~w7233;
assign w7415 = ~w7234 & ~w7235;
assign w7416 = ~w7236 & ~w7237;
assign w7417 = ~w7238 & ~w7239;
assign w7418 = ~w7240 & ~w7241;
assign w7419 = ~w7242 & ~w7243;
assign w7420 = ~w7244 & ~w7245;
assign w7421 = ~w7246 & ~w7247;
assign w7422 = ~w7248 & ~w7249;
assign w7423 = ~w7250 & ~w7251;
assign w7424 = ~w7252 & ~w7253;
assign w7425 = ~w7254 & ~w7255;
assign w7426 = ~w7256 & ~w7257;
assign w7427 = ~w7258 & ~w7259;
assign w7428 = ~w7260 & ~w7261;
assign w7429 = ~w7262 & ~w7263;
assign w7430 = ~w7264 & ~w7265;
assign w7431 = ~w7266 & ~w7267;
assign w7432 = ~w7268 & ~w7269;
assign w7433 = ~w7270 & ~w7271;
assign w7434 = ~w7272 & ~w7273;
assign w7435 = ~w7274 & ~w7275;
assign w7436 = ~w7276 & ~w7277;
assign w7437 = ~w7278 & ~w7279;
assign w7438 = ~w7280 & ~w7281;
assign w7439 = ~w7282 & ~w7283;
assign w7440 = ~w7284 & ~w7285;
assign w7441 = ~w7286 & ~w7287;
assign w7442 = ~w7288 & ~w7289;
assign w7443 = ~w7290 & ~w7291;
assign w7444 = ~w7292 & ~w7293;
assign w7445 = ~w7294 & ~w7295;
assign w7446 = ~w7296 & ~w7297;
assign w7447 = ~w7298 & ~w7299;
assign w7448 = ~w7300 & ~w7301;
assign w7449 = ~w7302 & ~w7303;
assign w7450 = ~w7304 & ~w7305;
assign w7451 = ~w7306 & ~w7307;
assign w7452 = ~w7308 & ~w7309;
assign w7453 = ~w7310 & ~w7311;
assign w7454 = ~w7312 & ~w7313;
assign w7455 = ~w7314 & ~w7315;
assign w7456 = ~w7316 & ~w7317;
assign w7457 = ~w7318 & ~w7319;
assign w7458 = ~w7320 & ~w7321;
assign w7459 = ~w7322 & ~w7323;
assign w7460 = ~w7324 & ~w7325;
assign w7461 = ~w7326 & ~w7327;
assign w7462 = ~w7328 & ~w7329;
assign w7463 = ~w7330 & ~w7331;
assign w7464 = ~w7332 & ~w7333;
assign w7465 = ~w7334 & ~w7335;
assign w7466 = ~w7336 & ~w7337;
assign w7467 = ~w7338 & ~w7339;
assign w7468 = w7466 & w7467;
assign w7469 = w7464 & w7465;
assign w7470 = w7462 & w7463;
assign w7471 = w7460 & w7461;
assign w7472 = w7458 & w7459;
assign w7473 = w7456 & w7457;
assign w7474 = w7454 & w7455;
assign w7475 = w7452 & w7453;
assign w7476 = w7450 & w7451;
assign w7477 = w7448 & w7449;
assign w7478 = w7446 & w7447;
assign w7479 = w7444 & w7445;
assign w7480 = w7442 & w7443;
assign w7481 = w7440 & w7441;
assign w7482 = w7438 & w7439;
assign w7483 = w7436 & w7437;
assign w7484 = w7434 & w7435;
assign w7485 = w7432 & w7433;
assign w7486 = w7430 & w7431;
assign w7487 = w7428 & w7429;
assign w7488 = w7426 & w7427;
assign w7489 = w7424 & w7425;
assign w7490 = w7422 & w7423;
assign w7491 = w7420 & w7421;
assign w7492 = w7418 & w7419;
assign w7493 = w7416 & w7417;
assign w7494 = w7414 & w7415;
assign w7495 = w7412 & w7413;
assign w7496 = w7410 & w7411;
assign w7497 = w7408 & w7409;
assign w7498 = w7406 & w7407;
assign w7499 = w7404 & w7405;
assign w7500 = w7402 & w7403;
assign w7501 = w7400 & w7401;
assign w7502 = w7398 & w7399;
assign w7503 = w7396 & w7397;
assign w7504 = w7394 & w7395;
assign w7505 = w7392 & w7393;
assign w7506 = w7390 & w7391;
assign w7507 = w7388 & w7389;
assign w7508 = w7386 & w7387;
assign w7509 = w7384 & w7385;
assign w7510 = w7382 & w7383;
assign w7511 = w7380 & w7381;
assign w7512 = w7378 & w7379;
assign w7513 = w7376 & w7377;
assign w7514 = w7374 & w7375;
assign w7515 = w7372 & w7373;
assign w7516 = w7370 & w7371;
assign w7517 = w7368 & w7369;
assign w7518 = w7366 & w7367;
assign w7519 = w7364 & w7365;
assign w7520 = w7362 & w7363;
assign w7521 = w7360 & w7361;
assign w7522 = w7358 & w7359;
assign w7523 = w7356 & w7357;
assign w7524 = w7354 & w7355;
assign w7525 = w7352 & w7353;
assign w7526 = w7350 & w7351;
assign w7527 = w7348 & w7349;
assign w7528 = w7346 & w7347;
assign w7529 = w7344 & w7345;
assign w7530 = w7342 & w7343;
assign w7531 = w7340 & w7341;
assign w7532 = w7530 & w7531;
assign w7533 = w7528 & w7529;
assign w7534 = w7526 & w7527;
assign w7535 = w7524 & w7525;
assign w7536 = w7522 & w7523;
assign w7537 = w7520 & w7521;
assign w7538 = w7518 & w7519;
assign w7539 = w7516 & w7517;
assign w7540 = w7514 & w7515;
assign w7541 = w7512 & w7513;
assign w7542 = w7510 & w7511;
assign w7543 = w7508 & w7509;
assign w7544 = w7506 & w7507;
assign w7545 = w7504 & w7505;
assign w7546 = w7502 & w7503;
assign w7547 = w7500 & w7501;
assign w7548 = w7498 & w7499;
assign w7549 = w7496 & w7497;
assign w7550 = w7494 & w7495;
assign w7551 = w7492 & w7493;
assign w7552 = w7490 & w7491;
assign w7553 = w7488 & w7489;
assign w7554 = w7486 & w7487;
assign w7555 = w7484 & w7485;
assign w7556 = w7482 & w7483;
assign w7557 = w7480 & w7481;
assign w7558 = w7478 & w7479;
assign w7559 = w7476 & w7477;
assign w7560 = w7474 & w7475;
assign w7561 = w7472 & w7473;
assign w7562 = w7470 & w7471;
assign w7563 = w7468 & w7469;
assign w7564 = w7562 & w7563;
assign w7565 = w7560 & w7561;
assign w7566 = w7558 & w7559;
assign w7567 = w7556 & w7557;
assign w7568 = w7554 & w7555;
assign w7569 = w7552 & w7553;
assign w7570 = w7550 & w7551;
assign w7571 = w7548 & w7549;
assign w7572 = w7546 & w7547;
assign w7573 = w7544 & w7545;
assign w7574 = w7542 & w7543;
assign w7575 = w7540 & w7541;
assign w7576 = w7538 & w7539;
assign w7577 = w7536 & w7537;
assign w7578 = w7534 & w7535;
assign w7579 = w7532 & w7533;
assign w7580 = w7578 & w7579;
assign w7581 = w7576 & w7577;
assign w7582 = w7574 & w7575;
assign w7583 = w7572 & w7573;
assign w7584 = w7570 & w7571;
assign w7585 = w7568 & w7569;
assign w7586 = w7566 & w7567;
assign w7587 = w7564 & w7565;
assign w7588 = w7586 & w7587;
assign w7589 = w7584 & w7585;
assign w7590 = w7582 & w7583;
assign w7591 = w7580 & w7581;
assign w7592 = w7590 & w7591;
assign w7593 = w7588 & w7589;
assign w7594 = w7592 & w7593;
assign w7595 = ~pi10577 & ~w7594;
assign w7596 = ~pi00365 & ~w6004;
assign w7597 = w6005 & ~w7596;
assign w7598 = ~pi00105 & w1121;
assign w7599 = ~w7597 & ~w7598;
assign w7600 = pi00465 & w1081;
assign w7601 = (w76 & w1081) | (w76 & w55707) | (w1081 & w55707);
assign w7602 = ~w7600 & w7601;
assign w7603 = pi05092 & w3232;
assign w7604 = pi03024 & w3310;
assign w7605 = pi09684 & w3398;
assign w7606 = pi02859 & w3336;
assign w7607 = pi09619 & w3286;
assign w7608 = pi05671 & w3508;
assign w7609 = pi09531 & w3188;
assign w7610 = pi02405 & w3606;
assign w7611 = pi02872 & w3500;
assign w7612 = pi06465 & w3242;
assign w7613 = pi02375 & w3612;
assign w7614 = pi05906 & w3238;
assign w7615 = pi06189 & w3096;
assign w7616 = pi02978 & w3424;
assign w7617 = pi05198 & w3528;
assign w7618 = pi05533 & w3340;
assign w7619 = pi03474 & w3211;
assign w7620 = pi05624 & w3272;
assign w7621 = pi05663 & w3434;
assign w7622 = pi02731 & w3620;
assign w7623 = pi02118 & w3258;
assign w7624 = pi05125 & w3436;
assign w7625 = pi03031 & w3244;
assign w7626 = pi03070 & w3209;
assign w7627 = pi05768 & w3171;
assign w7628 = pi05962 & w3175;
assign w7629 = pi06228 & w3580;
assign w7630 = pi05461 & w3384;
assign w7631 = pi03010 & w3260;
assign w7632 = pi05411 & w3514;
assign w7633 = pi03448 & w3177;
assign w7634 = pi02918 & w3530;
assign w7635 = pi06047 & w3468;
assign w7636 = pi05185 & w3554;
assign w7637 = pi03282 & w3115;
assign w7638 = pi06066 & w3584;
assign w7639 = pi03329 & w3618;
assign w7640 = pi06105 & w3320;
assign w7641 = pi05371 & w3304;
assign w7642 = pi06267 & w3294;
assign w7643 = pi05919 & w3516;
assign w7644 = pi02108 & w3162;
assign w7645 = pi05224 & w3480;
assign w7646 = pi05481 & w3300;
assign w7647 = pi05119 & w3308;
assign w7648 = pi02997 & w3262;
assign w7649 = pi06364 & w3160;
assign w7650 = pi06314 & w3602;
assign w7651 = pi06445 & w3408;
assign w7652 = pi05893 & w3125;
assign w7653 = pi05702 & w3165;
assign w7654 = pi05105 & w3266;
assign w7655 = pi06019 & w3608;
assign w7656 = pi03484 & w3582;
assign w7657 = pi05419 & w3186;
assign w7658 = pi05650 & w3566;
assign w7659 = pi03156 & w3428;
assign w7660 = pi02820 & w3614;
assign w7661 = pi06234 & w3229;
assign w7662 = pi03321 & w3370;
assign w7663 = pi06393 & w3418;
assign w7664 = pi06037 & w3594;
assign w7665 = pi05178 & w3219;
assign w7666 = pi09659 & w3466;
assign w7667 = pi02384 & w3446;
assign w7668 = pi05494 & w3234;
assign w7669 = pi05309 & w3236;
assign w7670 = pi05940 & w3532;
assign w7671 = pi03096 & w3592;
assign w7672 = pi06012 & w3440;
assign w7673 = pi02878 & w3268;
assign w7674 = pi05243 & w3378;
assign w7675 = pi02957 & w3103;
assign w7676 = pi05546 & w3552;
assign w7677 = pi03017 & w3610;
assign w7678 = pi03256 & w3214;
assign w7679 = pi09557 & w3318;
assign w7680 = pi05351 & w3199;
assign w7681 = pi06307 & w3158;
assign w7682 = pi01847 & w3129;
assign w7683 = pi06241 & w3560;
assign w7684 = pi05572 & w3364;
assign w7685 = pi05269 & w3414;
assign w7686 = pi06172 & w3280;
assign w7687 = pi05237 & w3112;
assign w7688 = pi02079 & w3396;
assign w7689 = pi05379 & w3462;
assign w7690 = pi02965 & w3274;
assign w7691 = pi03362 & w3562;
assign w7692 = pi03381 & w3302;
assign w7693 = pi02984 & w3296;
assign w7694 = pi02931 & w3064;
assign w7695 = pi06418 & w3110;
assign w7696 = pi06057 & w3173;
assign w7697 = pi05598 & w3225;
assign w7698 = pi09550 & w3135;
assign w7699 = pi05217 & w3288;
assign w7700 = pi05716 & w3372;
assign w7701 = pi05585 & w3205;
assign w7702 = pi03434 & w3556;
assign w7703 = pi03249 & w3334;
assign w7704 = pi05741 & w3600;
assign w7705 = pi09536 & w3474;
assign w7706 = pi06405 & w3246;
assign w7707 = pi02826 & w3306;
assign w7708 = pi05191 & w3452;
assign w7709 = pi03176 & w3181;
assign w7710 = pi09520 & w3156;
assign w7711 = pi03037 & w3548;
assign w7712 = pi02539 & w3616;
assign w7713 = pi02371 & w3148;
assign w7714 = pi03050 & w3526;
assign w7715 = pi06095 & w3444;
assign w7716 = pi03124 & w3071;
assign w7717 = pi02991 & w3137;
assign w7718 = pi05755 & w3590;
assign w7719 = pi05132 & w3248;
assign w7720 = pi03057 & w3350;
assign w7721 = pi05111 & w3143;
assign w7722 = pi03137 & w3574;
assign w7723 = pi05425 & w3284;
assign w7724 = pi05637 & w3358;
assign w7725 = pi05406 & w3278;
assign w7726 = pi03295 & w3328;
assign w7727 = pi03144 & w3494;
assign w7728 = pi05845 & w3270;
assign w7729 = pi05085 & w3486;
assign w7730 = pi05786 & w3458;
assign w7731 = pi01934 & w3392;
assign w7732 = pi03242 & w3326;
assign w7733 = pi05230 & w3217;
assign w7734 = pi02304 & w3324;
assign w7735 = pi02522 & w3448;
assign w7736 = pi03308 & w3146;
assign w7737 = pi09646 & w3572;
assign w7738 = pi03076 & w3338;
assign w7739 = pi02951 & w3322;
assign w7740 = pi02388 & w3344;
assign w7741 = pi06439 & w3558;
assign w7742 = pi05323 & w3354;
assign w7743 = pi03342 & w3412;
assign w7744 = pi03460 & w3588;
assign w7745 = pi02454 & w3276;
assign w7746 = pi02745 & w3472;
assign w7747 = pi05433 & w3078;
assign w7748 = pi01888 & w3430;
assign w7749 = pi06080 & w3106;
assign w7750 = pi05211 & w3568;
assign w7751 = pi03102 & w3498;
assign w7752 = pi05145 & w3604;
assign w7753 = pi05364 & w3227;
assign w7754 = pi05776 & w3476;
assign w7755 = pi05454 & w3442;
assign w7756 = pi02846 & w3520;
assign w7757 = pi05467 & w3432;
assign w7758 = pi06353 & w3368;
assign w7759 = pi05336 & w3203;
assign w7760 = pi03130 & w3118;
assign w7761 = pi05611 & w3221;
assign w7762 = pi03273 & w3086;
assign w7763 = pi02971 & w3536;
assign w7764 = pi02912 & w3330;
assign w7765 = pi02938 & w3534;
assign w7766 = pi05303 & w3450;
assign w7767 = pi05855 & w3386;
assign w7768 = pi06347 & w3438;
assign w7769 = pi02295 & w3201;
assign w7770 = pi06276 & w3316;
assign w7771 = pi05507 & w3127;
assign w7772 = pi06378 & w3524;
assign w7773 = pi05827 & w3464;
assign w7774 = pi05447 & w3518;
assign w7775 = pi02833 & w3380;
assign w7776 = pi05797 & w3192;
assign w7777 = pi05815 & w3390;
assign w7778 = pi03206 & w3454;
assign w7779 = pi05836 & w3207;
assign w7780 = pi09591 & w3410;
assign w7781 = pi05138 & w3598;
assign w7782 = pi09703 & w3506;
assign w7783 = pi06163 & w3542;
assign w7784 = pi06452 & w3510;
assign w7785 = pi05385 & w3496;
assign w7786 = pi03063 & w3576;
assign w7787 = pi05865 & w3382;
assign w7788 = pi05689 & w3312;
assign w7789 = pi02852 & w3197;
assign w7790 = pi05256 & w3460;
assign w7791 = pi02944 & w3400;
assign w7792 = pi03044 & w3490;
assign w7793 = pi03301 & w3484;
assign w7794 = pi02839 & w3346;
assign w7795 = pi05913 & w3426;
assign w7796 = pi06134 & w3264;
assign w7797 = pi06147 & w3546;
assign w7798 = pi05204 & w3550;
assign w7799 = pi02100 & w3184;
assign w7800 = pi06025 & w3366;
assign w7801 = pi03089 & w3456;
assign w7802 = pi05250 & w3356;
assign w7803 = pi05440 & w3256;
assign w7804 = pi06005 & w3570;
assign w7805 = pi02743 & w3254;
assign w7806 = pi03004 & w3292;
assign w7807 = pi05520 & w3406;
assign w7808 = pi03500 & w3488;
assign w7809 = pi06221 & w3402;
assign w7810 = pi03314 & w3564;
assign w7811 = pi06340 & w3179;
assign w7812 = pi06296 & w3332;
assign w7813 = pi03229 & w3290;
assign w7814 = pi02865 & w3544;
assign w7815 = pi02925 & w3250;
assign w7816 = pi02137 & w3512;
assign w7817 = pi05399 & w3082;
assign w7818 = pi02095 & w3388;
assign w7819 = pi05098 & w3240;
assign w7820 = pi06329 & w3578;
assign w7821 = pi01565 & w3376;
assign w7822 = pi03109 & w3132;
assign w7823 = pi06247 & w3342;
assign w7824 = pi06125 & w3282;
assign w7825 = pi05559 & w3420;
assign w7826 = pi02359 & w3252;
assign w7827 = pi05975 & w3223;
assign w7828 = pi05289 & w3314;
assign w7829 = pi03396 & w3122;
assign w7830 = pi05296 & w3538;
assign w7831 = pi02904 & w3404;
assign w7832 = pi02885 & w3416;
assign w7833 = pi05806 & w3360;
assign w7834 = pi05874 & w3352;
assign w7835 = pi02377 & w3492;
assign w7836 = pi03421 & w3504;
assign w7837 = pi05392 & w3153;
assign w7838 = pi05316 & w3298;
assign w7839 = pi03169 & w3522;
assign w7840 = pi05263 & w3586;
assign w7841 = pi05282 & w3482;
assign w7842 = pi05884 & w3596;
assign w7843 = pi06115 & w3478;
assign w7844 = pi03288 & w3190;
assign w7845 = pi09656 & w3139;
assign w7846 = pi02898 & w3362;
assign w7847 = pi05276 & w3540;
assign w7848 = pi05900 & w3093;
assign w7849 = pi05729 & w3374;
assign w7850 = pi03083 & w3348;
assign w7851 = pi03374 & w3169;
assign w7852 = pi01900 & w3194;
assign w7853 = pi02891 & w3470;
assign w7854 = pi03117 & w3394;
assign w7855 = pi05357 & w3422;
assign w7856 = pi05680 & w3167;
assign w7857 = pi03197 & w3502;
assign w7858 = pi06429 & w3150;
assign w7859 = ~w7603 & ~w7604;
assign w7860 = ~w7605 & ~w7606;
assign w7861 = ~w7607 & ~w7608;
assign w7862 = ~w7609 & ~w7610;
assign w7863 = ~w7611 & ~w7612;
assign w7864 = ~w7613 & ~w7614;
assign w7865 = ~w7615 & ~w7616;
assign w7866 = ~w7617 & ~w7618;
assign w7867 = ~w7619 & ~w7620;
assign w7868 = ~w7621 & ~w7622;
assign w7869 = ~w7623 & ~w7624;
assign w7870 = ~w7625 & ~w7626;
assign w7871 = ~w7627 & ~w7628;
assign w7872 = ~w7629 & ~w7630;
assign w7873 = ~w7631 & ~w7632;
assign w7874 = ~w7633 & ~w7634;
assign w7875 = ~w7635 & ~w7636;
assign w7876 = ~w7637 & ~w7638;
assign w7877 = ~w7639 & ~w7640;
assign w7878 = ~w7641 & ~w7642;
assign w7879 = ~w7643 & ~w7644;
assign w7880 = ~w7645 & ~w7646;
assign w7881 = ~w7647 & ~w7648;
assign w7882 = ~w7649 & ~w7650;
assign w7883 = ~w7651 & ~w7652;
assign w7884 = ~w7653 & ~w7654;
assign w7885 = ~w7655 & ~w7656;
assign w7886 = ~w7657 & ~w7658;
assign w7887 = ~w7659 & ~w7660;
assign w7888 = ~w7661 & ~w7662;
assign w7889 = ~w7663 & ~w7664;
assign w7890 = ~w7665 & ~w7666;
assign w7891 = ~w7667 & ~w7668;
assign w7892 = ~w7669 & ~w7670;
assign w7893 = ~w7671 & ~w7672;
assign w7894 = ~w7673 & ~w7674;
assign w7895 = ~w7675 & ~w7676;
assign w7896 = ~w7677 & ~w7678;
assign w7897 = ~w7679 & ~w7680;
assign w7898 = ~w7681 & ~w7682;
assign w7899 = ~w7683 & ~w7684;
assign w7900 = ~w7685 & ~w7686;
assign w7901 = ~w7687 & ~w7688;
assign w7902 = ~w7689 & ~w7690;
assign w7903 = ~w7691 & ~w7692;
assign w7904 = ~w7693 & ~w7694;
assign w7905 = ~w7695 & ~w7696;
assign w7906 = ~w7697 & ~w7698;
assign w7907 = ~w7699 & ~w7700;
assign w7908 = ~w7701 & ~w7702;
assign w7909 = ~w7703 & ~w7704;
assign w7910 = ~w7705 & ~w7706;
assign w7911 = ~w7707 & ~w7708;
assign w7912 = ~w7709 & ~w7710;
assign w7913 = ~w7711 & ~w7712;
assign w7914 = ~w7713 & ~w7714;
assign w7915 = ~w7715 & ~w7716;
assign w7916 = ~w7717 & ~w7718;
assign w7917 = ~w7719 & ~w7720;
assign w7918 = ~w7721 & ~w7722;
assign w7919 = ~w7723 & ~w7724;
assign w7920 = ~w7725 & ~w7726;
assign w7921 = ~w7727 & ~w7728;
assign w7922 = ~w7729 & ~w7730;
assign w7923 = ~w7731 & ~w7732;
assign w7924 = ~w7733 & ~w7734;
assign w7925 = ~w7735 & ~w7736;
assign w7926 = ~w7737 & ~w7738;
assign w7927 = ~w7739 & ~w7740;
assign w7928 = ~w7741 & ~w7742;
assign w7929 = ~w7743 & ~w7744;
assign w7930 = ~w7745 & ~w7746;
assign w7931 = ~w7747 & ~w7748;
assign w7932 = ~w7749 & ~w7750;
assign w7933 = ~w7751 & ~w7752;
assign w7934 = ~w7753 & ~w7754;
assign w7935 = ~w7755 & ~w7756;
assign w7936 = ~w7757 & ~w7758;
assign w7937 = ~w7759 & ~w7760;
assign w7938 = ~w7761 & ~w7762;
assign w7939 = ~w7763 & ~w7764;
assign w7940 = ~w7765 & ~w7766;
assign w7941 = ~w7767 & ~w7768;
assign w7942 = ~w7769 & ~w7770;
assign w7943 = ~w7771 & ~w7772;
assign w7944 = ~w7773 & ~w7774;
assign w7945 = ~w7775 & ~w7776;
assign w7946 = ~w7777 & ~w7778;
assign w7947 = ~w7779 & ~w7780;
assign w7948 = ~w7781 & ~w7782;
assign w7949 = ~w7783 & ~w7784;
assign w7950 = ~w7785 & ~w7786;
assign w7951 = ~w7787 & ~w7788;
assign w7952 = ~w7789 & ~w7790;
assign w7953 = ~w7791 & ~w7792;
assign w7954 = ~w7793 & ~w7794;
assign w7955 = ~w7795 & ~w7796;
assign w7956 = ~w7797 & ~w7798;
assign w7957 = ~w7799 & ~w7800;
assign w7958 = ~w7801 & ~w7802;
assign w7959 = ~w7803 & ~w7804;
assign w7960 = ~w7805 & ~w7806;
assign w7961 = ~w7807 & ~w7808;
assign w7962 = ~w7809 & ~w7810;
assign w7963 = ~w7811 & ~w7812;
assign w7964 = ~w7813 & ~w7814;
assign w7965 = ~w7815 & ~w7816;
assign w7966 = ~w7817 & ~w7818;
assign w7967 = ~w7819 & ~w7820;
assign w7968 = ~w7821 & ~w7822;
assign w7969 = ~w7823 & ~w7824;
assign w7970 = ~w7825 & ~w7826;
assign w7971 = ~w7827 & ~w7828;
assign w7972 = ~w7829 & ~w7830;
assign w7973 = ~w7831 & ~w7832;
assign w7974 = ~w7833 & ~w7834;
assign w7975 = ~w7835 & ~w7836;
assign w7976 = ~w7837 & ~w7838;
assign w7977 = ~w7839 & ~w7840;
assign w7978 = ~w7841 & ~w7842;
assign w7979 = ~w7843 & ~w7844;
assign w7980 = ~w7845 & ~w7846;
assign w7981 = ~w7847 & ~w7848;
assign w7982 = ~w7849 & ~w7850;
assign w7983 = ~w7851 & ~w7852;
assign w7984 = ~w7853 & ~w7854;
assign w7985 = ~w7855 & ~w7856;
assign w7986 = ~w7857 & ~w7858;
assign w7987 = w7985 & w7986;
assign w7988 = w7983 & w7984;
assign w7989 = w7981 & w7982;
assign w7990 = w7979 & w7980;
assign w7991 = w7977 & w7978;
assign w7992 = w7975 & w7976;
assign w7993 = w7973 & w7974;
assign w7994 = w7971 & w7972;
assign w7995 = w7969 & w7970;
assign w7996 = w7967 & w7968;
assign w7997 = w7965 & w7966;
assign w7998 = w7963 & w7964;
assign w7999 = w7961 & w7962;
assign w8000 = w7959 & w7960;
assign w8001 = w7957 & w7958;
assign w8002 = w7955 & w7956;
assign w8003 = w7953 & w7954;
assign w8004 = w7951 & w7952;
assign w8005 = w7949 & w7950;
assign w8006 = w7947 & w7948;
assign w8007 = w7945 & w7946;
assign w8008 = w7943 & w7944;
assign w8009 = w7941 & w7942;
assign w8010 = w7939 & w7940;
assign w8011 = w7937 & w7938;
assign w8012 = w7935 & w7936;
assign w8013 = w7933 & w7934;
assign w8014 = w7931 & w7932;
assign w8015 = w7929 & w7930;
assign w8016 = w7927 & w7928;
assign w8017 = w7925 & w7926;
assign w8018 = w7923 & w7924;
assign w8019 = w7921 & w7922;
assign w8020 = w7919 & w7920;
assign w8021 = w7917 & w7918;
assign w8022 = w7915 & w7916;
assign w8023 = w7913 & w7914;
assign w8024 = w7911 & w7912;
assign w8025 = w7909 & w7910;
assign w8026 = w7907 & w7908;
assign w8027 = w7905 & w7906;
assign w8028 = w7903 & w7904;
assign w8029 = w7901 & w7902;
assign w8030 = w7899 & w7900;
assign w8031 = w7897 & w7898;
assign w8032 = w7895 & w7896;
assign w8033 = w7893 & w7894;
assign w8034 = w7891 & w7892;
assign w8035 = w7889 & w7890;
assign w8036 = w7887 & w7888;
assign w8037 = w7885 & w7886;
assign w8038 = w7883 & w7884;
assign w8039 = w7881 & w7882;
assign w8040 = w7879 & w7880;
assign w8041 = w7877 & w7878;
assign w8042 = w7875 & w7876;
assign w8043 = w7873 & w7874;
assign w8044 = w7871 & w7872;
assign w8045 = w7869 & w7870;
assign w8046 = w7867 & w7868;
assign w8047 = w7865 & w7866;
assign w8048 = w7863 & w7864;
assign w8049 = w7861 & w7862;
assign w8050 = w7859 & w7860;
assign w8051 = w8049 & w8050;
assign w8052 = w8047 & w8048;
assign w8053 = w8045 & w8046;
assign w8054 = w8043 & w8044;
assign w8055 = w8041 & w8042;
assign w8056 = w8039 & w8040;
assign w8057 = w8037 & w8038;
assign w8058 = w8035 & w8036;
assign w8059 = w8033 & w8034;
assign w8060 = w8031 & w8032;
assign w8061 = w8029 & w8030;
assign w8062 = w8027 & w8028;
assign w8063 = w8025 & w8026;
assign w8064 = w8023 & w8024;
assign w8065 = w8021 & w8022;
assign w8066 = w8019 & w8020;
assign w8067 = w8017 & w8018;
assign w8068 = w8015 & w8016;
assign w8069 = w8013 & w8014;
assign w8070 = w8011 & w8012;
assign w8071 = w8009 & w8010;
assign w8072 = w8007 & w8008;
assign w8073 = w8005 & w8006;
assign w8074 = w8003 & w8004;
assign w8075 = w8001 & w8002;
assign w8076 = w7999 & w8000;
assign w8077 = w7997 & w7998;
assign w8078 = w7995 & w7996;
assign w8079 = w7993 & w7994;
assign w8080 = w7991 & w7992;
assign w8081 = w7989 & w7990;
assign w8082 = w7987 & w7988;
assign w8083 = w8081 & w8082;
assign w8084 = w8079 & w8080;
assign w8085 = w8077 & w8078;
assign w8086 = w8075 & w8076;
assign w8087 = w8073 & w8074;
assign w8088 = w8071 & w8072;
assign w8089 = w8069 & w8070;
assign w8090 = w8067 & w8068;
assign w8091 = w8065 & w8066;
assign w8092 = w8063 & w8064;
assign w8093 = w8061 & w8062;
assign w8094 = w8059 & w8060;
assign w8095 = w8057 & w8058;
assign w8096 = w8055 & w8056;
assign w8097 = w8053 & w8054;
assign w8098 = w8051 & w8052;
assign w8099 = w8097 & w8098;
assign w8100 = w8095 & w8096;
assign w8101 = w8093 & w8094;
assign w8102 = w8091 & w8092;
assign w8103 = w8089 & w8090;
assign w8104 = w8087 & w8088;
assign w8105 = w8085 & w8086;
assign w8106 = w8083 & w8084;
assign w8107 = w8105 & w8106;
assign w8108 = w8103 & w8104;
assign w8109 = w8101 & w8102;
assign w8110 = w8099 & w8100;
assign w8111 = w8109 & w8110;
assign w8112 = w8107 & w8108;
assign w8113 = w8111 & w8112;
assign w8114 = ~pi10577 & ~w8113;
assign w8115 = pi06235 & w3229;
assign w8116 = pi05605 & w3472;
assign w8117 = pi02992 & w3137;
assign w8118 = pi01489 & w3284;
assign w8119 = pi03131 & w3118;
assign w8120 = pi03336 & w3512;
assign w8121 = pi02966 & w3274;
assign w8122 = pi05579 & w3156;
assign w8123 = pi02979 & w3424;
assign w8124 = pi03415 & w3162;
assign w8125 = pi02214 & w3181;
assign w8126 = pi05199 & w3528;
assign w8127 = pi02190 & w3290;
assign w8128 = pi02827 & w3306;
assign w8129 = pi06430 & w3150;
assign w8130 = pi02932 & w3064;
assign w8131 = pi06173 & w3280;
assign w8132 = pi06308 & w3158;
assign w8133 = pi05749 & w3194;
assign w8134 = pi05152 & w3344;
assign w8135 = pi06466 & w3242;
assign w8136 = pi05159 & w3492;
assign w8137 = pi05212 & w3568;
assign w8138 = pi05644 & w3448;
assign w8139 = pi05468 & w3432;
assign w8140 = pi05372 & w3304;
assign w8141 = pi02985 & w3296;
assign w8142 = pi02461 & w3490;
assign w8143 = pi05756 & w3590;
assign w8144 = pi05310 & w3236;
assign w8145 = pi03011 & w3260;
assign w8146 = pi02401 & w3350;
assign w8147 = pi03441 & w3388;
assign w8148 = pi06096 & w3444;
assign w8149 = pi05251 & w3356;
assign w8150 = pi02130 & w3370;
assign w8151 = pi02148 & w3146;
assign w8152 = pi02860 & w3336;
assign w8153 = pi05534 & w3340;
assign w8154 = pi02316 & w3316;
assign w8155 = pi05930 & w3474;
assign w8156 = pi03018 & w3610;
assign w8157 = pi02399 & w3604;
assign w8158 = pi06453 & w3510;
assign w8159 = pi05816 & w3390;
assign w8160 = pi03467 & w3396;
assign w8161 = pi05337 & w3203;
assign w8162 = pi06287 & w3324;
assign w8163 = pi05651 & w3566;
assign w8164 = pi05270 & w3414;
assign w8165 = pi05172 & w3252;
assign w8166 = pi02305 & w3348;
assign w8167 = pi03157 & w3428;
assign w8168 = pi05901 & w3093;
assign w8169 = pi05553 & w3410;
assign w8170 = pi05672 & w3508;
assign w8171 = pi06190 & w3096;
assign w8172 = pi03388 & w3258;
assign w8173 = pi05488 & w3398;
assign w8174 = pi02343 & w3209;
assign w8175 = pi06394 & w3418;
assign w8176 = pi02734 & w3232;
assign w8177 = pi05482 & w3300;
assign w8178 = pi02840 & w3346;
assign w8179 = pi02905 & w3404;
assign w8180 = pi05238 & w3112;
assign w8181 = pi05331 & w3392;
assign w8182 = pi05742 & w3600;
assign w8183 = pi03501 & w3488;
assign w8184 = pi02919 & w3530;
assign w8185 = pi02517 & w3143;
assign w8186 = pi06211 & w3188;
assign w8187 = pi02240 & w3592;
assign w8188 = pi05573 & w3364;
assign w8189 = pi05995 & w3446;
assign w8190 = pi05777 & w3476;
assign w8191 = pi05218 & w3288;
assign w8192 = pi05638 & w3358;
assign w8193 = pi06135 & w3264;
assign w8194 = pi06365 & w3160;
assign w8195 = pi05304 & w3450;
assign w8196 = pi03475 & w3211;
assign w8197 = pi05283 & w3482;
assign w8198 = pi06058 & w3173;
assign w8199 = pi05769 & w3171;
assign w8200 = pi05441 & w3256;
assign w8201 = pi03198 & w3502;
assign w8202 = pi02181 & w3214;
assign w8203 = pi03051 & w3526;
assign w8204 = pi05894 & w3125;
assign w8205 = pi05501 & w3466;
assign w8206 = pi02415 & w3248;
assign w8207 = pi03330 & w3618;
assign w8208 = pi03103 & w3498;
assign w8209 = pi05186 & w3554;
assign w8210 = pi06348 & w3438;
assign w8211 = pi05179 & w3219;
assign w8212 = pi02847 & w3520;
assign w8213 = pi03274 & w3086;
assign w8214 = pi06026 & w3366;
assign w8215 = pi02737 & w3486;
assign w8216 = pi02420 & w3436;
assign w8217 = pi03025 & w3310;
assign w8218 = pi02263 & w3132;
assign w8219 = pi02879 & w3268;
assign w8220 = pi05941 & w3532;
assign w8221 = pi05976 & w3223;
assign w8222 = pi05875 & w3352;
assign w8223 = pi06406 & w3246;
assign w8224 = pi03302 & w3484;
assign w8225 = pi03207 & w3454;
assign w8226 = pi05586 & w3205;
assign w8227 = pi01633 & w3186;
assign w8228 = pi03461 & w3588;
assign w8229 = pi05787 & w3458;
assign w8230 = pi02547 & w3266;
assign w8231 = pi05514 & w3139;
assign w8232 = pi03077 & w3338;
assign w8233 = pi05365 & w3227;
assign w8234 = pi05244 & w3378;
assign w8235 = pi05914 & w3426;
assign w8236 = pi03449 & w3177;
assign w8237 = pi02866 & w3544;
assign w8238 = pi05475 & w3506;
assign w8239 = pi05625 & w3272;
assign w8240 = pi01733 & w3082;
assign w8241 = pi06067 & w3584;
assign w8242 = pi03485 & w3582;
assign w8243 = pi05448 & w3518;
assign w8244 = pi03397 & w3122;
assign w8245 = pi05866 & w3382;
assign w8246 = pi02972 & w3536;
assign w8247 = pi02939 & w3534;
assign w8248 = pi05592 & w3254;
assign w8249 = pi05527 & w3572;
assign w8250 = pi05717 & w3372;
assign w8251 = pi05920 & w3516;
assign w8252 = pi05690 & w3312;
assign w8253 = pi05324 & w3354;
assign w8254 = pi09713 & w3384;
assign w8255 = pi02124 & w3169;
assign w8256 = pi03289 & w3190;
assign w8257 = pi02892 & w3470;
assign w8258 = pi03038 & w3548;
assign w8259 = pi03422 & w3504;
assign w8260 = pi05257 & w3460;
assign w8261 = pi06198 & w3318;
assign w8262 = pi05434 & w3078;
assign w8263 = pi02352 & w3308;
assign w8264 = pi05703 & w3165;
assign w8265 = pi05949 & w3616;
assign w8266 = pi06164 & w3542;
assign w8267 = pi02886 & w3416;
assign w8268 = pi05264 & w3586;
assign w8269 = pi01745 & w3578;
assign w8270 = pi06268 & w3294;
assign w8271 = pi05599 & w3225;
assign w8272 = pi01863 & w3332;
assign w8273 = pi06248 & w3342;
assign w8274 = pi03064 & w3576;
assign w8275 = pi02998 & w3262;
assign w8276 = pi02958 & w3103;
assign w8277 = pi06229 & w3580;
assign w8278 = pi02913 & w3330;
assign w8279 = pi05521 & w3406;
assign w8280 = pi06341 & w3179;
assign w8281 = pi05508 & w3127;
assign w8282 = pi02251 & w3574;
assign w8283 = pi06006 & w3570;
assign w8284 = pi06446 & w3408;
assign w8285 = pi01903 & w3594;
assign w8286 = pi03428 & w3184;
assign w8287 = pi05165 & w3612;
assign w8288 = pi05837 & w3207;
assign w8289 = pi03343 & w3412;
assign w8290 = pi05231 & w3217;
assign w8291 = pi05566 & w3135;
assign w8292 = pi06148 & w3546;
assign w8293 = pi06419 & w3110;
assign w8294 = pi05455 & w3442;
assign w8295 = pi06315 & w3602;
assign w8296 = pi05380 & w3462;
assign w8297 = pi05358 & w3422;
assign w8298 = pi02899 & w3362;
assign w8299 = pi02257 & w3071;
assign w8300 = pi02408 & w3598;
assign w8301 = pi02834 & w3380;
assign w8302 = pi05612 & w3221;
assign w8303 = pi05225 & w3480;
assign w8304 = pi03250 & w3334;
assign w8305 = pi06257 & w3148;
assign w8306 = pi06106 & w3320;
assign w8307 = pi05664 & w3434;
assign w8308 = pi05856 & w3386;
assign w8309 = pi06242 & w3560;
assign w8310 = pi05297 & w3538;
assign w8311 = pi05807 & w3360;
assign w8312 = pi02952 & w3322;
assign w8313 = pi06116 & w3478;
assign w8314 = pi05985 & w3606;
assign w8315 = pi05317 & w3298;
assign w8316 = pi05412 & w3514;
assign w8317 = pi05540 & w3286;
assign w8318 = pi05495 & w3234;
assign w8319 = pi03170 & w3522;
assign w8320 = pi03435 & w3556;
assign w8321 = pi03118 & w3394;
assign w8322 = pi05205 & w3550;
assign w8323 = pi03145 & w3494;
assign w8324 = pi05631 & w3376;
assign w8325 = pi05709 & w3201;
assign w8326 = pi03315 & w3564;
assign w8327 = pi01703 & w3278;
assign w8328 = pi02527 & w3244;
assign w8329 = pi05393 & w3153;
assign w8330 = pi05192 & w3452;
assign w8331 = pi05618 & w3620;
assign w8332 = pi05846 & w3270;
assign w8333 = pi02873 & w3500;
assign w8334 = pi03090 & w3456;
assign w8335 = pi02150 & w3328;
assign w8336 = pi02945 & w3400;
assign w8337 = pi06440 & w3558;
assign w8338 = pi05560 & w3420;
assign w8339 = pi02821 & w3614;
assign w8340 = pi06222 & w3402;
assign w8341 = pi02613 & w3240;
assign w8342 = pi02163 & w3115;
assign w8343 = pi05344 & w3129;
assign w8344 = pi02926 & w3250;
assign w8345 = pi05386 & w3496;
assign w8346 = pi06126 & w3282;
assign w8347 = pi05730 & w3374;
assign w8348 = pi05963 & w3175;
assign w8349 = pi05352 & w3199;
assign w8350 = pi01794 & w3106;
assign w8351 = pi05657 & w3276;
assign w8352 = pi05907 & w3238;
assign w8353 = pi06020 & w3608;
assign w8354 = pi03005 & w3292;
assign w8355 = pi05885 & w3596;
assign w8356 = pi02853 & w3197;
assign w8357 = pi05290 & w3314;
assign w8358 = pi05798 & w3192;
assign w8359 = pi01608 & w3464;
assign w8360 = pi01894 & w3468;
assign w8361 = pi03382 & w3302;
assign w8362 = pi01686 & w3524;
assign w8363 = pi03363 & w3562;
assign w8364 = pi06013 & w3440;
assign w8365 = pi05547 & w3552;
assign w8366 = pi05277 & w3540;
assign w8367 = pi05681 & w3167;
assign w8368 = pi02186 & w3326;
assign w8369 = pi05762 & w3430;
assign w8370 = pi06354 & w3368;
assign w8371 = ~w8115 & ~w8116;
assign w8372 = ~w8117 & ~w8118;
assign w8373 = ~w8119 & ~w8120;
assign w8374 = ~w8121 & ~w8122;
assign w8375 = ~w8123 & ~w8124;
assign w8376 = ~w8125 & ~w8126;
assign w8377 = ~w8127 & ~w8128;
assign w8378 = ~w8129 & ~w8130;
assign w8379 = ~w8131 & ~w8132;
assign w8380 = ~w8133 & ~w8134;
assign w8381 = ~w8135 & ~w8136;
assign w8382 = ~w8137 & ~w8138;
assign w8383 = ~w8139 & ~w8140;
assign w8384 = ~w8141 & ~w8142;
assign w8385 = ~w8143 & ~w8144;
assign w8386 = ~w8145 & ~w8146;
assign w8387 = ~w8147 & ~w8148;
assign w8388 = ~w8149 & ~w8150;
assign w8389 = ~w8151 & ~w8152;
assign w8390 = ~w8153 & ~w8154;
assign w8391 = ~w8155 & ~w8156;
assign w8392 = ~w8157 & ~w8158;
assign w8393 = ~w8159 & ~w8160;
assign w8394 = ~w8161 & ~w8162;
assign w8395 = ~w8163 & ~w8164;
assign w8396 = ~w8165 & ~w8166;
assign w8397 = ~w8167 & ~w8168;
assign w8398 = ~w8169 & ~w8170;
assign w8399 = ~w8171 & ~w8172;
assign w8400 = ~w8173 & ~w8174;
assign w8401 = ~w8175 & ~w8176;
assign w8402 = ~w8177 & ~w8178;
assign w8403 = ~w8179 & ~w8180;
assign w8404 = ~w8181 & ~w8182;
assign w8405 = ~w8183 & ~w8184;
assign w8406 = ~w8185 & ~w8186;
assign w8407 = ~w8187 & ~w8188;
assign w8408 = ~w8189 & ~w8190;
assign w8409 = ~w8191 & ~w8192;
assign w8410 = ~w8193 & ~w8194;
assign w8411 = ~w8195 & ~w8196;
assign w8412 = ~w8197 & ~w8198;
assign w8413 = ~w8199 & ~w8200;
assign w8414 = ~w8201 & ~w8202;
assign w8415 = ~w8203 & ~w8204;
assign w8416 = ~w8205 & ~w8206;
assign w8417 = ~w8207 & ~w8208;
assign w8418 = ~w8209 & ~w8210;
assign w8419 = ~w8211 & ~w8212;
assign w8420 = ~w8213 & ~w8214;
assign w8421 = ~w8215 & ~w8216;
assign w8422 = ~w8217 & ~w8218;
assign w8423 = ~w8219 & ~w8220;
assign w8424 = ~w8221 & ~w8222;
assign w8425 = ~w8223 & ~w8224;
assign w8426 = ~w8225 & ~w8226;
assign w8427 = ~w8227 & ~w8228;
assign w8428 = ~w8229 & ~w8230;
assign w8429 = ~w8231 & ~w8232;
assign w8430 = ~w8233 & ~w8234;
assign w8431 = ~w8235 & ~w8236;
assign w8432 = ~w8237 & ~w8238;
assign w8433 = ~w8239 & ~w8240;
assign w8434 = ~w8241 & ~w8242;
assign w8435 = ~w8243 & ~w8244;
assign w8436 = ~w8245 & ~w8246;
assign w8437 = ~w8247 & ~w8248;
assign w8438 = ~w8249 & ~w8250;
assign w8439 = ~w8251 & ~w8252;
assign w8440 = ~w8253 & ~w8254;
assign w8441 = ~w8255 & ~w8256;
assign w8442 = ~w8257 & ~w8258;
assign w8443 = ~w8259 & ~w8260;
assign w8444 = ~w8261 & ~w8262;
assign w8445 = ~w8263 & ~w8264;
assign w8446 = ~w8265 & ~w8266;
assign w8447 = ~w8267 & ~w8268;
assign w8448 = ~w8269 & ~w8270;
assign w8449 = ~w8271 & ~w8272;
assign w8450 = ~w8273 & ~w8274;
assign w8451 = ~w8275 & ~w8276;
assign w8452 = ~w8277 & ~w8278;
assign w8453 = ~w8279 & ~w8280;
assign w8454 = ~w8281 & ~w8282;
assign w8455 = ~w8283 & ~w8284;
assign w8456 = ~w8285 & ~w8286;
assign w8457 = ~w8287 & ~w8288;
assign w8458 = ~w8289 & ~w8290;
assign w8459 = ~w8291 & ~w8292;
assign w8460 = ~w8293 & ~w8294;
assign w8461 = ~w8295 & ~w8296;
assign w8462 = ~w8297 & ~w8298;
assign w8463 = ~w8299 & ~w8300;
assign w8464 = ~w8301 & ~w8302;
assign w8465 = ~w8303 & ~w8304;
assign w8466 = ~w8305 & ~w8306;
assign w8467 = ~w8307 & ~w8308;
assign w8468 = ~w8309 & ~w8310;
assign w8469 = ~w8311 & ~w8312;
assign w8470 = ~w8313 & ~w8314;
assign w8471 = ~w8315 & ~w8316;
assign w8472 = ~w8317 & ~w8318;
assign w8473 = ~w8319 & ~w8320;
assign w8474 = ~w8321 & ~w8322;
assign w8475 = ~w8323 & ~w8324;
assign w8476 = ~w8325 & ~w8326;
assign w8477 = ~w8327 & ~w8328;
assign w8478 = ~w8329 & ~w8330;
assign w8479 = ~w8331 & ~w8332;
assign w8480 = ~w8333 & ~w8334;
assign w8481 = ~w8335 & ~w8336;
assign w8482 = ~w8337 & ~w8338;
assign w8483 = ~w8339 & ~w8340;
assign w8484 = ~w8341 & ~w8342;
assign w8485 = ~w8343 & ~w8344;
assign w8486 = ~w8345 & ~w8346;
assign w8487 = ~w8347 & ~w8348;
assign w8488 = ~w8349 & ~w8350;
assign w8489 = ~w8351 & ~w8352;
assign w8490 = ~w8353 & ~w8354;
assign w8491 = ~w8355 & ~w8356;
assign w8492 = ~w8357 & ~w8358;
assign w8493 = ~w8359 & ~w8360;
assign w8494 = ~w8361 & ~w8362;
assign w8495 = ~w8363 & ~w8364;
assign w8496 = ~w8365 & ~w8366;
assign w8497 = ~w8367 & ~w8368;
assign w8498 = ~w8369 & ~w8370;
assign w8499 = w8497 & w8498;
assign w8500 = w8495 & w8496;
assign w8501 = w8493 & w8494;
assign w8502 = w8491 & w8492;
assign w8503 = w8489 & w8490;
assign w8504 = w8487 & w8488;
assign w8505 = w8485 & w8486;
assign w8506 = w8483 & w8484;
assign w8507 = w8481 & w8482;
assign w8508 = w8479 & w8480;
assign w8509 = w8477 & w8478;
assign w8510 = w8475 & w8476;
assign w8511 = w8473 & w8474;
assign w8512 = w8471 & w8472;
assign w8513 = w8469 & w8470;
assign w8514 = w8467 & w8468;
assign w8515 = w8465 & w8466;
assign w8516 = w8463 & w8464;
assign w8517 = w8461 & w8462;
assign w8518 = w8459 & w8460;
assign w8519 = w8457 & w8458;
assign w8520 = w8455 & w8456;
assign w8521 = w8453 & w8454;
assign w8522 = w8451 & w8452;
assign w8523 = w8449 & w8450;
assign w8524 = w8447 & w8448;
assign w8525 = w8445 & w8446;
assign w8526 = w8443 & w8444;
assign w8527 = w8441 & w8442;
assign w8528 = w8439 & w8440;
assign w8529 = w8437 & w8438;
assign w8530 = w8435 & w8436;
assign w8531 = w8433 & w8434;
assign w8532 = w8431 & w8432;
assign w8533 = w8429 & w8430;
assign w8534 = w8427 & w8428;
assign w8535 = w8425 & w8426;
assign w8536 = w8423 & w8424;
assign w8537 = w8421 & w8422;
assign w8538 = w8419 & w8420;
assign w8539 = w8417 & w8418;
assign w8540 = w8415 & w8416;
assign w8541 = w8413 & w8414;
assign w8542 = w8411 & w8412;
assign w8543 = w8409 & w8410;
assign w8544 = w8407 & w8408;
assign w8545 = w8405 & w8406;
assign w8546 = w8403 & w8404;
assign w8547 = w8401 & w8402;
assign w8548 = w8399 & w8400;
assign w8549 = w8397 & w8398;
assign w8550 = w8395 & w8396;
assign w8551 = w8393 & w8394;
assign w8552 = w8391 & w8392;
assign w8553 = w8389 & w8390;
assign w8554 = w8387 & w8388;
assign w8555 = w8385 & w8386;
assign w8556 = w8383 & w8384;
assign w8557 = w8381 & w8382;
assign w8558 = w8379 & w8380;
assign w8559 = w8377 & w8378;
assign w8560 = w8375 & w8376;
assign w8561 = w8373 & w8374;
assign w8562 = w8371 & w8372;
assign w8563 = w8561 & w8562;
assign w8564 = w8559 & w8560;
assign w8565 = w8557 & w8558;
assign w8566 = w8555 & w8556;
assign w8567 = w8553 & w8554;
assign w8568 = w8551 & w8552;
assign w8569 = w8549 & w8550;
assign w8570 = w8547 & w8548;
assign w8571 = w8545 & w8546;
assign w8572 = w8543 & w8544;
assign w8573 = w8541 & w8542;
assign w8574 = w8539 & w8540;
assign w8575 = w8537 & w8538;
assign w8576 = w8535 & w8536;
assign w8577 = w8533 & w8534;
assign w8578 = w8531 & w8532;
assign w8579 = w8529 & w8530;
assign w8580 = w8527 & w8528;
assign w8581 = w8525 & w8526;
assign w8582 = w8523 & w8524;
assign w8583 = w8521 & w8522;
assign w8584 = w8519 & w8520;
assign w8585 = w8517 & w8518;
assign w8586 = w8515 & w8516;
assign w8587 = w8513 & w8514;
assign w8588 = w8511 & w8512;
assign w8589 = w8509 & w8510;
assign w8590 = w8507 & w8508;
assign w8591 = w8505 & w8506;
assign w8592 = w8503 & w8504;
assign w8593 = w8501 & w8502;
assign w8594 = w8499 & w8500;
assign w8595 = w8593 & w8594;
assign w8596 = w8591 & w8592;
assign w8597 = w8589 & w8590;
assign w8598 = w8587 & w8588;
assign w8599 = w8585 & w8586;
assign w8600 = w8583 & w8584;
assign w8601 = w8581 & w8582;
assign w8602 = w8579 & w8580;
assign w8603 = w8577 & w8578;
assign w8604 = w8575 & w8576;
assign w8605 = w8573 & w8574;
assign w8606 = w8571 & w8572;
assign w8607 = w8569 & w8570;
assign w8608 = w8567 & w8568;
assign w8609 = w8565 & w8566;
assign w8610 = w8563 & w8564;
assign w8611 = w8609 & w8610;
assign w8612 = w8607 & w8608;
assign w8613 = w8605 & w8606;
assign w8614 = w8603 & w8604;
assign w8615 = w8601 & w8602;
assign w8616 = w8599 & w8600;
assign w8617 = w8597 & w8598;
assign w8618 = w8595 & w8596;
assign w8619 = w8617 & w8618;
assign w8620 = w8615 & w8616;
assign w8621 = w8613 & w8614;
assign w8622 = w8611 & w8612;
assign w8623 = w8621 & w8622;
assign w8624 = w8619 & w8620;
assign w8625 = w8623 & w8624;
assign w8626 = ~pi10577 & ~w8625;
assign w8627 = pi02391 & w3606;
assign w8628 = pi06101 & w3320;
assign w8629 = pi02916 & w3530;
assign w8630 = pi02929 & w3064;
assign w8631 = pi05369 & w3304;
assign w8632 = pi03015 & w3610;
assign w8633 = pi02342 & w3490;
assign w8634 = pi03418 & w3504;
assign w8635 = pi02411 & w3598;
assign w8636 = pi03497 & w3488;
assign w8637 = pi05517 & w3406;
assign w8638 = pi05667 & w3508;
assign w8639 = pi06262 & w3294;
assign w8640 = pi05602 & w3472;
assign w8641 = pi05320 & w3354;
assign w8642 = pi02808 & w3310;
assign w8643 = pi05677 & w3167;
assign w8644 = pi02949 & w3322;
assign w8645 = pi09505 & w3242;
assign w8646 = pi03333 & w3512;
assign w8647 = pi05990 & w3446;
assign w8648 = pi02227 & w3522;
assign w8649 = pi03152 & w3428;
assign w8650 = pi03326 & w3618;
assign w8651 = pi06292 & w3332;
assign w8652 = pi05129 & w3248;
assign w8653 = pi06245 & w3342;
assign w8654 = pi02252 & w3118;
assign w8655 = pi05792 & w3192;
assign w8656 = pi05196 & w3528;
assign w8657 = pi05543 & w3552;
assign w8658 = pi02390 & w3223;
assign w8659 = pi02265 & w3132;
assign w8660 = pi05334 & w3203;
assign w8661 = pi03392 & w3122;
assign w8662 = pi06361 & w3160;
assign w8663 = pi05485 & w3398;
assign w8664 = pi03369 & w3169;
assign w8665 = pi05802 & w3360;
assign w8666 = pi01624 & w3284;
assign w8667 = pi05403 & w3278;
assign w8668 = pi03425 & w3184;
assign w8669 = pi05280 & w3482;
assign w8670 = pi05176 & w3219;
assign w8671 = pi02824 & w3306;
assign w8672 = pi02844 & w3520;
assign w8673 = pi05089 & w3232;
assign w8674 = pi06121 & w3282;
assign w8675 = pi09693 & w3318;
assign w8676 = pi02902 & w3404;
assign w8677 = pi05116 & w3308;
assign w8678 = pi05530 & w3340;
assign w8679 = pi03238 & w3326;
assign w8680 = pi05621 & w3272;
assign w8681 = pi02270 & w3592;
assign w8682 = pi02386 & w3526;
assign w8683 = pi05880 & w3596;
assign w8684 = pi02378 & w3338;
assign w8685 = pi03008 & w3260;
assign w8686 = pi05478 & w3300;
assign w8687 = pi02923 & w3250;
assign w8688 = pi02146 & w3370;
assign w8689 = pi06273 & w3316;
assign w8690 = pi05615 & w3620;
assign w8691 = pi02183 & w3334;
assign w8692 = pi06338 & w3179;
assign w8693 = pi03339 & w3412;
assign w8694 = pi02182 & w3214;
assign w8695 = pi03385 & w3258;
assign w8696 = pi02155 & w3484;
assign w8697 = pi06351 & w3368;
assign w8698 = pi02254 & w3574;
assign w8699 = pi02889 & w3470;
assign w8700 = pi05383 & w3496;
assign w8701 = pi06373 & w3524;
assign w8702 = pi03002 & w3292;
assign w8703 = pi05438 & w3256;
assign w8704 = pi03431 & w3556;
assign w8705 = pi02225 & w3181;
assign w8706 = pi06217 & w3402;
assign w8707 = pi05287 & w3314;
assign w8708 = pi05862 & w3382;
assign w8709 = pi05248 & w3356;
assign w8710 = pi05294 & w3538;
assign w8711 = pi09662 & w3280;
assign w8712 = pi06232 & w3229;
assign w8713 = pi02818 & w3614;
assign w8714 = pi05222 & w3480;
assign w8715 = pi02736 & w3240;
assign w8716 = pi05812 & w3390;
assign w8717 = pi05537 & w3286;
assign w8718 = pi03203 & w3454;
assign w8719 = pi06143 & w3546;
assign w8720 = pi05832 & w3207;
assign w8721 = pi02262 & w3394;
assign w8722 = pi05608 & w3221;
assign w8723 = pi02962 & w3274;
assign w8724 = pi02161 & w3328;
assign w8725 = pi05389 & w3153;
assign w8726 = pi02172 & w3086;
assign w8727 = pi02614 & w3616;
assign w8728 = pi05189 & w3452;
assign w8729 = pi02247 & w3494;
assign w8730 = pi09717 & w3384;
assign w8731 = pi02955 & w3103;
assign w8732 = pi03464 & w3396;
assign w8733 = pi02896 & w3362;
assign w8734 = pi05156 & w3492;
assign w8735 = pi05267 & w3414;
assign w8736 = pi05738 & w3600;
assign w8737 = pi05307 & w3236;
assign w8738 = pi05576 & w3156;
assign w8739 = pi05773 & w3476;
assign w8740 = pi06053 & w3173;
assign w8741 = pi02509 & w3175;
assign w8742 = pi02529 & w3143;
assign w8743 = pi06023 & w3366;
assign w8744 = pi03457 & w3588;
assign w8745 = pi05261 & w3586;
assign w8746 = pi05498 & w3466;
assign w8747 = pi03193 & w3502;
assign w8748 = pi05209 & w3568;
assign w8749 = pi02396 & w3576;
assign w8750 = pi09710 & w3432;
assign w8751 = pi02909 & w3330;
assign w8752 = pi02268 & w3498;
assign w8753 = pi02506 & w3548;
assign w8754 = pi02936 & w3534;
assign w8755 = pi05149 & w3344;
assign w8756 = pi02166 & w3115;
assign w8757 = pi05235 & w3112;
assign w8758 = pi06435 & w3558;
assign w8759 = pi02942 & w3400;
assign w8760 = pi05183 & w3554;
assign w8761 = pi06283 & w3324;
assign w8762 = pi05162 & w3612;
assign w8763 = pi05822 & w3464;
assign w8764 = pi05582 & w3205;
assign w8765 = pi05556 & w3420;
assign w8766 = pi05713 & w3372;
assign w8767 = pi03378 & w3302;
assign w8768 = pi05314 & w3298;
assign w8769 = pi09665 & w3096;
assign w8770 = pi02162 & w3190;
assign w8771 = pi05871 & w3352;
assign w8772 = pi05634 & w3358;
assign w8773 = pi03470 & w3211;
assign w8774 = pi06010 & w3440;
assign w8775 = pi05890 & w3125;
assign w8776 = pi06449 & w3510;
assign w8777 = pi05228 & w3217;
assign w8778 = pi02326 & w3456;
assign w8779 = pi02870 & w3500;
assign w8780 = pi02153 & w3146;
assign w8781 = pi02740 & w3486;
assign w8782 = pi05169 & w3252;
assign w8783 = pi06092 & w3444;
assign w8784 = pi06416 & w3110;
assign w8785 = pi05241 & w3378;
assign w8786 = pi05725 & w3374;
assign w8787 = pi06131 & w3264;
assign w8788 = pi02976 & w3424;
assign w8789 = pi06344 & w3438;
assign w8790 = pi05746 & w3194;
assign w8791 = pi02995 & w3262;
assign w8792 = pi03438 & w3388;
assign w8793 = pi02850 & w3197;
assign w8794 = pi02195 & w3290;
assign w8795 = pi06312 & w3602;
assign w8796 = pi05563 & w3135;
assign w8797 = pi05917 & w3516;
assign w8798 = pi02857 & w3336;
assign w8799 = pi05660 & w3434;
assign w8800 = pi06326 & w3578;
assign w8801 = pi01739 & w3082;
assign w8802 = pi02147 & w3564;
assign w8803 = pi05910 & w3426;
assign w8804 = pi05504 & w3127;
assign w8805 = pi05511 & w3139;
assign w8806 = pi06238 & w3560;
assign w8807 = pi05852 & w3386;
assign w8808 = pi02863 & w3544;
assign w8809 = pi05102 & w3266;
assign w8810 = pi05647 & w3566;
assign w8811 = pi06252 & w3148;
assign w8812 = pi05589 & w3254;
assign w8813 = pi02883 & w3416;
assign w8814 = pi05254 & w3460;
assign w8815 = pi09723 & w3442;
assign w8816 = pi05491 & w3234;
assign w8817 = pi02362 & w3570;
assign w8818 = pi05752 & w3590;
assign w8819 = pi05641 & w3448;
assign w8820 = pi05569 & w3364;
assign w8821 = pi05904 & w3238;
assign w8822 = pi06443 & w3408;
assign w8823 = pi06225 & w3580;
assign w8824 = pi05142 & w3604;
assign w8825 = pi05355 & w3422;
assign w8826 = pi05202 & w3550;
assign w8827 = pi02540 & w3244;
assign w8828 = pi02989 & w3137;
assign w8829 = pi05759 & w3430;
assign w8830 = pi05328 & w3392;
assign w8831 = pi06042 & w3468;
assign w8832 = pi05524 & w3572;
assign w8833 = pi05361 & w3227;
assign w8834 = pi05445 & w3518;
assign w8835 = pi03359 & w3562;
assign w8836 = pi06076 & w3106;
assign w8837 = pi02831 & w3380;
assign w8838 = pi01651 & w3514;
assign w8839 = pi09525 & w3188;
assign w8840 = pi02982 & w3296;
assign w8841 = pi05654 & w3276;
assign w8842 = pi05628 & w3376;
assign w8843 = pi05550 & w3410;
assign w8844 = pi06425 & w3150;
assign w8845 = pi05301 & w3450;
assign w8846 = pi02969 & w3536;
assign w8847 = pi02876 & w3268;
assign w8848 = pi02394 & w3209;
assign w8849 = pi02837 & w3346;
assign w8850 = pi03444 & w3177;
assign w8851 = pi06403 & w3246;
assign w8852 = pi05274 & w3540;
assign w8853 = pi05376 & w3462;
assign w8854 = pi05765 & w3171;
assign w8855 = pi09694 & w3506;
assign w8856 = pi02434 & w3436;
assign w8857 = pi06112 & w3478;
assign w8858 = pi05595 & w3225;
assign w8859 = pi02353 & w3348;
assign w8860 = pi02407 & w3350;
assign w8861 = pi05341 & w3129;
assign w8862 = pi05897 & w3093;
assign w8863 = pi05347 & w3199;
assign w8864 = pi05430 & w3078;
assign w8865 = pi05215 & w3288;
assign w8866 = pi05841 & w3270;
assign w8867 = pi02578 & w3542;
assign w8868 = pi03412 & w3162;
assign w8869 = pi02258 & w3071;
assign w8870 = pi02070 & w3582;
assign w8871 = pi05926 & w3474;
assign w8872 = pi05937 & w3532;
assign w8873 = pi02381 & w3312;
assign w8874 = pi05706 & w3201;
assign w8875 = pi06063 & w3584;
assign w8876 = pi06016 & w3608;
assign w8877 = pi06390 & w3418;
assign w8878 = pi06034 & w3594;
assign w8879 = pi05699 & w3165;
assign w8880 = pi05782 & w3458;
assign w8881 = pi06303 & w3158;
assign w8882 = pi05416 & w3186;
assign w8883 = ~w8627 & ~w8628;
assign w8884 = ~w8629 & ~w8630;
assign w8885 = ~w8631 & ~w8632;
assign w8886 = ~w8633 & ~w8634;
assign w8887 = ~w8635 & ~w8636;
assign w8888 = ~w8637 & ~w8638;
assign w8889 = ~w8639 & ~w8640;
assign w8890 = ~w8641 & ~w8642;
assign w8891 = ~w8643 & ~w8644;
assign w8892 = ~w8645 & ~w8646;
assign w8893 = ~w8647 & ~w8648;
assign w8894 = ~w8649 & ~w8650;
assign w8895 = ~w8651 & ~w8652;
assign w8896 = ~w8653 & ~w8654;
assign w8897 = ~w8655 & ~w8656;
assign w8898 = ~w8657 & ~w8658;
assign w8899 = ~w8659 & ~w8660;
assign w8900 = ~w8661 & ~w8662;
assign w8901 = ~w8663 & ~w8664;
assign w8902 = ~w8665 & ~w8666;
assign w8903 = ~w8667 & ~w8668;
assign w8904 = ~w8669 & ~w8670;
assign w8905 = ~w8671 & ~w8672;
assign w8906 = ~w8673 & ~w8674;
assign w8907 = ~w8675 & ~w8676;
assign w8908 = ~w8677 & ~w8678;
assign w8909 = ~w8679 & ~w8680;
assign w8910 = ~w8681 & ~w8682;
assign w8911 = ~w8683 & ~w8684;
assign w8912 = ~w8685 & ~w8686;
assign w8913 = ~w8687 & ~w8688;
assign w8914 = ~w8689 & ~w8690;
assign w8915 = ~w8691 & ~w8692;
assign w8916 = ~w8693 & ~w8694;
assign w8917 = ~w8695 & ~w8696;
assign w8918 = ~w8697 & ~w8698;
assign w8919 = ~w8699 & ~w8700;
assign w8920 = ~w8701 & ~w8702;
assign w8921 = ~w8703 & ~w8704;
assign w8922 = ~w8705 & ~w8706;
assign w8923 = ~w8707 & ~w8708;
assign w8924 = ~w8709 & ~w8710;
assign w8925 = ~w8711 & ~w8712;
assign w8926 = ~w8713 & ~w8714;
assign w8927 = ~w8715 & ~w8716;
assign w8928 = ~w8717 & ~w8718;
assign w8929 = ~w8719 & ~w8720;
assign w8930 = ~w8721 & ~w8722;
assign w8931 = ~w8723 & ~w8724;
assign w8932 = ~w8725 & ~w8726;
assign w8933 = ~w8727 & ~w8728;
assign w8934 = ~w8729 & ~w8730;
assign w8935 = ~w8731 & ~w8732;
assign w8936 = ~w8733 & ~w8734;
assign w8937 = ~w8735 & ~w8736;
assign w8938 = ~w8737 & ~w8738;
assign w8939 = ~w8739 & ~w8740;
assign w8940 = ~w8741 & ~w8742;
assign w8941 = ~w8743 & ~w8744;
assign w8942 = ~w8745 & ~w8746;
assign w8943 = ~w8747 & ~w8748;
assign w8944 = ~w8749 & ~w8750;
assign w8945 = ~w8751 & ~w8752;
assign w8946 = ~w8753 & ~w8754;
assign w8947 = ~w8755 & ~w8756;
assign w8948 = ~w8757 & ~w8758;
assign w8949 = ~w8759 & ~w8760;
assign w8950 = ~w8761 & ~w8762;
assign w8951 = ~w8763 & ~w8764;
assign w8952 = ~w8765 & ~w8766;
assign w8953 = ~w8767 & ~w8768;
assign w8954 = ~w8769 & ~w8770;
assign w8955 = ~w8771 & ~w8772;
assign w8956 = ~w8773 & ~w8774;
assign w8957 = ~w8775 & ~w8776;
assign w8958 = ~w8777 & ~w8778;
assign w8959 = ~w8779 & ~w8780;
assign w8960 = ~w8781 & ~w8782;
assign w8961 = ~w8783 & ~w8784;
assign w8962 = ~w8785 & ~w8786;
assign w8963 = ~w8787 & ~w8788;
assign w8964 = ~w8789 & ~w8790;
assign w8965 = ~w8791 & ~w8792;
assign w8966 = ~w8793 & ~w8794;
assign w8967 = ~w8795 & ~w8796;
assign w8968 = ~w8797 & ~w8798;
assign w8969 = ~w8799 & ~w8800;
assign w8970 = ~w8801 & ~w8802;
assign w8971 = ~w8803 & ~w8804;
assign w8972 = ~w8805 & ~w8806;
assign w8973 = ~w8807 & ~w8808;
assign w8974 = ~w8809 & ~w8810;
assign w8975 = ~w8811 & ~w8812;
assign w8976 = ~w8813 & ~w8814;
assign w8977 = ~w8815 & ~w8816;
assign w8978 = ~w8817 & ~w8818;
assign w8979 = ~w8819 & ~w8820;
assign w8980 = ~w8821 & ~w8822;
assign w8981 = ~w8823 & ~w8824;
assign w8982 = ~w8825 & ~w8826;
assign w8983 = ~w8827 & ~w8828;
assign w8984 = ~w8829 & ~w8830;
assign w8985 = ~w8831 & ~w8832;
assign w8986 = ~w8833 & ~w8834;
assign w8987 = ~w8835 & ~w8836;
assign w8988 = ~w8837 & ~w8838;
assign w8989 = ~w8839 & ~w8840;
assign w8990 = ~w8841 & ~w8842;
assign w8991 = ~w8843 & ~w8844;
assign w8992 = ~w8845 & ~w8846;
assign w8993 = ~w8847 & ~w8848;
assign w8994 = ~w8849 & ~w8850;
assign w8995 = ~w8851 & ~w8852;
assign w8996 = ~w8853 & ~w8854;
assign w8997 = ~w8855 & ~w8856;
assign w8998 = ~w8857 & ~w8858;
assign w8999 = ~w8859 & ~w8860;
assign w9000 = ~w8861 & ~w8862;
assign w9001 = ~w8863 & ~w8864;
assign w9002 = ~w8865 & ~w8866;
assign w9003 = ~w8867 & ~w8868;
assign w9004 = ~w8869 & ~w8870;
assign w9005 = ~w8871 & ~w8872;
assign w9006 = ~w8873 & ~w8874;
assign w9007 = ~w8875 & ~w8876;
assign w9008 = ~w8877 & ~w8878;
assign w9009 = ~w8879 & ~w8880;
assign w9010 = ~w8881 & ~w8882;
assign w9011 = w9009 & w9010;
assign w9012 = w9007 & w9008;
assign w9013 = w9005 & w9006;
assign w9014 = w9003 & w9004;
assign w9015 = w9001 & w9002;
assign w9016 = w8999 & w9000;
assign w9017 = w8997 & w8998;
assign w9018 = w8995 & w8996;
assign w9019 = w8993 & w8994;
assign w9020 = w8991 & w8992;
assign w9021 = w8989 & w8990;
assign w9022 = w8987 & w8988;
assign w9023 = w8985 & w8986;
assign w9024 = w8983 & w8984;
assign w9025 = w8981 & w8982;
assign w9026 = w8979 & w8980;
assign w9027 = w8977 & w8978;
assign w9028 = w8975 & w8976;
assign w9029 = w8973 & w8974;
assign w9030 = w8971 & w8972;
assign w9031 = w8969 & w8970;
assign w9032 = w8967 & w8968;
assign w9033 = w8965 & w8966;
assign w9034 = w8963 & w8964;
assign w9035 = w8961 & w8962;
assign w9036 = w8959 & w8960;
assign w9037 = w8957 & w8958;
assign w9038 = w8955 & w8956;
assign w9039 = w8953 & w8954;
assign w9040 = w8951 & w8952;
assign w9041 = w8949 & w8950;
assign w9042 = w8947 & w8948;
assign w9043 = w8945 & w8946;
assign w9044 = w8943 & w8944;
assign w9045 = w8941 & w8942;
assign w9046 = w8939 & w8940;
assign w9047 = w8937 & w8938;
assign w9048 = w8935 & w8936;
assign w9049 = w8933 & w8934;
assign w9050 = w8931 & w8932;
assign w9051 = w8929 & w8930;
assign w9052 = w8927 & w8928;
assign w9053 = w8925 & w8926;
assign w9054 = w8923 & w8924;
assign w9055 = w8921 & w8922;
assign w9056 = w8919 & w8920;
assign w9057 = w8917 & w8918;
assign w9058 = w8915 & w8916;
assign w9059 = w8913 & w8914;
assign w9060 = w8911 & w8912;
assign w9061 = w8909 & w8910;
assign w9062 = w8907 & w8908;
assign w9063 = w8905 & w8906;
assign w9064 = w8903 & w8904;
assign w9065 = w8901 & w8902;
assign w9066 = w8899 & w8900;
assign w9067 = w8897 & w8898;
assign w9068 = w8895 & w8896;
assign w9069 = w8893 & w8894;
assign w9070 = w8891 & w8892;
assign w9071 = w8889 & w8890;
assign w9072 = w8887 & w8888;
assign w9073 = w8885 & w8886;
assign w9074 = w8883 & w8884;
assign w9075 = w9073 & w9074;
assign w9076 = w9071 & w9072;
assign w9077 = w9069 & w9070;
assign w9078 = w9067 & w9068;
assign w9079 = w9065 & w9066;
assign w9080 = w9063 & w9064;
assign w9081 = w9061 & w9062;
assign w9082 = w9059 & w9060;
assign w9083 = w9057 & w9058;
assign w9084 = w9055 & w9056;
assign w9085 = w9053 & w9054;
assign w9086 = w9051 & w9052;
assign w9087 = w9049 & w9050;
assign w9088 = w9047 & w9048;
assign w9089 = w9045 & w9046;
assign w9090 = w9043 & w9044;
assign w9091 = w9041 & w9042;
assign w9092 = w9039 & w9040;
assign w9093 = w9037 & w9038;
assign w9094 = w9035 & w9036;
assign w9095 = w9033 & w9034;
assign w9096 = w9031 & w9032;
assign w9097 = w9029 & w9030;
assign w9098 = w9027 & w9028;
assign w9099 = w9025 & w9026;
assign w9100 = w9023 & w9024;
assign w9101 = w9021 & w9022;
assign w9102 = w9019 & w9020;
assign w9103 = w9017 & w9018;
assign w9104 = w9015 & w9016;
assign w9105 = w9013 & w9014;
assign w9106 = w9011 & w9012;
assign w9107 = w9105 & w9106;
assign w9108 = w9103 & w9104;
assign w9109 = w9101 & w9102;
assign w9110 = w9099 & w9100;
assign w9111 = w9097 & w9098;
assign w9112 = w9095 & w9096;
assign w9113 = w9093 & w9094;
assign w9114 = w9091 & w9092;
assign w9115 = w9089 & w9090;
assign w9116 = w9087 & w9088;
assign w9117 = w9085 & w9086;
assign w9118 = w9083 & w9084;
assign w9119 = w9081 & w9082;
assign w9120 = w9079 & w9080;
assign w9121 = w9077 & w9078;
assign w9122 = w9075 & w9076;
assign w9123 = w9121 & w9122;
assign w9124 = w9119 & w9120;
assign w9125 = w9117 & w9118;
assign w9126 = w9115 & w9116;
assign w9127 = w9113 & w9114;
assign w9128 = w9111 & w9112;
assign w9129 = w9109 & w9110;
assign w9130 = w9107 & w9108;
assign w9131 = w9129 & w9130;
assign w9132 = w9127 & w9128;
assign w9133 = w9125 & w9126;
assign w9134 = w9123 & w9124;
assign w9135 = w9133 & w9134;
assign w9136 = w9131 & w9132;
assign w9137 = w9135 & w9136;
assign w9138 = ~pi10577 & ~w9137;
assign w9139 = pi06161 & w3542;
assign w9140 = pi06218 & w3402;
assign w9141 = pi03299 & w3484;
assign w9142 = pi06002 & w3570;
assign w9143 = pi03312 & w3564;
assign w9144 = pi03141 & w3494;
assign w9145 = pi05833 & w3207;
assign w9146 = pi01756 & w3160;
assign w9147 = pi03081 & w3348;
assign w9148 = pi03035 & w3548;
assign w9149 = pi03029 & w3244;
assign w9150 = pi05452 & w3442;
assign w9151 = pi05616 & w3620;
assign w9152 = pi05130 & w3248;
assign w9153 = pi06391 & w3418;
assign w9154 = pi05190 & w3452;
assign w9155 = pi02877 & w3268;
assign w9156 = pi06293 & w3332;
assign w9157 = pi06352 & w3368;
assign w9158 = pi05774 & w3476;
assign w9159 = pi05853 & w3386;
assign w9160 = pi02832 & w3380;
assign w9161 = pi05177 & w3219;
assign w9162 = pi05223 & w3480;
assign w9163 = pi06462 & w3242;
assign w9164 = pi09579 & w3296;
assign w9165 = pi02858 & w3336;
assign w9166 = pi03498 & w3488;
assign w9167 = pi02838 & w3346;
assign w9168 = pi05262 & w3586;
assign w9169 = pi05242 & w3378;
assign w9170 = pi06246 & w3342;
assign w9171 = pi05960 & w3175;
assign w9172 = pi05512 & w3139;
assign w9173 = pi05281 & w3482;
assign w9174 = pi05275 & w3540;
assign w9175 = pi02903 & w3404;
assign w9176 = pi05700 & w3165;
assign w9177 = pi03340 & w3412;
assign w9178 = pi05793 & w3192;
assign w9179 = pi05669 & w3508;
assign w9180 = pi05928 & w3474;
assign w9181 = pi09586 & w3536;
assign w9182 = pi05109 & w3143;
assign w9183 = pi05982 & w3606;
assign w9184 = pi05117 & w3308;
assign w9185 = pi02825 & w3306;
assign w9186 = pi03094 & w3592;
assign w9187 = pi02890 & w3470;
assign w9188 = pi03413 & w3162;
assign w9189 = pi05947 & w3616;
assign w9190 = pi05726 & w3374;
assign w9191 = pi05655 & w3276;
assign w9192 = pi05577 & w3156;
assign w9193 = pi01865 & w3594;
assign w9194 = pi05824 & w3464;
assign w9195 = pi03042 & w3490;
assign w9196 = pi05622 & w3272;
assign w9197 = pi05417 & w3186;
assign w9198 = pi05197 & w3528;
assign w9199 = pi03386 & w3258;
assign w9200 = pi05492 & w3234;
assign w9201 = pi09535 & w3260;
assign w9202 = pi05629 & w3376;
assign w9203 = pi09566 & w3262;
assign w9204 = pi05918 & w3516;
assign w9205 = pi09705 & w3596;
assign w9206 = pi02008 & w3538;
assign w9207 = pi05096 & w3240;
assign w9208 = pi06284 & w3324;
assign w9209 = pi05410 & w3514;
assign w9210 = pi05157 & w3492;
assign w9211 = pi05163 & w3612;
assign w9212 = pi05590 & w3254;
assign w9213 = pi03371 & w3169;
assign w9214 = pi03379 & w3302;
assign w9215 = pi06103 & w3320;
assign w9216 = pi03471 & w3211;
assign w9217 = pi06132 & w3264;
assign w9218 = pi03458 & w3588;
assign w9219 = pi05551 & w3410;
assign w9220 = pi03135 & w3574;
assign w9221 = pi03061 & w3576;
assign w9222 = pi06404 & w3246;
assign w9223 = pi05362 & w3227;
assign w9224 = pi03174 & w3181;
assign w9225 = pi05505 & w3127;
assign w9226 = pi06417 & w3110;
assign w9227 = pi05583 & w3205;
assign w9228 = pi02884 & w3416;
assign w9229 = pi03194 & w3502;
assign w9230 = pi06444 & w3408;
assign w9231 = pi05570 & w3364;
assign w9232 = pi03115 & w3394;
assign w9233 = pi02864 & w3544;
assign w9234 = pi03254 & w3214;
assign w9235 = pi05564 & w3135;
assign w9236 = pi02819 & w3614;
assign w9237 = pi01881 & w3584;
assign w9238 = pi05973 & w3223;
assign w9239 = pi01867 & w3578;
assign w9240 = pi03293 & w3328;
assign w9241 = pi03100 & w3498;
assign w9242 = pi03360 & w3562;
assign w9243 = pi05707 & w3201;
assign w9244 = pi05538 & w3286;
assign w9245 = pi05397 & w3082;
assign w9246 = pi05249 & w3356;
assign w9247 = pi05898 & w3093;
assign w9248 = pi02845 & w3520;
assign w9249 = pi05635 & w3358;
assign w9250 = pi02937 & w3534;
assign w9251 = pi05150 & w3344;
assign w9252 = pi05911 & w3426;
assign w9253 = pi05083 & w3486;
assign w9254 = pi05479 & w3300;
assign w9255 = pi06017 & w3608;
assign w9256 = pi06233 & w3229;
assign w9257 = pi05473 & w3506;
assign w9258 = pi01972 & w3236;
assign w9259 = pi02323 & w3316;
assign w9260 = pi06264 & w3294;
assign w9261 = pi01501 & w3106;
assign w9262 = pi06024 & w3366;
assign w9263 = pi06450 & w3510;
assign w9264 = pi05747 & w3194;
assign w9265 = pi05377 & w3462;
assign w9266 = pi05216 & w3288;
assign w9267 = pi03426 & w3184;
assign w9268 = pi01893 & w3173;
assign w9269 = pi06436 & w3558;
assign w9270 = pi03445 & w3177;
assign w9271 = pi01952 & w3298;
assign w9272 = pi03247 & w3334;
assign w9273 = pi09660 & w3518;
assign w9274 = pi05661 & w3434;
assign w9275 = pi05356 & w3422;
assign w9276 = pi03465 & w3396;
assign w9277 = pi01783 & w3496;
assign w9278 = pi05268 & w3414;
assign w9279 = pi05557 & w3420;
assign w9280 = pi03439 & w3388;
assign w9281 = pi03074 & w3338;
assign w9282 = pi05170 & w3252;
assign w9283 = pi06011 & w3440;
assign w9284 = pi05229 & w3217;
assign w9285 = pi05766 & w3171;
assign w9286 = pi01693 & w3524;
assign w9287 = pi06054 & w3610;
assign w9288 = pi05609 & w3221;
assign w9289 = pi05465 & w3432;
assign w9290 = pi03128 & w3118;
assign w9291 = pi09585 & w3274;
assign w9292 = pi05210 & w3568;
assign w9293 = pi02943 & w3400;
assign w9294 = pi05784 & w3458;
assign w9295 = pi03107 & w3132;
assign w9296 = pi03022 & w3310;
assign w9297 = pi09546 & w3137;
assign w9298 = pi03068 & w3209;
assign w9299 = pi05872 & w3352;
assign w9300 = pi03481 & w3582;
assign w9301 = pi06170 & w3280;
assign w9302 = pi03167 & w3522;
assign w9303 = pi05518 & w3406;
assign w9304 = pi02930 & w3064;
assign w9305 = pi06427 & w3150;
assign w9306 = pi02950 & w3322;
assign w9307 = pi05390 & w3153;
assign w9308 = pi05938 & w3532;
assign w9309 = pi01806 & w3304;
assign w9310 = pi03087 & w3456;
assign w9311 = pi05123 & w3436;
assign w9312 = pi05753 & w3590;
assign w9313 = pi05678 & w3167;
assign w9314 = pi06345 & w3438;
assign w9315 = pi06304 & w3158;
assign w9316 = pi05459 & w3384;
assign w9317 = pi05136 & w3598;
assign w9318 = pi09559 & w3292;
assign w9319 = pi06186 & w3096;
assign w9320 = pi05525 & w3572;
assign w9321 = pi05648 & w3566;
assign w9322 = pi03122 & w3071;
assign w9323 = pi05804 & w3360;
assign w9324 = pi02188 & w3326;
assign w9325 = pi06339 & w3179;
assign w9326 = pi01889 & w3602;
assign w9327 = pi06144 & w3546;
assign w9328 = pi03048 & w3526;
assign w9329 = pi02871 & w3500;
assign w9330 = pi05432 & w3078;
assign w9331 = pi05486 & w3398;
assign w9332 = pi02234 & w3428;
assign w9333 = pi05891 & w3125;
assign w9334 = pi05760 & w3430;
assign w9335 = pi03055 & w3350;
assign w9336 = pi05603 & w3472;
assign w9337 = pi05342 & w3129;
assign w9338 = pi06208 & w3188;
assign w9339 = pi03419 & w3504;
assign w9340 = pi05714 & w3372;
assign w9341 = pi02897 & w3362;
assign w9342 = pi05203 & w3550;
assign w9343 = pi05687 & w3312;
assign w9344 = pi05531 & w3340;
assign w9345 = pi05992 & w3446;
assign w9346 = pi02917 & w3530;
assign w9347 = pi03306 & w3146;
assign w9348 = pi03334 & w3512;
assign w9349 = pi02924 & w3250;
assign w9350 = pi06226 & w3580;
assign w9351 = pi05184 & w3554;
assign w9352 = pi05905 & w3238;
assign w9353 = pi05255 & w3460;
assign w9354 = pi03393 & w3122;
assign w9355 = pi05236 & w3112;
assign w9356 = pi06093 & w3444;
assign w9357 = pi05499 & w3466;
assign w9358 = pi03319 & w3370;
assign w9359 = pi05843 & w3270;
assign w9360 = pi02851 & w3197;
assign w9361 = pi03327 & w3618;
assign w9362 = pi06044 & w3468;
assign w9363 = pi03227 & w3290;
assign w9364 = pi05143 & w3604;
assign w9365 = pi05596 & w3225;
assign w9366 = pi03271 & w3086;
assign w9367 = pi09582 & w3424;
assign w9368 = pi09739 & w3256;
assign w9369 = pi01948 & w3354;
assign w9370 = pi05642 & w3448;
assign w9371 = pi06253 & w3148;
assign w9372 = pi05404 & w3278;
assign w9373 = pi05349 & w3199;
assign w9374 = pi05813 & w3390;
assign w9375 = pi06122 & w3282;
assign w9376 = pi03286 & w3190;
assign w9377 = pi01992 & w3450;
assign w9378 = pi06195 & w3318;
assign w9379 = pi05863 & w3382;
assign w9380 = pi06239 & w3560;
assign w9381 = pi01975 & w3600;
assign w9382 = pi03432 & w3556;
assign w9383 = pi05329 & w3392;
assign w9384 = pi03280 & w3115;
assign w9385 = pi03204 & w3454;
assign w9386 = pi06113 & w3478;
assign w9387 = pi05544 & w3552;
assign w9388 = pi05423 & w3284;
assign w9389 = pi05288 & w3314;
assign w9390 = pi05090 & w3232;
assign w9391 = pi05103 & w3266;
assign w9392 = pi02910 & w3330;
assign w9393 = pi05335 & w3203;
assign w9394 = pi02956 & w3103;
assign w9395 = ~w9139 & ~w9140;
assign w9396 = ~w9141 & ~w9142;
assign w9397 = ~w9143 & ~w9144;
assign w9398 = ~w9145 & ~w9146;
assign w9399 = ~w9147 & ~w9148;
assign w9400 = ~w9149 & ~w9150;
assign w9401 = ~w9151 & ~w9152;
assign w9402 = ~w9153 & ~w9154;
assign w9403 = ~w9155 & ~w9156;
assign w9404 = ~w9157 & ~w9158;
assign w9405 = ~w9159 & ~w9160;
assign w9406 = ~w9161 & ~w9162;
assign w9407 = ~w9163 & ~w9164;
assign w9408 = ~w9165 & ~w9166;
assign w9409 = ~w9167 & ~w9168;
assign w9410 = ~w9169 & ~w9170;
assign w9411 = ~w9171 & ~w9172;
assign w9412 = ~w9173 & ~w9174;
assign w9413 = ~w9175 & ~w9176;
assign w9414 = ~w9177 & ~w9178;
assign w9415 = ~w9179 & ~w9180;
assign w9416 = ~w9181 & ~w9182;
assign w9417 = ~w9183 & ~w9184;
assign w9418 = ~w9185 & ~w9186;
assign w9419 = ~w9187 & ~w9188;
assign w9420 = ~w9189 & ~w9190;
assign w9421 = ~w9191 & ~w9192;
assign w9422 = ~w9193 & ~w9194;
assign w9423 = ~w9195 & ~w9196;
assign w9424 = ~w9197 & ~w9198;
assign w9425 = ~w9199 & ~w9200;
assign w9426 = ~w9201 & ~w9202;
assign w9427 = ~w9203 & ~w9204;
assign w9428 = ~w9205 & ~w9206;
assign w9429 = ~w9207 & ~w9208;
assign w9430 = ~w9209 & ~w9210;
assign w9431 = ~w9211 & ~w9212;
assign w9432 = ~w9213 & ~w9214;
assign w9433 = ~w9215 & ~w9216;
assign w9434 = ~w9217 & ~w9218;
assign w9435 = ~w9219 & ~w9220;
assign w9436 = ~w9221 & ~w9222;
assign w9437 = ~w9223 & ~w9224;
assign w9438 = ~w9225 & ~w9226;
assign w9439 = ~w9227 & ~w9228;
assign w9440 = ~w9229 & ~w9230;
assign w9441 = ~w9231 & ~w9232;
assign w9442 = ~w9233 & ~w9234;
assign w9443 = ~w9235 & ~w9236;
assign w9444 = ~w9237 & ~w9238;
assign w9445 = ~w9239 & ~w9240;
assign w9446 = ~w9241 & ~w9242;
assign w9447 = ~w9243 & ~w9244;
assign w9448 = ~w9245 & ~w9246;
assign w9449 = ~w9247 & ~w9248;
assign w9450 = ~w9249 & ~w9250;
assign w9451 = ~w9251 & ~w9252;
assign w9452 = ~w9253 & ~w9254;
assign w9453 = ~w9255 & ~w9256;
assign w9454 = ~w9257 & ~w9258;
assign w9455 = ~w9259 & ~w9260;
assign w9456 = ~w9261 & ~w9262;
assign w9457 = ~w9263 & ~w9264;
assign w9458 = ~w9265 & ~w9266;
assign w9459 = ~w9267 & ~w9268;
assign w9460 = ~w9269 & ~w9270;
assign w9461 = ~w9271 & ~w9272;
assign w9462 = ~w9273 & ~w9274;
assign w9463 = ~w9275 & ~w9276;
assign w9464 = ~w9277 & ~w9278;
assign w9465 = ~w9279 & ~w9280;
assign w9466 = ~w9281 & ~w9282;
assign w9467 = ~w9283 & ~w9284;
assign w9468 = ~w9285 & ~w9286;
assign w9469 = ~w9287 & ~w9288;
assign w9470 = ~w9289 & ~w9290;
assign w9471 = ~w9291 & ~w9292;
assign w9472 = ~w9293 & ~w9294;
assign w9473 = ~w9295 & ~w9296;
assign w9474 = ~w9297 & ~w9298;
assign w9475 = ~w9299 & ~w9300;
assign w9476 = ~w9301 & ~w9302;
assign w9477 = ~w9303 & ~w9304;
assign w9478 = ~w9305 & ~w9306;
assign w9479 = ~w9307 & ~w9308;
assign w9480 = ~w9309 & ~w9310;
assign w9481 = ~w9311 & ~w9312;
assign w9482 = ~w9313 & ~w9314;
assign w9483 = ~w9315 & ~w9316;
assign w9484 = ~w9317 & ~w9318;
assign w9485 = ~w9319 & ~w9320;
assign w9486 = ~w9321 & ~w9322;
assign w9487 = ~w9323 & ~w9324;
assign w9488 = ~w9325 & ~w9326;
assign w9489 = ~w9327 & ~w9328;
assign w9490 = ~w9329 & ~w9330;
assign w9491 = ~w9331 & ~w9332;
assign w9492 = ~w9333 & ~w9334;
assign w9493 = ~w9335 & ~w9336;
assign w9494 = ~w9337 & ~w9338;
assign w9495 = ~w9339 & ~w9340;
assign w9496 = ~w9341 & ~w9342;
assign w9497 = ~w9343 & ~w9344;
assign w9498 = ~w9345 & ~w9346;
assign w9499 = ~w9347 & ~w9348;
assign w9500 = ~w9349 & ~w9350;
assign w9501 = ~w9351 & ~w9352;
assign w9502 = ~w9353 & ~w9354;
assign w9503 = ~w9355 & ~w9356;
assign w9504 = ~w9357 & ~w9358;
assign w9505 = ~w9359 & ~w9360;
assign w9506 = ~w9361 & ~w9362;
assign w9507 = ~w9363 & ~w9364;
assign w9508 = ~w9365 & ~w9366;
assign w9509 = ~w9367 & ~w9368;
assign w9510 = ~w9369 & ~w9370;
assign w9511 = ~w9371 & ~w9372;
assign w9512 = ~w9373 & ~w9374;
assign w9513 = ~w9375 & ~w9376;
assign w9514 = ~w9377 & ~w9378;
assign w9515 = ~w9379 & ~w9380;
assign w9516 = ~w9381 & ~w9382;
assign w9517 = ~w9383 & ~w9384;
assign w9518 = ~w9385 & ~w9386;
assign w9519 = ~w9387 & ~w9388;
assign w9520 = ~w9389 & ~w9390;
assign w9521 = ~w9391 & ~w9392;
assign w9522 = ~w9393 & ~w9394;
assign w9523 = w9521 & w9522;
assign w9524 = w9519 & w9520;
assign w9525 = w9517 & w9518;
assign w9526 = w9515 & w9516;
assign w9527 = w9513 & w9514;
assign w9528 = w9511 & w9512;
assign w9529 = w9509 & w9510;
assign w9530 = w9507 & w9508;
assign w9531 = w9505 & w9506;
assign w9532 = w9503 & w9504;
assign w9533 = w9501 & w9502;
assign w9534 = w9499 & w9500;
assign w9535 = w9497 & w9498;
assign w9536 = w9495 & w9496;
assign w9537 = w9493 & w9494;
assign w9538 = w9491 & w9492;
assign w9539 = w9489 & w9490;
assign w9540 = w9487 & w9488;
assign w9541 = w9485 & w9486;
assign w9542 = w9483 & w9484;
assign w9543 = w9481 & w9482;
assign w9544 = w9479 & w9480;
assign w9545 = w9477 & w9478;
assign w9546 = w9475 & w9476;
assign w9547 = w9473 & w9474;
assign w9548 = w9471 & w9472;
assign w9549 = w9469 & w9470;
assign w9550 = w9467 & w9468;
assign w9551 = w9465 & w9466;
assign w9552 = w9463 & w9464;
assign w9553 = w9461 & w9462;
assign w9554 = w9459 & w9460;
assign w9555 = w9457 & w9458;
assign w9556 = w9455 & w9456;
assign w9557 = w9453 & w9454;
assign w9558 = w9451 & w9452;
assign w9559 = w9449 & w9450;
assign w9560 = w9447 & w9448;
assign w9561 = w9445 & w9446;
assign w9562 = w9443 & w9444;
assign w9563 = w9441 & w9442;
assign w9564 = w9439 & w9440;
assign w9565 = w9437 & w9438;
assign w9566 = w9435 & w9436;
assign w9567 = w9433 & w9434;
assign w9568 = w9431 & w9432;
assign w9569 = w9429 & w9430;
assign w9570 = w9427 & w9428;
assign w9571 = w9425 & w9426;
assign w9572 = w9423 & w9424;
assign w9573 = w9421 & w9422;
assign w9574 = w9419 & w9420;
assign w9575 = w9417 & w9418;
assign w9576 = w9415 & w9416;
assign w9577 = w9413 & w9414;
assign w9578 = w9411 & w9412;
assign w9579 = w9409 & w9410;
assign w9580 = w9407 & w9408;
assign w9581 = w9405 & w9406;
assign w9582 = w9403 & w9404;
assign w9583 = w9401 & w9402;
assign w9584 = w9399 & w9400;
assign w9585 = w9397 & w9398;
assign w9586 = w9395 & w9396;
assign w9587 = w9585 & w9586;
assign w9588 = w9583 & w9584;
assign w9589 = w9581 & w9582;
assign w9590 = w9579 & w9580;
assign w9591 = w9577 & w9578;
assign w9592 = w9575 & w9576;
assign w9593 = w9573 & w9574;
assign w9594 = w9571 & w9572;
assign w9595 = w9569 & w9570;
assign w9596 = w9567 & w9568;
assign w9597 = w9565 & w9566;
assign w9598 = w9563 & w9564;
assign w9599 = w9561 & w9562;
assign w9600 = w9559 & w9560;
assign w9601 = w9557 & w9558;
assign w9602 = w9555 & w9556;
assign w9603 = w9553 & w9554;
assign w9604 = w9551 & w9552;
assign w9605 = w9549 & w9550;
assign w9606 = w9547 & w9548;
assign w9607 = w9545 & w9546;
assign w9608 = w9543 & w9544;
assign w9609 = w9541 & w9542;
assign w9610 = w9539 & w9540;
assign w9611 = w9537 & w9538;
assign w9612 = w9535 & w9536;
assign w9613 = w9533 & w9534;
assign w9614 = w9531 & w9532;
assign w9615 = w9529 & w9530;
assign w9616 = w9527 & w9528;
assign w9617 = w9525 & w9526;
assign w9618 = w9523 & w9524;
assign w9619 = w9617 & w9618;
assign w9620 = w9615 & w9616;
assign w9621 = w9613 & w9614;
assign w9622 = w9611 & w9612;
assign w9623 = w9609 & w9610;
assign w9624 = w9607 & w9608;
assign w9625 = w9605 & w9606;
assign w9626 = w9603 & w9604;
assign w9627 = w9601 & w9602;
assign w9628 = w9599 & w9600;
assign w9629 = w9597 & w9598;
assign w9630 = w9595 & w9596;
assign w9631 = w9593 & w9594;
assign w9632 = w9591 & w9592;
assign w9633 = w9589 & w9590;
assign w9634 = w9587 & w9588;
assign w9635 = w9633 & w9634;
assign w9636 = w9631 & w9632;
assign w9637 = w9629 & w9630;
assign w9638 = w9627 & w9628;
assign w9639 = w9625 & w9626;
assign w9640 = w9623 & w9624;
assign w9641 = w9621 & w9622;
assign w9642 = w9619 & w9620;
assign w9643 = w9641 & w9642;
assign w9644 = w9639 & w9640;
assign w9645 = w9637 & w9638;
assign w9646 = w9635 & w9636;
assign w9647 = w9645 & w9646;
assign w9648 = w9643 & w9644;
assign w9649 = w9647 & w9648;
assign w9650 = ~pi10577 & ~w9649;
assign w9651 = pi02980 & w3296;
assign w9652 = pi05477 & w3300;
assign w9653 = pi05523 & w3572;
assign w9654 = pi05878 & w3596;
assign w9655 = pi03020 & w3310;
assign w9656 = pi01890 & w3602;
assign w9657 = pi06388 & w3418;
assign w9658 = pi06358 & w3160;
assign w9659 = pi03139 & w3494;
assign w9660 = pi02478 & w3229;
assign w9661 = pi03496 & w3488;
assign w9662 = pi03384 & w3258;
assign w9663 = pi05436 & w3256;
assign w9664 = pi03013 & w3610;
assign w9665 = pi05394 & w3082;
assign w9666 = pi09631 & w3530;
assign w9667 = pi05161 & w3612;
assign w9668 = pi03252 & w3214;
assign w9669 = pi09629 & w3404;
assign w9670 = pi03443 & w3177;
assign w9671 = pi05167 & w3252;
assign w9672 = pi09628 & w3426;
assign w9673 = pi03277 & w3115;
assign w9674 = pi09601 & w3400;
assign w9675 = pi03463 & w3396;
assign w9676 = pi05299 & w3450;
assign w9677 = pi06280 & w3324;
assign w9678 = pi06128 & w3264;
assign w9679 = pi02855 & w3336;
assign w9680 = pi05555 & w3420;
assign w9681 = pi02842 & w3520;
assign w9682 = pi03291 & w3328;
assign w9683 = pi02141 & w3460;
assign w9684 = pi02455 & w3223;
assign w9685 = pi05312 & w3298;
assign w9686 = pi03310 & w3564;
assign w9687 = pi05620 & w3272;
assign w9688 = pi05387 & w3153;
assign w9689 = pi05568 & w3364;
assign w9690 = pi05536 & w3286;
assign w9691 = pi05542 & w3552;
assign w9692 = pi05081 & w3486;
assign w9693 = pi05114 & w3308;
assign w9694 = pi02233 & w3217;
assign w9695 = pi05653 & w3276;
assign w9696 = pi02960 & w3274;
assign w9697 = pi02115 & w3122;
assign w9698 = pi05428 & w3078;
assign w9699 = pi05601 & w3472;
assign w9700 = pi03454 & w3588;
assign w9701 = pi05220 & w3480;
assign w9702 = pi05318 & w3354;
assign w9703 = pi02369 & w3570;
assign w9704 = pi05705 & w3201;
assign w9705 = pi05421 & w3284;
assign w9706 = pi02416 & w3342;
assign w9707 = pi03332 & w3512;
assign w9708 = pi05367 & w3304;
assign w9709 = pi02360 & w3219;
assign w9710 = pi05381 & w3496;
assign w9711 = pi09595 & w3103;
assign w9712 = pi05850 & w3386;
assign w9713 = pi02011 & w3538;
assign w9714 = pi05819 & w3464;
assign w9715 = pi06458 & w3242;
assign w9716 = pi03437 & w3388;
assign w9717 = pi05207 & w3568;
assign w9718 = pi02048 & w3482;
assign w9719 = pi05549 & w3410;
assign w9720 = pi02816 & w3614;
assign w9721 = pi05790 & w3192;
assign w9722 = pi03072 & w3338;
assign w9723 = pi05246 & w3356;
assign w9724 = pi03267 & w3086;
assign w9725 = pi05923 & w3474;
assign w9726 = pi05107 & w3143;
assign w9727 = pi05408 & w3514;
assign w9728 = pi03244 & w3334;
assign w9729 = pi03304 & w3146;
assign w9730 = pi05087 & w3232;
assign w9731 = pi02261 & w3288;
assign w9732 = pi03165 & w3522;
assign w9733 = pi06205 & w3188;
assign w9734 = pi03192 & w3502;
assign w9735 = pi05810 & w3390;
assign w9736 = pi05457 & w3384;
assign w9737 = pi05659 & w3434;
assign w9738 = pi05745 & w3194;
assign w9739 = pi03200 & w3454;
assign w9740 = pi01820 & w3227;
assign w9741 = pi02868 & w3500;
assign w9742 = pi05722 & w3374;
assign w9743 = pi03225 & w3290;
assign w9744 = pi02934 & w3534;
assign w9745 = pi05698 & w3165;
assign w9746 = pi05333 & w3203;
assign w9747 = pi02075 & w3582;
assign w9748 = pi03235 & w3326;
assign w9749 = pi03172 & w3181;
assign w9750 = pi03469 & w3211;
assign w9751 = pi06100 & w3320;
assign w9752 = pi03006 & w3260;
assign w9753 = pi06302 & w3158;
assign w9754 = pi02829 & w3380;
assign w9755 = pi09733 & w3408;
assign w9756 = pi02921 & w3250;
assign w9757 = pi01487 & w3346;
assign w9758 = pi06422 & w3150;
assign w9759 = pi09753 & w3544;
assign w9760 = pi01514 & w3608;
assign w9761 = pi02336 & w3550;
assign w9762 = pi05516 & w3406;
assign w9763 = pi02987 & w3137;
assign w9764 = pi06166 & w3280;
assign w9765 = pi03059 & w3576;
assign w9766 = pi05305 & w3236;
assign w9767 = pi06370 & w3524;
assign w9768 = pi05450 & w3442;
assign w9769 = pi05148 & w3344;
assign w9770 = pi05340 & w3129;
assign w9771 = pi05956 & w3175;
assign w9772 = pi02358 & w3440;
assign w9773 = pi03105 & w3132;
assign w9774 = pi01839 & w3179;
assign w9775 = pi05374 & w3462;
assign w9776 = pi05127 & w3248;
assign w9777 = pi05285 & w3314;
assign w9778 = pi01664 & w3246;
assign w9779 = pi03079 & w3348;
assign w9780 = pi05529 & w3340;
assign w9781 = pi02387 & w3446;
assign w9782 = pi05735 & w3600;
assign w9783 = pi03297 & w3484;
assign w9784 = pi05272 & w3540;
assign w9785 = pi03120 & w3071;
assign w9786 = pi03085 & w3456;
assign w9787 = pi03126 & w3118;
assign w9788 = pi02974 & w3424;
assign w9789 = pi09655 & w3238;
assign w9790 = pi01482 & w3306;
assign w9791 = pi03284 & w3190;
assign w9792 = pi05627 & w3376;
assign w9793 = pi05463 & w3432;
assign w9794 = pi03092 & w3592;
assign w9795 = pi06156 & w3542;
assign w9796 = pi05562 & w3135;
assign w9797 = pi06030 & w3594;
assign w9798 = pi06214 & w3402;
assign w9799 = pi01883 & w3173;
assign w9800 = pi05181 & w3554;
assign w9801 = pi02993 & w3262;
assign w9802 = pi09668 & w3093;
assign w9803 = pi03323 & w3618;
assign w9804 = pi06090 & w3444;
assign w9805 = pi03066 & w3209;
assign w9806 = pi02513 & w3580;
assign w9807 = pi05839 & w3270;
assign w9808 = pi03111 & w3394;
assign w9809 = pi03046 & w3526;
assign w9810 = pi03424 & w3184;
assign w9811 = pi02296 & w3332;
assign w9812 = pi05751 & w3590;
assign w9813 = pi05470 & w3506;
assign w9814 = pi05646 & w3566;
assign w9815 = pi05666 & w3508;
assign w9816 = pi03338 & w3412;
assign w9817 = pi05121 & w3436;
assign w9818 = pi02328 & w3316;
assign w9819 = pi09740 & w3510;
assign w9820 = pi02340 & w3366;
assign w9821 = pi02402 & w3148;
assign w9822 = pi02463 & w3560;
assign w9823 = pi05194 & w3528;
assign w9824 = pi05764 & w3171;
assign w9825 = pi01836 & w3422;
assign w9826 = pi01819 & w3438;
assign w9827 = pi01790 & w3368;
assign w9828 = pi09621 & w3516;
assign w9829 = pi06433 & w3558;
assign w9830 = pi09624 & w3064;
assign w9831 = pi06182 & w3096;
assign w9832 = pi09687 & w3470;
assign w9833 = pi06141 & w3546;
assign w9834 = pi05633 & w3358;
assign w9835 = pi05233 & w3112;
assign w9836 = pi02372 & w3294;
assign w9837 = pi05614 & w3620;
assign w9838 = pi05497 & w3466;
assign w9839 = pi05134 & w3598;
assign w9840 = pi06118 & w3282;
assign w9841 = pi05327 & w3392;
assign w9842 = pi05979 & w3606;
assign w9843 = pi03366 & w3169;
assign w9844 = pi06074 & w3106;
assign w9845 = pi03358 & w3562;
assign w9846 = pi02092 & w3414;
assign w9847 = pi05674 & w3167;
assign w9848 = pi05594 & w3225;
assign w9849 = pi05758 & w3430;
assign w9850 = pi05094 & w3240;
assign w9851 = pi03033 & w3548;
assign w9852 = pi05414 & w3186;
assign w9853 = pi03150 & w3428;
assign w9854 = pi05346 & w3199;
assign w9855 = pi05943 & w3616;
assign w9856 = pi05829 & w3207;
assign w9857 = pi05490 & w3234;
assign w9858 = pi05503 & w3127;
assign w9859 = pi09521 & w3532;
assign w9860 = pi05588 & w3254;
assign w9861 = pi02187 & w3378;
assign w9862 = pi03377 & w3302;
assign w9863 = pi05779 & w3458;
assign w9864 = pi03133 & w3574;
assign w9865 = pi02947 & w3322;
assign w9866 = pi05771 & w3476;
assign w9867 = pi06061 & w3584;
assign w9868 = pi03317 & w3370;
assign w9869 = pi01505 & w3197;
assign w9870 = pi02881 & w3416;
assign w9871 = pi05800 & w3360;
assign w9872 = pi06108 & w3478;
assign w9873 = pi05868 & w3352;
assign w9874 = pi03000 & w3292;
assign w9875 = pi02967 & w3536;
assign w9876 = pi03098 & w3498;
assign w9877 = pi02894 & w3362;
assign w9878 = pi03417 & w3504;
assign w9879 = pi05640 & w3448;
assign w9880 = pi05858 & w3382;
assign w9881 = pi03053 & w3350;
assign w9882 = pi06192 & w3318;
assign w9883 = pi05259 & w3586;
assign w9884 = pi05140 & w3604;
assign w9885 = pi05154 & w3492;
assign w9886 = pi06040 & w3468;
assign w9887 = pi05581 & w3205;
assign w9888 = pi01512 & w3110;
assign w9889 = pi02907 & w3330;
assign w9890 = pi02344 & w3452;
assign w9891 = pi03410 & w3162;
assign w9892 = pi05683 & w3312;
assign w9893 = pi05443 & w3518;
assign w9894 = pi05401 & w3278;
assign w9895 = pi05510 & w3139;
assign w9896 = pi05711 & w3372;
assign w9897 = pi05888 & w3125;
assign w9898 = pi01873 & w3578;
assign w9899 = pi05575 & w3156;
assign w9900 = pi03040 & w3490;
assign w9901 = pi05484 & w3398;
assign w9902 = pi05607 & w3221;
assign w9903 = pi03027 & w3244;
assign w9904 = pi03430 & w3556;
assign w9905 = pi05100 & w3266;
assign w9906 = pi09716 & w3268;
assign w9907 = ~w9651 & ~w9652;
assign w9908 = ~w9653 & ~w9654;
assign w9909 = ~w9655 & ~w9656;
assign w9910 = ~w9657 & ~w9658;
assign w9911 = ~w9659 & ~w9660;
assign w9912 = ~w9661 & ~w9662;
assign w9913 = ~w9663 & ~w9664;
assign w9914 = ~w9665 & ~w9666;
assign w9915 = ~w9667 & ~w9668;
assign w9916 = ~w9669 & ~w9670;
assign w9917 = ~w9671 & ~w9672;
assign w9918 = ~w9673 & ~w9674;
assign w9919 = ~w9675 & ~w9676;
assign w9920 = ~w9677 & ~w9678;
assign w9921 = ~w9679 & ~w9680;
assign w9922 = ~w9681 & ~w9682;
assign w9923 = ~w9683 & ~w9684;
assign w9924 = ~w9685 & ~w9686;
assign w9925 = ~w9687 & ~w9688;
assign w9926 = ~w9689 & ~w9690;
assign w9927 = ~w9691 & ~w9692;
assign w9928 = ~w9693 & ~w9694;
assign w9929 = ~w9695 & ~w9696;
assign w9930 = ~w9697 & ~w9698;
assign w9931 = ~w9699 & ~w9700;
assign w9932 = ~w9701 & ~w9702;
assign w9933 = ~w9703 & ~w9704;
assign w9934 = ~w9705 & ~w9706;
assign w9935 = ~w9707 & ~w9708;
assign w9936 = ~w9709 & ~w9710;
assign w9937 = ~w9711 & ~w9712;
assign w9938 = ~w9713 & ~w9714;
assign w9939 = ~w9715 & ~w9716;
assign w9940 = ~w9717 & ~w9718;
assign w9941 = ~w9719 & ~w9720;
assign w9942 = ~w9721 & ~w9722;
assign w9943 = ~w9723 & ~w9724;
assign w9944 = ~w9725 & ~w9726;
assign w9945 = ~w9727 & ~w9728;
assign w9946 = ~w9729 & ~w9730;
assign w9947 = ~w9731 & ~w9732;
assign w9948 = ~w9733 & ~w9734;
assign w9949 = ~w9735 & ~w9736;
assign w9950 = ~w9737 & ~w9738;
assign w9951 = ~w9739 & ~w9740;
assign w9952 = ~w9741 & ~w9742;
assign w9953 = ~w9743 & ~w9744;
assign w9954 = ~w9745 & ~w9746;
assign w9955 = ~w9747 & ~w9748;
assign w9956 = ~w9749 & ~w9750;
assign w9957 = ~w9751 & ~w9752;
assign w9958 = ~w9753 & ~w9754;
assign w9959 = ~w9755 & ~w9756;
assign w9960 = ~w9757 & ~w9758;
assign w9961 = ~w9759 & ~w9760;
assign w9962 = ~w9761 & ~w9762;
assign w9963 = ~w9763 & ~w9764;
assign w9964 = ~w9765 & ~w9766;
assign w9965 = ~w9767 & ~w9768;
assign w9966 = ~w9769 & ~w9770;
assign w9967 = ~w9771 & ~w9772;
assign w9968 = ~w9773 & ~w9774;
assign w9969 = ~w9775 & ~w9776;
assign w9970 = ~w9777 & ~w9778;
assign w9971 = ~w9779 & ~w9780;
assign w9972 = ~w9781 & ~w9782;
assign w9973 = ~w9783 & ~w9784;
assign w9974 = ~w9785 & ~w9786;
assign w9975 = ~w9787 & ~w9788;
assign w9976 = ~w9789 & ~w9790;
assign w9977 = ~w9791 & ~w9792;
assign w9978 = ~w9793 & ~w9794;
assign w9979 = ~w9795 & ~w9796;
assign w9980 = ~w9797 & ~w9798;
assign w9981 = ~w9799 & ~w9800;
assign w9982 = ~w9801 & ~w9802;
assign w9983 = ~w9803 & ~w9804;
assign w9984 = ~w9805 & ~w9806;
assign w9985 = ~w9807 & ~w9808;
assign w9986 = ~w9809 & ~w9810;
assign w9987 = ~w9811 & ~w9812;
assign w9988 = ~w9813 & ~w9814;
assign w9989 = ~w9815 & ~w9816;
assign w9990 = ~w9817 & ~w9818;
assign w9991 = ~w9819 & ~w9820;
assign w9992 = ~w9821 & ~w9822;
assign w9993 = ~w9823 & ~w9824;
assign w9994 = ~w9825 & ~w9826;
assign w9995 = ~w9827 & ~w9828;
assign w9996 = ~w9829 & ~w9830;
assign w9997 = ~w9831 & ~w9832;
assign w9998 = ~w9833 & ~w9834;
assign w9999 = ~w9835 & ~w9836;
assign w10000 = ~w9837 & ~w9838;
assign w10001 = ~w9839 & ~w9840;
assign w10002 = ~w9841 & ~w9842;
assign w10003 = ~w9843 & ~w9844;
assign w10004 = ~w9845 & ~w9846;
assign w10005 = ~w9847 & ~w9848;
assign w10006 = ~w9849 & ~w9850;
assign w10007 = ~w9851 & ~w9852;
assign w10008 = ~w9853 & ~w9854;
assign w10009 = ~w9855 & ~w9856;
assign w10010 = ~w9857 & ~w9858;
assign w10011 = ~w9859 & ~w9860;
assign w10012 = ~w9861 & ~w9862;
assign w10013 = ~w9863 & ~w9864;
assign w10014 = ~w9865 & ~w9866;
assign w10015 = ~w9867 & ~w9868;
assign w10016 = ~w9869 & ~w9870;
assign w10017 = ~w9871 & ~w9872;
assign w10018 = ~w9873 & ~w9874;
assign w10019 = ~w9875 & ~w9876;
assign w10020 = ~w9877 & ~w9878;
assign w10021 = ~w9879 & ~w9880;
assign w10022 = ~w9881 & ~w9882;
assign w10023 = ~w9883 & ~w9884;
assign w10024 = ~w9885 & ~w9886;
assign w10025 = ~w9887 & ~w9888;
assign w10026 = ~w9889 & ~w9890;
assign w10027 = ~w9891 & ~w9892;
assign w10028 = ~w9893 & ~w9894;
assign w10029 = ~w9895 & ~w9896;
assign w10030 = ~w9897 & ~w9898;
assign w10031 = ~w9899 & ~w9900;
assign w10032 = ~w9901 & ~w9902;
assign w10033 = ~w9903 & ~w9904;
assign w10034 = ~w9905 & ~w9906;
assign w10035 = w10033 & w10034;
assign w10036 = w10031 & w10032;
assign w10037 = w10029 & w10030;
assign w10038 = w10027 & w10028;
assign w10039 = w10025 & w10026;
assign w10040 = w10023 & w10024;
assign w10041 = w10021 & w10022;
assign w10042 = w10019 & w10020;
assign w10043 = w10017 & w10018;
assign w10044 = w10015 & w10016;
assign w10045 = w10013 & w10014;
assign w10046 = w10011 & w10012;
assign w10047 = w10009 & w10010;
assign w10048 = w10007 & w10008;
assign w10049 = w10005 & w10006;
assign w10050 = w10003 & w10004;
assign w10051 = w10001 & w10002;
assign w10052 = w9999 & w10000;
assign w10053 = w9997 & w9998;
assign w10054 = w9995 & w9996;
assign w10055 = w9993 & w9994;
assign w10056 = w9991 & w9992;
assign w10057 = w9989 & w9990;
assign w10058 = w9987 & w9988;
assign w10059 = w9985 & w9986;
assign w10060 = w9983 & w9984;
assign w10061 = w9981 & w9982;
assign w10062 = w9979 & w9980;
assign w10063 = w9977 & w9978;
assign w10064 = w9975 & w9976;
assign w10065 = w9973 & w9974;
assign w10066 = w9971 & w9972;
assign w10067 = w9969 & w9970;
assign w10068 = w9967 & w9968;
assign w10069 = w9965 & w9966;
assign w10070 = w9963 & w9964;
assign w10071 = w9961 & w9962;
assign w10072 = w9959 & w9960;
assign w10073 = w9957 & w9958;
assign w10074 = w9955 & w9956;
assign w10075 = w9953 & w9954;
assign w10076 = w9951 & w9952;
assign w10077 = w9949 & w9950;
assign w10078 = w9947 & w9948;
assign w10079 = w9945 & w9946;
assign w10080 = w9943 & w9944;
assign w10081 = w9941 & w9942;
assign w10082 = w9939 & w9940;
assign w10083 = w9937 & w9938;
assign w10084 = w9935 & w9936;
assign w10085 = w9933 & w9934;
assign w10086 = w9931 & w9932;
assign w10087 = w9929 & w9930;
assign w10088 = w9927 & w9928;
assign w10089 = w9925 & w9926;
assign w10090 = w9923 & w9924;
assign w10091 = w9921 & w9922;
assign w10092 = w9919 & w9920;
assign w10093 = w9917 & w9918;
assign w10094 = w9915 & w9916;
assign w10095 = w9913 & w9914;
assign w10096 = w9911 & w9912;
assign w10097 = w9909 & w9910;
assign w10098 = w9907 & w9908;
assign w10099 = w10097 & w10098;
assign w10100 = w10095 & w10096;
assign w10101 = w10093 & w10094;
assign w10102 = w10091 & w10092;
assign w10103 = w10089 & w10090;
assign w10104 = w10087 & w10088;
assign w10105 = w10085 & w10086;
assign w10106 = w10083 & w10084;
assign w10107 = w10081 & w10082;
assign w10108 = w10079 & w10080;
assign w10109 = w10077 & w10078;
assign w10110 = w10075 & w10076;
assign w10111 = w10073 & w10074;
assign w10112 = w10071 & w10072;
assign w10113 = w10069 & w10070;
assign w10114 = w10067 & w10068;
assign w10115 = w10065 & w10066;
assign w10116 = w10063 & w10064;
assign w10117 = w10061 & w10062;
assign w10118 = w10059 & w10060;
assign w10119 = w10057 & w10058;
assign w10120 = w10055 & w10056;
assign w10121 = w10053 & w10054;
assign w10122 = w10051 & w10052;
assign w10123 = w10049 & w10050;
assign w10124 = w10047 & w10048;
assign w10125 = w10045 & w10046;
assign w10126 = w10043 & w10044;
assign w10127 = w10041 & w10042;
assign w10128 = w10039 & w10040;
assign w10129 = w10037 & w10038;
assign w10130 = w10035 & w10036;
assign w10131 = w10129 & w10130;
assign w10132 = w10127 & w10128;
assign w10133 = w10125 & w10126;
assign w10134 = w10123 & w10124;
assign w10135 = w10121 & w10122;
assign w10136 = w10119 & w10120;
assign w10137 = w10117 & w10118;
assign w10138 = w10115 & w10116;
assign w10139 = w10113 & w10114;
assign w10140 = w10111 & w10112;
assign w10141 = w10109 & w10110;
assign w10142 = w10107 & w10108;
assign w10143 = w10105 & w10106;
assign w10144 = w10103 & w10104;
assign w10145 = w10101 & w10102;
assign w10146 = w10099 & w10100;
assign w10147 = w10145 & w10146;
assign w10148 = w10143 & w10144;
assign w10149 = w10141 & w10142;
assign w10150 = w10139 & w10140;
assign w10151 = w10137 & w10138;
assign w10152 = w10135 & w10136;
assign w10153 = w10133 & w10134;
assign w10154 = w10131 & w10132;
assign w10155 = w10153 & w10154;
assign w10156 = w10151 & w10152;
assign w10157 = w10149 & w10150;
assign w10158 = w10147 & w10148;
assign w10159 = w10157 & w10158;
assign w10160 = w10155 & w10156;
assign w10161 = w10159 & w10160;
assign w10162 = ~pi10577 & ~w10161;
assign w10163 = pi06237 & w3560;
assign w10164 = pi06142 & w3546;
assign w10165 = pi05382 & w3496;
assign w10166 = pi03014 & w3610;
assign w10167 = pi05945 & w3616;
assign w10168 = pi06324 & w3578;
assign w10169 = pi02065 & w3177;
assign w10170 = pi06290 & w3332;
assign w10171 = pi03391 & w3122;
assign w10172 = pi02882 & w3416;
assign w10173 = pi02142 & w3618;
assign w10174 = pi05260 & w3586;
assign w10175 = pi05234 & w3112;
assign w10176 = pi05415 & w3186;
assign w10177 = pi02975 & w3424;
assign w10178 = pi02954 & w3103;
assign w10179 = pi01717 & w3264;
assign w10180 = pi03093 & w3592;
assign w10181 = pi02081 & w3396;
assign w10182 = pi05313 & w3298;
assign w10183 = pi01841 & w3444;
assign w10184 = pi06167 & w3280;
assign w10185 = pi03060 & w3576;
assign w10186 = pi01704 & w3207;
assign w10187 = pi03411 & w3162;
assign w10188 = pi05266 & w3414;
assign w10189 = pi02119 & w3258;
assign w10190 = pi06022 & w3366;
assign w10191 = pi09664 & w3127;
assign w10192 = pi05999 & w3570;
assign w10193 = pi01875 & w3194;
assign w10194 = pi02981 & w3296;
assign w10195 = pi05409 & w3514;
assign w10196 = pi05723 & w3374;
assign w10197 = pi05182 & w3554;
assign w10198 = pi03279 & w3115;
assign w10199 = pi01937 & w3392;
assign w10200 = pi05122 & w3436;
assign w10201 = pi05458 & w3384;
assign w10202 = pi05388 & w3153;
assign w10203 = pi05128 & w3248;
assign w10204 = pi02862 & w3544;
assign w10205 = pi06402 & w3246;
assign w10206 = pi05903 & w3238;
assign w10207 = pi09602 & w3552;
assign w10208 = pi05936 & w3532;
assign w10209 = pi02206 & w3454;
assign w10210 = pi05737 & w3600;
assign w10211 = pi06448 & w3510;
assign w10212 = pi02403 & w3344;
assign w10213 = pi05368 & w3304;
assign w10214 = pi06310 & w3602;
assign w10215 = pi03455 & w3588;
assign w10216 = pi02747 & w3472;
assign w10217 = pi02428 & w3276;
assign w10218 = pi02337 & w3372;
assign w10219 = pi02750 & w3225;
assign w10220 = pi05221 & w3480;
assign w10221 = pi05300 & w3450;
assign w10222 = pi02409 & w3434;
assign w10223 = pi05471 & w3506;
assign w10224 = pi03269 & w3086;
assign w10225 = pi03041 & w3490;
assign w10226 = pi06184 & w3096;
assign w10227 = pi06442 & w3408;
assign w10228 = pi06051 & w3173;
assign w10229 = pi01825 & w3192;
assign w10230 = pi03285 & w3190;
assign w10231 = pi05293 & w3538;
assign w10232 = pi02732 & w3254;
assign w10233 = pi09648 & w3572;
assign w10234 = pi05082 & w3486;
assign w10235 = pi02843 & w3520;
assign w10236 = pi02632 & w3358;
assign w10237 = pi02948 & w3322;
assign w10238 = pi01880 & w3171;
assign w10239 = pi06001 & w3205;
assign w10240 = pi06337 & w3179;
assign w10241 = pi02093 & w3302;
assign w10242 = pi05464 & w3432;
assign w10243 = pi03368 & w3169;
assign w10244 = pi05141 & w3604;
assign w10245 = pi05909 & w3426;
assign w10246 = pi09683 & w3596;
assign w10247 = pi03106 & w3132;
assign w10248 = pi05971 & w3223;
assign w10249 = pi05208 & w3568;
assign w10250 = pi02915 & w3530;
assign w10251 = pi01781 & w3282;
assign w10252 = pi05188 & w3452;
assign w10253 = pi06015 & w3608;
assign w10254 = pi06282 & w3324;
assign w10255 = pi09672 & w3466;
assign w10256 = pi03292 & w3328;
assign w10257 = pi05896 & w3093;
assign w10258 = pi03073 & w3338;
assign w10259 = pi02413 & w3508;
assign w10260 = pi03021 & w3310;
assign w10261 = pi05437 & w3256;
assign w10262 = pi09593 & w3410;
assign w10263 = pi03478 & w3582;
assign w10264 = pi02994 & w3262;
assign w10265 = pi09552 & w3386;
assign w10266 = pi03166 & w3522;
assign w10267 = pi05155 & w3492;
assign w10268 = pi05115 & w3308;
assign w10269 = pi02875 & w3268;
assign w10270 = pi05286 & w3314;
assign w10271 = pi05214 & w3288;
assign w10272 = pi03121 & w3071;
assign w10273 = pi05201 & w3550;
assign w10274 = pi03298 & w3484;
assign w10275 = pi01892 & w3430;
assign w10276 = pi02888 & w3470;
assign w10277 = pi05429 & w3078;
assign w10278 = pi03226 & w3290;
assign w10279 = pi05395 & w3082;
assign w10280 = pi05279 & w3482;
assign w10281 = pi05227 & w3217;
assign w10282 = pi02136 & w3412;
assign w10283 = pi09532 & w3364;
assign w10284 = pi05360 & w3227;
assign w10285 = pi02516 & w3448;
assign w10286 = pi03173 & w3181;
assign w10287 = pi05095 & w3240;
assign w10288 = pi02830 & w3380;
assign w10289 = pi05247 & w3356;
assign w10290 = pi06158 & w3542;
assign w10291 = pi09645 & w3139;
assign w10292 = pi05422 & w3284;
assign w10293 = pi02105 & w3504;
assign w10294 = pi02836 & w3346;
assign w10295 = pi09690 & w3398;
assign w10296 = pi02849 & w3197;
assign w10297 = pi06424 & w3150;
assign w10298 = pi03245 & w3334;
assign w10299 = pi02139 & w3512;
assign w10300 = pi06224 & w3580;
assign w10301 = pi03134 & w3574;
assign w10302 = pi03318 & w3370;
assign w10303 = pi05101 & w3266;
assign w10304 = pi03054 & w3350;
assign w10305 = pi02504 & w3566;
assign w10306 = pi02077 & w3211;
assign w10307 = pi06360 & w3160;
assign w10308 = pi01853 & w3199;
assign w10309 = pi03112 & w3394;
assign w10310 = pi02357 & w3165;
assign w10311 = pi06110 & w3478;
assign w10312 = pi02908 & w3330;
assign w10313 = pi02739 & w3620;
assign w10314 = pi06261 & w3294;
assign w10315 = pi03001 & w3292;
assign w10316 = pi05980 & w3606;
assign w10317 = pi05306 & w3236;
assign w10318 = pi02089 & w3556;
assign w10319 = pi05781 & w3458;
assign w10320 = pi06206 & w3188;
assign w10321 = pi05402 & w3278;
assign w10322 = pi09673 & w3234;
assign w10323 = pi05168 & w3252;
assign w10324 = pi01647 & w3270;
assign w10325 = pi06372 & w3524;
assign w10326 = pi05175 & w3219;
assign w10327 = pi02941 & w3400;
assign w10328 = pi02213 & w3502;
assign w10329 = pi05958 & w3175;
assign w10330 = pi06032 & w3594;
assign w10331 = pi05821 & w3464;
assign w10332 = pi06193 & w3318;
assign w10333 = pi03236 & w3326;
assign w10334 = pi05135 & w3598;
assign w10335 = pi05240 & w3378;
assign w10336 = pi06434 & w3558;
assign w10337 = pi01678 & w3418;
assign w10338 = pi02126 & w3562;
assign w10339 = pi01898 & w3590;
assign w10340 = pi03034 & w3548;
assign w10341 = pi09636 & w3340;
assign w10342 = pi02099 & w3184;
assign w10343 = pi09571 & w3420;
assign w10344 = pi03311 & w3564;
assign w10345 = pi03086 & w3456;
assign w10346 = pi02069 & w3488;
assign w10347 = pi03028 & w3244;
assign w10348 = pi03151 & w3428;
assign w10349 = pi09569 & w3135;
assign w10350 = pi06415 & w3110;
assign w10351 = pi03099 & w3498;
assign w10352 = pi05253 & w3460;
assign w10353 = pi02901 & w3404;
assign w10354 = pi01727 & w3129;
assign w10355 = pi02968 & w3536;
assign w10356 = pi06343 & w3438;
assign w10357 = pi01793 & w3360;
assign w10358 = pi06250 & w3148;
assign w10359 = pi09727 & w3352;
assign w10360 = pi02988 & w3137;
assign w10361 = pi03047 & w3526;
assign w10362 = pi02345 & w3201;
assign w10363 = pi01907 & w3203;
assign w10364 = pi05925 & w3474;
assign w10365 = pi05108 & w3143;
assign w10366 = pi05811 & w3390;
assign w10367 = pi06459 & w3242;
assign w10368 = pi03007 & w3260;
assign w10369 = pi05451 & w3442;
assign w10370 = pi05916 & w3516;
assign w10371 = pi02856 & w3336;
assign w10372 = pi09622 & w3286;
assign w10373 = pi05375 & w3462;
assign w10374 = pi02817 & w3614;
assign w10375 = pi02928 & w3064;
assign w10376 = pi03080 & w3348;
assign w10377 = pi05685 & w3312;
assign w10378 = pi02961 & w3274;
assign w10379 = pi06244 & w3342;
assign w10380 = pi05675 & w3167;
assign w10381 = pi05273 & w3540;
assign w10382 = pi06216 & w3402;
assign w10383 = pi05088 & w3232;
assign w10384 = pi03067 & w3209;
assign w10385 = pi06062 & w3584;
assign w10386 = pi02647 & w3376;
assign w10387 = pi01901 & w3158;
assign w10388 = pi05195 & w3528;
assign w10389 = pi05444 & w3518;
assign w10390 = pi05861 & w3382;
assign w10391 = pi03253 & w3214;
assign w10392 = pi02869 & w3500;
assign w10393 = pi06075 & w3106;
assign w10394 = pi06009 & w3440;
assign w10395 = pi09654 & w3406;
assign w10396 = pi01821 & w3320;
assign w10397 = pi03140 & w3494;
assign w10398 = pi05989 & w3446;
assign w10399 = pi06231 & w3229;
assign w10400 = pi02383 & w3612;
assign w10401 = pi09539 & w3156;
assign w10402 = pi09697 & w3300;
assign w10403 = pi02823 & w3306;
assign w10404 = pi03127 & w3118;
assign w10405 = pi02738 & w3221;
assign w10406 = pi06041 & w3468;
assign w10407 = pi02935 & w3534;
assign w10408 = pi02735 & w3272;
assign w10409 = pi02097 & w3388;
assign w10410 = pi05889 & w3125;
assign w10411 = pi06271 & w3316;
assign w10412 = pi02922 & w3250;
assign w10413 = pi03305 & w3146;
assign w10414 = pi02895 & w3362;
assign w10415 = pi05354 & w3422;
assign w10416 = pi01866 & w3476;
assign w10417 = pi05319 & w3354;
assign w10418 = pi06350 & w3368;
assign w10419 = ~w10163 & ~w10164;
assign w10420 = ~w10165 & ~w10166;
assign w10421 = ~w10167 & ~w10168;
assign w10422 = ~w10169 & ~w10170;
assign w10423 = ~w10171 & ~w10172;
assign w10424 = ~w10173 & ~w10174;
assign w10425 = ~w10175 & ~w10176;
assign w10426 = ~w10177 & ~w10178;
assign w10427 = ~w10179 & ~w10180;
assign w10428 = ~w10181 & ~w10182;
assign w10429 = ~w10183 & ~w10184;
assign w10430 = ~w10185 & ~w10186;
assign w10431 = ~w10187 & ~w10188;
assign w10432 = ~w10189 & ~w10190;
assign w10433 = ~w10191 & ~w10192;
assign w10434 = ~w10193 & ~w10194;
assign w10435 = ~w10195 & ~w10196;
assign w10436 = ~w10197 & ~w10198;
assign w10437 = ~w10199 & ~w10200;
assign w10438 = ~w10201 & ~w10202;
assign w10439 = ~w10203 & ~w10204;
assign w10440 = ~w10205 & ~w10206;
assign w10441 = ~w10207 & ~w10208;
assign w10442 = ~w10209 & ~w10210;
assign w10443 = ~w10211 & ~w10212;
assign w10444 = ~w10213 & ~w10214;
assign w10445 = ~w10215 & ~w10216;
assign w10446 = ~w10217 & ~w10218;
assign w10447 = ~w10219 & ~w10220;
assign w10448 = ~w10221 & ~w10222;
assign w10449 = ~w10223 & ~w10224;
assign w10450 = ~w10225 & ~w10226;
assign w10451 = ~w10227 & ~w10228;
assign w10452 = ~w10229 & ~w10230;
assign w10453 = ~w10231 & ~w10232;
assign w10454 = ~w10233 & ~w10234;
assign w10455 = ~w10235 & ~w10236;
assign w10456 = ~w10237 & ~w10238;
assign w10457 = ~w10239 & ~w10240;
assign w10458 = ~w10241 & ~w10242;
assign w10459 = ~w10243 & ~w10244;
assign w10460 = ~w10245 & ~w10246;
assign w10461 = ~w10247 & ~w10248;
assign w10462 = ~w10249 & ~w10250;
assign w10463 = ~w10251 & ~w10252;
assign w10464 = ~w10253 & ~w10254;
assign w10465 = ~w10255 & ~w10256;
assign w10466 = ~w10257 & ~w10258;
assign w10467 = ~w10259 & ~w10260;
assign w10468 = ~w10261 & ~w10262;
assign w10469 = ~w10263 & ~w10264;
assign w10470 = ~w10265 & ~w10266;
assign w10471 = ~w10267 & ~w10268;
assign w10472 = ~w10269 & ~w10270;
assign w10473 = ~w10271 & ~w10272;
assign w10474 = ~w10273 & ~w10274;
assign w10475 = ~w10275 & ~w10276;
assign w10476 = ~w10277 & ~w10278;
assign w10477 = ~w10279 & ~w10280;
assign w10478 = ~w10281 & ~w10282;
assign w10479 = ~w10283 & ~w10284;
assign w10480 = ~w10285 & ~w10286;
assign w10481 = ~w10287 & ~w10288;
assign w10482 = ~w10289 & ~w10290;
assign w10483 = ~w10291 & ~w10292;
assign w10484 = ~w10293 & ~w10294;
assign w10485 = ~w10295 & ~w10296;
assign w10486 = ~w10297 & ~w10298;
assign w10487 = ~w10299 & ~w10300;
assign w10488 = ~w10301 & ~w10302;
assign w10489 = ~w10303 & ~w10304;
assign w10490 = ~w10305 & ~w10306;
assign w10491 = ~w10307 & ~w10308;
assign w10492 = ~w10309 & ~w10310;
assign w10493 = ~w10311 & ~w10312;
assign w10494 = ~w10313 & ~w10314;
assign w10495 = ~w10315 & ~w10316;
assign w10496 = ~w10317 & ~w10318;
assign w10497 = ~w10319 & ~w10320;
assign w10498 = ~w10321 & ~w10322;
assign w10499 = ~w10323 & ~w10324;
assign w10500 = ~w10325 & ~w10326;
assign w10501 = ~w10327 & ~w10328;
assign w10502 = ~w10329 & ~w10330;
assign w10503 = ~w10331 & ~w10332;
assign w10504 = ~w10333 & ~w10334;
assign w10505 = ~w10335 & ~w10336;
assign w10506 = ~w10337 & ~w10338;
assign w10507 = ~w10339 & ~w10340;
assign w10508 = ~w10341 & ~w10342;
assign w10509 = ~w10343 & ~w10344;
assign w10510 = ~w10345 & ~w10346;
assign w10511 = ~w10347 & ~w10348;
assign w10512 = ~w10349 & ~w10350;
assign w10513 = ~w10351 & ~w10352;
assign w10514 = ~w10353 & ~w10354;
assign w10515 = ~w10355 & ~w10356;
assign w10516 = ~w10357 & ~w10358;
assign w10517 = ~w10359 & ~w10360;
assign w10518 = ~w10361 & ~w10362;
assign w10519 = ~w10363 & ~w10364;
assign w10520 = ~w10365 & ~w10366;
assign w10521 = ~w10367 & ~w10368;
assign w10522 = ~w10369 & ~w10370;
assign w10523 = ~w10371 & ~w10372;
assign w10524 = ~w10373 & ~w10374;
assign w10525 = ~w10375 & ~w10376;
assign w10526 = ~w10377 & ~w10378;
assign w10527 = ~w10379 & ~w10380;
assign w10528 = ~w10381 & ~w10382;
assign w10529 = ~w10383 & ~w10384;
assign w10530 = ~w10385 & ~w10386;
assign w10531 = ~w10387 & ~w10388;
assign w10532 = ~w10389 & ~w10390;
assign w10533 = ~w10391 & ~w10392;
assign w10534 = ~w10393 & ~w10394;
assign w10535 = ~w10395 & ~w10396;
assign w10536 = ~w10397 & ~w10398;
assign w10537 = ~w10399 & ~w10400;
assign w10538 = ~w10401 & ~w10402;
assign w10539 = ~w10403 & ~w10404;
assign w10540 = ~w10405 & ~w10406;
assign w10541 = ~w10407 & ~w10408;
assign w10542 = ~w10409 & ~w10410;
assign w10543 = ~w10411 & ~w10412;
assign w10544 = ~w10413 & ~w10414;
assign w10545 = ~w10415 & ~w10416;
assign w10546 = ~w10417 & ~w10418;
assign w10547 = w10545 & w10546;
assign w10548 = w10543 & w10544;
assign w10549 = w10541 & w10542;
assign w10550 = w10539 & w10540;
assign w10551 = w10537 & w10538;
assign w10552 = w10535 & w10536;
assign w10553 = w10533 & w10534;
assign w10554 = w10531 & w10532;
assign w10555 = w10529 & w10530;
assign w10556 = w10527 & w10528;
assign w10557 = w10525 & w10526;
assign w10558 = w10523 & w10524;
assign w10559 = w10521 & w10522;
assign w10560 = w10519 & w10520;
assign w10561 = w10517 & w10518;
assign w10562 = w10515 & w10516;
assign w10563 = w10513 & w10514;
assign w10564 = w10511 & w10512;
assign w10565 = w10509 & w10510;
assign w10566 = w10507 & w10508;
assign w10567 = w10505 & w10506;
assign w10568 = w10503 & w10504;
assign w10569 = w10501 & w10502;
assign w10570 = w10499 & w10500;
assign w10571 = w10497 & w10498;
assign w10572 = w10495 & w10496;
assign w10573 = w10493 & w10494;
assign w10574 = w10491 & w10492;
assign w10575 = w10489 & w10490;
assign w10576 = w10487 & w10488;
assign w10577 = w10485 & w10486;
assign w10578 = w10483 & w10484;
assign w10579 = w10481 & w10482;
assign w10580 = w10479 & w10480;
assign w10581 = w10477 & w10478;
assign w10582 = w10475 & w10476;
assign w10583 = w10473 & w10474;
assign w10584 = w10471 & w10472;
assign w10585 = w10469 & w10470;
assign w10586 = w10467 & w10468;
assign w10587 = w10465 & w10466;
assign w10588 = w10463 & w10464;
assign w10589 = w10461 & w10462;
assign w10590 = w10459 & w10460;
assign w10591 = w10457 & w10458;
assign w10592 = w10455 & w10456;
assign w10593 = w10453 & w10454;
assign w10594 = w10451 & w10452;
assign w10595 = w10449 & w10450;
assign w10596 = w10447 & w10448;
assign w10597 = w10445 & w10446;
assign w10598 = w10443 & w10444;
assign w10599 = w10441 & w10442;
assign w10600 = w10439 & w10440;
assign w10601 = w10437 & w10438;
assign w10602 = w10435 & w10436;
assign w10603 = w10433 & w10434;
assign w10604 = w10431 & w10432;
assign w10605 = w10429 & w10430;
assign w10606 = w10427 & w10428;
assign w10607 = w10425 & w10426;
assign w10608 = w10423 & w10424;
assign w10609 = w10421 & w10422;
assign w10610 = w10419 & w10420;
assign w10611 = w10609 & w10610;
assign w10612 = w10607 & w10608;
assign w10613 = w10605 & w10606;
assign w10614 = w10603 & w10604;
assign w10615 = w10601 & w10602;
assign w10616 = w10599 & w10600;
assign w10617 = w10597 & w10598;
assign w10618 = w10595 & w10596;
assign w10619 = w10593 & w10594;
assign w10620 = w10591 & w10592;
assign w10621 = w10589 & w10590;
assign w10622 = w10587 & w10588;
assign w10623 = w10585 & w10586;
assign w10624 = w10583 & w10584;
assign w10625 = w10581 & w10582;
assign w10626 = w10579 & w10580;
assign w10627 = w10577 & w10578;
assign w10628 = w10575 & w10576;
assign w10629 = w10573 & w10574;
assign w10630 = w10571 & w10572;
assign w10631 = w10569 & w10570;
assign w10632 = w10567 & w10568;
assign w10633 = w10565 & w10566;
assign w10634 = w10563 & w10564;
assign w10635 = w10561 & w10562;
assign w10636 = w10559 & w10560;
assign w10637 = w10557 & w10558;
assign w10638 = w10555 & w10556;
assign w10639 = w10553 & w10554;
assign w10640 = w10551 & w10552;
assign w10641 = w10549 & w10550;
assign w10642 = w10547 & w10548;
assign w10643 = w10641 & w10642;
assign w10644 = w10639 & w10640;
assign w10645 = w10637 & w10638;
assign w10646 = w10635 & w10636;
assign w10647 = w10633 & w10634;
assign w10648 = w10631 & w10632;
assign w10649 = w10629 & w10630;
assign w10650 = w10627 & w10628;
assign w10651 = w10625 & w10626;
assign w10652 = w10623 & w10624;
assign w10653 = w10621 & w10622;
assign w10654 = w10619 & w10620;
assign w10655 = w10617 & w10618;
assign w10656 = w10615 & w10616;
assign w10657 = w10613 & w10614;
assign w10658 = w10611 & w10612;
assign w10659 = w10657 & w10658;
assign w10660 = w10655 & w10656;
assign w10661 = w10653 & w10654;
assign w10662 = w10651 & w10652;
assign w10663 = w10649 & w10650;
assign w10664 = w10647 & w10648;
assign w10665 = w10645 & w10646;
assign w10666 = w10643 & w10644;
assign w10667 = w10665 & w10666;
assign w10668 = w10663 & w10664;
assign w10669 = w10661 & w10662;
assign w10670 = w10659 & w10660;
assign w10671 = w10669 & w10670;
assign w10672 = w10667 & w10668;
assign w10673 = w10671 & w10672;
assign w10674 = ~pi10577 & ~w10673;
assign w10675 = w76 & w1084;
assign w10676 = ~w2275 & w55708;
assign w10677 = ~pi09872 & ~pi10586;
assign w10678 = ~pi01606 & pi09872;
assign w10679 = ~w10677 & ~w10678;
assign w10680 = w145 & w10679;
assign w10681 = ~w10676 & w10680;
assign w10682 = ~pi10581 & ~pi10582;
assign w10683 = ~pi00441 & pi00460;
assign w10684 = ~w10682 & ~w10683;
assign w10685 = ~pi00461 & w10682;
assign w10686 = ~pi01216 & ~pi01450;
assign w10687 = ~pi01454 & w10686;
assign w10688 = w10686 & w55709;
assign w10689 = ~pi01274 & w10688;
assign w10690 = pi00441 & ~pi00460;
assign w10691 = ~w10683 & ~w10690;
assign w10692 = (w10685 & ~w10689) | (w10685 & w55710) | (~w10689 & w55710);
assign w10693 = pi00461 & ~w10690;
assign w10694 = ~pi02348 & pi10352;
assign w10695 = pi00442 & w10694;
assign w10696 = ~w10684 & ~w10693;
assign w10697 = w10695 & w10696;
assign w10698 = ~w10692 & w10697;
assign w10699 = (~pi00461 & ~w10688) | (~pi00461 & w55711) | (~w10688 & w55711);
assign w10700 = pi00441 & w10682;
assign w10701 = ~pi00460 & pi00461;
assign w10702 = pi00460 & ~pi00461;
assign w10703 = ~w10701 & ~w10702;
assign w10704 = w10700 & ~w10703;
assign w10705 = w10685 & ~w10690;
assign w10706 = w10685 & w55712;
assign w10707 = ~w10704 & ~w10706;
assign w10708 = ~pi00442 & w10694;
assign w10709 = ~w10699 & w10708;
assign w10710 = ~w10707 & w10709;
assign w10711 = ~w10698 & ~w10710;
assign w10712 = ~pi00441 & ~w10682;
assign w10713 = ~w10700 & ~w10712;
assign w10714 = w10682 & w10694;
assign w10715 = w10701 & ~w10714;
assign w10716 = ~w10713 & w10715;
assign w10717 = (~w10688 & w55714) | (~w10688 & w55715) | (w55714 & w55715);
assign w10718 = (w10717 & w10716) | (w10717 & w55716) | (w10716 & w55716);
assign w10719 = (~pi00474 & ~w10694) | (~pi00474 & w55717) | (~w10694 & w55717);
assign w10720 = ~w10689 & w10719;
assign w10721 = ~w10707 & w10720;
assign w10722 = ~w10718 & ~w10721;
assign w10723 = w10711 & w10722;
assign w10724 = pi00375 & w10723;
assign w10725 = ~pi00488 & ~pi00540;
assign w10726 = ~pi00643 & w10725;
assign w10727 = w10718 & ~w10726;
assign w10728 = ~w10722 & ~w10727;
assign w10729 = pi00095 & w10728;
assign w10730 = ~pi00457 & ~pi00458;
assign w10731 = ~pi00459 & w10730;
assign w10732 = w10698 & ~w10731;
assign w10733 = ~w10727 & ~w10732;
assign w10734 = ~pi00375 & ~w10733;
assign w10735 = w10698 & w10731;
assign w10736 = ~w10710 & ~w10735;
assign w10737 = (pi00098 & w10735) | (pi00098 & w55718) | (w10735 & w55718);
assign w10738 = ~w10724 & ~w10729;
assign w10739 = ~w10734 & ~w10737;
assign w10740 = w10738 & w10739;
assign w10741 = ~pi00376 & ~pi10516;
assign w10742 = ~w3014 & ~w10741;
assign w10743 = ~w1122 & ~w1128;
assign w10744 = ~pi00320 & ~w10743;
assign w10745 = ~pi01272 & w2425;
assign w10746 = pi00203 & ~pi00230;
assign w10747 = pi01272 & w10746;
assign w10748 = ~w10745 & ~w10747;
assign w10749 = (pi00377 & ~w10744) | (pi00377 & w55719) | (~w10744 & w55719);
assign w10750 = w10744 & w55720;
assign w10751 = ~w10749 & ~w10750;
assign w10752 = (pi00378 & ~w10744) | (pi00378 & w55721) | (~w10744 & w55721);
assign w10753 = w10744 & w55722;
assign w10754 = ~w10752 & ~w10753;
assign w10755 = (pi00379 & ~w10744) | (pi00379 & w55723) | (~w10744 & w55723);
assign w10756 = w10744 & w55724;
assign w10757 = ~w10755 & ~w10756;
assign w10758 = (pi00380 & ~w10744) | (pi00380 & w55725) | (~w10744 & w55725);
assign w10759 = w10744 & w55726;
assign w10760 = ~w10758 & ~w10759;
assign w10761 = (pi00381 & ~w10744) | (pi00381 & w55727) | (~w10744 & w55727);
assign w10762 = w10744 & w55728;
assign w10763 = ~w10761 & ~w10762;
assign w10764 = (pi00382 & ~w10744) | (pi00382 & w55729) | (~w10744 & w55729);
assign w10765 = w10744 & w55730;
assign w10766 = ~w10764 & ~w10765;
assign w10767 = w10744 & w10748;
assign w10768 = ~w2429 & w10767;
assign w10769 = pi00383 & ~w10768;
assign w10770 = pi10511 & w10768;
assign w10771 = ~w10769 & ~w10770;
assign w10772 = pi00384 & ~w10768;
assign w10773 = ~pi10489 & w10768;
assign w10774 = ~w10772 & ~w10773;
assign w10775 = pi00385 & ~w10768;
assign w10776 = ~pi10520 & w10768;
assign w10777 = ~w10775 & ~w10776;
assign w10778 = pi00386 & ~w10768;
assign w10779 = pi10486 & w10768;
assign w10780 = ~w10778 & ~w10779;
assign w10781 = pi00387 & ~w10768;
assign w10782 = ~pi10495 & w10768;
assign w10783 = ~w10781 & ~w10782;
assign w10784 = pi00388 & ~w10768;
assign w10785 = ~pi10492 & w10768;
assign w10786 = ~w10784 & ~w10785;
assign w10787 = pi00389 & ~w10768;
assign w10788 = ~pi10505 & w10768;
assign w10789 = ~w10787 & ~w10788;
assign w10790 = pi00390 & ~w10768;
assign w10791 = pi10483 & w10768;
assign w10792 = ~w10790 & ~w10791;
assign w10793 = w2585 & w10767;
assign w10794 = pi00391 & ~w10793;
assign w10795 = pi10511 & w10793;
assign w10796 = ~w10794 & ~w10795;
assign w10797 = pi00392 & ~w10793;
assign w10798 = ~pi10489 & w10793;
assign w10799 = ~w10797 & ~w10798;
assign w10800 = pi00393 & ~w10793;
assign w10801 = ~pi10520 & w10793;
assign w10802 = ~w10800 & ~w10801;
assign w10803 = pi00394 & ~w10793;
assign w10804 = pi10486 & w10793;
assign w10805 = ~w10803 & ~w10804;
assign w10806 = pi00395 & ~w10793;
assign w10807 = ~pi10495 & w10793;
assign w10808 = ~w10806 & ~w10807;
assign w10809 = pi00396 & ~w10793;
assign w10810 = ~pi10492 & w10793;
assign w10811 = ~w10809 & ~w10810;
assign w10812 = pi00397 & ~w10793;
assign w10813 = ~pi10505 & w10793;
assign w10814 = ~w10812 & ~w10813;
assign w10815 = pi00398 & ~w10793;
assign w10816 = pi10483 & w10793;
assign w10817 = ~w10815 & ~w10816;
assign w10818 = (pi00399 & ~w10744) | (pi00399 & w55731) | (~w10744 & w55731);
assign w10819 = w10744 & w55732;
assign w10820 = ~w10818 & ~w10819;
assign w10821 = (pi00400 & ~w10744) | (pi00400 & w55733) | (~w10744 & w55733);
assign w10822 = w10744 & w55734;
assign w10823 = ~w10821 & ~w10822;
assign w10824 = w799 & w55736;
assign w10825 = (w799 & w55737) | (w799 & w55738) | (w55737 & w55738);
assign w10826 = ~w10824 & w10825;
assign w10827 = ~pi00536 & w6048;
assign w10828 = (w671 & w6048) | (w671 & w55739) | (w6048 & w55739);
assign w10829 = ~w10827 & w10828;
assign w10830 = pi00375 & pi00414;
assign w10831 = pi00432 & w10830;
assign w10832 = w10830 & w54698;
assign w10833 = pi00424 & w10832;
assign w10834 = w10832 & w54699;
assign w10835 = w10832 & w54718;
assign w10836 = pi00427 & w10835;
assign w10837 = w10835 & w54741;
assign w10838 = w10835 & w54742;
assign w10839 = w10835 & w54768;
assign w10840 = pi00404 & pi00407;
assign w10841 = pi00408 & pi00409;
assign w10842 = pi00410 & pi00411;
assign w10843 = pi00412 & pi00431;
assign w10844 = w10842 & w10843;
assign w10845 = w10840 & w10841;
assign w10846 = w10844 & w10845;
assign w10847 = w10839 & w10846;
assign w10848 = w10839 & w54796;
assign w10849 = pi00415 & w10848;
assign w10850 = w10848 & w54826;
assign w10851 = pi00417 & pi00418;
assign w10852 = w10848 & w55740;
assign w10853 = w10848 & w55741;
assign w10854 = w10848 & w55742;
assign w10855 = pi00420 & pi00421;
assign w10856 = w10848 & w55743;
assign w10857 = ~pi00403 & ~w10733;
assign w10858 = ~w10733 & w55744;
assign w10859 = ~w10733 & ~w10856;
assign w10860 = ~w10723 & ~w10859;
assign w10861 = (pi00403 & w10859) | (pi00403 & w55745) | (w10859 & w55745);
assign w10862 = ~pi00251 & w10728;
assign w10863 = (~pi00252 & w10735) | (~pi00252 & w55746) | (w10735 & w55746);
assign w10864 = ~w10862 & ~w10863;
assign w10865 = ~w10858 & w10864;
assign w10866 = ~w10861 & w10865;
assign w10867 = (pi00293 & w10735) | (pi00293 & w55747) | (w10735 & w55747);
assign w10868 = pi00407 & w10839;
assign w10869 = w10839 & w55748;
assign w10870 = w10839 & w55749;
assign w10871 = w10839 & w55750;
assign w10872 = w10839 & w55751;
assign w10873 = pi00404 & w10872;
assign w10874 = ~w10733 & ~w10873;
assign w10875 = ~w10723 & ~w10874;
assign w10876 = (pi00404 & w10874) | (pi00404 & w55752) | (w10874 & w55752);
assign w10877 = ~w10733 & w55753;
assign w10878 = pi00290 & w10728;
assign w10879 = ~w10867 & ~w10878;
assign w10880 = ~w10877 & w10879;
assign w10881 = ~w10876 & w10880;
assign w10882 = ~w10733 & w55754;
assign w10883 = ~pi00405 & w10851;
assign w10884 = w10882 & w10883;
assign w10885 = ~w10733 & ~w10852;
assign w10886 = (pi00405 & w10885) | (pi00405 & w55755) | (w10885 & w55755);
assign w10887 = (pi00225 & w10735) | (pi00225 & w55756) | (w10735 & w55756);
assign w10888 = pi00221 & w10728;
assign w10889 = ~w10887 & ~w10888;
assign w10890 = ~w10884 & w10889;
assign w10891 = ~w10886 & w10890;
assign w10892 = pi00117 & w10728;
assign w10893 = ~w10733 & ~w10839;
assign w10894 = ~w10723 & ~w10893;
assign w10895 = (pi00406 & w10893) | (pi00406 & w55757) | (w10893 & w55757);
assign w10896 = ~w10733 & w55758;
assign w10897 = (pi00123 & w10735) | (pi00123 & w55759) | (w10735 & w55759);
assign w10898 = ~w10892 & ~w10897;
assign w10899 = ~w10896 & w10898;
assign w10900 = ~w10895 & w10899;
assign w10901 = (pi00407 & w10893) | (pi00407 & w55760) | (w10893 & w55760);
assign w10902 = pi00129 & w10728;
assign w10903 = (pi00135 & w10735) | (pi00135 & w55761) | (w10735 & w55761);
assign w10904 = ~w10733 & w55762;
assign w10905 = ~w10902 & ~w10903;
assign w10906 = ~w10904 & w10905;
assign w10907 = ~w10901 & w10906;
assign w10908 = ~w10733 & w55763;
assign w10909 = ~w10733 & ~w10869;
assign w10910 = (pi00408 & w10909) | (pi00408 & w55764) | (w10909 & w55764);
assign w10911 = pi00182 & w10728;
assign w10912 = (pi00183 & w10735) | (pi00183 & w55765) | (w10735 & w55765);
assign w10913 = ~w10911 & ~w10912;
assign w10914 = ~w10908 & w10913;
assign w10915 = ~w10910 & w10914;
assign w10916 = pi00304 & w10728;
assign w10917 = ~w10733 & ~w10871;
assign w10918 = ~w10723 & ~w10917;
assign w10919 = (pi00409 & w10917) | (pi00409 & w55766) | (w10917 & w55766);
assign w10920 = ~w10733 & w55767;
assign w10921 = (pi00306 & w10735) | (pi00306 & w55768) | (w10735 & w55768);
assign w10922 = ~w10916 & ~w10921;
assign w10923 = ~w10920 & w10922;
assign w10924 = ~w10919 & w10923;
assign w10925 = ~w10733 & w55769;
assign w10926 = pi00410 & ~w10918;
assign w10927 = pi00305 & w10728;
assign w10928 = (pi00307 & w10735) | (pi00307 & w55770) | (w10735 & w55770);
assign w10929 = ~w10927 & ~w10928;
assign w10930 = ~w10925 & w10929;
assign w10931 = ~w10926 & w10930;
assign w10932 = ~w10733 & w55771;
assign w10933 = pi00411 & ~w10875;
assign w10934 = (pi00287 & w10735) | (pi00287 & w55772) | (w10735 & w55772);
assign w10935 = pi00284 & w10728;
assign w10936 = ~w10934 & ~w10935;
assign w10937 = ~w10932 & w10936;
assign w10938 = ~w10933 & w10937;
assign w10939 = ~w10733 & ~w10846;
assign w10940 = ~w10733 & w55774;
assign w10941 = (pi00412 & ~w10894) | (pi00412 & w55775) | (~w10894 & w55775);
assign w10942 = pi00261 & w10728;
assign w10943 = (pi00264 & w10735) | (pi00264 & w55776) | (w10735 & w55776);
assign w10944 = ~w10942 & ~w10943;
assign w10945 = ~w10941 & w10944;
assign w10946 = ~w10940 & w10945;
assign w10947 = pi00285 & w10728;
assign w10948 = (pi00413 & ~w10894) | (pi00413 & w55777) | (~w10894 & w55777);
assign w10949 = pi00289 & ~w10736;
assign w10950 = ~w10733 & w55778;
assign w10951 = ~w10947 & ~w10949;
assign w10952 = ~w10950 & w10951;
assign w10953 = ~w10948 & w10952;
assign w10954 = pi00096 & w10728;
assign w10955 = (pi00414 & w10734) | (pi00414 & w55779) | (w10734 & w55779);
assign w10956 = pi00099 & ~w10736;
assign w10957 = pi00375 & ~pi00414;
assign w10958 = ~w10733 & w10957;
assign w10959 = ~w10954 & ~w10956;
assign w10960 = ~w10958 & w10959;
assign w10961 = ~w10955 & w10960;
assign w10962 = (pi00288 & w10735) | (pi00288 & w55780) | (w10735 & w55780);
assign w10963 = ~pi00415 & ~w10848;
assign w10964 = ~w10733 & w55781;
assign w10965 = pi00286 & w10728;
assign w10966 = pi00415 & w10723;
assign w10967 = ~w10962 & ~w10965;
assign w10968 = ~w10966 & w10967;
assign w10969 = ~w10964 & w10968;
assign w10970 = pi00262 & w10728;
assign w10971 = ~w10733 & ~w10850;
assign w10972 = ~w10723 & ~w10971;
assign w10973 = (~pi00416 & w10733) | (~pi00416 & w55782) | (w10733 & w55782);
assign w10974 = ~w10972 & ~w10973;
assign w10975 = (pi00265 & w10735) | (pi00265 & w55783) | (w10735 & w55783);
assign w10976 = ~w10970 & ~w10975;
assign w10977 = ~w10974 & w10976;
assign w10978 = (pi00227 & w10735) | (pi00227 & w55784) | (w10735 & w55784);
assign w10979 = (pi00417 & w10971) | (pi00417 & w55785) | (w10971 & w55785);
assign w10980 = ~pi00417 & w10882;
assign w10981 = pi00219 & w10728;
assign w10982 = ~w10978 & ~w10981;
assign w10983 = ~w10980 & w10982;
assign w10984 = ~w10979 & w10983;
assign w10985 = w10848 & w55786;
assign w10986 = ~w10733 & w55787;
assign w10987 = (pi00418 & w10885) | (pi00418 & w55788) | (w10885 & w55788);
assign w10988 = pi00220 & w10728;
assign w10989 = (pi00228 & w10735) | (pi00228 & w55789) | (w10735 & w55789);
assign w10990 = ~w10988 & ~w10989;
assign w10991 = ~w10986 & w10990;
assign w10992 = ~w10987 & w10991;
assign w10993 = (pi00224 & w10735) | (pi00224 & w55790) | (w10735 & w55790);
assign w10994 = ~w10733 & ~w10854;
assign w10995 = (pi00419 & w10994) | (pi00419 & w55791) | (w10994 & w55791);
assign w10996 = ~w10733 & w55792;
assign w10997 = pi00222 & w10728;
assign w10998 = ~w10993 & ~w10997;
assign w10999 = ~w10996 & w10998;
assign w11000 = ~w10995 & w10999;
assign w11001 = (pi00200 & w10735) | (pi00200 & w55793) | (w10735 & w55793);
assign w11002 = (pi00420 & w10994) | (pi00420 & w55794) | (w10994 & w55794);
assign w11003 = ~w10733 & w55795;
assign w11004 = pi00199 & w10728;
assign w11005 = ~w11001 & ~w11004;
assign w11006 = ~w11003 & w11005;
assign w11007 = ~w11002 & w11006;
assign w11008 = (pi00421 & w10859) | (pi00421 & w55796) | (w10859 & w55796);
assign w11009 = (pi00266 & w10735) | (pi00266 & w55797) | (w10735 & w55797);
assign w11010 = pi00263 & w10728;
assign w11011 = pi00420 & ~pi00421;
assign w11012 = ~w10733 & w55798;
assign w11013 = ~w11009 & ~w11010;
assign w11014 = ~w11012 & w11013;
assign w11015 = ~w11008 & w11014;
assign w11016 = (pi00422 & ~w10860) | (pi00422 & w55799) | (~w10860 & w55799);
assign w11017 = ~pi00226 & ~w10736;
assign w11018 = ~pi00223 & w10728;
assign w11019 = pi00403 & ~pi00422;
assign w11020 = ~w10733 & w55800;
assign w11021 = ~w11017 & ~w11018;
assign w11022 = ~w11020 & w11021;
assign w11023 = ~w11016 & w11022;
assign w11024 = pi00120 & w10728;
assign w11025 = ~w10733 & ~w10831;
assign w11026 = (pi00423 & w11025) | (pi00423 & w55801) | (w11025 & w55801);
assign w11027 = (pi00126 & w10735) | (pi00126 & w55802) | (w10735 & w55802);
assign w11028 = w10830 & w55803;
assign w11029 = ~w10733 & w11028;
assign w11030 = ~w11024 & ~w11027;
assign w11031 = ~w11029 & w11030;
assign w11032 = ~w11026 & w11031;
assign w11033 = (pi00181 & w10735) | (pi00181 & w55804) | (w10735 & w55804);
assign w11034 = ~w10733 & ~w10833;
assign w11035 = (pi00424 & w11034) | (pi00424 & w55805) | (w11034 & w55805);
assign w11036 = ~w10733 & w55806;
assign w11037 = pi00180 & w10728;
assign w11038 = ~w11033 & ~w11037;
assign w11039 = ~w11036 & w11038;
assign w11040 = ~w11035 & w11039;
assign w11041 = pi00121 & w10728;
assign w11042 = (pi00425 & w11034) | (pi00425 & w55807) | (w11034 & w55807);
assign w11043 = pi00127 & ~w10736;
assign w11044 = w10832 & w55808;
assign w11045 = ~w10733 & w11044;
assign w11046 = ~w11041 & ~w11043;
assign w11047 = ~w11045 & w11046;
assign w11048 = ~w11042 & w11047;
assign w11049 = (pi00136 & w10735) | (pi00136 & w55809) | (w10735 & w55809);
assign w11050 = ~w10733 & ~w10835;
assign w11051 = (pi00426 & w11050) | (pi00426 & w55810) | (w11050 & w55810);
assign w11052 = ~w10733 & w55811;
assign w11053 = pi00131 & w10728;
assign w11054 = ~w11049 & ~w11053;
assign w11055 = ~w11052 & w11054;
assign w11056 = ~w11051 & w11055;
assign w11057 = pi00115 & w10728;
assign w11058 = (pi00427 & w11050) | (pi00427 & w55812) | (w11050 & w55812);
assign w11059 = pi00130 & ~w10736;
assign w11060 = ~pi00427 & w10835;
assign w11061 = ~w10733 & w11060;
assign w11062 = ~w11057 & ~w11059;
assign w11063 = ~w11061 & w11062;
assign w11064 = ~w11058 & w11063;
assign w11065 = (pi00097 & w10735) | (pi00097 & w55813) | (w10735 & w55813);
assign w11066 = ~w10733 & ~w10837;
assign w11067 = (pi00428 & w11066) | (pi00428 & w55814) | (w11066 & w55814);
assign w11068 = ~w10733 & w55815;
assign w11069 = pi00094 & w10728;
assign w11070 = ~w11065 & ~w11069;
assign w11071 = ~w11068 & w11070;
assign w11072 = ~w11067 & w11071;
assign w11073 = w10835 & w55816;
assign w11074 = ~w10733 & w11073;
assign w11075 = (pi00429 & w11066) | (pi00429 & w55817) | (w11066 & w55817);
assign w11076 = pi00134 & ~w10736;
assign w11077 = pi00128 & w10728;
assign w11078 = ~w11074 & ~w11076;
assign w11079 = ~w11077 & w11078;
assign w11080 = ~w11075 & w11079;
assign w11081 = pi00430 & w10711;
assign w11082 = w10722 & ~w11081;
assign w11083 = (pi00122 & w10735) | (pi00122 & w55818) | (w10735 & w55818);
assign w11084 = (pi00431 & w10909) | (pi00431 & w55819) | (w10909 & w55819);
assign w11085 = w10868 & w10909;
assign w11086 = pi00125 & w10728;
assign w11087 = ~w11083 & ~w11086;
assign w11088 = ~w11085 & w11087;
assign w11089 = ~w11084 & w11088;
assign w11090 = (pi00124 & w10735) | (pi00124 & w55820) | (w10735 & w55820);
assign w11091 = (pi00432 & w11025) | (pi00432 & w55821) | (w11025 & w55821);
assign w11092 = w10830 & w11025;
assign w11093 = pi00119 & w10728;
assign w11094 = ~w11090 & ~w11093;
assign w11095 = ~w11092 & w11094;
assign w11096 = ~w11091 & w11095;
assign w11097 = ~pi00433 & w10723;
assign w11098 = pi00434 & ~pi00869;
assign w11099 = ~w149 & ~w158;
assign w11100 = ~w642 & w749;
assign w11101 = w11099 & w11100;
assign w11102 = w10680 & w11101;
assign w11103 = ~w11098 & ~w11102;
assign w11104 = w10688 & w55822;
assign w11105 = w10706 & w11104;
assign w11106 = ~w10703 & w10712;
assign w11107 = ~w10713 & w11104;
assign w11108 = w10707 & ~w11107;
assign w11109 = ~w11106 & w11108;
assign w11110 = (~w11105 & ~w11108) | (~w11105 & w55823) | (~w11108 & w55823);
assign w11111 = ~pi00435 & ~w11110;
assign w11112 = w10711 & ~w11111;
assign w11113 = pi09926 & pi09963;
assign w11114 = ~pi09819 & ~pi09912;
assign w11115 = ~w11113 & w11114;
assign w11116 = (pi00250 & ~w25) | (pi00250 & w55825) | (~w25 & w55825);
assign w11117 = ~w11116 & w55826;
assign w11118 = pi00812 & w11116;
assign w11119 = ~w11117 & ~w11118;
assign w11120 = pi00437 & pi10546;
assign w11121 = ~pi10345 & w1121;
assign w11122 = ~w11120 & ~w11121;
assign w11123 = w830 & w55827;
assign w11124 = pi10006 & ~w11123;
assign w11125 = w830 & w55828;
assign w11126 = pi02665 & ~pi10418;
assign w11127 = w2041 & w2049;
assign w11128 = pi00870 & ~pi01209;
assign w11129 = ~pi01217 & ~pi01262;
assign w11130 = ~pi01463 & w11129;
assign w11131 = w11126 & w11128;
assign w11132 = w11130 & w11131;
assign w11133 = w2041 & w55829;
assign w11134 = ~w11125 & ~w11133;
assign w11135 = pi00440 & ~w11110;
assign w11136 = w10723 & ~w11135;
assign w11137 = w10694 & w55830;
assign w11138 = (~w10688 & w55831) | (~w10688 & w55832) | (w55831 & w55832);
assign w11139 = w11106 & ~w11137;
assign w11140 = w11139 & w55833;
assign w11141 = ~pi00441 & ~w11140;
assign w11142 = w11108 & ~w11141;
assign w11143 = ~w11105 & ~w11140;
assign w11144 = pi00457 & w10698;
assign w11145 = w10698 & w55834;
assign w11146 = w11143 & ~w11145;
assign w11147 = pi00442 & w11146;
assign w11148 = pi00459 & w10698;
assign w11149 = pi01217 & pi01262;
assign w11150 = (~pi00268 & w2049) | (~pi00268 & w55835) | (w2049 & w55835);
assign w11151 = pi00209 & ~w11150;
assign w11152 = ~pi01209 & ~w11149;
assign w11153 = (w11152 & ~w2040) | (w11152 & w55836) | (~w2040 & w55836);
assign w11154 = ~w11143 & w11153;
assign w11155 = ~w11148 & ~w11154;
assign w11156 = ~w11147 & w11155;
assign w11157 = ~pi00443 & w2927;
assign w11158 = w25 & w55837;
assign w11159 = ~w11157 & ~w11158;
assign w11160 = ~pi00025 & pi10543;
assign w11161 = pi00444 & ~w11160;
assign w11162 = pi00535 & w11160;
assign w11163 = ~w11161 & ~w11162;
assign w11164 = pi10047 & pi10360;
assign w11165 = pi00445 & ~w11164;
assign w11166 = w832 & w11165;
assign w11167 = pi00292 & w11164;
assign w11168 = w2041 & w11167;
assign w11169 = ~w11166 & ~w11168;
assign w11170 = pi00446 & ~w11164;
assign w11171 = w832 & w11170;
assign w11172 = pi00291 & w11164;
assign w11173 = w2041 & w11172;
assign w11174 = ~w11171 & ~w11173;
assign w11175 = ~pi00845 & pi10445;
assign w11176 = ~pi00113 & ~pi00177;
assign w11177 = pi00845 & w11126;
assign w11178 = w11176 & w11177;
assign w11179 = (~w11175 & ~w11177) | (~w11175 & w55838) | (~w11177 & w55838);
assign w11180 = pi10000 & w11126;
assign w11181 = w11179 & w55839;
assign w11182 = pi00113 & pi00177;
assign w11183 = w11175 & w11182;
assign w11184 = (pi01187 & w11178) | (pi01187 & w55840) | (w11178 & w55840);
assign w11185 = w11175 & w11176;
assign w11186 = pi01171 & w11185;
assign w11187 = pi00113 & ~pi00177;
assign w11188 = w11175 & w11187;
assign w11189 = pi01178 & w11188;
assign w11190 = ~pi00113 & pi00177;
assign w11191 = w11175 & w11190;
assign w11192 = pi01201 & w11191;
assign w11193 = w11126 & w55841;
assign w11194 = pi01271 & w11193;
assign w11195 = w11179 & w11194;
assign w11196 = pi00611 & w11195;
assign w11197 = w11179 & w11180;
assign w11198 = ~pi01270 & ~pi01271;
assign w11199 = pi00627 & w11198;
assign w11200 = ~pi01270 & pi01271;
assign w11201 = pi00639 & w11200;
assign w11202 = pi01270 & ~pi01271;
assign w11203 = pi00618 & w11202;
assign w11204 = ~w11199 & ~w11201;
assign w11205 = ~w11203 & w11204;
assign w11206 = w11197 & ~w11205;
assign w11207 = ~w11186 & ~w11189;
assign w11208 = ~w11192 & w11207;
assign w11209 = w11208 & w55842;
assign w11210 = ~w11196 & ~w11206;
assign w11211 = w11209 & w11210;
assign w11212 = w11179 & w55843;
assign w11213 = (pi01188 & w11178) | (pi01188 & w55844) | (w11178 & w55844);
assign w11214 = pi01179 & w11188;
assign w11215 = pi01182 & w11185;
assign w11216 = pi01202 & w11191;
assign w11217 = pi00622 & w11195;
assign w11218 = pi00628 & w11198;
assign w11219 = pi00641 & w11200;
assign w11220 = pi00619 & w11202;
assign w11221 = ~w11218 & ~w11219;
assign w11222 = ~w11220 & w11221;
assign w11223 = w11197 & ~w11222;
assign w11224 = ~w11214 & ~w11215;
assign w11225 = ~w11216 & w11224;
assign w11226 = w11225 & w55845;
assign w11227 = ~w11217 & ~w11223;
assign w11228 = w11226 & w11227;
assign w11229 = w11179 & w55846;
assign w11230 = (pi01189 & w11178) | (pi01189 & w55847) | (w11178 & w55847);
assign w11231 = pi01172 & w11191;
assign w11232 = pi01180 & w11188;
assign w11233 = pi01193 & w11185;
assign w11234 = pi00633 & w11195;
assign w11235 = pi00620 & w11202;
assign w11236 = pi00629 & w11198;
assign w11237 = pi00612 & w11200;
assign w11238 = ~w11235 & ~w11236;
assign w11239 = ~w11237 & w11238;
assign w11240 = w11197 & ~w11239;
assign w11241 = ~w11231 & ~w11232;
assign w11242 = ~w11233 & w11241;
assign w11243 = w11242 & w55848;
assign w11244 = ~w11234 & ~w11240;
assign w11245 = w11243 & w11244;
assign w11246 = w11179 & w55849;
assign w11247 = (pi01190 & w11178) | (pi01190 & w55850) | (w11178 & w55850);
assign w11248 = pi01173 & w11191;
assign w11249 = pi01181 & w11188;
assign w11250 = pi01196 & w11185;
assign w11251 = pi00642 & w11195;
assign w11252 = pi00613 & w11200;
assign w11253 = pi00621 & w11202;
assign w11254 = pi00630 & w11198;
assign w11255 = ~w11252 & ~w11253;
assign w11256 = ~w11254 & w11255;
assign w11257 = w11197 & ~w11256;
assign w11258 = ~w11248 & ~w11249;
assign w11259 = ~w11250 & w11258;
assign w11260 = w11259 & w55851;
assign w11261 = ~w11251 & ~w11257;
assign w11262 = w11260 & w11261;
assign w11263 = pi00636 & w11195;
assign w11264 = (pi01191 & w11178) | (pi01191 & w55852) | (w11178 & w55852);
assign w11265 = pi01174 & w11191;
assign w11266 = pi01183 & w11188;
assign w11267 = pi01197 & w11185;
assign w11268 = w11179 & w55853;
assign w11269 = pi00614 & w11200;
assign w11270 = pi00623 & w11202;
assign w11271 = pi00631 & w11198;
assign w11272 = ~w11269 & ~w11270;
assign w11273 = ~w11271 & w11272;
assign w11274 = w11197 & ~w11273;
assign w11275 = ~w11265 & ~w11266;
assign w11276 = ~w11267 & w11275;
assign w11277 = ~w11264 & w11276;
assign w11278 = ~w11263 & w11277;
assign w11279 = ~w11268 & ~w11274;
assign w11280 = w11278 & w11279;
assign w11281 = pi00640 & w11195;
assign w11282 = (pi01195 & w11178) | (pi01195 & w55854) | (w11178 & w55854);
assign w11283 = pi01177 & w11191;
assign w11284 = pi01186 & w11188;
assign w11285 = pi01200 & w11185;
assign w11286 = w11179 & w55855;
assign w11287 = pi00626 & w11202;
assign w11288 = pi00635 & w11198;
assign w11289 = pi00617 & w11200;
assign w11290 = ~w11287 & ~w11288;
assign w11291 = ~w11289 & w11290;
assign w11292 = w11197 & ~w11291;
assign w11293 = ~w11283 & ~w11284;
assign w11294 = ~w11285 & w11293;
assign w11295 = ~w11282 & w11294;
assign w11296 = ~w11281 & w11295;
assign w11297 = ~w11286 & ~w11292;
assign w11298 = w11296 & w11297;
assign w11299 = pi00637 & w11195;
assign w11300 = (pi01194 & w11178) | (pi01194 & w55856) | (w11178 & w55856);
assign w11301 = pi01176 & w11191;
assign w11302 = pi01185 & w11188;
assign w11303 = pi01199 & w11185;
assign w11304 = w11179 & w55857;
assign w11305 = pi00625 & w11202;
assign w11306 = pi00634 & w11198;
assign w11307 = pi00616 & w11200;
assign w11308 = ~w11305 & ~w11306;
assign w11309 = ~w11307 & w11308;
assign w11310 = w11197 & ~w11309;
assign w11311 = ~w11301 & ~w11302;
assign w11312 = ~w11303 & w11311;
assign w11313 = ~w11300 & w11312;
assign w11314 = ~w11299 & w11313;
assign w11315 = ~w11304 & ~w11310;
assign w11316 = w11314 & w11315;
assign w11317 = pi00638 & w11195;
assign w11318 = (pi01192 & w11178) | (pi01192 & w55858) | (w11178 & w55858);
assign w11319 = pi01175 & w11191;
assign w11320 = pi01184 & w11188;
assign w11321 = pi01198 & w11185;
assign w11322 = w11179 & w55859;
assign w11323 = pi00632 & w11198;
assign w11324 = pi00615 & w11200;
assign w11325 = pi00624 & w11202;
assign w11326 = ~w11323 & ~w11324;
assign w11327 = ~w11325 & w11326;
assign w11328 = w11197 & ~w11327;
assign w11329 = ~w11319 & ~w11320;
assign w11330 = ~w11321 & w11329;
assign w11331 = ~w11318 & w11330;
assign w11332 = ~w11317 & w11331;
assign w11333 = ~w11322 & ~w11328;
assign w11334 = w11332 & w11333;
assign w11335 = ~pi10031 & ~pi10356;
assign w11336 = ~pi02648 & w11335;
assign w11337 = w11335 & w54827;
assign w11338 = ~pi01204 & w11337;
assign w11339 = w11337 & w55860;
assign w11340 = w11337 & w55861;
assign w11341 = ~pi01205 & w11340;
assign w11342 = w11340 & w55862;
assign w11343 = (~pi00455 & ~w11340) | (~pi00455 & w55863) | (~w11340 & w55863);
assign w11344 = pi00962 & ~pi01306;
assign w11345 = pi01309 & w11344;
assign w11346 = ~pi01213 & ~pi01275;
assign w11347 = ~pi01308 & w11346;
assign w11348 = pi00957 & pi01305;
assign w11349 = w11345 & w11348;
assign w11350 = w11347 & w11349;
assign w11351 = w11349 & w55864;
assign w11352 = ~pi01309 & pi09863;
assign w11353 = pi01309 & ~pi09863;
assign w11354 = ~w11352 & ~w11353;
assign w11355 = w11346 & w55865;
assign w11356 = ~pi01306 & ~pi01307;
assign w11357 = w11355 & w11356;
assign w11358 = pi00962 & ~w11354;
assign w11359 = w11357 & w11358;
assign w11360 = pi09851 & w11359;
assign w11361 = w11344 & w55866;
assign w11362 = w11355 & w11361;
assign w11363 = w11349 & w55867;
assign w11364 = pi09827 & w11363;
assign w11365 = (~w11362 & ~w11351) | (~w11362 & w55868) | (~w11351 & w55868);
assign w11366 = ~w11360 & ~w11364;
assign w11367 = (w11342 & ~w11366) | (w11342 & w55869) | (~w11366 & w55869);
assign w11368 = w11342 & ~w11359;
assign w11369 = ~w11350 & ~w11362;
assign w11370 = w11368 & w11369;
assign w11371 = ~pi00485 & w11370;
assign w11372 = ~w11343 & ~w11367;
assign w11373 = ~w11371 & w11372;
assign w11374 = ~pi00469 & w11370;
assign w11375 = (pi00456 & ~w11340) | (pi00456 & w55870) | (~w11340 & w55870);
assign w11376 = pi09810 & w11362;
assign w11377 = ~pi09836 & w11351;
assign w11378 = pi09831 & w11363;
assign w11379 = ~w11376 & ~w11377;
assign w11380 = w11379 & w55871;
assign w11381 = ~w11375 & ~w11380;
assign w11382 = ~w11374 & ~w11381;
assign w11383 = ~pi00457 & ~w10698;
assign w11384 = w11143 & ~w11144;
assign w11385 = ~w11383 & w11384;
assign w11386 = ~w11140 & w55872;
assign w11387 = ~w11144 & ~w11386;
assign w11388 = ~w11145 & ~w11387;
assign w11389 = (~pi00459 & ~w10698) | (~pi00459 & w55873) | (~w10698 & w55873);
assign w11390 = pi00459 & ~w11146;
assign w11391 = ~w11389 & ~w11390;
assign w11392 = (pi00460 & w11109) | (pi00460 & w55874) | (w11109 & w55874);
assign w11393 = w10711 & ~w11392;
assign w11394 = (pi00461 & w11109) | (pi00461 & w55875) | (w11109 & w55875);
assign w11395 = w10722 & ~w11394;
assign w11396 = pi00462 & w10723;
assign w11397 = ~pi00089 & ~w10722;
assign w11398 = w10711 & ~w11397;
assign w11399 = ~pi00105 & ~w10722;
assign w11400 = ~w11396 & ~w11399;
assign w11401 = w11398 & w11400;
assign w11402 = (pi00824 & ~w799) | (pi00824 & w55876) | (~w799 & w55876);
assign w11403 = w799 & w55877;
assign w11404 = w671 & ~w11402;
assign w11405 = ~w11403 & w11404;
assign w11406 = ~pi00825 & w6042;
assign w11407 = (w671 & w6042) | (w671 & w55878) | (w6042 & w55878);
assign w11408 = ~w11406 & w11407;
assign w11409 = pi00610 & w76;
assign w11410 = (~pi00466 & ~w11340) | (~pi00466 & w55879) | (~w11340 & w55879);
assign w11411 = pi09829 & w11363;
assign w11412 = ~pi09853 & w11359;
assign w11413 = ~pi09835 & w11351;
assign w11414 = pi09811 & w11362;
assign w11415 = ~w11411 & ~w11414;
assign w11416 = ~w11412 & ~w11413;
assign w11417 = w11415 & w11416;
assign w11418 = ~pi00468 & w11370;
assign w11419 = (~w11410 & w11417) | (~w11410 & w55880) | (w11417 & w55880);
assign w11420 = ~w11418 & w11419;
assign w11421 = (~pi00467 & ~w11340) | (~pi00467 & w55881) | (~w11340 & w55881);
assign w11422 = pi09817 & w11363;
assign w11423 = ~pi09815 & w11351;
assign w11424 = pi00957 & w11359;
assign w11425 = pi09858 & w11362;
assign w11426 = ~w11422 & ~w11425;
assign w11427 = ~w11423 & ~w11424;
assign w11428 = w11426 & w11427;
assign w11429 = ~pi00466 & w11370;
assign w11430 = (~w11421 & w11428) | (~w11421 & w55882) | (w11428 & w55882);
assign w11431 = ~w11429 & w11430;
assign w11432 = (~pi00468 & ~w11340) | (~pi00468 & w55883) | (~w11340 & w55883);
assign w11433 = pi09828 & w11363;
assign w11434 = ~pi09852 & w11359;
assign w11435 = ~pi09834 & w11351;
assign w11436 = pi09854 & w11362;
assign w11437 = ~w11433 & ~w11436;
assign w11438 = ~w11434 & ~w11435;
assign w11439 = w11437 & w11438;
assign w11440 = ~pi00455 & w11370;
assign w11441 = (~w11432 & w11439) | (~w11432 & w55884) | (w11439 & w55884);
assign w11442 = ~w11440 & w11441;
assign w11443 = (~pi00469 & ~w11340) | (~pi00469 & w55885) | (~w11340 & w55885);
assign w11444 = pi09830 & w11363;
assign w11445 = ~pi00957 & w11359;
assign w11446 = ~pi09838 & w11351;
assign w11447 = pi09857 & w11362;
assign w11448 = ~w11444 & ~w11447;
assign w11449 = ~w11445 & ~w11446;
assign w11450 = w11448 & w11449;
assign w11451 = ~pi00467 & w11370;
assign w11452 = (~w11443 & w11450) | (~w11443 & w55886) | (w11450 & w55886);
assign w11453 = ~w11451 & w11452;
assign w11454 = pi00470 & w10722;
assign w11455 = w11398 & ~w11454;
assign w11456 = pi00471 & w10722;
assign w11457 = ~w10722 & w55887;
assign w11458 = w10711 & ~w11456;
assign w11459 = ~w11457 & w11458;
assign w11460 = ~pi01167 & w664;
assign w11461 = (w76 & w664) | (w76 & w55888) | (w664 & w55888);
assign w11462 = ~w11460 & w11461;
assign w11463 = ~w11116 & w55889;
assign w11464 = pi00886 & w11116;
assign w11465 = ~w11463 & ~w11464;
assign w11466 = pi00643 & w10718;
assign w11467 = ~pi01274 & ~pi01312;
assign w11468 = (pi01454 & ~w10686) | (pi01454 & w55890) | (~w10686 & w55890);
assign w11469 = w11467 & ~w11468;
assign w11470 = w11140 & ~w11469;
assign w11471 = ~w11107 & ~w11140;
assign w11472 = pi00540 & w10718;
assign w11473 = w10718 & w55891;
assign w11474 = w11471 & ~w11473;
assign w11475 = pi00474 & w11474;
assign w11476 = ~w11466 & ~w11470;
assign w11477 = ~w11475 & w11476;
assign w11478 = pi00475 & ~w11160;
assign w11479 = ~pi00036 & w11160;
assign w11480 = pi00034 & pi00035;
assign w11481 = pi00881 & ~w11480;
assign w11482 = w11479 & w11481;
assign w11483 = ~w11478 & ~w11482;
assign w11484 = w1209 & w55892;
assign w11485 = w1209 & w55893;
assign w11486 = ~pi10590 & ~pi10591;
assign w11487 = ~pi10592 & ~pi10593;
assign w11488 = ~pi10594 & ~pi10595;
assign w11489 = ~pi10596 & w11488;
assign w11490 = w11486 & w11487;
assign w11491 = w11489 & w11490;
assign w11492 = pi10597 & ~w11491;
assign w11493 = ~pi10598 & ~pi10599;
assign w11494 = ~pi10600 & ~pi10601;
assign w11495 = ~pi10602 & ~pi10603;
assign w11496 = ~pi10604 & ~pi10605;
assign w11497 = ~pi10606 & ~pi10607;
assign w11498 = ~pi10608 & ~pi10609;
assign w11499 = ~pi10610 & ~pi10611;
assign w11500 = ~pi10612 & ~pi10613;
assign w11501 = ~pi10614 & ~pi10615;
assign w11502 = ~pi10616 & ~pi10617;
assign w11503 = ~pi10618 & ~pi10619;
assign w11504 = ~pi10620 & ~pi10621;
assign w11505 = w11503 & w11504;
assign w11506 = w11501 & w11502;
assign w11507 = w11499 & w11500;
assign w11508 = w11497 & w11498;
assign w11509 = w11495 & w11496;
assign w11510 = w11493 & w11494;
assign w11511 = w11509 & w11510;
assign w11512 = w11507 & w11508;
assign w11513 = w11505 & w11506;
assign w11514 = w11512 & w11513;
assign w11515 = w11511 & w11514;
assign w11516 = w1277 & ~w11492;
assign w11517 = w11515 & w11516;
assign w11518 = (pi00477 & ~w11517) | (pi00477 & w55894) | (~w11517 & w55894);
assign w11519 = w11517 & w55895;
assign w11520 = ~w11518 & ~w11519;
assign w11521 = (pi00478 & ~w11517) | (pi00478 & w55896) | (~w11517 & w55896);
assign w11522 = w11517 & w55897;
assign w11523 = ~w11521 & ~w11522;
assign w11524 = (pi00479 & ~w11517) | (pi00479 & w55898) | (~w11517 & w55898);
assign w11525 = w11517 & w55899;
assign w11526 = ~w11524 & ~w11525;
assign w11527 = (pi00480 & ~w11517) | (pi00480 & w55900) | (~w11517 & w55900);
assign w11528 = w11517 & w55901;
assign w11529 = ~w11527 & ~w11528;
assign w11530 = (pi00481 & ~w11517) | (pi00481 & w55902) | (~w11517 & w55902);
assign w11531 = w11517 & w55903;
assign w11532 = ~w11530 & ~w11531;
assign w11533 = (pi00482 & ~w11517) | (pi00482 & w55904) | (~w11517 & w55904);
assign w11534 = w11517 & w55905;
assign w11535 = ~w11533 & ~w11534;
assign w11536 = (pi00483 & ~w11517) | (pi00483 & w55906) | (~w11517 & w55906);
assign w11537 = w11517 & w55907;
assign w11538 = ~w11536 & ~w11537;
assign w11539 = (pi00484 & ~w11517) | (pi00484 & w55908) | (~w11517 & w55908);
assign w11540 = w11517 & w55909;
assign w11541 = ~w11539 & ~w11540;
assign w11542 = (~pi00485 & ~w11340) | (~pi00485 & w55910) | (~w11340 & w55910);
assign w11543 = pi09850 & w11359;
assign w11544 = pi09826 & w11363;
assign w11545 = pi09832 & w11351;
assign w11546 = ~w11543 & ~w11544;
assign w11547 = (w11342 & ~w11546) | (w11342 & w55911) | (~w11546 & w55911);
assign w11548 = pi10589 & w11370;
assign w11549 = ~w11542 & ~w11547;
assign w11550 = ~w11548 & w11549;
assign w11551 = (~pi00486 & ~w11340) | (~pi00486 & w55912) | (~w11340 & w55912);
assign w11552 = pi09816 & w11363;
assign w11553 = ~pi09837 & w11351;
assign w11554 = pi09849 & w11362;
assign w11555 = ~w11552 & ~w11554;
assign w11556 = (w11342 & ~w11555) | (w11342 & w55913) | (~w11555 & w55913);
assign w11557 = ~pi00456 & w11370;
assign w11558 = ~w11551 & ~w11556;
assign w11559 = ~w11557 & w11558;
assign w11560 = ~pi00443 & pi09931;
assign w11561 = pi00487 & ~w11560;
assign w11562 = pi00875 & ~pi00877;
assign w11563 = ~pi00875 & pi00877;
assign w11564 = pi09991 & w11563;
assign w11565 = pi00875 & pi00877;
assign w11566 = pi10011 & w11565;
assign w11567 = ~pi00875 & ~pi00877;
assign w11568 = pi09913 & w11567;
assign w11569 = (pi00876 & ~w11562) | (pi00876 & w55914) | (~w11562 & w55914);
assign w11570 = ~w11564 & ~w11566;
assign w11571 = w11570 & w55915;
assign w11572 = pi09983 & w11563;
assign w11573 = pi10249 & w11565;
assign w11574 = pi09904 & w11567;
assign w11575 = (~pi00876 & ~w11562) | (~pi00876 & w55916) | (~w11562 & w55916);
assign w11576 = ~w11572 & ~w11573;
assign w11577 = w11576 & w55917;
assign w11578 = ~pi00005 & ~w11571;
assign w11579 = ~w11577 & w11578;
assign w11580 = pi00005 & pi00876;
assign w11581 = pi09914 & w11567;
assign w11582 = pi09936 & w11563;
assign w11583 = pi10259 & w11565;
assign w11584 = pi10014 & w11562;
assign w11585 = ~w11581 & ~w11582;
assign w11586 = ~w11583 & ~w11584;
assign w11587 = w11585 & w11586;
assign w11588 = pi00005 & ~pi00876;
assign w11589 = pi09905 & w11567;
assign w11590 = pi09940 & w11563;
assign w11591 = pi10250 & w11565;
assign w11592 = pi10244 & w11562;
assign w11593 = ~w11589 & ~w11590;
assign w11594 = ~w11591 & ~w11592;
assign w11595 = w11593 & w11594;
assign w11596 = w11588 & ~w11595;
assign w11597 = (pi00874 & w11587) | (pi00874 & w55918) | (w11587 & w55918);
assign w11598 = ~w11596 & w11597;
assign w11599 = ~w11579 & w11598;
assign w11600 = pi09938 & w11563;
assign w11601 = pi09908 & w11567;
assign w11602 = pi10246 & w11562;
assign w11603 = (~pi00876 & ~w11565) | (~pi00876 & w55919) | (~w11565 & w55919);
assign w11604 = ~w11600 & ~w11601;
assign w11605 = w11604 & w55920;
assign w11606 = pi10257 & w11562;
assign w11607 = pi10009 & w11565;
assign w11608 = pi09993 & w11563;
assign w11609 = (pi00876 & ~w11567) | (pi00876 & w55921) | (~w11567 & w55921);
assign w11610 = ~w11606 & ~w11607;
assign w11611 = w11610 & w55922;
assign w11612 = ~pi00005 & ~w11605;
assign w11613 = ~w11611 & w11612;
assign w11614 = pi09909 & w11567;
assign w11615 = pi09989 & w11563;
assign w11616 = pi10247 & w11562;
assign w11617 = pi10017 & w11565;
assign w11618 = ~w11614 & ~w11615;
assign w11619 = ~w11616 & ~w11617;
assign w11620 = w11618 & w11619;
assign w11621 = pi09798 & w11567;
assign w11622 = pi09934 & w11563;
assign w11623 = pi10233 & w11562;
assign w11624 = pi10007 & w11565;
assign w11625 = ~w11621 & ~w11622;
assign w11626 = ~w11623 & ~w11624;
assign w11627 = w11625 & w11626;
assign w11628 = w11580 & ~w11627;
assign w11629 = (~pi00874 & w11620) | (~pi00874 & w55923) | (w11620 & w55923);
assign w11630 = ~w11628 & w11629;
assign w11631 = ~w11613 & w11630;
assign w11632 = ~pi00001 & ~w11599;
assign w11633 = pi09992 & w11563;
assign w11634 = pi10010 & w11565;
assign w11635 = pi10255 & w11562;
assign w11636 = (pi00876 & ~w11567) | (pi00876 & w55924) | (~w11567 & w55924);
assign w11637 = ~w11633 & ~w11634;
assign w11638 = w11637 & w55925;
assign w11639 = pi10245 & w11562;
assign w11640 = pi09986 & w11563;
assign w11641 = pi10013 & w11565;
assign w11642 = (~pi00876 & ~w11567) | (~pi00876 & w55926) | (~w11567 & w55926);
assign w11643 = ~w11639 & ~w11640;
assign w11644 = w11643 & w55927;
assign w11645 = ~pi00005 & ~w11638;
assign w11646 = ~w11644 & w11645;
assign w11647 = pi09916 & w11567;
assign w11648 = pi09935 & w11563;
assign w11649 = pi10260 & w11565;
assign w11650 = pi10256 & w11562;
assign w11651 = ~w11647 & ~w11648;
assign w11652 = ~w11649 & ~w11650;
assign w11653 = w11651 & w11652;
assign w11654 = pi09907 & w11567;
assign w11655 = pi09987 & w11563;
assign w11656 = pi10251 & w11565;
assign w11657 = pi10019 & w11562;
assign w11658 = ~w11654 & ~w11655;
assign w11659 = ~w11656 & ~w11657;
assign w11660 = w11658 & w11659;
assign w11661 = w11588 & ~w11660;
assign w11662 = (pi00874 & w11653) | (pi00874 & w55918) | (w11653 & w55918);
assign w11663 = ~w11661 & w11662;
assign w11664 = ~w11646 & w11663;
assign w11665 = pi09910 & w11567;
assign w11666 = pi10015 & w11565;
assign w11667 = pi09990 & w11563;
assign w11668 = (~pi00876 & ~w11562) | (~pi00876 & w55928) | (~w11562 & w55928);
assign w11669 = ~w11665 & ~w11666;
assign w11670 = w11669 & w55929;
assign w11671 = pi10012 & w11562;
assign w11672 = pi10261 & w11565;
assign w11673 = pi09918 & w11567;
assign w11674 = (pi00876 & ~w11563) | (pi00876 & w55930) | (~w11563 & w55930);
assign w11675 = ~w11671 & ~w11672;
assign w11676 = w11675 & w55931;
assign w11677 = ~pi00005 & ~w11670;
assign w11678 = ~w11676 & w11677;
assign w11679 = pi09911 & w11567;
assign w11680 = pi09937 & w11563;
assign w11681 = pi10253 & w11565;
assign w11682 = pi10248 & w11562;
assign w11683 = ~w11679 & ~w11680;
assign w11684 = ~w11681 & ~w11682;
assign w11685 = w11683 & w11684;
assign w11686 = pi09919 & w11567;
assign w11687 = pi09995 & w11563;
assign w11688 = pi10258 & w11562;
assign w11689 = pi10008 & w11565;
assign w11690 = ~w11686 & ~w11687;
assign w11691 = ~w11688 & ~w11689;
assign w11692 = w11690 & w11691;
assign w11693 = w11580 & ~w11692;
assign w11694 = (~pi00874 & w11685) | (~pi00874 & w55923) | (w11685 & w55923);
assign w11695 = ~w11693 & w11694;
assign w11696 = ~w11678 & w11695;
assign w11697 = pi00001 & ~w11664;
assign w11698 = ~w11696 & w11697;
assign w11699 = (w11560 & ~w11632) | (w11560 & w55932) | (~w11632 & w55932);
assign w11700 = ~w11698 & w11699;
assign w11701 = w2927 & ~w11561;
assign w11702 = ~w11700 & w11701;
assign w11703 = (~pi00488 & ~w10718) | (~pi00488 & w10725) | (~w10718 & w10725);
assign w11704 = w11474 & ~w11703;
assign w11705 = pi00808 & ~pi00809;
assign w11706 = pi10469 & pi10510;
assign w11707 = pi10468 & pi10496;
assign w11708 = pi01274 & w10688;
assign w11709 = (w11707 & ~w10688) | (w11707 & w55933) | (~w10688 & w55933);
assign w11710 = pi00810 & ~w11706;
assign w11711 = w11709 & w55934;
assign w11712 = (pi00489 & ~w11711) | (pi00489 & w55935) | (~w11711 & w55935);
assign w11713 = w11711 & w55936;
assign w11714 = ~w11712 & ~w11713;
assign w11715 = (pi00490 & ~w11711) | (pi00490 & w55937) | (~w11711 & w55937);
assign w11716 = w11711 & w55938;
assign w11717 = ~w11715 & ~w11716;
assign w11718 = (pi00491 & ~w11711) | (pi00491 & w55939) | (~w11711 & w55939);
assign w11719 = w11711 & w55940;
assign w11720 = ~w11718 & ~w11719;
assign w11721 = (pi00492 & ~w11711) | (pi00492 & w55941) | (~w11711 & w55941);
assign w11722 = w11711 & w55942;
assign w11723 = ~w11721 & ~w11722;
assign w11724 = (pi00493 & ~w11711) | (pi00493 & w55943) | (~w11711 & w55943);
assign w11725 = w11711 & w55944;
assign w11726 = ~w11724 & ~w11725;
assign w11727 = (pi00494 & ~w11711) | (pi00494 & w55945) | (~w11711 & w55945);
assign w11728 = w11711 & w55946;
assign w11729 = ~w11727 & ~w11728;
assign w11730 = (pi00495 & ~w11711) | (pi00495 & w55947) | (~w11711 & w55947);
assign w11731 = w11711 & w55948;
assign w11732 = ~w11730 & ~w11731;
assign w11733 = ~pi00808 & pi00809;
assign w11734 = (pi00496 & ~w11711) | (pi00496 & w55949) | (~w11711 & w55949);
assign w11735 = w11711 & w55950;
assign w11736 = ~w11734 & ~w11735;
assign w11737 = (pi00497 & ~w11711) | (pi00497 & w55951) | (~w11711 & w55951);
assign w11738 = w11711 & w55952;
assign w11739 = ~w11737 & ~w11738;
assign w11740 = (pi00498 & ~w11711) | (pi00498 & w55953) | (~w11711 & w55953);
assign w11741 = w11711 & w55954;
assign w11742 = ~w11740 & ~w11741;
assign w11743 = (pi00499 & ~w11711) | (pi00499 & w55955) | (~w11711 & w55955);
assign w11744 = w11711 & w55956;
assign w11745 = ~w11743 & ~w11744;
assign w11746 = (pi00500 & ~w11711) | (pi00500 & w55957) | (~w11711 & w55957);
assign w11747 = w11711 & w55958;
assign w11748 = ~w11746 & ~w11747;
assign w11749 = (pi00501 & ~w11711) | (pi00501 & w55959) | (~w11711 & w55959);
assign w11750 = w11711 & w55960;
assign w11751 = ~w11749 & ~w11750;
assign w11752 = (pi00502 & ~w11711) | (pi00502 & w55961) | (~w11711 & w55961);
assign w11753 = w11711 & w55962;
assign w11754 = ~w11752 & ~w11753;
assign w11755 = (pi00503 & ~w11711) | (pi00503 & w55963) | (~w11711 & w55963);
assign w11756 = w11711 & w55964;
assign w11757 = ~w11755 & ~w11756;
assign w11758 = (pi00504 & ~w11711) | (pi00504 & w55965) | (~w11711 & w55965);
assign w11759 = w11711 & w55966;
assign w11760 = ~w11758 & ~w11759;
assign w11761 = ~pi00810 & ~w11706;
assign w11762 = w11709 & w55967;
assign w11763 = (pi00505 & ~w11762) | (pi00505 & w55968) | (~w11762 & w55968);
assign w11764 = w11762 & w55936;
assign w11765 = ~w11763 & ~w11764;
assign w11766 = (pi00506 & ~w11762) | (pi00506 & w55969) | (~w11762 & w55969);
assign w11767 = w11762 & w55938;
assign w11768 = ~w11766 & ~w11767;
assign w11769 = (pi00507 & ~w11762) | (pi00507 & w55970) | (~w11762 & w55970);
assign w11770 = w11762 & w55971;
assign w11771 = ~w11769 & ~w11770;
assign w11772 = (pi00508 & ~w11762) | (pi00508 & w55972) | (~w11762 & w55972);
assign w11773 = w11762 & w55973;
assign w11774 = ~w11772 & ~w11773;
assign w11775 = (pi00509 & ~w11762) | (pi00509 & w55974) | (~w11762 & w55974);
assign w11776 = w11762 & w55975;
assign w11777 = ~w11775 & ~w11776;
assign w11778 = (pi00510 & ~w11762) | (pi00510 & w55976) | (~w11762 & w55976);
assign w11779 = w11762 & w55977;
assign w11780 = ~w11778 & ~w11779;
assign w11781 = (pi00511 & ~w11762) | (pi00511 & w55978) | (~w11762 & w55978);
assign w11782 = w11762 & w55979;
assign w11783 = ~w11781 & ~w11782;
assign w11784 = (pi00512 & ~w11762) | (pi00512 & w55980) | (~w11762 & w55980);
assign w11785 = w11762 & w55944;
assign w11786 = ~w11784 & ~w11785;
assign w11787 = (pi00513 & ~w11762) | (pi00513 & w55981) | (~w11762 & w55981);
assign w11788 = w11762 & w55982;
assign w11789 = ~w11787 & ~w11788;
assign w11790 = (pi00514 & ~w11762) | (pi00514 & w55983) | (~w11762 & w55983);
assign w11791 = w11762 & w55984;
assign w11792 = ~w11790 & ~w11791;
assign w11793 = (pi00515 & ~w11762) | (pi00515 & w55985) | (~w11762 & w55985);
assign w11794 = w11762 & w55958;
assign w11795 = ~w11793 & ~w11794;
assign w11796 = (pi00516 & ~w11762) | (pi00516 & w55986) | (~w11762 & w55986);
assign w11797 = w11762 & w55987;
assign w11798 = ~w11796 & ~w11797;
assign w11799 = pi00808 & pi00809;
assign w11800 = w11709 & w55988;
assign w11801 = (pi00517 & ~w11800) | (pi00517 & w55989) | (~w11800 & w55989);
assign w11802 = w11800 & w55990;
assign w11803 = ~w11801 & ~w11802;
assign w11804 = (pi00518 & ~w11800) | (pi00518 & w55991) | (~w11800 & w55991);
assign w11805 = w11800 & w55992;
assign w11806 = ~w11804 & ~w11805;
assign w11807 = (pi00519 & ~w11800) | (pi00519 & w55993) | (~w11800 & w55993);
assign w11808 = w11800 & w55994;
assign w11809 = ~w11807 & ~w11808;
assign w11810 = (pi00520 & ~w11800) | (pi00520 & w55995) | (~w11800 & w55995);
assign w11811 = w11800 & w55996;
assign w11812 = ~w11810 & ~w11811;
assign w11813 = (pi00521 & ~w11800) | (pi00521 & w55997) | (~w11800 & w55997);
assign w11814 = w11800 & w55998;
assign w11815 = ~w11813 & ~w11814;
assign w11816 = (pi00522 & ~w11800) | (pi00522 & w55999) | (~w11800 & w55999);
assign w11817 = w11800 & w56000;
assign w11818 = ~w11816 & ~w11817;
assign w11819 = (pi00523 & ~w11800) | (pi00523 & w56001) | (~w11800 & w56001);
assign w11820 = w11800 & w56002;
assign w11821 = ~w11819 & ~w11820;
assign w11822 = (pi00524 & ~w11800) | (pi00524 & w56003) | (~w11800 & w56003);
assign w11823 = w11800 & w56004;
assign w11824 = ~w11822 & ~w11823;
assign w11825 = ~pi00808 & ~pi00809;
assign w11826 = pi00541 & ~w11706;
assign w11827 = w11709 & w11826;
assign w11828 = w11709 & w56005;
assign w11829 = (pi00525 & ~w11828) | (pi00525 & w56006) | (~w11828 & w56006);
assign w11830 = w11828 & w56007;
assign w11831 = ~w11829 & ~w11830;
assign w11832 = (pi00526 & ~w11828) | (pi00526 & w56008) | (~w11828 & w56008);
assign w11833 = w11828 & w56009;
assign w11834 = ~w11832 & ~w11833;
assign w11835 = (pi00527 & ~w11828) | (pi00527 & w56010) | (~w11828 & w56010);
assign w11836 = w11828 & w56011;
assign w11837 = ~w11835 & ~w11836;
assign w11838 = (pi00528 & ~w11828) | (pi00528 & w56012) | (~w11828 & w56012);
assign w11839 = w11828 & w56013;
assign w11840 = ~w11838 & ~w11839;
assign w11841 = (pi00529 & ~w11828) | (pi00529 & w56014) | (~w11828 & w56014);
assign w11842 = w11828 & w56015;
assign w11843 = ~w11841 & ~w11842;
assign w11844 = (pi00530 & ~w11828) | (pi00530 & w56016) | (~w11828 & w56016);
assign w11845 = w11828 & w56017;
assign w11846 = ~w11844 & ~w11845;
assign w11847 = (pi00531 & ~w11828) | (pi00531 & w56018) | (~w11828 & w56018);
assign w11848 = w11828 & w56019;
assign w11849 = ~w11847 & ~w11848;
assign w11850 = (pi00532 & ~w11828) | (pi00532 & w56020) | (~w11828 & w56020);
assign w11851 = w11828 & w56021;
assign w11852 = ~w11850 & ~w11851;
assign w11853 = (pi00533 & ~w11828) | (pi00533 & w56022) | (~w11828 & w56022);
assign w11854 = w11828 & w56023;
assign w11855 = ~w11853 & ~w11854;
assign w11856 = (pi00534 & ~w11828) | (pi00534 & w56024) | (~w11828 & w56024);
assign w11857 = w11828 & w56025;
assign w11858 = ~w11856 & ~w11857;
assign w11859 = ~pi00881 & ~pi10500;
assign w11860 = pi00881 & pi10500;
assign w11861 = ~w11859 & ~w11860;
assign w11862 = ~pi09821 & w6042;
assign w11863 = (w671 & w6042) | (w671 & w56026) | (w6042 & w56026);
assign w11864 = ~w11862 & w11863;
assign w11865 = ~pi01276 & w6048;
assign w11866 = (w671 & w6048) | (w671 & w56027) | (w6048 & w56027);
assign w11867 = ~w11865 & w11866;
assign w11868 = pi00833 & pi00834;
assign w11869 = pi00827 & pi00831;
assign w11870 = pi00832 & pi00835;
assign w11871 = pi00836 & pi00837;
assign w11872 = w11870 & w11871;
assign w11873 = w11868 & w11869;
assign w11874 = w11872 & w11873;
assign w11875 = pi00538 & pi00826;
assign w11876 = pi00828 & pi00829;
assign w11877 = pi00830 & pi00838;
assign w11878 = pi00839 & pi00840;
assign w11879 = w11877 & w11878;
assign w11880 = w11875 & w11876;
assign w11881 = w11879 & w11880;
assign w11882 = w11874 & w11881;
assign w11883 = w406 & w11882;
assign w11884 = (~pi09964 & w536) | (~pi09964 & w56028) | (w536 & w56028);
assign w11885 = ~w11882 & ~w11884;
assign w11886 = (w11874 & w11885) | (w11874 & w56029) | (w11885 & w56029);
assign w11887 = pi00838 & w11886;
assign w11888 = w11886 & w54828;
assign w11889 = w11886 & w56030;
assign w11890 = w11886 & w56031;
assign w11891 = w11886 & w56032;
assign w11892 = w11886 & w56033;
assign w11893 = w11886 & w56034;
assign w11894 = ~pi00538 & ~w11893;
assign w11895 = ~pi00037 & ~w573;
assign w11896 = (w11895 & ~w656) | (w11895 & w56035) | (~w656 & w56035);
assign w11897 = ~w11883 & w11896;
assign w11898 = ~w11894 & w11897;
assign w11899 = (~w789 & ~w762) | (~w789 & w56036) | (~w762 & w56036);
assign w11900 = ~w686 & ~w11899;
assign w11901 = ~w11140 & w56037;
assign w11902 = ~w10718 & ~w11901;
assign w11903 = ~w11472 & ~w11902;
assign w11904 = ~w11709 & ~w11826;
assign w11905 = ~w11827 & ~w11904;
assign w11906 = (pi00542 & ~w11711) | (pi00542 & w56038) | (~w11711 & w56038);
assign w11907 = w11711 & w56039;
assign w11908 = ~w11906 & ~w11907;
assign w11909 = (pi00543 & ~w11711) | (pi00543 & w56040) | (~w11711 & w56040);
assign w11910 = w11711 & w56041;
assign w11911 = ~w11909 & ~w11910;
assign w11912 = (pi00544 & ~w11711) | (pi00544 & w56042) | (~w11711 & w56042);
assign w11913 = w11711 & w56043;
assign w11914 = ~w11912 & ~w11913;
assign w11915 = (pi00545 & ~w11711) | (pi00545 & w56044) | (~w11711 & w56044);
assign w11916 = w11711 & w55975;
assign w11917 = ~w11915 & ~w11916;
assign w11918 = (pi00546 & ~w11711) | (pi00546 & w56045) | (~w11711 & w56045);
assign w11919 = w11711 & w55977;
assign w11920 = ~w11918 & ~w11919;
assign w11921 = (pi00547 & ~w11711) | (pi00547 & w56046) | (~w11711 & w56046);
assign w11922 = w11711 & w56047;
assign w11923 = ~w11921 & ~w11922;
assign w11924 = (pi00548 & ~w11711) | (pi00548 & w56048) | (~w11711 & w56048);
assign w11925 = w11711 & w55982;
assign w11926 = ~w11924 & ~w11925;
assign w11927 = (pi00549 & ~w11711) | (pi00549 & w56049) | (~w11711 & w56049);
assign w11928 = w11711 & w56050;
assign w11929 = ~w11927 & ~w11928;
assign w11930 = (pi00550 & ~w11711) | (pi00550 & w56051) | (~w11711 & w56051);
assign w11931 = w11711 & w56052;
assign w11932 = ~w11930 & ~w11931;
assign w11933 = (pi00551 & ~w11711) | (pi00551 & w56053) | (~w11711 & w56053);
assign w11934 = w11711 & w56054;
assign w11935 = ~w11933 & ~w11934;
assign w11936 = (pi00552 & ~w11711) | (pi00552 & w56055) | (~w11711 & w56055);
assign w11937 = w11711 & w56056;
assign w11938 = ~w11936 & ~w11937;
assign w11939 = (pi00553 & ~w11711) | (pi00553 & w56057) | (~w11711 & w56057);
assign w11940 = w11711 & w56058;
assign w11941 = ~w11939 & ~w11940;
assign w11942 = (pi00554 & ~w11711) | (pi00554 & w56059) | (~w11711 & w56059);
assign w11943 = w11711 & w56060;
assign w11944 = ~w11942 & ~w11943;
assign w11945 = (pi00555 & ~w11711) | (pi00555 & w56061) | (~w11711 & w56061);
assign w11946 = w11711 & w56062;
assign w11947 = ~w11945 & ~w11946;
assign w11948 = (pi00556 & ~w11762) | (pi00556 & w56063) | (~w11762 & w56063);
assign w11949 = w11762 & w56064;
assign w11950 = ~w11948 & ~w11949;
assign w11951 = (pi00557 & ~w11762) | (pi00557 & w56065) | (~w11762 & w56065);
assign w11952 = w11762 & w56041;
assign w11953 = ~w11951 & ~w11952;
assign w11954 = (pi00558 & ~w11762) | (pi00558 & w56066) | (~w11762 & w56066);
assign w11955 = w11762 & w56067;
assign w11956 = ~w11954 & ~w11955;
assign w11957 = (pi00559 & ~w11762) | (pi00559 & w56068) | (~w11762 & w56068);
assign w11958 = w11762 & w56069;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = (pi00560 & ~w11762) | (pi00560 & w56070) | (~w11762 & w56070);
assign w11961 = w11762 & w56071;
assign w11962 = ~w11960 & ~w11961;
assign w11963 = (pi00561 & ~w11762) | (pi00561 & w56072) | (~w11762 & w56072);
assign w11964 = w11762 & w55946;
assign w11965 = ~w11963 & ~w11964;
assign w11966 = (pi00562 & ~w11762) | (pi00562 & w56073) | (~w11762 & w56073);
assign w11967 = w11762 & w55948;
assign w11968 = ~w11966 & ~w11967;
assign w11969 = (pi00563 & ~w11762) | (pi00563 & w56074) | (~w11762 & w56074);
assign w11970 = w11762 & w56075;
assign w11971 = ~w11969 & ~w11970;
assign w11972 = (pi00564 & ~w11762) | (pi00564 & w56076) | (~w11762 & w56076);
assign w11973 = w11762 & w56077;
assign w11974 = ~w11972 & ~w11973;
assign w11975 = (pi00565 & ~w11762) | (pi00565 & w56078) | (~w11762 & w56078);
assign w11976 = w11762 & w55954;
assign w11977 = ~w11975 & ~w11976;
assign w11978 = (pi00566 & ~w11762) | (pi00566 & w56079) | (~w11762 & w56079);
assign w11979 = w11762 & w55960;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = (pi00567 & ~w11762) | (pi00567 & w56080) | (~w11762 & w56080);
assign w11982 = w11762 & w56081;
assign w11983 = ~w11981 & ~w11982;
assign w11984 = (pi00568 & ~w11762) | (pi00568 & w56082) | (~w11762 & w56082);
assign w11985 = w11762 & w56083;
assign w11986 = ~w11984 & ~w11985;
assign w11987 = (pi00569 & ~w11762) | (pi00569 & w56084) | (~w11762 & w56084);
assign w11988 = w11762 & w55962;
assign w11989 = ~w11987 & ~w11988;
assign w11990 = (pi00570 & ~w11762) | (pi00570 & w56085) | (~w11762 & w56085);
assign w11991 = w11762 & w56054;
assign w11992 = ~w11990 & ~w11991;
assign w11993 = (pi00571 & ~w11762) | (pi00571 & w56086) | (~w11762 & w56086);
assign w11994 = w11762 & w55964;
assign w11995 = ~w11993 & ~w11994;
assign w11996 = (pi00572 & ~w11762) | (pi00572 & w56087) | (~w11762 & w56087);
assign w11997 = w11762 & w56052;
assign w11998 = ~w11996 & ~w11997;
assign w11999 = (pi00573 & ~w11762) | (pi00573 & w56088) | (~w11762 & w56088);
assign w12000 = w11762 & w56060;
assign w12001 = ~w11999 & ~w12000;
assign w12002 = (pi00574 & ~w11762) | (pi00574 & w56089) | (~w11762 & w56089);
assign w12003 = w11762 & w56090;
assign w12004 = ~w12002 & ~w12003;
assign w12005 = (pi00575 & ~w11762) | (pi00575 & w56091) | (~w11762 & w56091);
assign w12006 = w11762 & w56092;
assign w12007 = ~w12005 & ~w12006;
assign w12008 = (pi00576 & ~w11800) | (pi00576 & w56093) | (~w11800 & w56093);
assign w12009 = w11800 & w56094;
assign w12010 = ~w12008 & ~w12009;
assign w12011 = (pi00577 & ~w11800) | (pi00577 & w56095) | (~w11800 & w56095);
assign w12012 = w11800 & w56096;
assign w12013 = ~w12011 & ~w12012;
assign w12014 = (pi00578 & ~w11800) | (pi00578 & w56097) | (~w11800 & w56097);
assign w12015 = w11800 & w56098;
assign w12016 = ~w12014 & ~w12015;
assign w12017 = (pi00579 & ~w11800) | (pi00579 & w56099) | (~w11800 & w56099);
assign w12018 = w11800 & w56100;
assign w12019 = ~w12017 & ~w12018;
assign w12020 = (pi00580 & ~w11800) | (pi00580 & w56101) | (~w11800 & w56101);
assign w12021 = w11800 & w56102;
assign w12022 = ~w12020 & ~w12021;
assign w12023 = (pi00581 & ~w11800) | (pi00581 & w56103) | (~w11800 & w56103);
assign w12024 = w11800 & w56104;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = (pi00582 & ~w11762) | (pi00582 & w56105) | (~w11762 & w56105);
assign w12027 = w11762 & w56106;
assign w12028 = ~w12026 & ~w12027;
assign w12029 = (pi00583 & ~w11800) | (pi00583 & w56107) | (~w11800 & w56107);
assign w12030 = w11800 & w56108;
assign w12031 = ~w12029 & ~w12030;
assign w12032 = (pi00584 & ~w11800) | (pi00584 & w56109) | (~w11800 & w56109);
assign w12033 = w11800 & w56110;
assign w12034 = ~w12032 & ~w12033;
assign w12035 = (pi00585 & ~w11800) | (pi00585 & w56111) | (~w11800 & w56111);
assign w12036 = w11800 & w56112;
assign w12037 = ~w12035 & ~w12036;
assign w12038 = (pi00586 & ~w11800) | (pi00586 & w56113) | (~w11800 & w56113);
assign w12039 = w11800 & w56114;
assign w12040 = ~w12038 & ~w12039;
assign w12041 = (pi00587 & ~w11800) | (pi00587 & w56115) | (~w11800 & w56115);
assign w12042 = w11800 & w56116;
assign w12043 = ~w12041 & ~w12042;
assign w12044 = (pi00588 & ~w11800) | (pi00588 & w56117) | (~w11800 & w56117);
assign w12045 = w11800 & w56118;
assign w12046 = ~w12044 & ~w12045;
assign w12047 = (pi00589 & ~w11800) | (pi00589 & w56119) | (~w11800 & w56119);
assign w12048 = w11800 & w56120;
assign w12049 = ~w12047 & ~w12048;
assign w12050 = (pi00590 & ~w11800) | (pi00590 & w56121) | (~w11800 & w56121);
assign w12051 = w11800 & w56122;
assign w12052 = ~w12050 & ~w12051;
assign w12053 = (pi00591 & ~w11800) | (pi00591 & w56123) | (~w11800 & w56123);
assign w12054 = w11800 & w56124;
assign w12055 = ~w12053 & ~w12054;
assign w12056 = (pi00592 & ~w11828) | (pi00592 & w56125) | (~w11828 & w56125);
assign w12057 = w11828 & w56126;
assign w12058 = ~w12056 & ~w12057;
assign w12059 = (pi00593 & ~w11828) | (pi00593 & w56127) | (~w11828 & w56127);
assign w12060 = w11828 & w56128;
assign w12061 = ~w12059 & ~w12060;
assign w12062 = (pi00594 & ~w11828) | (pi00594 & w56129) | (~w11828 & w56129);
assign w12063 = w11828 & w56130;
assign w12064 = ~w12062 & ~w12063;
assign w12065 = (pi00595 & ~w11828) | (pi00595 & w56131) | (~w11828 & w56131);
assign w12066 = w11828 & w56132;
assign w12067 = ~w12065 & ~w12066;
assign w12068 = (pi00596 & ~w11828) | (pi00596 & w56133) | (~w11828 & w56133);
assign w12069 = w11828 & w56134;
assign w12070 = ~w12068 & ~w12069;
assign w12071 = (pi00597 & ~w11828) | (pi00597 & w56135) | (~w11828 & w56135);
assign w12072 = w11828 & w56136;
assign w12073 = ~w12071 & ~w12072;
assign w12074 = (pi00598 & ~w11828) | (pi00598 & w56137) | (~w11828 & w56137);
assign w12075 = w11828 & w56138;
assign w12076 = ~w12074 & ~w12075;
assign w12077 = (pi00599 & ~w11828) | (pi00599 & w56139) | (~w11828 & w56139);
assign w12078 = w11828 & w56140;
assign w12079 = ~w12077 & ~w12078;
assign w12080 = (pi00600 & ~w11828) | (pi00600 & w56141) | (~w11828 & w56141);
assign w12081 = w11828 & w56142;
assign w12082 = ~w12080 & ~w12081;
assign w12083 = (pi00601 & ~w11828) | (pi00601 & w56143) | (~w11828 & w56143);
assign w12084 = w11828 & w56144;
assign w12085 = ~w12083 & ~w12084;
assign w12086 = (pi00602 & ~w11828) | (pi00602 & w56145) | (~w11828 & w56145);
assign w12087 = w11828 & w56146;
assign w12088 = ~w12086 & ~w12087;
assign w12089 = (pi00603 & ~w11828) | (pi00603 & w56147) | (~w11828 & w56147);
assign w12090 = w11828 & w56148;
assign w12091 = ~w12089 & ~w12090;
assign w12092 = (pi00604 & ~w11828) | (pi00604 & w56149) | (~w11828 & w56149);
assign w12093 = w11828 & w56150;
assign w12094 = ~w12092 & ~w12093;
assign w12095 = (pi00605 & ~w11828) | (pi00605 & w56151) | (~w11828 & w56151);
assign w12096 = w11828 & w56152;
assign w12097 = ~w12095 & ~w12096;
assign w12098 = (pi00606 & ~w11828) | (pi00606 & w56153) | (~w11828 & w56153);
assign w12099 = w11828 & w56154;
assign w12100 = ~w12098 & ~w12099;
assign w12101 = (pi00607 & ~w11800) | (pi00607 & w56155) | (~w11800 & w56155);
assign w12102 = w11800 & w55952;
assign w12103 = ~w12101 & ~w12102;
assign w12104 = w11762 & w11799;
assign w12105 = (pi00608 & ~w11762) | (pi00608 & w56156) | (~w11762 & w56156);
assign w12106 = w11762 & w56102;
assign w12107 = ~w12105 & ~w12106;
assign w12108 = pi00609 & ~w11160;
assign w12109 = pi00033 & w11480;
assign w12110 = w11160 & w56157;
assign w12111 = ~w12109 & w12110;
assign w12112 = ~w12108 & ~w12111;
assign w12113 = (~pi00064 & ~w146) | (~pi00064 & w56158) | (~w146 & w56158);
assign w12114 = w146 & w56159;
assign w12115 = w76 & ~w12113;
assign w12116 = ~w12114 & w12115;
assign w12117 = pi00845 & w11198;
assign w12118 = w11180 & w12117;
assign w12119 = ~w11175 & ~w12118;
assign w12120 = (pi01171 & ~w12119) | (pi01171 & w56160) | (~w12119 & w56160);
assign w12121 = w12119 & w56161;
assign w12122 = ~w12120 & ~w12121;
assign w12123 = (pi01172 & ~w12119) | (pi01172 & w56162) | (~w12119 & w56162);
assign w12124 = w12119 & w56163;
assign w12125 = ~w12123 & ~w12124;
assign w12126 = (pi01173 & ~w12119) | (pi01173 & w56164) | (~w12119 & w56164);
assign w12127 = w12119 & w56165;
assign w12128 = ~w12126 & ~w12127;
assign w12129 = (pi01174 & ~w12119) | (pi01174 & w56166) | (~w12119 & w56166);
assign w12130 = w12119 & w56167;
assign w12131 = ~w12129 & ~w12130;
assign w12132 = (pi01175 & ~w12119) | (pi01175 & w56168) | (~w12119 & w56168);
assign w12133 = w12119 & w56169;
assign w12134 = ~w12132 & ~w12133;
assign w12135 = (pi01176 & ~w12119) | (pi01176 & w56170) | (~w12119 & w56170);
assign w12136 = w12119 & w56171;
assign w12137 = ~w12135 & ~w12136;
assign w12138 = (pi01177 & ~w12119) | (pi01177 & w56172) | (~w12119 & w56172);
assign w12139 = w12119 & w56173;
assign w12140 = ~w12138 & ~w12139;
assign w12141 = (pi01178 & ~w12119) | (pi01178 & w56174) | (~w12119 & w56174);
assign w12142 = w12119 & w56175;
assign w12143 = ~w12141 & ~w12142;
assign w12144 = (pi01179 & ~w12119) | (pi01179 & w56176) | (~w12119 & w56176);
assign w12145 = w12119 & w56177;
assign w12146 = ~w12144 & ~w12145;
assign w12147 = (pi01180 & ~w12119) | (pi01180 & w56178) | (~w12119 & w56178);
assign w12148 = w12119 & w56179;
assign w12149 = ~w12147 & ~w12148;
assign w12150 = (pi01181 & ~w12119) | (pi01181 & w56180) | (~w12119 & w56180);
assign w12151 = w12119 & w56181;
assign w12152 = ~w12150 & ~w12151;
assign w12153 = (pi01182 & ~w12119) | (pi01182 & w56182) | (~w12119 & w56182);
assign w12154 = w12119 & w56183;
assign w12155 = ~w12153 & ~w12154;
assign w12156 = (pi01183 & ~w12119) | (pi01183 & w56184) | (~w12119 & w56184);
assign w12157 = w12119 & w56185;
assign w12158 = ~w12156 & ~w12157;
assign w12159 = (pi01184 & ~w12119) | (pi01184 & w56186) | (~w12119 & w56186);
assign w12160 = w12119 & w56187;
assign w12161 = ~w12159 & ~w12160;
assign w12162 = (pi01185 & ~w12119) | (pi01185 & w56188) | (~w12119 & w56188);
assign w12163 = w12119 & w56189;
assign w12164 = ~w12162 & ~w12163;
assign w12165 = (pi01186 & ~w12119) | (pi01186 & w56190) | (~w12119 & w56190);
assign w12166 = w12119 & w56191;
assign w12167 = ~w12165 & ~w12166;
assign w12168 = (pi01187 & ~w12119) | (pi01187 & w56192) | (~w12119 & w56192);
assign w12169 = w12119 & w56193;
assign w12170 = ~w12168 & ~w12169;
assign w12171 = (pi01188 & ~w12119) | (pi01188 & w56194) | (~w12119 & w56194);
assign w12172 = w12119 & w56195;
assign w12173 = ~w12171 & ~w12172;
assign w12174 = (pi01189 & ~w12119) | (pi01189 & w56196) | (~w12119 & w56196);
assign w12175 = w12119 & w56197;
assign w12176 = ~w12174 & ~w12175;
assign w12177 = (pi01190 & ~w12119) | (pi01190 & w56198) | (~w12119 & w56198);
assign w12178 = w12119 & w56199;
assign w12179 = ~w12177 & ~w12178;
assign w12180 = (pi01191 & ~w12119) | (pi01191 & w56200) | (~w12119 & w56200);
assign w12181 = w12119 & w56201;
assign w12182 = ~w12180 & ~w12181;
assign w12183 = (pi01192 & ~w12119) | (pi01192 & w56202) | (~w12119 & w56202);
assign w12184 = w12119 & w56203;
assign w12185 = ~w12183 & ~w12184;
assign w12186 = (pi01193 & ~w12119) | (pi01193 & w56204) | (~w12119 & w56204);
assign w12187 = w12119 & w56205;
assign w12188 = ~w12186 & ~w12187;
assign w12189 = (pi01194 & ~w12119) | (pi01194 & w56206) | (~w12119 & w56206);
assign w12190 = w12119 & w56207;
assign w12191 = ~w12189 & ~w12190;
assign w12192 = (pi01195 & ~w12119) | (pi01195 & w56208) | (~w12119 & w56208);
assign w12193 = w12119 & w56209;
assign w12194 = ~w12192 & ~w12193;
assign w12195 = (pi01197 & ~w12119) | (pi01197 & w56210) | (~w12119 & w56210);
assign w12196 = w12119 & w56211;
assign w12197 = ~w12195 & ~w12196;
assign w12198 = (pi01199 & ~w12119) | (pi01199 & w56212) | (~w12119 & w56212);
assign w12199 = w12119 & w56213;
assign w12200 = ~w12198 & ~w12199;
assign w12201 = (pi01198 & ~w12119) | (pi01198 & w56214) | (~w12119 & w56214);
assign w12202 = w12119 & w56215;
assign w12203 = ~w12201 & ~w12202;
assign w12204 = (pi01201 & ~w12119) | (pi01201 & w56216) | (~w12119 & w56216);
assign w12205 = w12119 & w56217;
assign w12206 = ~w12204 & ~w12205;
assign w12207 = (pi01200 & ~w12119) | (pi01200 & w56218) | (~w12119 & w56218);
assign w12208 = w12119 & w56219;
assign w12209 = ~w12207 & ~w12208;
assign w12210 = (pi01202 & ~w12119) | (pi01202 & w56220) | (~w12119 & w56220);
assign w12211 = w12119 & w56221;
assign w12212 = ~w12210 & ~w12211;
assign w12213 = (pi01196 & ~w12119) | (pi01196 & w56222) | (~w12119 & w56222);
assign w12214 = w12119 & w56223;
assign w12215 = ~w12213 & ~w12214;
assign w12216 = (~pi00643 & ~w10718) | (~pi00643 & w56224) | (~w10718 & w56224);
assign w12217 = pi00643 & ~w11474;
assign w12218 = ~w12216 & ~w12217;
assign w12219 = w11706 & w11709;
assign w12220 = w11800 & w11825;
assign w12221 = (pi00087 & w12220) | (pi00087 & w56225) | (w12220 & w56225);
assign w12222 = ~w12220 & w56226;
assign w12223 = ~w12221 & ~w12222;
assign w12224 = (pi00074 & w12220) | (pi00074 & w56227) | (w12220 & w56227);
assign w12225 = ~w12220 & w56228;
assign w12226 = ~w12224 & ~w12225;
assign w12227 = (pi00075 & w12220) | (pi00075 & w56229) | (w12220 & w56229);
assign w12228 = ~w12220 & w56230;
assign w12229 = ~w12227 & ~w12228;
assign w12230 = (pi00080 & w12220) | (pi00080 & w56231) | (w12220 & w56231);
assign w12231 = ~w12220 & w56232;
assign w12232 = ~w12230 & ~w12231;
assign w12233 = (pi00076 & w12220) | (pi00076 & w56233) | (w12220 & w56233);
assign w12234 = ~w12220 & w56234;
assign w12235 = ~w12233 & ~w12234;
assign w12236 = (pi00077 & w12220) | (pi00077 & w56235) | (w12220 & w56235);
assign w12237 = ~w12220 & w56236;
assign w12238 = ~w12236 & ~w12237;
assign w12239 = (pi00078 & w12220) | (pi00078 & w56237) | (w12220 & w56237);
assign w12240 = ~w12220 & w56238;
assign w12241 = ~w12239 & ~w12240;
assign w12242 = (pi00165 & w12220) | (pi00165 & w56239) | (w12220 & w56239);
assign w12243 = ~w12220 & w56240;
assign w12244 = ~w12242 & ~w12243;
assign w12245 = (pi00166 & w12220) | (pi00166 & w56241) | (w12220 & w56241);
assign w12246 = ~w12220 & w56242;
assign w12247 = ~w12245 & ~w12246;
assign w12248 = (pi00172 & w12220) | (pi00172 & w56243) | (w12220 & w56243);
assign w12249 = ~w12220 & w56244;
assign w12250 = ~w12248 & ~w12249;
assign w12251 = (pi00167 & w12220) | (pi00167 & w56245) | (w12220 & w56245);
assign w12252 = ~w12220 & w56246;
assign w12253 = ~w12251 & ~w12252;
assign w12254 = (pi00079 & w12220) | (pi00079 & w56247) | (w12220 & w56247);
assign w12255 = ~w12220 & w56248;
assign w12256 = ~w12254 & ~w12255;
assign w12257 = (pi00168 & w12220) | (pi00168 & w56249) | (w12220 & w56249);
assign w12258 = ~w12220 & w56250;
assign w12259 = ~w12257 & ~w12258;
assign w12260 = (pi00169 & w12220) | (pi00169 & w56251) | (w12220 & w56251);
assign w12261 = ~w12220 & w56252;
assign w12262 = ~w12260 & ~w12261;
assign w12263 = (pi00170 & w12220) | (pi00170 & w56253) | (w12220 & w56253);
assign w12264 = ~w12220 & w56254;
assign w12265 = ~w12263 & ~w12264;
assign w12266 = (pi00171 & w12220) | (pi00171 & w56255) | (w12220 & w56255);
assign w12267 = ~w12220 & w56256;
assign w12268 = ~w12266 & ~w12267;
assign w12269 = (pi00157 & w12220) | (pi00157 & w56257) | (w12220 & w56257);
assign w12270 = ~w12220 & w56258;
assign w12271 = ~w12269 & ~w12270;
assign w12272 = (pi00158 & w12220) | (pi00158 & w56259) | (w12220 & w56259);
assign w12273 = ~w12220 & w56260;
assign w12274 = ~w12272 & ~w12273;
assign w12275 = (pi00159 & w12220) | (pi00159 & w56261) | (w12220 & w56261);
assign w12276 = ~w12220 & w56262;
assign w12277 = ~w12275 & ~w12276;
assign w12278 = (pi00160 & w12220) | (pi00160 & w56263) | (w12220 & w56263);
assign w12279 = ~w12220 & w56264;
assign w12280 = ~w12278 & ~w12279;
assign w12281 = (pi00161 & w12220) | (pi00161 & w56265) | (w12220 & w56265);
assign w12282 = ~w12220 & w56266;
assign w12283 = ~w12281 & ~w12282;
assign w12284 = (pi00162 & w12220) | (pi00162 & w56267) | (w12220 & w56267);
assign w12285 = ~w12220 & w56268;
assign w12286 = ~w12284 & ~w12285;
assign w12287 = (pi00081 & w12220) | (pi00081 & w56269) | (w12220 & w56269);
assign w12288 = ~w12220 & w56270;
assign w12289 = ~w12287 & ~w12288;
assign w12290 = (pi00163 & w12220) | (pi00163 & w56271) | (w12220 & w56271);
assign w12291 = ~w12220 & w56272;
assign w12292 = ~w12290 & ~w12291;
assign w12293 = (pi00164 & w12220) | (pi00164 & w56273) | (w12220 & w56273);
assign w12294 = ~w12220 & w56274;
assign w12295 = ~w12293 & ~w12294;
assign w12296 = (pi00088 & w12220) | (pi00088 & w56275) | (w12220 & w56275);
assign w12297 = ~w12220 & w56276;
assign w12298 = ~w12296 & ~w12297;
assign w12299 = (pi00082 & w12220) | (pi00082 & w56277) | (w12220 & w56277);
assign w12300 = ~w12220 & w56278;
assign w12301 = ~w12299 & ~w12300;
assign w12302 = (pi00083 & w12220) | (pi00083 & w56279) | (w12220 & w56279);
assign w12303 = ~w12220 & w56280;
assign w12304 = ~w12302 & ~w12303;
assign w12305 = (pi00084 & w12220) | (pi00084 & w56281) | (w12220 & w56281);
assign w12306 = ~w12220 & w56282;
assign w12307 = ~w12305 & ~w12306;
assign w12308 = (pi00085 & w12220) | (pi00085 & w56283) | (w12220 & w56283);
assign w12309 = ~w12220 & w56284;
assign w12310 = ~w12308 & ~w12309;
assign w12311 = (pi00086 & w12220) | (pi00086 & w56285) | (w12220 & w56285);
assign w12312 = ~w12220 & w56286;
assign w12313 = ~w12311 & ~w12312;
assign w12314 = (pi00072 & w12220) | (pi00072 & w56287) | (w12220 & w56287);
assign w12315 = ~w12220 & w56288;
assign w12316 = ~w12314 & ~w12315;
assign w12317 = (pi00676 & ~w11828) | (pi00676 & w56289) | (~w11828 & w56289);
assign w12318 = w11828 & w56290;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = (pi00677 & ~w11828) | (pi00677 & w56291) | (~w11828 & w56291);
assign w12321 = w11828 & w56292;
assign w12322 = ~w12320 & ~w12321;
assign w12323 = (pi00678 & ~w11828) | (pi00678 & w56293) | (~w11828 & w56293);
assign w12324 = w11828 & w56064;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = (pi00679 & ~w11828) | (pi00679 & w56294) | (~w11828 & w56294);
assign w12327 = w11828 & w56295;
assign w12328 = ~w12326 & ~w12327;
assign w12329 = (pi00680 & ~w11828) | (pi00680 & w56296) | (~w11828 & w56296);
assign w12330 = w11828 & w56039;
assign w12331 = ~w12329 & ~w12330;
assign w12332 = (pi00681 & ~w11828) | (pi00681 & w56297) | (~w11828 & w56297);
assign w12333 = w11828 & w56067;
assign w12334 = ~w12332 & ~w12333;
assign w12335 = (pi00682 & ~w11828) | (pi00682 & w56298) | (~w11828 & w56298);
assign w12336 = w11828 & w55971;
assign w12337 = ~w12335 & ~w12336;
assign w12338 = (pi00683 & ~w11828) | (pi00683 & w56299) | (~w11828 & w56299);
assign w12339 = w11828 & w56300;
assign w12340 = ~w12338 & ~w12339;
assign w12341 = (pi00684 & ~w11828) | (pi00684 & w56301) | (~w11828 & w56301);
assign w12342 = w11828 & w56302;
assign w12343 = ~w12341 & ~w12342;
assign w12344 = (pi00685 & ~w11828) | (pi00685 & w56303) | (~w11828 & w56303);
assign w12345 = w11828 & w56069;
assign w12346 = ~w12344 & ~w12345;
assign w12347 = (pi00686 & ~w11828) | (pi00686 & w56304) | (~w11828 & w56304);
assign w12348 = w11828 & w56071;
assign w12349 = ~w12347 & ~w12348;
assign w12350 = (pi00687 & ~w11828) | (pi00687 & w56305) | (~w11828 & w56305);
assign w12351 = w11828 & w55944;
assign w12352 = ~w12350 & ~w12351;
assign w12353 = (pi00688 & ~w11828) | (pi00688 & w56306) | (~w11828 & w56306);
assign w12354 = w11828 & w55946;
assign w12355 = ~w12353 & ~w12354;
assign w12356 = (pi00689 & ~w11828) | (pi00689 & w56307) | (~w11828 & w56307);
assign w12357 = w11828 & w56047;
assign w12358 = ~w12356 & ~w12357;
assign w12359 = (pi00690 & ~w11828) | (pi00690 & w56308) | (~w11828 & w56308);
assign w12360 = w11828 & w55948;
assign w12361 = ~w12359 & ~w12360;
assign w12362 = (pi00691 & ~w11828) | (pi00691 & w56309) | (~w11828 & w56309);
assign w12363 = w11828 & w56310;
assign w12364 = ~w12362 & ~w12363;
assign w12365 = (pi00692 & ~w11828) | (pi00692 & w56311) | (~w11828 & w56311);
assign w12366 = w11828 & w56077;
assign w12367 = ~w12365 & ~w12366;
assign w12368 = (pi00693 & ~w11828) | (pi00693 & w56312) | (~w11828 & w56312);
assign w12369 = w11828 & w55952;
assign w12370 = ~w12368 & ~w12369;
assign w12371 = (pi00694 & ~w11828) | (pi00694 & w56313) | (~w11828 & w56313);
assign w12372 = w11828 & w55984;
assign w12373 = ~w12371 & ~w12372;
assign w12374 = (pi00695 & ~w11828) | (pi00695 & w56314) | (~w11828 & w56314);
assign w12375 = w11828 & w55958;
assign w12376 = ~w12374 & ~w12375;
assign w12377 = (pi00696 & ~w11828) | (pi00696 & w56315) | (~w11828 & w56315);
assign w12378 = w11828 & w56316;
assign w12379 = ~w12377 & ~w12378;
assign w12380 = (pi00697 & ~w11828) | (pi00697 & w56317) | (~w11828 & w56317);
assign w12381 = w11828 & w56081;
assign w12382 = ~w12380 & ~w12381;
assign w12383 = (pi00698 & ~w11828) | (pi00698 & w56318) | (~w11828 & w56318);
assign w12384 = w11828 & w56083;
assign w12385 = ~w12383 & ~w12384;
assign w12386 = (pi00699 & ~w11828) | (pi00699 & w56319) | (~w11828 & w56319);
assign w12387 = w11828 & w55950;
assign w12388 = ~w12386 & ~w12387;
assign w12389 = (pi00700 & ~w11828) | (pi00700 & w56320) | (~w11828 & w56320);
assign w12390 = w11828 & w56058;
assign w12391 = ~w12389 & ~w12390;
assign w12392 = (pi00701 & ~w11828) | (pi00701 & w56321) | (~w11828 & w56321);
assign w12393 = w11828 & w56106;
assign w12394 = ~w12392 & ~w12393;
assign w12395 = (pi00702 & ~w11828) | (pi00702 & w56322) | (~w11828 & w56322);
assign w12396 = w11828 & w56323;
assign w12397 = ~w12395 & ~w12396;
assign w12398 = (pi00703 & ~w11711) | (pi00703 & w56324) | (~w11711 & w56324);
assign w12399 = w11711 & w56096;
assign w12400 = ~w12398 & ~w12399;
assign w12401 = (pi00704 & ~w11711) | (pi00704 & w56325) | (~w11711 & w56325);
assign w12402 = w11711 & w56326;
assign w12403 = ~w12401 & ~w12402;
assign w12404 = (pi00705 & ~w11711) | (pi00705 & w56327) | (~w11711 & w56327);
assign w12405 = w11711 & w55994;
assign w12406 = ~w12404 & ~w12405;
assign w12407 = (pi00706 & ~w11711) | (pi00706 & w56328) | (~w11711 & w56328);
assign w12408 = w11711 & w56002;
assign w12409 = ~w12407 & ~w12408;
assign w12410 = (pi00707 & ~w11711) | (pi00707 & w56329) | (~w11711 & w56329);
assign w12411 = w11711 & w56110;
assign w12412 = ~w12410 & ~w12411;
assign w12413 = (pi00708 & ~w11711) | (pi00708 & w56330) | (~w11711 & w56330);
assign w12414 = w11711 & w56112;
assign w12415 = ~w12413 & ~w12414;
assign w12416 = (pi00709 & ~w11711) | (pi00709 & w56331) | (~w11711 & w56331);
assign w12417 = w11711 & w56118;
assign w12418 = ~w12416 & ~w12417;
assign w12419 = (pi00710 & ~w11711) | (pi00710 & w56332) | (~w11711 & w56332);
assign w12420 = w11711 & w56333;
assign w12421 = ~w12419 & ~w12420;
assign w12422 = (pi00711 & ~w11711) | (pi00711 & w56334) | (~w11711 & w56334);
assign w12423 = w11711 & w56335;
assign w12424 = ~w12422 & ~w12423;
assign w12425 = (pi00712 & ~w11711) | (pi00712 & w56336) | (~w11711 & w56336);
assign w12426 = w11711 & w56120;
assign w12427 = ~w12425 & ~w12426;
assign w12428 = (pi00713 & ~w11711) | (pi00713 & w56337) | (~w11711 & w56337);
assign w12429 = w11711 & w56122;
assign w12430 = ~w12428 & ~w12429;
assign w12431 = (pi00714 & ~w11711) | (pi00714 & w56338) | (~w11711 & w56338);
assign w12432 = w11711 & w56124;
assign w12433 = ~w12431 & ~w12432;
assign w12434 = (pi00715 & ~w11828) | (pi00715 & w56339) | (~w11828 & w56339);
assign w12435 = w11828 & w56096;
assign w12436 = ~w12434 & ~w12435;
assign w12437 = (pi00716 & ~w11828) | (pi00716 & w56340) | (~w11828 & w56340);
assign w12438 = w11828 & w56341;
assign w12439 = ~w12437 & ~w12438;
assign w12440 = (pi00717 & ~w11828) | (pi00717 & w56342) | (~w11828 & w56342);
assign w12441 = w11828 & w56098;
assign w12442 = ~w12440 & ~w12441;
assign w12443 = (pi00718 & ~w11828) | (pi00718 & w56343) | (~w11828 & w56343);
assign w12444 = w11828 & w56326;
assign w12445 = ~w12443 & ~w12444;
assign w12446 = (pi00719 & ~w11828) | (pi00719 & w56344) | (~w11828 & w56344);
assign w12447 = w11828 & w55996;
assign w12448 = ~w12446 & ~w12447;
assign w12449 = (pi00720 & ~w11828) | (pi00720 & w56345) | (~w11828 & w56345);
assign w12450 = w11828 & w56110;
assign w12451 = ~w12449 & ~w12450;
assign w12452 = (pi00721 & ~w11828) | (pi00721 & w56346) | (~w11828 & w56346);
assign w12453 = w11828 & w56114;
assign w12454 = ~w12452 & ~w12453;
assign w12455 = (pi00722 & ~w11828) | (pi00722 & w56347) | (~w11828 & w56347);
assign w12456 = w11828 & w56120;
assign w12457 = ~w12455 & ~w12456;
assign w12458 = (pi00723 & ~w11762) | (pi00723 & w56348) | (~w11762 & w56348);
assign w12459 = w11762 & w56128;
assign w12460 = ~w12458 & ~w12459;
assign w12461 = (pi00724 & ~w11762) | (pi00724 & w56349) | (~w11762 & w56349);
assign w12462 = w11762 & w56130;
assign w12463 = ~w12461 & ~w12462;
assign w12464 = (pi00725 & ~w11762) | (pi00725 & w56350) | (~w11762 & w56350);
assign w12465 = w11762 & w56351;
assign w12466 = ~w12464 & ~w12465;
assign w12467 = (pi00726 & ~w11762) | (pi00726 & w56352) | (~w11762 & w56352);
assign w12468 = w11762 & w56142;
assign w12469 = ~w12467 & ~w12468;
assign w12470 = (pi00727 & ~w11762) | (pi00727 & w56353) | (~w11762 & w56353);
assign w12471 = w11762 & w56011;
assign w12472 = ~w12470 & ~w12471;
assign w12473 = (pi00728 & ~w11762) | (pi00728 & w56354) | (~w11762 & w56354);
assign w12474 = w11762 & w56138;
assign w12475 = ~w12473 & ~w12474;
assign w12476 = (pi00729 & ~w11762) | (pi00729 & w56355) | (~w11762 & w56355);
assign w12477 = w11762 & w56013;
assign w12478 = ~w12476 & ~w12477;
assign w12479 = (pi00730 & ~w11762) | (pi00730 & w56356) | (~w11762 & w56356);
assign w12480 = w11762 & w56015;
assign w12481 = ~w12479 & ~w12480;
assign w12482 = (pi00731 & ~w11762) | (pi00731 & w56357) | (~w11762 & w56357);
assign w12483 = w11762 & w56140;
assign w12484 = ~w12482 & ~w12483;
assign w12485 = (pi00732 & ~w11762) | (pi00732 & w56358) | (~w11762 & w56358);
assign w12486 = w11762 & w56017;
assign w12487 = ~w12485 & ~w12486;
assign w12488 = (pi00733 & ~w11762) | (pi00733 & w56359) | (~w11762 & w56359);
assign w12489 = w11762 & w56144;
assign w12490 = ~w12488 & ~w12489;
assign w12491 = (pi00734 & ~w11762) | (pi00734 & w56360) | (~w11762 & w56360);
assign w12492 = w11762 & w56146;
assign w12493 = ~w12491 & ~w12492;
assign w12494 = (pi00735 & ~w11762) | (pi00735 & w56361) | (~w11762 & w56361);
assign w12495 = w11762 & w56362;
assign w12496 = ~w12494 & ~w12495;
assign w12497 = (pi00736 & ~w11800) | (pi00736 & w56363) | (~w11800 & w56363);
assign w12498 = w11800 & w56290;
assign w12499 = ~w12497 & ~w12498;
assign w12500 = (pi00737 & ~w11800) | (pi00737 & w56364) | (~w11800 & w56364);
assign w12501 = w11800 & w56295;
assign w12502 = ~w12500 & ~w12501;
assign w12503 = (pi00738 & ~w11762) | (pi00738 & w56365) | (~w11762 & w56365);
assign w12504 = w11762 & w56126;
assign w12505 = ~w12503 & ~w12504;
assign w12506 = (pi00739 & ~w11800) | (pi00739 & w56366) | (~w11800 & w56366);
assign w12507 = w11800 & w56067;
assign w12508 = ~w12506 & ~w12507;
assign w12509 = (pi00740 & ~w11800) | (pi00740 & w56367) | (~w11800 & w56367);
assign w12510 = w11800 & w55940;
assign w12511 = ~w12509 & ~w12510;
assign w12512 = (pi00741 & ~w11800) | (pi00741 & w56368) | (~w11800 & w56368);
assign w12513 = w11800 & w56369;
assign w12514 = ~w12512 & ~w12513;
assign w12515 = (pi00742 & ~w11800) | (pi00742 & w56370) | (~w11800 & w56370);
assign w12516 = w11800 & w56075;
assign w12517 = ~w12515 & ~w12516;
assign w12518 = (pi00743 & ~w11800) | (pi00743 & w56371) | (~w11800 & w56371);
assign w12519 = w11800 & w55982;
assign w12520 = ~w12518 & ~w12519;
assign w12521 = (pi00744 & ~w11800) | (pi00744 & w56372) | (~w11800 & w56372);
assign w12522 = w11800 & w55948;
assign w12523 = ~w12521 & ~w12522;
assign w12524 = (pi00745 & ~w11800) | (pi00745 & w56373) | (~w11800 & w56373);
assign w12525 = w11800 & w56310;
assign w12526 = ~w12524 & ~w12525;
assign w12527 = (pi00746 & ~w11800) | (pi00746 & w56374) | (~w11800 & w56374);
assign w12528 = w11800 & w56375;
assign w12529 = ~w12527 & ~w12528;
assign w12530 = (pi00747 & ~w11800) | (pi00747 & w56376) | (~w11800 & w56376);
assign w12531 = w11800 & w55984;
assign w12532 = ~w12530 & ~w12531;
assign w12533 = (pi00748 & ~w11800) | (pi00748 & w56377) | (~w11800 & w56377);
assign w12534 = w11800 & w55956;
assign w12535 = ~w12533 & ~w12534;
assign w12536 = (pi00749 & ~w11800) | (pi00749 & w56378) | (~w11800 & w56378);
assign w12537 = w11800 & w56316;
assign w12538 = ~w12536 & ~w12537;
assign w12539 = (pi00750 & ~w11800) | (pi00750 & w56379) | (~w11800 & w56379);
assign w12540 = w11800 & w55960;
assign w12541 = ~w12539 & ~w12540;
assign w12542 = (pi00751 & ~w11800) | (pi00751 & w56380) | (~w11800 & w56380);
assign w12543 = w11800 & w56081;
assign w12544 = ~w12542 & ~w12543;
assign w12545 = (pi00752 & ~w11800) | (pi00752 & w56381) | (~w11800 & w56381);
assign w12546 = w11800 & w56052;
assign w12547 = ~w12545 & ~w12546;
assign w12548 = (pi00753 & ~w11800) | (pi00753 & w56382) | (~w11800 & w56382);
assign w12549 = w11800 & w56054;
assign w12550 = ~w12548 & ~w12549;
assign w12551 = (pi00754 & ~w11800) | (pi00754 & w56383) | (~w11800 & w56383);
assign w12552 = w11800 & w55964;
assign w12553 = ~w12551 & ~w12552;
assign w12554 = (pi00755 & ~w11800) | (pi00755 & w56384) | (~w11800 & w56384);
assign w12555 = w11800 & w56385;
assign w12556 = ~w12554 & ~w12555;
assign w12557 = (pi00756 & ~w11800) | (pi00756 & w56386) | (~w11800 & w56386);
assign w12558 = w11800 & w56090;
assign w12559 = ~w12557 & ~w12558;
assign w12560 = (pi00757 & ~w11800) | (pi00757 & w56387) | (~w11800 & w56387);
assign w12561 = w11800 & w56060;
assign w12562 = ~w12560 & ~w12561;
assign w12563 = (pi00758 & ~w11800) | (pi00758 & w56388) | (~w11800 & w56388);
assign w12564 = w11800 & w56389;
assign w12565 = ~w12563 & ~w12564;
assign w12566 = (pi00759 & ~w11800) | (pi00759 & w56390) | (~w11800 & w56390);
assign w12567 = w11800 & w56391;
assign w12568 = ~w12566 & ~w12567;
assign w12569 = (pi00760 & ~w11800) | (pi00760 & w56392) | (~w11800 & w56392);
assign w12570 = w11800 & w56393;
assign w12571 = ~w12569 & ~w12570;
assign w12572 = (pi00761 & ~w11800) | (pi00761 & w56394) | (~w11800 & w56394);
assign w12573 = w11800 & w56058;
assign w12574 = ~w12572 & ~w12573;
assign w12575 = (pi00762 & ~w11800) | (pi00762 & w56395) | (~w11800 & w56395);
assign w12576 = w11800 & w55987;
assign w12577 = ~w12575 & ~w12576;
assign w12578 = (pi00763 & ~w11800) | (pi00763 & w56396) | (~w11800 & w56396);
assign w12579 = w11800 & w56062;
assign w12580 = ~w12578 & ~w12579;
assign w12581 = (pi00764 & ~w11800) | (pi00764 & w56397) | (~w11800 & w56397);
assign w12582 = w11800 & w56154;
assign w12583 = ~w12581 & ~w12582;
assign w12584 = (pi00765 & ~w11800) | (pi00765 & w56398) | (~w11800 & w56398);
assign w12585 = w11800 & w56323;
assign w12586 = ~w12584 & ~w12585;
assign w12587 = (pi00766 & ~w11800) | (pi00766 & w56399) | (~w11800 & w56399);
assign w12588 = w11800 & w55966;
assign w12589 = ~w12587 & ~w12588;
assign w12590 = (pi00767 & ~w11800) | (pi00767 & w56400) | (~w11800 & w56400);
assign w12591 = w11800 & w55950;
assign w12592 = ~w12590 & ~w12591;
assign w12593 = (pi00768 & ~w11762) | (pi00768 & w56401) | (~w11762 & w56401);
assign w12594 = w11762 & w55990;
assign w12595 = ~w12593 & ~w12594;
assign w12596 = (pi00769 & ~w11762) | (pi00769 & w56402) | (~w11762 & w56402);
assign w12597 = w11762 & w56341;
assign w12598 = ~w12596 & ~w12597;
assign w12599 = (pi00770 & ~w11762) | (pi00770 & w56403) | (~w11762 & w56403);
assign w12600 = w11762 & w56098;
assign w12601 = ~w12599 & ~w12600;
assign w12602 = (pi00771 & ~w11762) | (pi00771 & w56404) | (~w11762 & w56404);
assign w12603 = w11762 & w56100;
assign w12604 = ~w12602 & ~w12603;
assign w12605 = (pi00772 & ~w11762) | (pi00772 & w56405) | (~w11762 & w56405);
assign w12606 = w11762 & w56406;
assign w12607 = ~w12605 & ~w12606;
assign w12608 = (pi00773 & ~w11762) | (pi00773 & w56407) | (~w11762 & w56407);
assign w12609 = w11762 & w56104;
assign w12610 = ~w12608 & ~w12609;
assign w12611 = (pi00774 & ~w11762) | (pi00774 & w56408) | (~w11762 & w56408);
assign w12612 = w11762 & w55992;
assign w12613 = ~w12611 & ~w12612;
assign w12614 = (pi00775 & ~w11762) | (pi00775 & w56409) | (~w11762 & w56409);
assign w12615 = w11762 & w55994;
assign w12616 = ~w12614 & ~w12615;
assign w12617 = (pi00776 & ~w11762) | (pi00776 & w56410) | (~w11762 & w56410);
assign w12618 = w11762 & w55996;
assign w12619 = ~w12617 & ~w12618;
assign w12620 = (pi00777 & ~w11762) | (pi00777 & w56411) | (~w11762 & w56411);
assign w12621 = w11762 & w56000;
assign w12622 = ~w12620 & ~w12621;
assign w12623 = (pi00778 & ~w11762) | (pi00778 & w56412) | (~w11762 & w56412);
assign w12624 = w11762 & w56002;
assign w12625 = ~w12623 & ~w12624;
assign w12626 = (pi00779 & ~w11762) | (pi00779 & w56413) | (~w11762 & w56413);
assign w12627 = w11762 & w56110;
assign w12628 = ~w12626 & ~w12627;
assign w12629 = (pi00780 & ~w11762) | (pi00780 & w56414) | (~w11762 & w56414);
assign w12630 = w11762 & w56112;
assign w12631 = ~w12629 & ~w12630;
assign w12632 = (pi00781 & ~w11762) | (pi00781 & w56415) | (~w11762 & w56415);
assign w12633 = w11762 & w56118;
assign w12634 = ~w12632 & ~w12633;
assign w12635 = (pi00782 & ~w11762) | (pi00782 & w56416) | (~w11762 & w56416);
assign w12636 = w11762 & w56333;
assign w12637 = ~w12635 & ~w12636;
assign w12638 = (pi00783 & ~w11762) | (pi00783 & w56417) | (~w11762 & w56417);
assign w12639 = w11762 & w56418;
assign w12640 = ~w12638 & ~w12639;
assign w12641 = (pi00784 & ~w11762) | (pi00784 & w56419) | (~w11762 & w56419);
assign w12642 = w11762 & w56420;
assign w12643 = ~w12641 & ~w12642;
assign w12644 = (pi00785 & ~w11762) | (pi00785 & w56421) | (~w11762 & w56421);
assign w12645 = w11762 & w56004;
assign w12646 = ~w12644 & ~w12645;
assign w12647 = (pi00786 & ~w11762) | (pi00786 & w56422) | (~w11762 & w56422);
assign w12648 = w11762 & w56120;
assign w12649 = ~w12647 & ~w12648;
assign w12650 = (pi00787 & ~w11762) | (pi00787 & w56423) | (~w11762 & w56423);
assign w12651 = w11762 & w56122;
assign w12652 = ~w12650 & ~w12651;
assign w12653 = (pi00788 & ~w11762) | (pi00788 & w56424) | (~w11762 & w56424);
assign w12654 = w11762 & w56124;
assign w12655 = ~w12653 & ~w12654;
assign w12656 = (pi00789 & ~w11711) | (pi00789 & w56425) | (~w11711 & w56425);
assign w12657 = w11711 & w56007;
assign w12658 = ~w12656 & ~w12657;
assign w12659 = (pi00790 & ~w11711) | (pi00790 & w56426) | (~w11711 & w56426);
assign w12660 = w11711 & w56126;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = (pi00791 & ~w11711) | (pi00791 & w56427) | (~w11711 & w56427);
assign w12663 = w11711 & w56428;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = (pi00792 & ~w11711) | (pi00792 & w56429) | (~w11711 & w56429);
assign w12666 = w11711 & w56130;
assign w12667 = ~w12665 & ~w12666;
assign w12668 = (pi00793 & ~w11711) | (pi00793 & w56430) | (~w11711 & w56430);
assign w12669 = w11711 & w56351;
assign w12670 = ~w12668 & ~w12669;
assign w12671 = (pi00794 & ~w11711) | (pi00794 & w56431) | (~w11711 & w56431);
assign w12672 = w11711 & w56134;
assign w12673 = ~w12671 & ~w12672;
assign w12674 = (pi00795 & ~w11711) | (pi00795 & w56432) | (~w11711 & w56432);
assign w12675 = w11711 & w56009;
assign w12676 = ~w12674 & ~w12675;
assign w12677 = (pi00796 & ~w11711) | (pi00796 & w56433) | (~w11711 & w56433);
assign w12678 = w11711 & w56142;
assign w12679 = ~w12677 & ~w12678;
assign w12680 = (pi00797 & ~w11711) | (pi00797 & w56434) | (~w11711 & w56434);
assign w12681 = w11711 & w56138;
assign w12682 = ~w12680 & ~w12681;
assign w12683 = (pi00798 & ~w11711) | (pi00798 & w56435) | (~w11711 & w56435);
assign w12684 = w11711 & w56140;
assign w12685 = ~w12683 & ~w12684;
assign w12686 = (pi00799 & ~w11711) | (pi00799 & w56436) | (~w11711 & w56436);
assign w12687 = w11711 & w56017;
assign w12688 = ~w12686 & ~w12687;
assign w12689 = (pi00800 & ~w11762) | (pi00800 & w56437) | (~w11762 & w56437);
assign w12690 = w11762 & w56335;
assign w12691 = ~w12689 & ~w12690;
assign w12692 = (pi00801 & ~w11711) | (pi00801 & w56438) | (~w11711 & w56438);
assign w12693 = w11711 & w56148;
assign w12694 = ~w12692 & ~w12693;
assign w12695 = (pi00802 & ~w11711) | (pi00802 & w56439) | (~w11711 & w56439);
assign w12696 = w11711 & w56019;
assign w12697 = ~w12695 & ~w12696;
assign w12698 = (pi00803 & ~w11711) | (pi00803 & w56440) | (~w11711 & w56440);
assign w12699 = w11711 & w56441;
assign w12700 = ~w12698 & ~w12699;
assign w12701 = (pi00804 & ~w11711) | (pi00804 & w56442) | (~w11711 & w56442);
assign w12702 = w11711 & w56443;
assign w12703 = ~w12701 & ~w12702;
assign w12704 = (pi00805 & ~w11711) | (pi00805 & w56444) | (~w11711 & w56444);
assign w12705 = w11711 & w56445;
assign w12706 = ~w12704 & ~w12705;
assign w12707 = (pi00806 & ~w11711) | (pi00806 & w56446) | (~w11711 & w56446);
assign w12708 = w11711 & w56362;
assign w12709 = ~w12707 & ~w12708;
assign w12710 = (pi00807 & ~w11711) | (pi00807 & w56447) | (~w11711 & w56447);
assign w12711 = w11711 & w56144;
assign w12712 = ~w12710 & ~w12711;
assign w12713 = w11709 & w56448;
assign w12714 = (~pi00808 & ~w11709) | (~pi00808 & w56449) | (~w11709 & w56449);
assign w12715 = ~w11706 & ~w12713;
assign w12716 = ~w12714 & w12715;
assign w12717 = (~pi00809 & ~w11709) | (~pi00809 & w56450) | (~w11709 & w56450);
assign w12718 = (~w11706 & ~w11709) | (~w11706 & w56452) | (~w11709 & w56452);
assign w12719 = ~w12717 & w12718;
assign w12720 = pi00810 & w12718;
assign w12721 = ~w12104 & ~w12720;
assign w12722 = (pi00460 & w10682) | (pi00460 & w55830) | (w10682 & w55830);
assign w12723 = ~pi00816 & pi10020;
assign w12724 = ~w12722 & w12723;
assign w12725 = (~pi00811 & w12722) | (~pi00811 & w56453) | (w12722 & w56453);
assign w12726 = pi00811 & w826;
assign w12727 = ~w12725 & ~w12726;
assign w12728 = ~pi00274 & pi00815;
assign w12729 = pi09842 & ~w1435;
assign w12730 = ~pi09842 & w1435;
assign w12731 = ~pi00233 & pi09845;
assign w12732 = pi00233 & ~pi09845;
assign w12733 = ~w12731 & ~w12732;
assign w12734 = ~pi00240 & pi09840;
assign w12735 = pi00240 & ~pi09840;
assign w12736 = ~w12734 & ~w12735;
assign w12737 = ~pi09841 & ~w1432;
assign w12738 = pi09844 & ~w1429;
assign w12739 = ~pi09844 & w1429;
assign w12740 = ~w12738 & ~w12739;
assign w12741 = pi09841 & w1432;
assign w12742 = ~pi09843 & ~w1448;
assign w12743 = pi09843 & w1448;
assign w12744 = pi00249 & ~pi10587;
assign w12745 = ~w12733 & w12744;
assign w12746 = ~w12736 & w12745;
assign w12747 = ~w12737 & ~w12741;
assign w12748 = w12746 & w12747;
assign w12749 = ~w12729 & ~w12730;
assign w12750 = w12748 & w12749;
assign w12751 = ~w12742 & ~w12743;
assign w12752 = w12750 & w12751;
assign w12753 = ~w12740 & w12752;
assign w12754 = ~w12728 & ~w12753;
assign w12755 = ~pi00816 & ~pi00880;
assign w12756 = pi01481 & ~pi10020;
assign w12757 = ~w12755 & ~w12756;
assign w12758 = w11160 & w56454;
assign w12759 = pi00817 & ~w11160;
assign w12760 = ~w12758 & ~w12759;
assign w12761 = ~w11116 & w56455;
assign w12762 = pi10367 & w11116;
assign w12763 = ~w12761 & ~w12762;
assign w12764 = ~w11116 & w56456;
assign w12765 = pi10427 & w11116;
assign w12766 = ~w12764 & ~w12765;
assign w12767 = ~w11116 & w56457;
assign w12768 = pi10383 & w11116;
assign w12769 = ~w12767 & ~w12768;
assign w12770 = ~w11116 & w56458;
assign w12771 = pi10429 & w11116;
assign w12772 = ~w12770 & ~w12771;
assign w12773 = ~w11116 & w56459;
assign w12774 = pi10534 & w11116;
assign w12775 = ~w12773 & ~w12774;
assign w12776 = ~w11116 & w56460;
assign w12777 = pi10464 & w11116;
assign w12778 = ~w12776 & ~w12777;
assign w12779 = w671 & ~w2917;
assign w12780 = w671 & w2923;
assign w12781 = (~pi00826 & ~w11886) | (~pi00826 & w56461) | (~w11886 & w56461);
assign w12782 = ~w11890 & w11896;
assign w12783 = ~w12781 & w12782;
assign w12784 = ~w11885 & w56462;
assign w12785 = (pi00827 & w11885) | (pi00827 & w56463) | (w11885 & w56463);
assign w12786 = w11896 & ~w12784;
assign w12787 = ~w12785 & w12786;
assign w12788 = (~pi00828 & ~w11886) | (~pi00828 & w56464) | (~w11886 & w56464);
assign w12789 = ~w11889 & w11896;
assign w12790 = ~w12788 & w12789;
assign w12791 = (~pi00829 & ~w11886) | (~pi00829 & w56465) | (~w11886 & w56465);
assign w12792 = ~w11891 & w11896;
assign w12793 = ~w12791 & w12792;
assign w12794 = (~pi00830 & ~w11886) | (~pi00830 & w56466) | (~w11886 & w56466);
assign w12795 = ~w11892 & w11896;
assign w12796 = ~w12794 & w12795;
assign w12797 = ~pi00831 & ~w12785;
assign w12798 = pi00831 & w12785;
assign w12799 = w11896 & ~w12797;
assign w12800 = ~w12798 & w12799;
assign w12801 = (~pi00832 & ~w12785) | (~pi00832 & w56467) | (~w12785 & w56467);
assign w12802 = w12785 & w56468;
assign w12803 = w11896 & ~w12801;
assign w12804 = ~w12802 & w12803;
assign w12805 = (~pi00833 & ~w12785) | (~pi00833 & w56469) | (~w12785 & w56469);
assign w12806 = w12785 & w56470;
assign w12807 = w11896 & ~w12805;
assign w12808 = ~w12806 & w12807;
assign w12809 = (~pi00834 & ~w12785) | (~pi00834 & w56471) | (~w12785 & w56471);
assign w12810 = w12785 & w56472;
assign w12811 = w11896 & ~w12810;
assign w12812 = ~w12809 & w12811;
assign w12813 = (~pi00835 & ~w12785) | (~pi00835 & w56473) | (~w12785 & w56473);
assign w12814 = w12785 & w56474;
assign w12815 = w11896 & ~w12813;
assign w12816 = ~w12814 & w12815;
assign w12817 = (~pi00836 & ~w12785) | (~pi00836 & w56475) | (~w12785 & w56475);
assign w12818 = w12785 & w56476;
assign w12819 = w11896 & ~w12817;
assign w12820 = ~w12818 & w12819;
assign w12821 = (~pi00837 & ~w12785) | (~pi00837 & w56477) | (~w12785 & w56477);
assign w12822 = ~w11886 & w11896;
assign w12823 = ~w12821 & w12822;
assign w12824 = ~pi00838 & ~w11886;
assign w12825 = ~w11887 & w11896;
assign w12826 = ~w12824 & w12825;
assign w12827 = (~pi00839 & ~w11886) | (~pi00839 & w56478) | (~w11886 & w56478);
assign w12828 = ~w11888 & w11896;
assign w12829 = ~w12827 & w12828;
assign w12830 = (~pi00840 & ~w11886) | (~pi00840 & w56479) | (~w11886 & w56479);
assign w12831 = ~w11893 & w11896;
assign w12832 = ~w12830 & w12831;
assign w12833 = w25 & w56480;
assign w12834 = w2431 & ~w12833;
assign w12835 = pi01277 & ~w12834;
assign w12836 = (~pi00842 & ~w11485) | (~pi00842 & w56481) | (~w11485 & w56481);
assign w12837 = w11485 & w56482;
assign w12838 = ~pi10001 & ~w12836;
assign w12839 = ~w12837 & w12838;
assign w12840 = (~pi00843 & ~w11485) | (~pi00843 & w56483) | (~w11485 & w56483);
assign w12841 = w11485 & w56484;
assign w12842 = ~pi10357 & ~w12840;
assign w12843 = ~w12841 & w12842;
assign w12844 = pi00053 & pi00539;
assign w12845 = (~pi10577 & w12844) | (~pi10577 & w56485) | (w12844 & w56485);
assign w12846 = pi10381 & pi10552;
assign w12847 = pi02665 & w12846;
assign w12848 = (~pi00857 & ~w12846) | (~pi00857 & w56486) | (~w12846 & w56486);
assign w12849 = pi09930 & pi10002;
assign w12850 = pi09969 & ~w12849;
assign w12851 = ~pi00844 & ~pi00857;
assign w12852 = ~pi00868 & w12851;
assign w12853 = w12851 & w54829;
assign w12854 = w12853 & w56487;
assign w12855 = (pi02665 & ~w12853) | (pi02665 & w56488) | (~w12853 & w56488);
assign w12856 = (pi10418 & w12849) | (pi10418 & w56489) | (w12849 & w56489);
assign w12857 = (w12856 & w12855) | (w12856 & w56490) | (w12855 & w56490);
assign w12858 = w12857 & w56491;
assign w12859 = (~pi00844 & ~w12857) | (~pi00844 & w56492) | (~w12857 & w56492);
assign w12860 = w12857 & w56493;
assign w12861 = w12845 & ~w12859;
assign w12862 = ~w12860 & w12861;
assign w12863 = ~pi01170 & pi10518;
assign w12864 = pi00845 & pi10474;
assign w12865 = ~w12863 & w12864;
assign w12866 = ~pi10445 & ~w12865;
assign w12867 = ~pi02123 & pi02661;
assign w12868 = (pi00848 & ~w11370) | (pi00848 & w56494) | (~w11370 & w56494);
assign w12869 = w11370 & w56495;
assign w12870 = ~w12868 & ~w12869;
assign w12871 = pi00007 & pi00849;
assign w12872 = ~w686 & w12871;
assign w12873 = ~w523 & ~w12872;
assign w12874 = ~pi00483 & pi09868;
assign w12875 = ~pi10527 & w12874;
assign w12876 = (pi00132 & ~w12874) | (pi00132 & w56496) | (~w12874 & w56496);
assign w12877 = pi09519 & w1193;
assign w12878 = ~w12875 & ~w12877;
assign w12879 = ~w12876 & ~w12878;
assign w12880 = ~w12878 & w56497;
assign w12881 = w1193 & w56498;
assign w12882 = pi10374 & w12881;
assign w12883 = pi01304 & w12876;
assign w12884 = w12882 & w12883;
assign w12885 = pi01207 & w12884;
assign w12886 = w12884 & w56499;
assign w12887 = w12884 & w56500;
assign w12888 = w12884 & w56501;
assign w12889 = (pi00850 & w12878) | (pi00850 & w56502) | (w12878 & w56502);
assign w12890 = ~w12887 & w12889;
assign w12891 = ~w12880 & ~w12888;
assign w12892 = ~w12890 & w12891;
assign w12893 = ~pi00851 & pi00857;
assign w12894 = pi00852 & ~pi00858;
assign w12895 = pi00844 & ~pi00857;
assign w12896 = ~pi00868 & w12895;
assign w12897 = w12896 & w56503;
assign w12898 = pi02787 & w12897;
assign w12899 = ~pi00852 & ~pi00858;
assign w12900 = pi00867 & w12899;
assign w12901 = pi00868 & w12851;
assign w12902 = w12900 & w12901;
assign w12903 = pi00844 & pi00868;
assign w12904 = ~pi00857 & w12903;
assign w12905 = ~pi00867 & w12899;
assign w12906 = w12904 & w12905;
assign w12907 = pi09874 & w12906;
assign w12908 = w12901 & w12905;
assign w12909 = pi09981 & w12908;
assign w12910 = w12900 & w12904;
assign w12911 = pi02797 & w12910;
assign w12912 = w12853 & w56504;
assign w12913 = w12853 & w56505;
assign w12914 = w12853 & w56506;
assign w12915 = w12896 & w56507;
assign w12916 = pi01475 & w12915;
assign w12917 = (pi00852 & w12852) | (pi00852 & w56508) | (w12852 & w56508);
assign w12918 = ~w12850 & w12853;
assign w12919 = ~pi00867 & ~w12918;
assign w12920 = (~pi00858 & w12917) | (~pi00858 & w56509) | (w12917 & w56509);
assign w12921 = ~w12919 & w12920;
assign w12922 = (~pi00857 & ~w12902) | (~pi00857 & w56510) | (~w12902 & w56510);
assign w12923 = ~w12907 & ~w12909;
assign w12924 = ~w12898 & w12922;
assign w12925 = ~w12916 & w12924;
assign w12926 = w12923 & w56511;
assign w12927 = ~w12914 & w12926;
assign w12928 = ~w12921 & w12925;
assign w12929 = w12927 & w12928;
assign w12930 = ~w12893 & ~w12929;
assign w12931 = pi00852 & w12860;
assign w12932 = (w12845 & w12860) | (w12845 & w56512) | (w12860 & w56512);
assign w12933 = ~w12931 & w12932;
assign w12934 = w11485 & w56513;
assign w12935 = pi00853 & ~w12934;
assign w12936 = pi10349 & ~w12935;
assign w12937 = w11485 & w56514;
assign w12938 = pi00854 & ~w12937;
assign w12939 = pi10421 & ~w12938;
assign w12940 = w11485 & w56515;
assign w12941 = pi00855 & ~w12940;
assign w12942 = pi10348 & ~w12941;
assign w12943 = w11485 & w56516;
assign w12944 = pi00856 & ~w12943;
assign w12945 = pi10547 & pi10550;
assign w12946 = ~w12944 & ~w12945;
assign w12947 = (~pi00857 & ~w12857) | (~pi00857 & w56517) | (~w12857 & w56517);
assign w12948 = w12857 & w56518;
assign w12949 = w12845 & ~w12947;
assign w12950 = ~w12948 & w12949;
assign w12951 = w12860 & w56521;
assign w12952 = (w12860 & w56522) | (w12860 & w56523) | (w56522 & w56523);
assign w12953 = ~w12951 & w12952;
assign w12954 = (pi00859 & ~w11370) | (pi00859 & w56524) | (~w11370 & w56524);
assign w12955 = w11370 & w56525;
assign w12956 = ~w12954 & ~w12955;
assign w12957 = (pi00860 & ~w11370) | (pi00860 & w56526) | (~w11370 & w56526);
assign w12958 = w11370 & w56527;
assign w12959 = ~w12957 & ~w12958;
assign w12960 = (pi00861 & ~w11370) | (pi00861 & w56528) | (~w11370 & w56528);
assign w12961 = w11370 & w56529;
assign w12962 = ~w12960 & ~w12961;
assign w12963 = (pi00862 & ~w11370) | (pi00862 & w56530) | (~w11370 & w56530);
assign w12964 = w11370 & w56531;
assign w12965 = ~w12963 & ~w12964;
assign w12966 = (pi00863 & ~w11370) | (pi00863 & w56532) | (~w11370 & w56532);
assign w12967 = w11370 & w56533;
assign w12968 = ~w12966 & ~w12967;
assign w12969 = (pi00864 & ~w11370) | (pi00864 & w56534) | (~w11370 & w56534);
assign w12970 = w11370 & w56535;
assign w12971 = ~w12969 & ~w12970;
assign w12972 = (pi00865 & ~w11370) | (pi00865 & w56536) | (~w11370 & w56536);
assign w12973 = w11370 & w56537;
assign w12974 = ~w12972 & ~w12973;
assign w12975 = (pi00869 & w1480) | (pi00869 & w56538) | (w1480 & w56538);
assign w12976 = pi00866 & ~pi00869;
assign w12977 = ~w12975 & ~w12976;
assign w12978 = (~pi00867 & ~w12857) | (~pi00867 & w56539) | (~w12857 & w56539);
assign w12979 = w12845 & ~w12858;
assign w12980 = ~w12978 & w12979;
assign w12981 = (~pi00868 & ~w12860) | (~pi00868 & w54829) | (~w12860 & w54829);
assign w12982 = (w12845 & ~w12860) | (w12845 & w56540) | (~w12860 & w56540);
assign w12983 = ~w12981 & w12982;
assign w12984 = pi10442 & pi10517;
assign w12985 = ~pi00870 & ~pi01463;
assign w12986 = ~pi01262 & w12985;
assign w12987 = w12985 & w11129;
assign w12988 = ~pi01209 & w12987;
assign w12989 = (w12984 & ~w12987) | (w12984 & w56541) | (~w12987 & w56541);
assign w12990 = ~w1789 & w12989;
assign w12991 = w1789 & ~w12989;
assign w12992 = ~w12990 & ~w12991;
assign w12993 = ~pi10362 & ~pi10373;
assign w12994 = pi00870 & w12993;
assign w12995 = w12992 & w12994;
assign w12996 = ~w12992 & ~w12994;
assign w12997 = ~w12995 & ~w12996;
assign w12998 = pi00869 & w1491;
assign w12999 = ~pi00869 & pi00871;
assign w13000 = ~w12998 & ~w12999;
assign w13001 = (pi00872 & ~w11485) | (pi00872 & w56542) | (~w11485 & w56542);
assign w13002 = w11485 & w56543;
assign w13003 = ~w13001 & ~w13002;
assign w13004 = (pi00869 & w1467) | (pi00869 & w56544) | (w1467 & w56544);
assign w13005 = ~pi00869 & pi00873;
assign w13006 = ~w13004 & ~w13005;
assign w13007 = ~pi00874 & w67;
assign w13008 = pi00004 & w69;
assign w13009 = ~w13007 & ~w13008;
assign w13010 = pi00875 & w67;
assign w13011 = pi00026 & w69;
assign w13012 = ~w13010 & ~w13011;
assign w13013 = pi00876 & w67;
assign w13014 = pi00002 & w69;
assign w13015 = ~w13013 & ~w13014;
assign w13016 = pi00877 & w67;
assign w13017 = pi00205 & w69;
assign w13018 = ~w13016 & ~w13017;
assign w13019 = pi00878 & ~w11160;
assign w13020 = pi00035 & pi00036;
assign w13021 = w11160 & ~w13020;
assign w13022 = pi00036 & ~w693;
assign w13023 = ~pi10350 & w13021;
assign w13024 = ~w13022 & w13023;
assign w13025 = ~w13019 & ~w13024;
assign w13026 = w76 & ~w649;
assign w13027 = ~pi02810 & ~w11706;
assign w13028 = ~w11706 & w56545;
assign w13029 = pi01164 & pi01477;
assign w13030 = w13028 & w13029;
assign w13031 = w13028 & w56546;
assign w13032 = ~pi01164 & ~pi01477;
assign w13033 = w13028 & w13032;
assign w13034 = w13028 & w56547;
assign w13035 = ~pi01164 & pi01477;
assign w13036 = ~w11706 & w56548;
assign w13037 = w13036 & w56549;
assign w13038 = pi01164 & ~pi01477;
assign w13039 = ~w11706 & w56550;
assign w13040 = w13039 & w56551;
assign w13041 = w13028 & w56552;
assign w13042 = ~pi02810 & ~pi02812;
assign w13043 = w13032 & w13042;
assign w13044 = (~pi00666 & w13043) | (~pi00666 & w56553) | (w13043 & w56553);
assign w13045 = ~w11706 & w13042;
assign w13046 = w13038 & w13045;
assign w13047 = w13045 & w56554;
assign w13048 = w13028 & w13035;
assign w13049 = w13028 & w56555;
assign w13050 = w13035 & w13045;
assign w13051 = w13045 & w56556;
assign w13052 = w13036 & w56557;
assign w13053 = w13029 & w13045;
assign w13054 = w13045 & w56558;
assign w13055 = w13039 & w56559;
assign w13056 = w13039 & w56560;
assign w13057 = w13036 & w13038;
assign w13058 = w13036 & w56561;
assign w13059 = w13032 & w13039;
assign w13060 = w13039 & w56562;
assign w13061 = w13036 & w56563;
assign w13062 = ~w13044 & ~w13047;
assign w13063 = ~w13051 & ~w13054;
assign w13064 = w13062 & w13063;
assign w13065 = ~w13031 & ~w13034;
assign w13066 = ~w13037 & ~w13040;
assign w13067 = ~w13041 & ~w13049;
assign w13068 = ~w13052 & ~w13055;
assign w13069 = ~w13056 & ~w13058;
assign w13070 = ~w13060 & ~w13061;
assign w13071 = w13069 & w13070;
assign w13072 = w13067 & w13068;
assign w13073 = w13065 & w13066;
assign w13074 = w13064 & w13073;
assign w13075 = w13071 & w13072;
assign w13076 = w13074 & w13075;
assign w13077 = w13039 & w56564;
assign w13078 = w13036 & w56565;
assign w13079 = w13039 & w56566;
assign w13080 = w13039 & w56567;
assign w13081 = w13028 & w56568;
assign w13082 = (~pi00649 & w13043) | (~pi00649 & w56569) | (w13043 & w56569);
assign w13083 = w13045 & w56570;
assign w13084 = w13036 & w56571;
assign w13085 = w13045 & w56572;
assign w13086 = w13028 & w56573;
assign w13087 = w13045 & w56574;
assign w13088 = w13039 & w56575;
assign w13089 = w13028 & w56576;
assign w13090 = w13036 & w56577;
assign w13091 = w13028 & w56578;
assign w13092 = w13036 & w56579;
assign w13093 = ~w13082 & ~w13083;
assign w13094 = ~w13085 & ~w13087;
assign w13095 = w13093 & w13094;
assign w13096 = ~w13077 & ~w13078;
assign w13097 = ~w13079 & ~w13080;
assign w13098 = ~w13081 & ~w13084;
assign w13099 = ~w13086 & ~w13088;
assign w13100 = ~w13089 & ~w13090;
assign w13101 = ~w13091 & ~w13092;
assign w13102 = w13100 & w13101;
assign w13103 = w13098 & w13099;
assign w13104 = w13096 & w13097;
assign w13105 = w13095 & w13104;
assign w13106 = w13102 & w13103;
assign w13107 = w13105 & w13106;
assign w13108 = w13028 & w56580;
assign w13109 = w13036 & w56581;
assign w13110 = w13028 & w56582;
assign w13111 = w13036 & w56583;
assign w13112 = w13039 & w56584;
assign w13113 = (~pi00645 & w13043) | (~pi00645 & w56585) | (w13043 & w56585);
assign w13114 = w13045 & w56586;
assign w13115 = w13028 & w56587;
assign w13116 = w13045 & w56588;
assign w13117 = w13039 & w56589;
assign w13118 = w13045 & w56590;
assign w13119 = w13039 & w56591;
assign w13120 = w13036 & w56592;
assign w13121 = w13039 & w56593;
assign w13122 = w13028 & w56594;
assign w13123 = w13036 & w56595;
assign w13124 = ~w13113 & ~w13114;
assign w13125 = ~w13116 & ~w13118;
assign w13126 = w13124 & w13125;
assign w13127 = ~w13108 & ~w13109;
assign w13128 = ~w13110 & ~w13111;
assign w13129 = ~w13112 & ~w13115;
assign w13130 = ~w13117 & ~w13119;
assign w13131 = ~w13120 & ~w13121;
assign w13132 = ~w13122 & ~w13123;
assign w13133 = w13131 & w13132;
assign w13134 = w13129 & w13130;
assign w13135 = w13127 & w13128;
assign w13136 = w13126 & w13135;
assign w13137 = w13133 & w13134;
assign w13138 = w13136 & w13137;
assign w13139 = w13039 & w56596;
assign w13140 = w13036 & w56597;
assign w13141 = w13039 & w56598;
assign w13142 = w13028 & w56599;
assign w13143 = w13028 & w56600;
assign w13144 = (~pi00653 & w13043) | (~pi00653 & w56601) | (w13043 & w56601);
assign w13145 = w13045 & w56602;
assign w13146 = w13028 & w56603;
assign w13147 = w13045 & w56604;
assign w13148 = w13036 & w56605;
assign w13149 = w13045 & w56606;
assign w13150 = w13036 & w56607;
assign w13151 = w13028 & w56608;
assign w13152 = w13036 & w56609;
assign w13153 = w13039 & w56610;
assign w13154 = w13039 & w56611;
assign w13155 = ~w13144 & ~w13145;
assign w13156 = ~w13147 & ~w13149;
assign w13157 = w13155 & w13156;
assign w13158 = ~w13139 & ~w13140;
assign w13159 = ~w13141 & ~w13142;
assign w13160 = ~w13143 & ~w13146;
assign w13161 = ~w13148 & ~w13150;
assign w13162 = ~w13151 & ~w13152;
assign w13163 = ~w13153 & ~w13154;
assign w13164 = w13162 & w13163;
assign w13165 = w13160 & w13161;
assign w13166 = w13158 & w13159;
assign w13167 = w13157 & w13166;
assign w13168 = w13164 & w13165;
assign w13169 = w13167 & w13168;
assign w13170 = (pi00887 & ~w11711) | (pi00887 & w56612) | (~w11711 & w56612);
assign w13171 = w11711 & w56613;
assign w13172 = ~w13170 & ~w13171;
assign w13173 = (pi00888 & ~w11828) | (pi00888 & w56614) | (~w11828 & w56614);
assign w13174 = w11828 & w56351;
assign w13175 = ~w13173 & ~w13174;
assign w13176 = (pi00889 & ~w11828) | (pi00889 & w56615) | (~w11828 & w56615);
assign w13177 = w11828 & w56445;
assign w13178 = ~w13176 & ~w13177;
assign w13179 = (pi00890 & ~w11711) | (pi00890 & w56616) | (~w11711 & w56616);
assign w13180 = w11711 & w56011;
assign w13181 = ~w13179 & ~w13180;
assign w13182 = (pi00891 & ~w11711) | (pi00891 & w56617) | (~w11711 & w56617);
assign w13183 = w11711 & w56128;
assign w13184 = ~w13182 & ~w13183;
assign w13185 = (pi00892 & ~w11762) | (pi00892 & w56618) | (~w11762 & w56618);
assign w13186 = w11762 & w56096;
assign w13187 = ~w13185 & ~w13186;
assign w13188 = (pi00893 & ~w11800) | (pi00893 & w56619) | (~w11800 & w56619);
assign w13189 = w11800 & w56406;
assign w13190 = ~w13188 & ~w13189;
assign w13191 = (pi00894 & ~w11800) | (pi00894 & w56620) | (~w11800 & w56620);
assign w13192 = w11800 & w56420;
assign w13193 = ~w13191 & ~w13192;
assign w13194 = (pi00895 & ~w11800) | (pi00895 & w56621) | (~w11800 & w56621);
assign w13195 = w11800 & w56039;
assign w13196 = ~w13194 & ~w13195;
assign w13197 = (pi00896 & ~w11762) | (pi00896 & w56622) | (~w11762 & w56622);
assign w13198 = w11762 & w55952;
assign w13199 = ~w13197 & ~w13198;
assign w13200 = (pi00897 & ~w11762) | (pi00897 & w56623) | (~w11762 & w56623);
assign w13201 = w11762 & w56391;
assign w13202 = ~w13200 & ~w13201;
assign w13203 = (pi00898 & ~w11762) | (pi00898 & w56624) | (~w11762 & w56624);
assign w13204 = w11762 & w56385;
assign w13205 = ~w13203 & ~w13204;
assign w13206 = (pi00899 & ~w11762) | (pi00899 & w56625) | (~w11762 & w56625);
assign w13207 = w11762 & w56626;
assign w13208 = ~w13206 & ~w13207;
assign w13209 = (pi00900 & ~w11800) | (pi00900 & w56627) | (~w11800 & w56627);
assign w13210 = w11800 & w55958;
assign w13211 = ~w13209 & ~w13210;
assign w13212 = (pi00901 & ~w11762) | (pi00901 & w56628) | (~w11762 & w56628);
assign w13213 = w11762 & w56302;
assign w13214 = ~w13212 & ~w13213;
assign w13215 = (pi00902 & ~w11762) | (pi00902 & w56629) | (~w11762 & w56629);
assign w13216 = w11762 & w56295;
assign w13217 = ~w13215 & ~w13216;
assign w13218 = (pi00903 & ~w11800) | (pi00903 & w56630) | (~w11800 & w56630);
assign w13219 = w11800 & w56047;
assign w13220 = ~w13218 & ~w13219;
assign w13221 = (pi00904 & ~w11800) | (pi00904 & w56631) | (~w11800 & w56631);
assign w13222 = w11800 & w55979;
assign w13223 = ~w13221 & ~w13222;
assign w13224 = (pi00905 & ~w11800) | (pi00905 & w56632) | (~w11800 & w56632);
assign w13225 = w11800 & w56633;
assign w13226 = ~w13224 & ~w13225;
assign w13227 = (pi00906 & ~w11800) | (pi00906 & w56634) | (~w11800 & w56634);
assign w13228 = w11800 & w56292;
assign w13229 = ~w13227 & ~w13228;
assign w13230 = (pi00907 & ~w11762) | (pi00907 & w56635) | (~w11762 & w56635);
assign w13231 = w11762 & w56441;
assign w13232 = ~w13230 & ~w13231;
assign w13233 = (pi00908 & ~w11762) | (pi00908 & w56636) | (~w11762 & w56636);
assign w13234 = w11762 & w56613;
assign w13235 = ~w13233 & ~w13234;
assign w13236 = (pi00909 & ~w11762) | (pi00909 & w56637) | (~w11762 & w56637);
assign w13237 = w11762 & w56134;
assign w13238 = ~w13236 & ~w13237;
assign w13239 = (pi00910 & ~w11828) | (pi00910 & w56638) | (~w11828 & w56638);
assign w13240 = w11828 & w56335;
assign w13241 = ~w13239 & ~w13240;
assign w13242 = (pi00911 & ~w11711) | (pi00911 & w56639) | (~w11711 & w56639);
assign w13243 = w11711 & w56418;
assign w13244 = ~w13242 & ~w13243;
assign w13245 = (pi00912 & ~w11828) | (pi00912 & w56640) | (~w11828 & w56640);
assign w13246 = w11828 & w56333;
assign w13247 = ~w13245 & ~w13246;
assign w13248 = (pi00913 & ~w11828) | (pi00913 & w56641) | (~w11828 & w56641);
assign w13249 = w11828 & w56000;
assign w13250 = ~w13248 & ~w13249;
assign w13251 = (pi00914 & ~w11828) | (pi00914 & w56642) | (~w11828 & w56642);
assign w13252 = w11828 & w56100;
assign w13253 = ~w13251 & ~w13252;
assign w13254 = (pi00915 & ~w11711) | (pi00915 & w56643) | (~w11711 & w56643);
assign w13255 = w11711 & w56644;
assign w13256 = ~w13254 & ~w13255;
assign w13257 = (pi00916 & ~w11828) | (pi00916 & w56645) | (~w11828 & w56645);
assign w13258 = w11828 & w56054;
assign w13259 = ~w13257 & ~w13258;
assign w13260 = (pi00917 & ~w11711) | (pi00917 & w56646) | (~w11711 & w56646);
assign w13261 = w11711 & w56341;
assign w13262 = ~w13260 & ~w13261;
assign w13263 = (pi00918 & ~w11711) | (pi00918 & w56647) | (~w11711 & w56647);
assign w13264 = w11711 & w56098;
assign w13265 = ~w13263 & ~w13264;
assign w13266 = (pi00919 & ~w11828) | (pi00919 & w56648) | (~w11828 & w56648);
assign w13267 = w11828 & w56056;
assign w13268 = ~w13266 & ~w13267;
assign w13269 = (pi00920 & ~w11828) | (pi00920 & w56649) | (~w11828 & w56649);
assign w13270 = w11828 & w55956;
assign w13271 = ~w13269 & ~w13270;
assign w13272 = (pi00921 & ~w11711) | (pi00921 & w56650) | (~w11711 & w56650);
assign w13273 = w11711 & w56385;
assign w13274 = ~w13272 & ~w13273;
assign w13275 = (pi00922 & ~w11711) | (pi00922 & w56651) | (~w11711 & w56651);
assign w13276 = w11711 & w56391;
assign w13277 = ~w13275 & ~w13276;
assign w13278 = (pi00923 & ~w11711) | (pi00923 & w56652) | (~w11711 & w56652);
assign w13279 = w11711 & w55984;
assign w13280 = ~w13278 & ~w13279;
assign w13281 = (pi00924 & ~w11828) | (pi00924 & w56653) | (~w11828 & w56653);
assign w13282 = w11828 & w56633;
assign w13283 = ~w13281 & ~w13282;
assign w13284 = (pi00925 & ~w11828) | (pi00925 & w56654) | (~w11828 & w56654);
assign w13285 = w11828 & w55977;
assign w13286 = ~w13284 & ~w13285;
assign w13287 = (pi00926 & ~w11828) | (pi00926 & w56655) | (~w11828 & w56655);
assign w13288 = w11828 & w56375;
assign w13289 = ~w13287 & ~w13288;
assign w13290 = (pi00927 & ~w11711) | (pi00927 & w56656) | (~w11711 & w56656);
assign w13291 = w11711 & w55979;
assign w13292 = ~w13290 & ~w13291;
assign w13293 = (pi00928 & ~w11711) | (pi00928 & w56657) | (~w11711 & w56657);
assign w13294 = w11711 & w56633;
assign w13295 = ~w13293 & ~w13294;
assign w13296 = (~pi00929 & ~w518) | (~pi00929 & w56658) | (~w518 & w56658);
assign w13297 = ~w523 & ~w13296;
assign w13298 = w13028 & w56659;
assign w13299 = w13039 & w56660;
assign w13300 = w13039 & w56661;
assign w13301 = w13036 & w56662;
assign w13302 = w13036 & w56663;
assign w13303 = (~pi00668 & w13043) | (~pi00668 & w56664) | (w13043 & w56664);
assign w13304 = w13045 & w56665;
assign w13305 = w13028 & w56666;
assign w13306 = w13045 & w56667;
assign w13307 = w13039 & w56668;
assign w13308 = w13045 & w56669;
assign w13309 = w13036 & w56670;
assign w13310 = w13036 & w56671;
assign w13311 = w13028 & w56672;
assign w13312 = w13039 & w56673;
assign w13313 = w13028 & w56674;
assign w13314 = ~w13303 & ~w13304;
assign w13315 = ~w13306 & ~w13308;
assign w13316 = w13314 & w13315;
assign w13317 = ~w13298 & ~w13299;
assign w13318 = ~w13300 & ~w13301;
assign w13319 = ~w13302 & ~w13305;
assign w13320 = ~w13307 & ~w13309;
assign w13321 = ~w13310 & ~w13311;
assign w13322 = ~w13312 & ~w13313;
assign w13323 = w13321 & w13322;
assign w13324 = w13319 & w13320;
assign w13325 = w13317 & w13318;
assign w13326 = w13316 & w13325;
assign w13327 = w13323 & w13324;
assign w13328 = w13326 & w13327;
assign w13329 = w13036 & w56675;
assign w13330 = w13028 & w56676;
assign w13331 = w13039 & w56677;
assign w13332 = w13036 & w56678;
assign w13333 = w13036 & w56679;
assign w13334 = (~pi00667 & w13043) | (~pi00667 & w56680) | (w13043 & w56680);
assign w13335 = w13045 & w56681;
assign w13336 = w13028 & w56682;
assign w13337 = w13045 & w56683;
assign w13338 = w13039 & w56684;
assign w13339 = w13045 & w56685;
assign w13340 = w13039 & w56686;
assign w13341 = w13028 & w56687;
assign w13342 = w13028 & w56688;
assign w13343 = w13039 & w56689;
assign w13344 = w13036 & w56690;
assign w13345 = ~w13334 & ~w13335;
assign w13346 = ~w13337 & ~w13339;
assign w13347 = w13345 & w13346;
assign w13348 = ~w13329 & ~w13330;
assign w13349 = ~w13331 & ~w13332;
assign w13350 = ~w13333 & ~w13336;
assign w13351 = ~w13338 & ~w13340;
assign w13352 = ~w13341 & ~w13342;
assign w13353 = ~w13343 & ~w13344;
assign w13354 = w13352 & w13353;
assign w13355 = w13350 & w13351;
assign w13356 = w13348 & w13349;
assign w13357 = w13347 & w13356;
assign w13358 = w13354 & w13355;
assign w13359 = w13357 & w13358;
assign w13360 = w13036 & w56691;
assign w13361 = w13039 & w56692;
assign w13362 = w13039 & w56693;
assign w13363 = w13039 & w56694;
assign w13364 = w13028 & w56695;
assign w13365 = (~pi00665 & w13043) | (~pi00665 & w56696) | (w13043 & w56696);
assign w13366 = w13045 & w56697;
assign w13367 = w13028 & w56698;
assign w13368 = w13045 & w56699;
assign w13369 = w13036 & w56700;
assign w13370 = w13045 & w56701;
assign w13371 = w13036 & w56702;
assign w13372 = w13036 & w56703;
assign w13373 = w13028 & w56704;
assign w13374 = w13028 & w56705;
assign w13375 = w13039 & w56706;
assign w13376 = ~w13365 & ~w13366;
assign w13377 = ~w13368 & ~w13370;
assign w13378 = w13376 & w13377;
assign w13379 = ~w13360 & ~w13361;
assign w13380 = ~w13362 & ~w13363;
assign w13381 = ~w13364 & ~w13367;
assign w13382 = ~w13369 & ~w13371;
assign w13383 = ~w13372 & ~w13373;
assign w13384 = ~w13374 & ~w13375;
assign w13385 = w13383 & w13384;
assign w13386 = w13381 & w13382;
assign w13387 = w13379 & w13380;
assign w13388 = w13378 & w13387;
assign w13389 = w13385 & w13386;
assign w13390 = w13388 & w13389;
assign w13391 = w13028 & w56707;
assign w13392 = w13036 & w56708;
assign w13393 = w13028 & w56709;
assign w13394 = w13036 & w56710;
assign w13395 = w13036 & w56711;
assign w13396 = (~pi00664 & w13043) | (~pi00664 & w56712) | (w13043 & w56712);
assign w13397 = w13045 & w56713;
assign w13398 = w13039 & w56714;
assign w13399 = w13045 & w56715;
assign w13400 = w13036 & w56716;
assign w13401 = w13045 & w56717;
assign w13402 = w13028 & w56718;
assign w13403 = w13039 & w56719;
assign w13404 = w13028 & w56720;
assign w13405 = w13039 & w56721;
assign w13406 = w13039 & w56722;
assign w13407 = ~w13396 & ~w13397;
assign w13408 = ~w13399 & ~w13401;
assign w13409 = w13407 & w13408;
assign w13410 = ~w13391 & ~w13392;
assign w13411 = ~w13393 & ~w13394;
assign w13412 = ~w13395 & ~w13398;
assign w13413 = ~w13400 & ~w13402;
assign w13414 = ~w13403 & ~w13404;
assign w13415 = ~w13405 & ~w13406;
assign w13416 = w13414 & w13415;
assign w13417 = w13412 & w13413;
assign w13418 = w13410 & w13411;
assign w13419 = w13409 & w13418;
assign w13420 = w13416 & w13417;
assign w13421 = w13419 & w13420;
assign w13422 = w13028 & w56723;
assign w13423 = w13028 & w56724;
assign w13424 = w13039 & w56725;
assign w13425 = w13036 & w56726;
assign w13426 = w13039 & w56727;
assign w13427 = (~pi00663 & w13043) | (~pi00663 & w56728) | (w13043 & w56728);
assign w13428 = w13045 & w56729;
assign w13429 = w13028 & w56730;
assign w13430 = w13045 & w56731;
assign w13431 = w13036 & w56732;
assign w13432 = w13045 & w56733;
assign w13433 = w13036 & w56734;
assign w13434 = w13039 & w56735;
assign w13435 = w13036 & w56736;
assign w13436 = w13028 & w56737;
assign w13437 = w13039 & w56738;
assign w13438 = ~w13427 & ~w13428;
assign w13439 = ~w13430 & ~w13432;
assign w13440 = w13438 & w13439;
assign w13441 = ~w13422 & ~w13423;
assign w13442 = ~w13424 & ~w13425;
assign w13443 = ~w13426 & ~w13429;
assign w13444 = ~w13431 & ~w13433;
assign w13445 = ~w13434 & ~w13435;
assign w13446 = ~w13436 & ~w13437;
assign w13447 = w13445 & w13446;
assign w13448 = w13443 & w13444;
assign w13449 = w13441 & w13442;
assign w13450 = w13440 & w13449;
assign w13451 = w13447 & w13448;
assign w13452 = w13450 & w13451;
assign w13453 = w13039 & w56739;
assign w13454 = w13036 & w56740;
assign w13455 = w13036 & w56741;
assign w13456 = w13039 & w56742;
assign w13457 = w13036 & w56743;
assign w13458 = (~pi00662 & w13043) | (~pi00662 & w56744) | (w13043 & w56744);
assign w13459 = w13045 & w56745;
assign w13460 = w13028 & w56746;
assign w13461 = w13045 & w56747;
assign w13462 = w13036 & w56748;
assign w13463 = w13045 & w56749;
assign w13464 = w13028 & w56750;
assign w13465 = w13039 & w56751;
assign w13466 = w13028 & w56752;
assign w13467 = w13028 & w56753;
assign w13468 = w13039 & w56754;
assign w13469 = ~w13458 & ~w13459;
assign w13470 = ~w13461 & ~w13463;
assign w13471 = w13469 & w13470;
assign w13472 = ~w13453 & ~w13454;
assign w13473 = ~w13455 & ~w13456;
assign w13474 = ~w13457 & ~w13460;
assign w13475 = ~w13462 & ~w13464;
assign w13476 = ~w13465 & ~w13466;
assign w13477 = ~w13467 & ~w13468;
assign w13478 = w13476 & w13477;
assign w13479 = w13474 & w13475;
assign w13480 = w13472 & w13473;
assign w13481 = w13471 & w13480;
assign w13482 = w13478 & w13479;
assign w13483 = w13481 & w13482;
assign w13484 = w13039 & w56755;
assign w13485 = w13036 & w56756;
assign w13486 = w13036 & w56757;
assign w13487 = w13039 & w56758;
assign w13488 = w13028 & w56759;
assign w13489 = (~pi00661 & w13043) | (~pi00661 & w56760) | (w13043 & w56760);
assign w13490 = w13045 & w56761;
assign w13491 = w13039 & w56762;
assign w13492 = w13045 & w56763;
assign w13493 = w13036 & w56764;
assign w13494 = w13045 & w56765;
assign w13495 = w13028 & w56766;
assign w13496 = w13036 & w56767;
assign w13497 = w13028 & w56768;
assign w13498 = w13028 & w56769;
assign w13499 = w13039 & w56770;
assign w13500 = ~w13489 & ~w13490;
assign w13501 = ~w13492 & ~w13494;
assign w13502 = w13500 & w13501;
assign w13503 = ~w13484 & ~w13485;
assign w13504 = ~w13486 & ~w13487;
assign w13505 = ~w13488 & ~w13491;
assign w13506 = ~w13493 & ~w13495;
assign w13507 = ~w13496 & ~w13497;
assign w13508 = ~w13498 & ~w13499;
assign w13509 = w13507 & w13508;
assign w13510 = w13505 & w13506;
assign w13511 = w13503 & w13504;
assign w13512 = w13502 & w13511;
assign w13513 = w13509 & w13510;
assign w13514 = w13512 & w13513;
assign w13515 = w13028 & w56771;
assign w13516 = w13039 & w56772;
assign w13517 = w13036 & w56773;
assign w13518 = w13039 & w56774;
assign w13519 = w13039 & w56775;
assign w13520 = (~pi00659 & w13043) | (~pi00659 & w56776) | (w13043 & w56776);
assign w13521 = w13045 & w56777;
assign w13522 = w13028 & w56778;
assign w13523 = w13045 & w56779;
assign w13524 = w13036 & w56780;
assign w13525 = w13045 & w56781;
assign w13526 = w13036 & w56782;
assign w13527 = w13036 & w56783;
assign w13528 = w13028 & w56784;
assign w13529 = w13028 & w56785;
assign w13530 = w13039 & w56786;
assign w13531 = ~w13520 & ~w13521;
assign w13532 = ~w13523 & ~w13525;
assign w13533 = w13531 & w13532;
assign w13534 = ~w13515 & ~w13516;
assign w13535 = ~w13517 & ~w13518;
assign w13536 = ~w13519 & ~w13522;
assign w13537 = ~w13524 & ~w13526;
assign w13538 = ~w13527 & ~w13528;
assign w13539 = ~w13529 & ~w13530;
assign w13540 = w13538 & w13539;
assign w13541 = w13536 & w13537;
assign w13542 = w13534 & w13535;
assign w13543 = w13533 & w13542;
assign w13544 = w13540 & w13541;
assign w13545 = w13543 & w13544;
assign w13546 = w13036 & w56787;
assign w13547 = w13028 & w56788;
assign w13548 = w13039 & w56789;
assign w13549 = w13028 & w56790;
assign w13550 = w13028 & w56791;
assign w13551 = (~pi00660 & w13043) | (~pi00660 & w56792) | (w13043 & w56792);
assign w13552 = w13045 & w56793;
assign w13553 = w13039 & w56794;
assign w13554 = w13045 & w56795;
assign w13555 = w13028 & w56796;
assign w13556 = w13045 & w56797;
assign w13557 = w13039 & w56798;
assign w13558 = w13036 & w56799;
assign w13559 = w13036 & w56800;
assign w13560 = w13039 & w56801;
assign w13561 = w13036 & w56802;
assign w13562 = ~w13551 & ~w13552;
assign w13563 = ~w13554 & ~w13556;
assign w13564 = w13562 & w13563;
assign w13565 = ~w13546 & ~w13547;
assign w13566 = ~w13548 & ~w13549;
assign w13567 = ~w13550 & ~w13553;
assign w13568 = ~w13555 & ~w13557;
assign w13569 = ~w13558 & ~w13559;
assign w13570 = ~w13560 & ~w13561;
assign w13571 = w13569 & w13570;
assign w13572 = w13567 & w13568;
assign w13573 = w13565 & w13566;
assign w13574 = w13564 & w13573;
assign w13575 = w13571 & w13572;
assign w13576 = w13574 & w13575;
assign w13577 = w13039 & w56803;
assign w13578 = w13028 & w56804;
assign w13579 = w13039 & w56805;
assign w13580 = w13039 & w56806;
assign w13581 = w13036 & w56807;
assign w13582 = (~pi00658 & w13043) | (~pi00658 & w56808) | (w13043 & w56808);
assign w13583 = w13045 & w56809;
assign w13584 = w13036 & w56810;
assign w13585 = w13045 & w56811;
assign w13586 = w13036 & w56812;
assign w13587 = w13045 & w56813;
assign w13588 = w13028 & w56814;
assign w13589 = w13036 & w56815;
assign w13590 = w13039 & w56816;
assign w13591 = w13028 & w56817;
assign w13592 = w13028 & w56818;
assign w13593 = ~w13582 & ~w13583;
assign w13594 = ~w13585 & ~w13587;
assign w13595 = w13593 & w13594;
assign w13596 = ~w13577 & ~w13578;
assign w13597 = ~w13579 & ~w13580;
assign w13598 = ~w13581 & ~w13584;
assign w13599 = ~w13586 & ~w13588;
assign w13600 = ~w13589 & ~w13590;
assign w13601 = ~w13591 & ~w13592;
assign w13602 = w13600 & w13601;
assign w13603 = w13598 & w13599;
assign w13604 = w13596 & w13597;
assign w13605 = w13595 & w13604;
assign w13606 = w13602 & w13603;
assign w13607 = w13605 & w13606;
assign w13608 = w13036 & w56819;
assign w13609 = w13039 & w56820;
assign w13610 = w13028 & w56821;
assign w13611 = w13036 & w56822;
assign w13612 = w13028 & w56823;
assign w13613 = (~pi00657 & w13043) | (~pi00657 & w56824) | (w13043 & w56824);
assign w13614 = w13045 & w56825;
assign w13615 = w13039 & w56826;
assign w13616 = w13045 & w56827;
assign w13617 = w13028 & w56828;
assign w13618 = w13045 & w56829;
assign w13619 = w13039 & w56830;
assign w13620 = w13036 & w56831;
assign w13621 = w13028 & w56832;
assign w13622 = w13036 & w56833;
assign w13623 = w13039 & w56834;
assign w13624 = ~w13613 & ~w13614;
assign w13625 = ~w13616 & ~w13618;
assign w13626 = w13624 & w13625;
assign w13627 = ~w13608 & ~w13609;
assign w13628 = ~w13610 & ~w13611;
assign w13629 = ~w13612 & ~w13615;
assign w13630 = ~w13617 & ~w13619;
assign w13631 = ~w13620 & ~w13621;
assign w13632 = ~w13622 & ~w13623;
assign w13633 = w13631 & w13632;
assign w13634 = w13629 & w13630;
assign w13635 = w13627 & w13628;
assign w13636 = w13626 & w13635;
assign w13637 = w13633 & w13634;
assign w13638 = w13636 & w13637;
assign w13639 = w13036 & w56835;
assign w13640 = w13036 & w56836;
assign w13641 = w13039 & w56837;
assign w13642 = w13039 & w56838;
assign w13643 = w13036 & w56839;
assign w13644 = (~pi00656 & w13043) | (~pi00656 & w56840) | (w13043 & w56840);
assign w13645 = w13045 & w56841;
assign w13646 = w13039 & w56842;
assign w13647 = w13045 & w56843;
assign w13648 = w13028 & w56844;
assign w13649 = w13045 & w56845;
assign w13650 = w13028 & w56846;
assign w13651 = w13028 & w56847;
assign w13652 = w13036 & w56848;
assign w13653 = w13039 & w56849;
assign w13654 = w13028 & w56850;
assign w13655 = ~w13644 & ~w13645;
assign w13656 = ~w13647 & ~w13649;
assign w13657 = w13655 & w13656;
assign w13658 = ~w13639 & ~w13640;
assign w13659 = ~w13641 & ~w13642;
assign w13660 = ~w13643 & ~w13646;
assign w13661 = ~w13648 & ~w13650;
assign w13662 = ~w13651 & ~w13652;
assign w13663 = ~w13653 & ~w13654;
assign w13664 = w13662 & w13663;
assign w13665 = w13660 & w13661;
assign w13666 = w13658 & w13659;
assign w13667 = w13657 & w13666;
assign w13668 = w13664 & w13665;
assign w13669 = w13667 & w13668;
assign w13670 = w13036 & w56851;
assign w13671 = w13039 & w56852;
assign w13672 = w13028 & w56853;
assign w13673 = w13036 & w56854;
assign w13674 = w13036 & w56855;
assign w13675 = (~pi00654 & w13043) | (~pi00654 & w56856) | (w13043 & w56856);
assign w13676 = w13045 & w56857;
assign w13677 = w13028 & w56858;
assign w13678 = w13045 & w56859;
assign w13679 = w13039 & w56860;
assign w13680 = w13045 & w56861;
assign w13681 = w13028 & w56862;
assign w13682 = w13028 & w56863;
assign w13683 = w13036 & w56864;
assign w13684 = w13039 & w56865;
assign w13685 = w13039 & w56866;
assign w13686 = ~w13675 & ~w13676;
assign w13687 = ~w13678 & ~w13680;
assign w13688 = w13686 & w13687;
assign w13689 = ~w13670 & ~w13671;
assign w13690 = ~w13672 & ~w13673;
assign w13691 = ~w13674 & ~w13677;
assign w13692 = ~w13679 & ~w13681;
assign w13693 = ~w13682 & ~w13683;
assign w13694 = ~w13684 & ~w13685;
assign w13695 = w13693 & w13694;
assign w13696 = w13691 & w13692;
assign w13697 = w13689 & w13690;
assign w13698 = w13688 & w13697;
assign w13699 = w13695 & w13696;
assign w13700 = w13698 & w13699;
assign w13701 = w13036 & w56867;
assign w13702 = w13036 & w56868;
assign w13703 = w13028 & w56869;
assign w13704 = w13039 & w56870;
assign w13705 = w13036 & w56871;
assign w13706 = (~pi00652 & w13043) | (~pi00652 & w56872) | (w13043 & w56872);
assign w13707 = w13045 & w56873;
assign w13708 = w13028 & w56874;
assign w13709 = w13045 & w56875;
assign w13710 = w13028 & w56876;
assign w13711 = w13045 & w56877;
assign w13712 = w13028 & w56878;
assign w13713 = w13039 & w56879;
assign w13714 = w13039 & w56880;
assign w13715 = w13039 & w56881;
assign w13716 = w13036 & w56882;
assign w13717 = ~w13706 & ~w13707;
assign w13718 = ~w13709 & ~w13711;
assign w13719 = w13717 & w13718;
assign w13720 = ~w13701 & ~w13702;
assign w13721 = ~w13703 & ~w13704;
assign w13722 = ~w13705 & ~w13708;
assign w13723 = ~w13710 & ~w13712;
assign w13724 = ~w13713 & ~w13714;
assign w13725 = ~w13715 & ~w13716;
assign w13726 = w13724 & w13725;
assign w13727 = w13722 & w13723;
assign w13728 = w13720 & w13721;
assign w13729 = w13719 & w13728;
assign w13730 = w13726 & w13727;
assign w13731 = w13729 & w13730;
assign w13732 = w13036 & w56883;
assign w13733 = w13039 & w56884;
assign w13734 = w13036 & w56885;
assign w13735 = w13036 & w56886;
assign w13736 = w13028 & w56887;
assign w13737 = (~pi00651 & w13043) | (~pi00651 & w56888) | (w13043 & w56888);
assign w13738 = w13045 & w56889;
assign w13739 = w13028 & w56890;
assign w13740 = w13045 & w56891;
assign w13741 = w13036 & w56892;
assign w13742 = w13045 & w56893;
assign w13743 = w13028 & w56894;
assign w13744 = w13039 & w56895;
assign w13745 = w13039 & w56896;
assign w13746 = w13028 & w56897;
assign w13747 = w13039 & w56898;
assign w13748 = ~w13737 & ~w13738;
assign w13749 = ~w13740 & ~w13742;
assign w13750 = w13748 & w13749;
assign w13751 = ~w13732 & ~w13733;
assign w13752 = ~w13734 & ~w13735;
assign w13753 = ~w13736 & ~w13739;
assign w13754 = ~w13741 & ~w13743;
assign w13755 = ~w13744 & ~w13745;
assign w13756 = ~w13746 & ~w13747;
assign w13757 = w13755 & w13756;
assign w13758 = w13753 & w13754;
assign w13759 = w13751 & w13752;
assign w13760 = w13750 & w13759;
assign w13761 = w13757 & w13758;
assign w13762 = w13760 & w13761;
assign w13763 = w13036 & w56899;
assign w13764 = w13028 & w56900;
assign w13765 = w13036 & w56901;
assign w13766 = w13039 & w56902;
assign w13767 = w13039 & w56903;
assign w13768 = (~pi00650 & w13043) | (~pi00650 & w56904) | (w13043 & w56904);
assign w13769 = w13045 & w56905;
assign w13770 = w13036 & w56906;
assign w13771 = w13045 & w56907;
assign w13772 = w13039 & w56908;
assign w13773 = w13045 & w56909;
assign w13774 = w13028 & w56910;
assign w13775 = w13036 & w56911;
assign w13776 = w13039 & w56912;
assign w13777 = w13028 & w56913;
assign w13778 = w13028 & w56914;
assign w13779 = ~w13768 & ~w13769;
assign w13780 = ~w13771 & ~w13773;
assign w13781 = w13779 & w13780;
assign w13782 = ~w13763 & ~w13764;
assign w13783 = ~w13765 & ~w13766;
assign w13784 = ~w13767 & ~w13770;
assign w13785 = ~w13772 & ~w13774;
assign w13786 = ~w13775 & ~w13776;
assign w13787 = ~w13777 & ~w13778;
assign w13788 = w13786 & w13787;
assign w13789 = w13784 & w13785;
assign w13790 = w13782 & w13783;
assign w13791 = w13781 & w13790;
assign w13792 = w13788 & w13789;
assign w13793 = w13791 & w13792;
assign w13794 = w13036 & w56915;
assign w13795 = w13039 & w56916;
assign w13796 = w13039 & w56917;
assign w13797 = w13036 & w56918;
assign w13798 = w13028 & w56919;
assign w13799 = (~pi00648 & w13043) | (~pi00648 & w56920) | (w13043 & w56920);
assign w13800 = w13045 & w56921;
assign w13801 = w13036 & w56922;
assign w13802 = w13045 & w56923;
assign w13803 = w13028 & w56924;
assign w13804 = w13045 & w56925;
assign w13805 = w13028 & w56926;
assign w13806 = w13039 & w56927;
assign w13807 = w13039 & w56928;
assign w13808 = w13028 & w56929;
assign w13809 = w13036 & w56930;
assign w13810 = ~w13799 & ~w13800;
assign w13811 = ~w13802 & ~w13804;
assign w13812 = w13810 & w13811;
assign w13813 = ~w13794 & ~w13795;
assign w13814 = ~w13796 & ~w13797;
assign w13815 = ~w13798 & ~w13801;
assign w13816 = ~w13803 & ~w13805;
assign w13817 = ~w13806 & ~w13807;
assign w13818 = ~w13808 & ~w13809;
assign w13819 = w13817 & w13818;
assign w13820 = w13815 & w13816;
assign w13821 = w13813 & w13814;
assign w13822 = w13812 & w13821;
assign w13823 = w13819 & w13820;
assign w13824 = w13822 & w13823;
assign w13825 = w13028 & w56931;
assign w13826 = w13028 & w56932;
assign w13827 = w13039 & w56933;
assign w13828 = w13039 & w56934;
assign w13829 = w13036 & w56935;
assign w13830 = (~pi00647 & w13043) | (~pi00647 & w56936) | (w13043 & w56936);
assign w13831 = w13045 & w56937;
assign w13832 = w13028 & w56938;
assign w13833 = w13045 & w56939;
assign w13834 = w13039 & w56940;
assign w13835 = w13045 & w56941;
assign w13836 = w13039 & w56942;
assign w13837 = w13036 & w56943;
assign w13838 = w13036 & w56944;
assign w13839 = w13036 & w56945;
assign w13840 = w13028 & w56946;
assign w13841 = ~w13830 & ~w13831;
assign w13842 = ~w13833 & ~w13835;
assign w13843 = w13841 & w13842;
assign w13844 = ~w13825 & ~w13826;
assign w13845 = ~w13827 & ~w13828;
assign w13846 = ~w13829 & ~w13832;
assign w13847 = ~w13834 & ~w13836;
assign w13848 = ~w13837 & ~w13838;
assign w13849 = ~w13839 & ~w13840;
assign w13850 = w13848 & w13849;
assign w13851 = w13846 & w13847;
assign w13852 = w13844 & w13845;
assign w13853 = w13843 & w13852;
assign w13854 = w13850 & w13851;
assign w13855 = w13853 & w13854;
assign w13856 = w13036 & w56947;
assign w13857 = w13028 & w56948;
assign w13858 = w13039 & w56949;
assign w13859 = w13028 & w56950;
assign w13860 = w13039 & w56951;
assign w13861 = (~pi00646 & w13043) | (~pi00646 & w56952) | (w13043 & w56952);
assign w13862 = w13045 & w56953;
assign w13863 = w13036 & w56954;
assign w13864 = w13045 & w56955;
assign w13865 = w13036 & w56956;
assign w13866 = w13045 & w56957;
assign w13867 = w13028 & w56958;
assign w13868 = w13036 & w56959;
assign w13869 = w13039 & w56960;
assign w13870 = w13028 & w56961;
assign w13871 = w13039 & w56962;
assign w13872 = ~w13861 & ~w13862;
assign w13873 = ~w13864 & ~w13866;
assign w13874 = w13872 & w13873;
assign w13875 = ~w13856 & ~w13857;
assign w13876 = ~w13858 & ~w13859;
assign w13877 = ~w13860 & ~w13863;
assign w13878 = ~w13865 & ~w13867;
assign w13879 = ~w13868 & ~w13869;
assign w13880 = ~w13870 & ~w13871;
assign w13881 = w13879 & w13880;
assign w13882 = w13877 & w13878;
assign w13883 = w13875 & w13876;
assign w13884 = w13874 & w13883;
assign w13885 = w13881 & w13882;
assign w13886 = w13884 & w13885;
assign w13887 = w13036 & w56963;
assign w13888 = w13039 & w56964;
assign w13889 = w13028 & w56965;
assign w13890 = w13036 & w56966;
assign w13891 = w13028 & w56967;
assign w13892 = (~pi00674 & w13043) | (~pi00674 & w56968) | (w13043 & w56968);
assign w13893 = w13045 & w56969;
assign w13894 = w13039 & w56970;
assign w13895 = w13045 & w56971;
assign w13896 = w13028 & w56972;
assign w13897 = w13045 & w56973;
assign w13898 = w13036 & w56974;
assign w13899 = w13039 & w56975;
assign w13900 = w13039 & w56976;
assign w13901 = w13028 & w56977;
assign w13902 = w13036 & w56978;
assign w13903 = ~w13892 & ~w13893;
assign w13904 = ~w13895 & ~w13897;
assign w13905 = w13903 & w13904;
assign w13906 = ~w13887 & ~w13888;
assign w13907 = ~w13889 & ~w13890;
assign w13908 = ~w13891 & ~w13894;
assign w13909 = ~w13896 & ~w13898;
assign w13910 = ~w13899 & ~w13900;
assign w13911 = ~w13901 & ~w13902;
assign w13912 = w13910 & w13911;
assign w13913 = w13908 & w13909;
assign w13914 = w13906 & w13907;
assign w13915 = w13905 & w13914;
assign w13916 = w13912 & w13913;
assign w13917 = w13915 & w13916;
assign w13918 = w13028 & w56979;
assign w13919 = w13036 & w56980;
assign w13920 = w13036 & w56981;
assign w13921 = w13028 & w56982;
assign w13922 = w13036 & w56983;
assign w13923 = (~pi00673 & w13043) | (~pi00673 & w56984) | (w13043 & w56984);
assign w13924 = w13045 & w56985;
assign w13925 = w13039 & w56986;
assign w13926 = w13045 & w56987;
assign w13927 = w13039 & w56988;
assign w13928 = w13045 & w56989;
assign w13929 = w13028 & w56990;
assign w13930 = w13036 & w56991;
assign w13931 = w13028 & w56992;
assign w13932 = w13039 & w56993;
assign w13933 = w13039 & w56994;
assign w13934 = ~w13923 & ~w13924;
assign w13935 = ~w13926 & ~w13928;
assign w13936 = w13934 & w13935;
assign w13937 = ~w13918 & ~w13919;
assign w13938 = ~w13920 & ~w13921;
assign w13939 = ~w13922 & ~w13925;
assign w13940 = ~w13927 & ~w13929;
assign w13941 = ~w13930 & ~w13931;
assign w13942 = ~w13932 & ~w13933;
assign w13943 = w13941 & w13942;
assign w13944 = w13939 & w13940;
assign w13945 = w13937 & w13938;
assign w13946 = w13936 & w13945;
assign w13947 = w13943 & w13944;
assign w13948 = w13946 & w13947;
assign w13949 = w13039 & w56995;
assign w13950 = w13036 & w56996;
assign w13951 = w13028 & w56997;
assign w13952 = w13036 & w56998;
assign w13953 = w13039 & w56999;
assign w13954 = (~pi00672 & w13043) | (~pi00672 & w57000) | (w13043 & w57000);
assign w13955 = w13045 & w57001;
assign w13956 = w13039 & w57002;
assign w13957 = w13045 & w57003;
assign w13958 = w13028 & w57004;
assign w13959 = w13045 & w57005;
assign w13960 = w13028 & w57006;
assign w13961 = w13028 & w57007;
assign w13962 = w13039 & w57008;
assign w13963 = w13036 & w57009;
assign w13964 = w13036 & w57010;
assign w13965 = ~w13954 & ~w13955;
assign w13966 = ~w13957 & ~w13959;
assign w13967 = w13965 & w13966;
assign w13968 = ~w13949 & ~w13950;
assign w13969 = ~w13951 & ~w13952;
assign w13970 = ~w13953 & ~w13956;
assign w13971 = ~w13958 & ~w13960;
assign w13972 = ~w13961 & ~w13962;
assign w13973 = ~w13963 & ~w13964;
assign w13974 = w13972 & w13973;
assign w13975 = w13970 & w13971;
assign w13976 = w13968 & w13969;
assign w13977 = w13967 & w13976;
assign w13978 = w13974 & w13975;
assign w13979 = w13977 & w13978;
assign w13980 = w13028 & w57011;
assign w13981 = w13039 & w57012;
assign w13982 = w13028 & w57013;
assign w13983 = w13036 & w57014;
assign w13984 = w13036 & w57015;
assign w13985 = (~pi00671 & w13043) | (~pi00671 & w57016) | (w13043 & w57016);
assign w13986 = w13045 & w57017;
assign w13987 = w13039 & w57018;
assign w13988 = w13045 & w57019;
assign w13989 = w13039 & w57020;
assign w13990 = w13045 & w57021;
assign w13991 = w13028 & w57022;
assign w13992 = w13039 & w57023;
assign w13993 = w13036 & w57024;
assign w13994 = w13028 & w57025;
assign w13995 = w13036 & w57026;
assign w13996 = ~w13985 & ~w13986;
assign w13997 = ~w13988 & ~w13990;
assign w13998 = w13996 & w13997;
assign w13999 = ~w13980 & ~w13981;
assign w14000 = ~w13982 & ~w13983;
assign w14001 = ~w13984 & ~w13987;
assign w14002 = ~w13989 & ~w13991;
assign w14003 = ~w13992 & ~w13993;
assign w14004 = ~w13994 & ~w13995;
assign w14005 = w14003 & w14004;
assign w14006 = w14001 & w14002;
assign w14007 = w13999 & w14000;
assign w14008 = w13998 & w14007;
assign w14009 = w14005 & w14006;
assign w14010 = w14008 & w14009;
assign w14011 = w13028 & w57027;
assign w14012 = w13028 & w57028;
assign w14013 = w13039 & w57029;
assign w14014 = w13039 & w57030;
assign w14015 = w13036 & w57031;
assign w14016 = (~pi00669 & w13043) | (~pi00669 & w57032) | (w13043 & w57032);
assign w14017 = w13045 & w57033;
assign w14018 = w13028 & w57034;
assign w14019 = w13045 & w57035;
assign w14020 = w13039 & w57036;
assign w14021 = w13045 & w57037;
assign w14022 = w13039 & w57038;
assign w14023 = w13036 & w57039;
assign w14024 = w13036 & w57040;
assign w14025 = w13028 & w57041;
assign w14026 = w13036 & w57042;
assign w14027 = ~w14016 & ~w14017;
assign w14028 = ~w14019 & ~w14021;
assign w14029 = w14027 & w14028;
assign w14030 = ~w14011 & ~w14012;
assign w14031 = ~w14013 & ~w14014;
assign w14032 = ~w14015 & ~w14018;
assign w14033 = ~w14020 & ~w14022;
assign w14034 = ~w14023 & ~w14024;
assign w14035 = ~w14025 & ~w14026;
assign w14036 = w14034 & w14035;
assign w14037 = w14032 & w14033;
assign w14038 = w14030 & w14031;
assign w14039 = w14029 & w14038;
assign w14040 = w14036 & w14037;
assign w14041 = w14039 & w14040;
assign w14042 = w13028 & w57043;
assign w14043 = w13039 & w57044;
assign w14044 = w13036 & w57045;
assign w14045 = w13039 & w57046;
assign w14046 = w13036 & w57047;
assign w14047 = (~pi00670 & w13043) | (~pi00670 & w57048) | (w13043 & w57048);
assign w14048 = w13045 & w57049;
assign w14049 = w13039 & w57050;
assign w14050 = w13045 & w57051;
assign w14051 = w13028 & w57052;
assign w14052 = w13045 & w57053;
assign w14053 = w13028 & w57054;
assign w14054 = w13028 & w57055;
assign w14055 = w13036 & w57056;
assign w14056 = w13039 & w57057;
assign w14057 = w13036 & w57058;
assign w14058 = ~w14047 & ~w14048;
assign w14059 = ~w14050 & ~w14052;
assign w14060 = w14058 & w14059;
assign w14061 = ~w14042 & ~w14043;
assign w14062 = ~w14044 & ~w14045;
assign w14063 = ~w14046 & ~w14049;
assign w14064 = ~w14051 & ~w14053;
assign w14065 = ~w14054 & ~w14055;
assign w14066 = ~w14056 & ~w14057;
assign w14067 = w14065 & w14066;
assign w14068 = w14063 & w14064;
assign w14069 = w14061 & w14062;
assign w14070 = w14060 & w14069;
assign w14071 = w14067 & w14068;
assign w14072 = w14070 & w14071;
assign w14073 = w13039 & w57059;
assign w14074 = w13028 & w57060;
assign w14075 = w13036 & w57061;
assign w14076 = w13036 & w57062;
assign w14077 = w13028 & w57063;
assign w14078 = (~pi00655 & w13043) | (~pi00655 & w57064) | (w13043 & w57064);
assign w14079 = w13045 & w57065;
assign w14080 = w13039 & w57066;
assign w14081 = w13045 & w57067;
assign w14082 = w13039 & w57068;
assign w14083 = w13045 & w57069;
assign w14084 = w13028 & w57070;
assign w14085 = w13036 & w57071;
assign w14086 = w13039 & w57072;
assign w14087 = w13036 & w57073;
assign w14088 = w13028 & w57074;
assign w14089 = ~w14078 & ~w14079;
assign w14090 = ~w14081 & ~w14083;
assign w14091 = w14089 & w14090;
assign w14092 = ~w14073 & ~w14074;
assign w14093 = ~w14075 & ~w14076;
assign w14094 = ~w14077 & ~w14080;
assign w14095 = ~w14082 & ~w14084;
assign w14096 = ~w14085 & ~w14086;
assign w14097 = ~w14087 & ~w14088;
assign w14098 = w14096 & w14097;
assign w14099 = w14094 & w14095;
assign w14100 = w14092 & w14093;
assign w14101 = w14091 & w14100;
assign w14102 = w14098 & w14099;
assign w14103 = w14101 & w14102;
assign w14104 = w13036 & w57075;
assign w14105 = w13036 & w57076;
assign w14106 = w13028 & w57077;
assign w14107 = w13028 & w57078;
assign w14108 = w13039 & w57079;
assign w14109 = (~pi00644 & w13043) | (~pi00644 & w57080) | (w13043 & w57080);
assign w14110 = w13045 & w57081;
assign w14111 = w13039 & w57082;
assign w14112 = w13045 & w57083;
assign w14113 = w13028 & w57084;
assign w14114 = w13045 & w57085;
assign w14115 = w13036 & w57086;
assign w14116 = w13039 & w57087;
assign w14117 = w13036 & w57088;
assign w14118 = w13028 & w57089;
assign w14119 = w13039 & w57090;
assign w14120 = ~w14109 & ~w14110;
assign w14121 = ~w14112 & ~w14114;
assign w14122 = w14120 & w14121;
assign w14123 = ~w14104 & ~w14105;
assign w14124 = ~w14106 & ~w14107;
assign w14125 = ~w14108 & ~w14111;
assign w14126 = ~w14113 & ~w14115;
assign w14127 = ~w14116 & ~w14117;
assign w14128 = ~w14118 & ~w14119;
assign w14129 = w14127 & w14128;
assign w14130 = w14125 & w14126;
assign w14131 = w14123 & w14124;
assign w14132 = w14122 & w14131;
assign w14133 = w14129 & w14130;
assign w14134 = w14132 & w14133;
assign w14135 = pi02341 & ~pi02662;
assign w14136 = w11340 & w57091;
assign w14137 = w11340 & w57092;
assign w14138 = w11340 & w57093;
assign w14139 = ~pi00962 & ~pi01310;
assign w14140 = ~pi02657 & pi02660;
assign w14141 = w14139 & w14140;
assign w14142 = ~pi02659 & pi02663;
assign w14143 = ~w14135 & ~w14142;
assign w14144 = ~w14141 & w14143;
assign w14145 = pi01275 & pi01307;
assign w14146 = pi01308 & w14145;
assign w14147 = pi01213 & pi01305;
assign w14148 = w14146 & w14147;
assign w14149 = w14136 & w14148;
assign w14150 = w14136 & w57094;
assign w14151 = ~pi01306 & w14144;
assign w14152 = w14150 & w14151;
assign w14153 = (pi00957 & ~w14137) | (pi00957 & w57095) | (~w14137 & w57095);
assign w14154 = ~w14152 & w14153;
assign w14155 = ~w14138 & ~w14154;
assign w14156 = w13039 & w57096;
assign w14157 = ~pi01000 & w13030;
assign w14158 = w13036 & w57097;
assign w14159 = w13039 & w57098;
assign w14160 = ~pi00765 & w13059;
assign w14161 = (~pi00675 & w13043) | (~pi00675 & w57099) | (w13043 & w57099);
assign w14162 = ~pi01157 & w13050;
assign w14163 = w13036 & w57100;
assign w14164 = ~pi00534 & w13053;
assign w14165 = w13036 & w57101;
assign w14166 = ~pi01080 & w13046;
assign w14167 = w13028 & w57102;
assign w14168 = ~pi00548 & w13048;
assign w14169 = w13039 & w57103;
assign w14170 = ~pi00743 & w13033;
assign w14171 = w13036 & w57104;
assign w14172 = ~w14161 & ~w14162;
assign w14173 = ~w14164 & ~w14166;
assign w14174 = w14172 & w14173;
assign w14175 = ~w14156 & ~w14157;
assign w14176 = ~w14158 & ~w14159;
assign w14177 = ~w14160 & ~w14163;
assign w14178 = ~w14165 & ~w14167;
assign w14179 = ~w14168 & ~w14169;
assign w14180 = ~w14170 & ~w14171;
assign w14181 = w14179 & w14180;
assign w14182 = w14177 & w14178;
assign w14183 = w14175 & w14176;
assign w14184 = w14174 & w14183;
assign w14185 = w14181 & w14182;
assign w14186 = w14184 & w14185;
assign w14187 = ~pi09805 & ~pi09808;
assign w14188 = ~pi09860 & ~pi09861;
assign w14189 = ~pi09862 & ~pi09864;
assign w14190 = w14188 & w14189;
assign w14191 = (~pi09809 & ~w14190) | (~pi09809 & w57105) | (~w14190 & w57105);
assign w14192 = ~pi09860 & w14191;
assign w14193 = w14191 & w57106;
assign w14194 = w14191 & w57107;
assign w14195 = w14191 & w57108;
assign w14196 = ~pi09808 & w14195;
assign w14197 = (w14195 & w57110) | (w14195 & w57111) | (w57110 & w57111);
assign w14198 = w11340 & ~w14197;
assign w14199 = (pi00959 & ~w11337) | (pi00959 & w57112) | (~w11337 & w57112);
assign w14200 = ~w14198 & ~w14199;
assign w14201 = pi00869 & ~w1462;
assign w14202 = ~pi00869 & pi00960;
assign w14203 = ~w14201 & ~w14202;
assign w14204 = ~pi00024 & w503;
assign w14205 = w503 & w57113;
assign w14206 = (pi00025 & ~w403) | (pi00025 & w43935) | (~w403 & w43935);
assign w14207 = w504 & ~w14206;
assign w14208 = w724 & ~w14205;
assign w14209 = ~w14207 & w14208;
assign w14210 = (~pi00962 & ~w14137) | (~pi00962 & w57114) | (~w14137 & w57114);
assign w14211 = ~w14152 & ~w14210;
assign w14212 = (~pi00963 & ~w573) | (~pi00963 & w57115) | (~w573 & w57115);
assign w14213 = pi09964 & w291;
assign w14214 = ~w502 & ~w14213;
assign w14215 = ~w288 & ~w14214;
assign w14216 = ~w14212 & ~w14215;
assign w14217 = w507 & w14216;
assign w14218 = w11485 & w57116;
assign w14219 = ~pi00964 & ~w14218;
assign w14220 = pi10431 & ~w14219;
assign w14221 = w11485 & w57117;
assign w14222 = ~pi00965 & ~w14221;
assign w14223 = pi10371 & ~w14222;
assign w14224 = w11485 & w57118;
assign w14225 = ~pi00966 & ~w14224;
assign w14226 = pi10358 & ~w14225;
assign w14227 = pi02792 & w12897;
assign w14228 = pi09988 & w12908;
assign w14229 = w12853 & w57119;
assign w14230 = w12894 & w12901;
assign w14231 = w12853 & w57120;
assign w14232 = ~w14230 & ~w14231;
assign w14233 = ~pi00867 & ~w14232;
assign w14234 = pi09895 & w12906;
assign w14235 = pi02804 & w12910;
assign w14236 = w12896 & w12905;
assign w14237 = pi00857 & pi00967;
assign w14238 = pi01474 & w12915;
assign w14239 = pi00868 & ~pi09903;
assign w14240 = w12851 & ~w14239;
assign w14241 = w12900 & w14240;
assign w14242 = ~w14236 & ~w14237;
assign w14243 = ~w14241 & w14242;
assign w14244 = ~w14228 & ~w14234;
assign w14245 = ~w14235 & w14244;
assign w14246 = w14243 & w57121;
assign w14247 = ~w14229 & w14245;
assign w14248 = w14246 & w14247;
assign w14249 = ~w14233 & w14248;
assign w14250 = pi02123 & w11370;
assign w14251 = w11370 & w57122;
assign w14252 = (pi00968 & ~w11370) | (pi00968 & w57123) | (~w11370 & w57123);
assign w14253 = ~w14251 & ~w14252;
assign w14254 = w11370 & w57124;
assign w14255 = (pi00969 & ~w11370) | (pi00969 & w57125) | (~w11370 & w57125);
assign w14256 = ~w14254 & ~w14255;
assign w14257 = (~pi00970 & ~w25) | (~pi00970 & w57127) | (~w25 & w57127);
assign w14258 = ~pi00299 & ~pi09803;
assign w14259 = pi00487 & ~w14258;
assign w14260 = w25 & w57128;
assign w14261 = pi00063 & pi01251;
assign w14262 = ~pi00300 & ~w14261;
assign w14263 = w14260 & w14262;
assign w14264 = ~w14257 & ~w14263;
assign w14265 = (pi00971 & ~w11711) | (pi00971 & w57129) | (~w11711 & w57129);
assign w14266 = w11711 & w56290;
assign w14267 = ~w14265 & ~w14266;
assign w14268 = (pi00972 & ~w11711) | (pi00972 & w57130) | (~w11711 & w57130);
assign w14269 = w11711 & w56292;
assign w14270 = ~w14268 & ~w14269;
assign w14271 = (pi00973 & ~w11711) | (pi00973 & w57131) | (~w11711 & w57131);
assign w14272 = w11711 & w56064;
assign w14273 = ~w14271 & ~w14272;
assign w14274 = (pi00974 & ~w11711) | (pi00974 & w57132) | (~w11711 & w57132);
assign w14275 = w11711 & w56295;
assign w14276 = ~w14274 & ~w14275;
assign w14277 = (pi00975 & ~w11711) | (pi00975 & w57133) | (~w11711 & w57133);
assign w14278 = w11711 & w56375;
assign w14279 = ~w14277 & ~w14278;
assign w14280 = (pi00976 & ~w11711) | (pi00976 & w57134) | (~w11711 & w57134);
assign w14281 = w11711 & w56067;
assign w14282 = ~w14280 & ~w14281;
assign w14283 = (pi00977 & ~w11711) | (pi00977 & w57135) | (~w11711 & w57135);
assign w14284 = w11711 & w55971;
assign w14285 = ~w14283 & ~w14284;
assign w14286 = (pi00978 & ~w11711) | (pi00978 & w57136) | (~w11711 & w57136);
assign w14287 = w11711 & w56369;
assign w14288 = ~w14286 & ~w14287;
assign w14289 = (pi00979 & ~w11711) | (pi00979 & w57137) | (~w11711 & w57137);
assign w14290 = w11711 & w56300;
assign w14291 = ~w14289 & ~w14290;
assign w14292 = (pi00980 & ~w11711) | (pi00980 & w57138) | (~w11711 & w57138);
assign w14293 = w11711 & w55973;
assign w14294 = ~w14292 & ~w14293;
assign w14295 = (pi00981 & ~w11711) | (pi00981 & w57139) | (~w11711 & w57139);
assign w14296 = w11711 & w56302;
assign w14297 = ~w14295 & ~w14296;
assign w14298 = (pi00982 & ~w11711) | (pi00982 & w57140) | (~w11711 & w57140);
assign w14299 = w11711 & w56069;
assign w14300 = ~w14298 & ~w14299;
assign w14301 = (pi00983 & ~w11711) | (pi00983 & w57141) | (~w11711 & w57141);
assign w14302 = w11711 & w56071;
assign w14303 = ~w14301 & ~w14302;
assign w14304 = (pi00984 & ~w11711) | (pi00984 & w57142) | (~w11711 & w57142);
assign w14305 = w11711 & w57143;
assign w14306 = ~w14304 & ~w14305;
assign w14307 = (pi00985 & ~w11711) | (pi00985 & w57144) | (~w11711 & w57144);
assign w14308 = w11711 & w56626;
assign w14309 = ~w14307 & ~w14308;
assign w14310 = (pi00986 & ~w11711) | (pi00986 & w57145) | (~w11711 & w57145);
assign w14311 = w11711 & w56075;
assign w14312 = ~w14310 & ~w14311;
assign w14313 = (pi00987 & ~w11828) | (pi00987 & w57146) | (~w11828 & w57146);
assign w14314 = w11828 & w55936;
assign w14315 = ~w14313 & ~w14314;
assign w14316 = (pi00988 & ~w11828) | (pi00988 & w57147) | (~w11828 & w57147);
assign w14317 = w11828 & w55938;
assign w14318 = ~w14316 & ~w14317;
assign w14319 = (pi00989 & ~w11828) | (pi00989 & w57148) | (~w11828 & w57148);
assign w14320 = w11828 & w56041;
assign w14321 = ~w14319 & ~w14320;
assign w14322 = (pi00990 & ~w11828) | (pi00990 & w57149) | (~w11828 & w57149);
assign w14323 = w11828 & w56043;
assign w14324 = ~w14322 & ~w14323;
assign w14325 = (pi00991 & ~w11828) | (pi00991 & w57150) | (~w11828 & w57150);
assign w14326 = w11828 & w56369;
assign w14327 = ~w14325 & ~w14326;
assign w14328 = (pi00992 & ~w11828) | (pi00992 & w57151) | (~w11828 & w57151);
assign w14329 = w11828 & w55940;
assign w14330 = ~w14328 & ~w14329;
assign w14331 = (pi00993 & ~w11828) | (pi00993 & w57152) | (~w11828 & w57152);
assign w14332 = w11828 & w55973;
assign w14333 = ~w14331 & ~w14332;
assign w14334 = (pi00994 & ~w11828) | (pi00994 & w57153) | (~w11828 & w57153);
assign w14335 = w11828 & w55942;
assign w14336 = ~w14334 & ~w14335;
assign w14337 = (pi00995 & ~w11828) | (pi00995 & w57154) | (~w11828 & w57154);
assign w14338 = w11828 & w55975;
assign w14339 = ~w14337 & ~w14338;
assign w14340 = (pi00996 & ~w11828) | (pi00996 & w57155) | (~w11828 & w57155);
assign w14341 = w11828 & w55979;
assign w14342 = ~w14340 & ~w14341;
assign w14343 = (pi00997 & ~w11828) | (pi00997 & w57156) | (~w11828 & w57156);
assign w14344 = w11828 & w57143;
assign w14345 = ~w14343 & ~w14344;
assign w14346 = (pi00998 & ~w11828) | (pi00998 & w57157) | (~w11828 & w57157);
assign w14347 = w11828 & w56626;
assign w14348 = ~w14346 & ~w14347;
assign w14349 = (pi00999 & ~w11828) | (pi00999 & w57158) | (~w11828 & w57158);
assign w14350 = w11828 & w56075;
assign w14351 = ~w14349 & ~w14350;
assign w14352 = (pi01000 & ~w11828) | (pi01000 & w57159) | (~w11828 & w57159);
assign w14353 = w11828 & w55982;
assign w14354 = ~w14352 & ~w14353;
assign w14355 = (pi01001 & ~w11711) | (pi01001 & w57160) | (~w11711 & w57160);
assign w14356 = w11711 & w56077;
assign w14357 = ~w14355 & ~w14356;
assign w14358 = (pi01002 & ~w11711) | (pi01002 & w57161) | (~w11711 & w57161);
assign w14359 = w11711 & w56310;
assign w14360 = ~w14358 & ~w14359;
assign w14361 = (pi01003 & ~w11711) | (pi01003 & w57162) | (~w11711 & w57162);
assign w14362 = w11711 & w56316;
assign w14363 = ~w14361 & ~w14362;
assign w14364 = (pi01004 & ~w11711) | (pi01004 & w57163) | (~w11711 & w57163);
assign w14365 = w11711 & w56081;
assign w14366 = ~w14364 & ~w14365;
assign w14367 = (pi01005 & ~w11711) | (pi01005 & w57164) | (~w11711 & w57164);
assign w14368 = w11711 & w56083;
assign w14369 = ~w14367 & ~w14368;
assign w14370 = (pi01006 & ~w11711) | (pi01006 & w57165) | (~w11711 & w57165);
assign w14371 = w11711 & w56090;
assign w14372 = ~w14370 & ~w14371;
assign w14373 = (pi01007 & ~w11711) | (pi01007 & w57166) | (~w11711 & w57166);
assign w14374 = w11711 & w56389;
assign w14375 = ~w14373 & ~w14374;
assign w14376 = (pi01008 & ~w11711) | (pi01008 & w57167) | (~w11711 & w57167);
assign w14377 = w11711 & w56393;
assign w14378 = ~w14376 & ~w14377;
assign w14379 = (pi01009 & ~w11711) | (pi01009 & w57168) | (~w11711 & w57168);
assign w14380 = w11711 & w55987;
assign w14381 = ~w14379 & ~w14380;
assign w14382 = (pi01010 & ~w11711) | (pi01010 & w57169) | (~w11711 & w57169);
assign w14383 = w11711 & w56154;
assign w14384 = ~w14382 & ~w14383;
assign w14385 = (pi01011 & ~w11711) | (pi01011 & w57170) | (~w11711 & w57170);
assign w14386 = w11711 & w56092;
assign w14387 = ~w14385 & ~w14386;
assign w14388 = (pi01012 & ~w11711) | (pi01012 & w57171) | (~w11711 & w57171);
assign w14389 = w11711 & w56106;
assign w14390 = ~w14388 & ~w14389;
assign w14391 = (pi01013 & ~w11711) | (pi01013 & w57172) | (~w11711 & w57172);
assign w14392 = w11711 & w56323;
assign w14393 = ~w14391 & ~w14392;
assign w14394 = (pi01014 & ~w11828) | (pi01014 & w57173) | (~w11828 & w57173);
assign w14395 = w11828 & w56050;
assign w14396 = ~w14394 & ~w14395;
assign w14397 = (pi01015 & ~w11828) | (pi01015 & w57174) | (~w11828 & w57174);
assign w14398 = w11828 & w55954;
assign w14399 = ~w14397 & ~w14398;
assign w14400 = (pi01016 & ~w11828) | (pi01016 & w57175) | (~w11828 & w57175);
assign w14401 = w11828 & w55960;
assign w14402 = ~w14400 & ~w14401;
assign w14403 = (pi01017 & ~w11828) | (pi01017 & w57176) | (~w11828 & w57176);
assign w14404 = w11828 & w56052;
assign w14405 = ~w14403 & ~w14404;
assign w14406 = (pi01018 & ~w11828) | (pi01018 & w57177) | (~w11828 & w57177);
assign w14407 = w11828 & w55962;
assign w14408 = ~w14406 & ~w14407;
assign w14409 = (pi01019 & ~w11828) | (pi01019 & w57178) | (~w11828 & w57178);
assign w14410 = w11828 & w55964;
assign w14411 = ~w14409 & ~w14410;
assign w14412 = (pi01020 & ~w11828) | (pi01020 & w57179) | (~w11828 & w57179);
assign w14413 = w11828 & w56385;
assign w14414 = ~w14412 & ~w14413;
assign w14415 = (pi01021 & ~w11828) | (pi01021 & w57180) | (~w11828 & w57180);
assign w14416 = w11828 & w56090;
assign w14417 = ~w14415 & ~w14416;
assign w14418 = (pi01022 & ~w11828) | (pi01022 & w57181) | (~w11828 & w57181);
assign w14419 = w11828 & w56060;
assign w14420 = ~w14418 & ~w14419;
assign w14421 = (pi01023 & ~w11828) | (pi01023 & w57182) | (~w11828 & w57182);
assign w14422 = w11828 & w56389;
assign w14423 = ~w14421 & ~w14422;
assign w14424 = (pi01024 & ~w11828) | (pi01024 & w57183) | (~w11828 & w57183);
assign w14425 = w11828 & w56391;
assign w14426 = ~w14424 & ~w14425;
assign w14427 = (pi01025 & ~w11828) | (pi01025 & w57184) | (~w11828 & w57184);
assign w14428 = w11828 & w56393;
assign w14429 = ~w14427 & ~w14428;
assign w14430 = (pi01026 & ~w11828) | (pi01026 & w57185) | (~w11828 & w57185);
assign w14431 = w11828 & w56062;
assign w14432 = ~w14430 & ~w14431;
assign w14433 = (pi01027 & ~w11828) | (pi01027 & w57186) | (~w11828 & w57186);
assign w14434 = w11828 & w55987;
assign w14435 = ~w14433 & ~w14434;
assign w14436 = (pi01028 & ~w11828) | (pi01028 & w57187) | (~w11828 & w57187);
assign w14437 = w11828 & w56092;
assign w14438 = ~w14436 & ~w14437;
assign w14439 = (pi01029 & ~w11828) | (pi01029 & w57188) | (~w11828 & w57188);
assign w14440 = w11828 & w55966;
assign w14441 = ~w14439 & ~w14440;
assign w14442 = (pi01030 & ~w11711) | (pi01030 & w57189) | (~w11711 & w57189);
assign w14443 = w11711 & w56094;
assign w14444 = ~w14442 & ~w14443;
assign w14445 = (pi01031 & ~w11711) | (pi01031 & w57190) | (~w11711 & w57190);
assign w14446 = w11711 & w55990;
assign w14447 = ~w14445 & ~w14446;
assign w14448 = (pi01032 & ~w11711) | (pi01032 & w57191) | (~w11711 & w57191);
assign w14449 = w11711 & w57192;
assign w14450 = ~w14448 & ~w14449;
assign w14451 = (pi01033 & ~w11711) | (pi01033 & w57193) | (~w11711 & w57193);
assign w14452 = w11711 & w56100;
assign w14453 = ~w14451 & ~w14452;
assign w14454 = (pi01034 & ~w11711) | (pi01034 & w57194) | (~w11711 & w57194);
assign w14455 = w11711 & w56102;
assign w14456 = ~w14454 & ~w14455;
assign w14457 = (pi01035 & ~w11711) | (pi01035 & w57195) | (~w11711 & w57195);
assign w14458 = w11711 & w56406;
assign w14459 = ~w14457 & ~w14458;
assign w14460 = (pi01036 & ~w11711) | (pi01036 & w57196) | (~w11711 & w57196);
assign w14461 = w11711 & w56108;
assign w14462 = ~w14460 & ~w14461;
assign w14463 = (pi01037 & ~w11711) | (pi01037 & w57197) | (~w11711 & w57197);
assign w14464 = w11711 & w56104;
assign w14465 = ~w14463 & ~w14464;
assign w14466 = (pi01038 & ~w11711) | (pi01038 & w57198) | (~w11711 & w57198);
assign w14467 = w11711 & w55992;
assign w14468 = ~w14466 & ~w14467;
assign w14469 = (pi01039 & ~w11711) | (pi01039 & w57199) | (~w11711 & w57199);
assign w14470 = w11711 & w55996;
assign w14471 = ~w14469 & ~w14470;
assign w14472 = (pi01040 & ~w11711) | (pi01040 & w57200) | (~w11711 & w57200);
assign w14473 = w11711 & w55998;
assign w14474 = ~w14472 & ~w14473;
assign w14475 = (pi01041 & ~w11711) | (pi01041 & w57201) | (~w11711 & w57201);
assign w14476 = w11711 & w56000;
assign w14477 = ~w14475 & ~w14476;
assign w14478 = (pi01042 & ~w11711) | (pi01042 & w57202) | (~w11711 & w57202);
assign w14479 = w11711 & w56114;
assign w14480 = ~w14478 & ~w14479;
assign w14481 = (pi01043 & ~w11711) | (pi01043 & w57203) | (~w11711 & w57203);
assign w14482 = w11711 & w56420;
assign w14483 = ~w14481 & ~w14482;
assign w14484 = (pi01044 & ~w11711) | (pi01044 & w57204) | (~w11711 & w57204);
assign w14485 = w11711 & w56116;
assign w14486 = ~w14484 & ~w14485;
assign w14487 = (pi01045 & ~w11711) | (pi01045 & w57205) | (~w11711 & w57205);
assign w14488 = w11711 & w56004;
assign w14489 = ~w14487 & ~w14488;
assign w14490 = (pi01046 & ~w11828) | (pi01046 & w57206) | (~w11828 & w57206);
assign w14491 = w11828 & w56094;
assign w14492 = ~w14490 & ~w14491;
assign w14493 = (pi01047 & ~w11828) | (pi01047 & w57207) | (~w11828 & w57207);
assign w14494 = w11828 & w55990;
assign w14495 = ~w14493 & ~w14494;
assign w14496 = (pi01048 & ~w11828) | (pi01048 & w57208) | (~w11828 & w57208);
assign w14497 = w11828 & w57192;
assign w14498 = ~w14496 & ~w14497;
assign w14499 = (pi01049 & ~w11828) | (pi01049 & w57209) | (~w11828 & w57209);
assign w14500 = w11828 & w56102;
assign w14501 = ~w14499 & ~w14500;
assign w14502 = (pi01050 & ~w11828) | (pi01050 & w57210) | (~w11828 & w57210);
assign w14503 = w11828 & w56406;
assign w14504 = ~w14502 & ~w14503;
assign w14505 = (pi01051 & ~w11828) | (pi01051 & w57211) | (~w11828 & w57211);
assign w14506 = w11828 & w56104;
assign w14507 = ~w14505 & ~w14506;
assign w14508 = (pi01052 & ~w11828) | (pi01052 & w57212) | (~w11828 & w57212);
assign w14509 = w11828 & w56108;
assign w14510 = ~w14508 & ~w14509;
assign w14511 = (pi01053 & ~w11828) | (pi01053 & w57213) | (~w11828 & w57213);
assign w14512 = w11828 & w55992;
assign w14513 = ~w14511 & ~w14512;
assign w14514 = (pi01054 & ~w11828) | (pi01054 & w57214) | (~w11828 & w57214);
assign w14515 = w11828 & w55994;
assign w14516 = ~w14514 & ~w14515;
assign w14517 = (pi01055 & ~w11828) | (pi01055 & w57215) | (~w11828 & w57215);
assign w14518 = w11828 & w55998;
assign w14519 = ~w14517 & ~w14518;
assign w14520 = (pi01056 & ~w11828) | (pi01056 & w57216) | (~w11828 & w57216);
assign w14521 = w11828 & w56002;
assign w14522 = ~w14520 & ~w14521;
assign w14523 = (pi01057 & ~w11828) | (pi01057 & w57217) | (~w11828 & w57217);
assign w14524 = w11828 & w56112;
assign w14525 = ~w14523 & ~w14524;
assign w14526 = (pi01058 & ~w11828) | (pi01058 & w57218) | (~w11828 & w57218);
assign w14527 = w11828 & w56118;
assign w14528 = ~w14526 & ~w14527;
assign w14529 = (pi01059 & ~w11828) | (pi01059 & w57219) | (~w11828 & w57219);
assign w14530 = w11828 & w56418;
assign w14531 = ~w14529 & ~w14530;
assign w14532 = (pi01060 & ~w11828) | (pi01060 & w57220) | (~w11828 & w57220);
assign w14533 = w11828 & w56116;
assign w14534 = ~w14532 & ~w14533;
assign w14535 = (pi01061 & ~w11828) | (pi01061 & w57221) | (~w11828 & w57221);
assign w14536 = w11828 & w56420;
assign w14537 = ~w14535 & ~w14536;
assign w14538 = (pi01062 & ~w11828) | (pi01062 & w57222) | (~w11828 & w57222);
assign w14539 = w11828 & w56004;
assign w14540 = ~w14538 & ~w14539;
assign w14541 = (pi01063 & ~w11828) | (pi01063 & w57223) | (~w11828 & w57223);
assign w14542 = w11828 & w56122;
assign w14543 = ~w14541 & ~w14542;
assign w14544 = (pi01064 & ~w11828) | (pi01064 & w57224) | (~w11828 & w57224);
assign w14545 = w11828 & w56644;
assign w14546 = ~w14544 & ~w14545;
assign w14547 = (pi01065 & ~w11828) | (pi01065 & w57225) | (~w11828 & w57225);
assign w14548 = w11828 & w56124;
assign w14549 = ~w14547 & ~w14548;
assign w14550 = (pi01066 & ~w11762) | (pi01066 & w57226) | (~w11762 & w57226);
assign w14551 = w11762 & w56007;
assign w14552 = ~w14550 & ~w14551;
assign w14553 = (pi01067 & ~w11762) | (pi01067 & w57227) | (~w11762 & w57227);
assign w14554 = w11762 & w56428;
assign w14555 = ~w14553 & ~w14554;
assign w14556 = (pi01068 & ~w11762) | (pi01068 & w57228) | (~w11762 & w57228);
assign w14557 = w11762 & w57229;
assign w14558 = ~w14556 & ~w14557;
assign w14559 = (pi01069 & ~w11762) | (pi01069 & w57230) | (~w11762 & w57230);
assign w14560 = w11762 & w56136;
assign w14561 = ~w14559 & ~w14560;
assign w14562 = (pi01070 & ~w11762) | (pi01070 & w57231) | (~w11762 & w57231);
assign w14563 = w11762 & w56132;
assign w14564 = ~w14562 & ~w14563;
assign w14565 = (pi01071 & ~w11762) | (pi01071 & w57232) | (~w11762 & w57232);
assign w14566 = w11762 & w56009;
assign w14567 = ~w14565 & ~w14566;
assign w14568 = (pi01072 & ~w11762) | (pi01072 & w57233) | (~w11762 & w57233);
assign w14569 = w11762 & w56148;
assign w14570 = ~w14568 & ~w14569;
assign w14571 = (pi01073 & ~w11762) | (pi01073 & w57234) | (~w11762 & w57234);
assign w14572 = w11762 & w56019;
assign w14573 = ~w14571 & ~w14572;
assign w14574 = (pi01074 & ~w11762) | (pi01074 & w57235) | (~w11762 & w57235);
assign w14575 = w11762 & w56150;
assign w14576 = ~w14574 & ~w14575;
assign w14577 = (pi01075 & ~w11762) | (pi01075 & w57236) | (~w11762 & w57236);
assign w14578 = w11762 & w56443;
assign w14579 = ~w14577 & ~w14578;
assign w14580 = (pi01076 & ~w11762) | (pi01076 & w57237) | (~w11762 & w57237);
assign w14581 = w11762 & w56152;
assign w14582 = ~w14580 & ~w14581;
assign w14583 = (pi01077 & ~w11762) | (pi01077 & w57238) | (~w11762 & w57238);
assign w14584 = w11762 & w56021;
assign w14585 = ~w14583 & ~w14584;
assign w14586 = (pi01078 & ~w11762) | (pi01078 & w57239) | (~w11762 & w57239);
assign w14587 = w11762 & w56445;
assign w14588 = ~w14586 & ~w14587;
assign w14589 = (pi01079 & ~w11762) | (pi01079 & w57240) | (~w11762 & w57240);
assign w14590 = w11762 & w56023;
assign w14591 = ~w14589 & ~w14590;
assign w14592 = (pi01080 & ~w11762) | (pi01080 & w57241) | (~w11762 & w57241);
assign w14593 = w11762 & w56025;
assign w14594 = ~w14592 & ~w14593;
assign w14595 = (pi01081 & ~w11800) | (pi01081 & w57242) | (~w11800 & w57242);
assign w14596 = w11800 & w55936;
assign w14597 = ~w14595 & ~w14596;
assign w14598 = (pi01082 & ~w11800) | (pi01082 & w57243) | (~w11800 & w57243);
assign w14599 = w11800 & w55938;
assign w14600 = ~w14598 & ~w14599;
assign w14601 = (pi01083 & ~w11800) | (pi01083 & w57244) | (~w11800 & w57244);
assign w14602 = w11800 & w56064;
assign w14603 = ~w14601 & ~w14602;
assign w14604 = (pi01084 & ~w11800) | (pi01084 & w57245) | (~w11800 & w57245);
assign w14605 = w11800 & w56041;
assign w14606 = ~w14604 & ~w14605;
assign w14607 = (pi01085 & ~w11800) | (pi01085 & w57246) | (~w11800 & w57246);
assign w14608 = w11800 & w55971;
assign w14609 = ~w14607 & ~w14608;
assign w14610 = (pi01086 & ~w11800) | (pi01086 & w57247) | (~w11800 & w57247);
assign w14611 = w11800 & w56043;
assign w14612 = ~w14610 & ~w14611;
assign w14613 = (pi01087 & ~w11800) | (pi01087 & w57248) | (~w11800 & w57248);
assign w14614 = w11800 & w56300;
assign w14615 = ~w14613 & ~w14614;
assign w14616 = (pi01088 & ~w11800) | (pi01088 & w57249) | (~w11800 & w57249);
assign w14617 = w11800 & w55973;
assign w14618 = ~w14616 & ~w14617;
assign w14619 = (pi01089 & ~w11800) | (pi01089 & w57250) | (~w11800 & w57250);
assign w14620 = w11800 & w56302;
assign w14621 = ~w14619 & ~w14620;
assign w14622 = (pi01090 & ~w11800) | (pi01090 & w57251) | (~w11800 & w57251);
assign w14623 = w11800 & w56069;
assign w14624 = ~w14622 & ~w14623;
assign w14625 = (pi01091 & ~w11800) | (pi01091 & w57252) | (~w11800 & w57252);
assign w14626 = w11800 & w55942;
assign w14627 = ~w14625 & ~w14626;
assign w14628 = (pi01092 & ~w11800) | (pi01092 & w57253) | (~w11800 & w57253);
assign w14629 = w11800 & w55975;
assign w14630 = ~w14628 & ~w14629;
assign w14631 = (pi01093 & ~w11800) | (pi01093 & w57254) | (~w11800 & w57254);
assign w14632 = w11800 & w55977;
assign w14633 = ~w14631 & ~w14632;
assign w14634 = (pi01094 & ~w11800) | (pi01094 & w57255) | (~w11800 & w57255);
assign w14635 = w11800 & w56071;
assign w14636 = ~w14634 & ~w14635;
assign w14637 = (pi01095 & ~w11800) | (pi01095 & w57256) | (~w11800 & w57256);
assign w14638 = w11800 & w55944;
assign w14639 = ~w14637 & ~w14638;
assign w14640 = (pi01096 & ~w11800) | (pi01096 & w57257) | (~w11800 & w57257);
assign w14641 = w11800 & w57143;
assign w14642 = ~w14640 & ~w14641;
assign w14643 = (pi01097 & ~w11800) | (pi01097 & w57258) | (~w11800 & w57258);
assign w14644 = w11800 & w55946;
assign w14645 = ~w14643 & ~w14644;
assign w14646 = (pi01098 & ~w11800) | (pi01098 & w57259) | (~w11800 & w57259);
assign w14647 = w11800 & w56626;
assign w14648 = ~w14646 & ~w14647;
assign w14649 = (pi01099 & ~w11762) | (pi01099 & w57260) | (~w11762 & w57260);
assign w14650 = w11762 & w56290;
assign w14651 = ~w14649 & ~w14650;
assign w14652 = (pi01100 & ~w11762) | (pi01100 & w57261) | (~w11762 & w57261);
assign w14653 = w11762 & w56292;
assign w14654 = ~w14652 & ~w14653;
assign w14655 = (pi01101 & ~w11762) | (pi01101 & w57262) | (~w11762 & w57262);
assign w14656 = w11762 & w56375;
assign w14657 = ~w14655 & ~w14656;
assign w14658 = (pi01102 & ~w11762) | (pi01102 & w57263) | (~w11762 & w57263);
assign w14659 = w11762 & w56039;
assign w14660 = ~w14658 & ~w14659;
assign w14661 = (pi01103 & ~w11762) | (pi01103 & w57264) | (~w11762 & w57264);
assign w14662 = w11762 & w55940;
assign w14663 = ~w14661 & ~w14662;
assign w14664 = (pi01104 & ~w11762) | (pi01104 & w57265) | (~w11762 & w57265);
assign w14665 = w11762 & w56369;
assign w14666 = ~w14664 & ~w14665;
assign w14667 = (pi01105 & ~w11762) | (pi01105 & w57266) | (~w11762 & w57266);
assign w14668 = w11762 & w56300;
assign w14669 = ~w14667 & ~w14668;
assign w14670 = (pi01106 & ~w11762) | (pi01106 & w57267) | (~w11762 & w57267);
assign w14671 = w11762 & w56633;
assign w14672 = ~w14670 & ~w14671;
assign w14673 = (pi01107 & ~w11762) | (pi01107 & w57268) | (~w11762 & w57268);
assign w14674 = w11762 & w56043;
assign w14675 = ~w14673 & ~w14674;
assign w14676 = (pi01108 & ~w11762) | (pi01108 & w57269) | (~w11762 & w57269);
assign w14677 = w11762 & w55942;
assign w14678 = ~w14676 & ~w14677;
assign w14679 = (pi01109 & ~w11762) | (pi01109 & w57270) | (~w11762 & w57270);
assign w14680 = w11762 & w57143;
assign w14681 = ~w14679 & ~w14680;
assign w14682 = (pi01110 & ~w11762) | (pi01110 & w57271) | (~w11762 & w57271);
assign w14683 = w11762 & w56047;
assign w14684 = ~w14682 & ~w14683;
assign w14685 = (pi01111 & ~w11800) | (pi01111 & w57272) | (~w11800 & w57272);
assign w14686 = w11800 & w56077;
assign w14687 = ~w14685 & ~w14686;
assign w14688 = (pi01112 & ~w11800) | (pi01112 & w57273) | (~w11800 & w57273);
assign w14689 = w11800 & w56050;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = (pi01113 & ~w11800) | (pi01113 & w57274) | (~w11800 & w57274);
assign w14692 = w11800 & w55954;
assign w14693 = ~w14691 & ~w14692;
assign w14694 = (pi01114 & ~w11800) | (pi01114 & w57275) | (~w11800 & w57275);
assign w14695 = w11800 & w56083;
assign w14696 = ~w14694 & ~w14695;
assign w14697 = (pi01115 & ~w11800) | (pi01115 & w57276) | (~w11800 & w57276);
assign w14698 = w11800 & w55962;
assign w14699 = ~w14697 & ~w14698;
assign w14700 = (pi01116 & ~w11800) | (pi01116 & w57277) | (~w11800 & w57277);
assign w14701 = w11800 & w56056;
assign w14702 = ~w14700 & ~w14701;
assign w14703 = (pi01117 & ~w11800) | (pi01117 & w57278) | (~w11800 & w57278);
assign w14704 = w11800 & w56092;
assign w14705 = ~w14703 & ~w14704;
assign w14706 = (pi01118 & ~w11800) | (pi01118 & w57279) | (~w11800 & w57279);
assign w14707 = w11800 & w56106;
assign w14708 = ~w14706 & ~w14707;
assign w14709 = (pi01119 & ~w11762) | (pi01119 & w57280) | (~w11762 & w57280);
assign w14710 = w11762 & w56310;
assign w14711 = ~w14709 & ~w14710;
assign w14712 = (pi01120 & ~w11762) | (pi01120 & w57281) | (~w11762 & w57281);
assign w14713 = w11762 & w55950;
assign w14714 = ~w14712 & ~w14713;
assign w14715 = (pi01121 & ~w11762) | (pi01121 & w57282) | (~w11762 & w57282);
assign w14716 = w11762 & w56050;
assign w14717 = ~w14715 & ~w14716;
assign w14718 = (pi01122 & ~w11762) | (pi01122 & w57283) | (~w11762 & w57283);
assign w14719 = w11762 & w55956;
assign w14720 = ~w14718 & ~w14719;
assign w14721 = (pi01123 & ~w11762) | (pi01123 & w57284) | (~w11762 & w57284);
assign w14722 = w11762 & w56316;
assign w14723 = ~w14721 & ~w14722;
assign w14724 = (pi01124 & ~w11762) | (pi01124 & w57285) | (~w11762 & w57285);
assign w14725 = w11762 & w56056;
assign w14726 = ~w14724 & ~w14725;
assign w14727 = (pi01125 & ~w11762) | (pi01125 & w57286) | (~w11762 & w57286);
assign w14728 = w11762 & w56389;
assign w14729 = ~w14727 & ~w14728;
assign w14730 = (pi01126 & ~w11762) | (pi01126 & w57287) | (~w11762 & w57287);
assign w14731 = w11762 & w56393;
assign w14732 = ~w14730 & ~w14731;
assign w14733 = (pi01127 & ~w11762) | (pi01127 & w57288) | (~w11762 & w57288);
assign w14734 = w11762 & w56058;
assign w14735 = ~w14733 & ~w14734;
assign w14736 = (pi01128 & ~w11762) | (pi01128 & w57289) | (~w11762 & w57289);
assign w14737 = w11762 & w55966;
assign w14738 = ~w14736 & ~w14737;
assign w14739 = (pi01129 & ~w11762) | (pi01129 & w57290) | (~w11762 & w57290);
assign w14740 = w11762 & w56323;
assign w14741 = ~w14739 & ~w14740;
assign w14742 = (pi01130 & ~w11762) | (pi01130 & w57291) | (~w11762 & w57291);
assign w14743 = w11762 & w56062;
assign w14744 = ~w14742 & ~w14743;
assign w14745 = (pi01131 & ~w11762) | (pi01131 & w57292) | (~w11762 & w57292);
assign w14746 = w11762 & w56154;
assign w14747 = ~w14745 & ~w14746;
assign w14748 = (pi01132 & ~w11800) | (pi01132 & w57293) | (~w11800 & w57293);
assign w14749 = w11800 & w57192;
assign w14750 = ~w14748 & ~w14749;
assign w14751 = (pi01133 & ~w11800) | (pi01133 & w57294) | (~w11800 & w57294);
assign w14752 = w11800 & w56341;
assign w14753 = ~w14751 & ~w14752;
assign w14754 = (pi01134 & ~w11800) | (pi01134 & w57295) | (~w11800 & w57295);
assign w14755 = w11800 & w56326;
assign w14756 = ~w14754 & ~w14755;
assign w14757 = (pi01135 & ~w11800) | (pi01135 & w57296) | (~w11800 & w57296);
assign w14758 = w11800 & w56333;
assign w14759 = ~w14757 & ~w14758;
assign w14760 = (pi01136 & ~w11800) | (pi01136 & w57297) | (~w11800 & w57297);
assign w14761 = w11800 & w56418;
assign w14762 = ~w14760 & ~w14761;
assign w14763 = (pi01137 & ~w11800) | (pi01137 & w57298) | (~w11800 & w57298);
assign w14764 = w11800 & w56335;
assign w14765 = ~w14763 & ~w14764;
assign w14766 = (pi01138 & ~w11800) | (pi01138 & w57299) | (~w11800 & w57299);
assign w14767 = w11800 & w56644;
assign w14768 = ~w14766 & ~w14767;
assign w14769 = (pi01139 & ~w11762) | (pi01139 & w57300) | (~w11762 & w57300);
assign w14770 = w11762 & w56094;
assign w14771 = ~w14769 & ~w14770;
assign w14772 = (pi01140 & ~w11762) | (pi01140 & w57301) | (~w11762 & w57301);
assign w14773 = w11762 & w57192;
assign w14774 = ~w14772 & ~w14773;
assign w14775 = (pi01141 & ~w11762) | (pi01141 & w57302) | (~w11762 & w57302);
assign w14776 = w11762 & w56108;
assign w14777 = ~w14775 & ~w14776;
assign w14778 = (pi01142 & ~w11762) | (pi01142 & w57303) | (~w11762 & w57303);
assign w14779 = w11762 & w56326;
assign w14780 = ~w14778 & ~w14779;
assign w14781 = (pi01143 & ~w11762) | (pi01143 & w57304) | (~w11762 & w57304);
assign w14782 = w11762 & w55998;
assign w14783 = ~w14781 & ~w14782;
assign w14784 = (pi01144 & ~w11762) | (pi01144 & w57305) | (~w11762 & w57305);
assign w14785 = w11762 & w56114;
assign w14786 = ~w14784 & ~w14785;
assign w14787 = (pi01145 & ~w11762) | (pi01145 & w57306) | (~w11762 & w57306);
assign w14788 = w11762 & w56116;
assign w14789 = ~w14787 & ~w14788;
assign w14790 = (pi01146 & ~w11762) | (pi01146 & w57307) | (~w11762 & w57307);
assign w14791 = w11762 & w56644;
assign w14792 = ~w14790 & ~w14791;
assign w14793 = (pi01147 & ~w11711) | (pi01147 & w57308) | (~w11711 & w57308);
assign w14794 = w11711 & w57229;
assign w14795 = ~w14793 & ~w14794;
assign w14796 = (pi01148 & ~w11711) | (pi01148 & w57309) | (~w11711 & w57309);
assign w14797 = w11711 & w56132;
assign w14798 = ~w14796 & ~w14797;
assign w14799 = (pi01149 & ~w11711) | (pi01149 & w57310) | (~w11711 & w57310);
assign w14800 = w11711 & w56136;
assign w14801 = ~w14799 & ~w14800;
assign w14802 = (pi01150 & ~w11711) | (pi01150 & w57311) | (~w11711 & w57311);
assign w14803 = w11711 & w56013;
assign w14804 = ~w14802 & ~w14803;
assign w14805 = (pi01151 & ~w11711) | (pi01151 & w57312) | (~w11711 & w57312);
assign w14806 = w11711 & w56015;
assign w14807 = ~w14805 & ~w14806;
assign w14808 = (pi01152 & ~w11711) | (pi01152 & w57313) | (~w11711 & w57313);
assign w14809 = w11711 & w56146;
assign w14810 = ~w14808 & ~w14809;
assign w14811 = (pi01153 & ~w11711) | (pi01153 & w57314) | (~w11711 & w57314);
assign w14812 = w11711 & w56150;
assign w14813 = ~w14811 & ~w14812;
assign w14814 = (pi01154 & ~w11711) | (pi01154 & w57315) | (~w11711 & w57315);
assign w14815 = w11711 & w56021;
assign w14816 = ~w14814 & ~w14815;
assign w14817 = (pi01155 & ~w11711) | (pi01155 & w57316) | (~w11711 & w57316);
assign w14818 = w11711 & w56152;
assign w14819 = ~w14817 & ~w14818;
assign w14820 = (pi01156 & ~w11711) | (pi01156 & w57317) | (~w11711 & w57317);
assign w14821 = w11711 & w56023;
assign w14822 = ~w14820 & ~w14821;
assign w14823 = (pi01157 & ~w11711) | (pi01157 & w57318) | (~w11711 & w57318);
assign w14824 = w11711 & w56025;
assign w14825 = ~w14823 & ~w14824;
assign w14826 = (pi01158 & ~w11828) | (pi01158 & w57319) | (~w11828 & w57319);
assign w14827 = w11828 & w56428;
assign w14828 = ~w14826 & ~w14827;
assign w14829 = (pi01159 & ~w11828) | (pi01159 & w57320) | (~w11828 & w57320);
assign w14830 = w11828 & w57229;
assign w14831 = ~w14829 & ~w14830;
assign w14832 = (pi01160 & ~w11828) | (pi01160 & w57321) | (~w11828 & w57321);
assign w14833 = w11828 & w56613;
assign w14834 = ~w14832 & ~w14833;
assign w14835 = (pi01161 & ~w11828) | (pi01161 & w57322) | (~w11828 & w57322);
assign w14836 = w11828 & w56441;
assign w14837 = ~w14835 & ~w14836;
assign w14838 = (pi01162 & ~w11828) | (pi01162 & w57323) | (~w11828 & w57323);
assign w14839 = w11828 & w56443;
assign w14840 = ~w14838 & ~w14839;
assign w14841 = (pi01163 & ~w11828) | (pi01163 & w57324) | (~w11828 & w57324);
assign w14842 = w11828 & w56362;
assign w14843 = ~w14841 & ~w14842;
assign w14844 = (w1192 & ~w10688) | (w1192 & w57325) | (~w10688 & w57325);
assign w14845 = pi01164 & w14844;
assign w14846 = pi01164 & ~w11706;
assign w14847 = ~w14844 & ~w14846;
assign w14848 = ~w14845 & ~w14847;
assign w14849 = w1192 & w11706;
assign w14850 = ~w14848 & ~w14849;
assign w14851 = pi01253 & pi10359;
assign w14852 = ~pi01165 & ~w14851;
assign w14853 = ~w290 & ~w14852;
assign w14854 = w76 & ~w810;
assign w14855 = w76 & w1100;
assign w14856 = ~pi10020 & ~pi10266;
assign w14857 = pi10030 & w826;
assign w14858 = ~w12726 & ~w14857;
assign w14859 = ~pi01168 & w14858;
assign w14860 = ~w14856 & ~w14859;
assign w14861 = pi09825 & pi09856;
assign w14862 = ~pi09855 & w12993;
assign w14863 = pi01209 & w12987;
assign w14864 = (w1789 & ~w12987) | (w1789 & w57326) | (~w12987 & w57326);
assign w14865 = w14864 & w57327;
assign w14866 = w14861 & w14865;
assign w14867 = (pi01169 & ~w14865) | (pi01169 & w57328) | (~w14865 & w57328);
assign w14868 = w14865 & w57329;
assign w14869 = ~w14867 & ~w14868;
assign w14870 = (pi01170 & ~w318) | (pi01170 & w57330) | (~w318 & w57330);
assign w14871 = ~w789 & ~w14870;
assign w14872 = ~pi09818 & ~pi09955;
assign w14873 = ~pi09958 & ~pi09960;
assign w14874 = w14872 & w14873;
assign w14875 = (~pi02670 & w14874) | (~pi02670 & w57331) | (w14874 & w57331);
assign w14876 = pi09818 & pi09955;
assign w14877 = pi09958 & ~pi09960;
assign w14878 = w12993 & w14876;
assign w14879 = w14877 & w14878;
assign w14880 = w14878 & w57332;
assign w14881 = w14872 & w14877;
assign w14882 = ~pi01415 & w14881;
assign w14883 = pi09818 & ~pi09955;
assign w14884 = w14877 & w14883;
assign w14885 = ~pi10171 & w14884;
assign w14886 = w14873 & w14876;
assign w14887 = ~pi10293 & w14886;
assign w14888 = ~pi09958 & pi09960;
assign w14889 = w14883 & w14888;
assign w14890 = ~pi10041 & w14889;
assign w14891 = w14876 & w14888;
assign w14892 = ~pi10338 & w14891;
assign w14893 = w14872 & w14888;
assign w14894 = ~pi10204 & w14893;
assign w14895 = pi09958 & pi09960;
assign w14896 = w14872 & w14895;
assign w14897 = ~pi10080 & w14896;
assign w14898 = ~pi09818 & pi09955;
assign w14899 = w14877 & w14898;
assign w14900 = ~pi10271 & w14899;
assign w14901 = w14883 & w14895;
assign w14902 = ~pi01359 & w14901;
assign w14903 = w14873 & w14898;
assign w14904 = ~pi10298 & w14903;
assign w14905 = w14895 & w14898;
assign w14906 = ~pi10313 & w14905;
assign w14907 = w14888 & w14898;
assign w14908 = ~pi10054 & w14907;
assign w14909 = w14876 & w14895;
assign w14910 = ~pi01289 & w14909;
assign w14911 = w14873 & w14883;
assign w14912 = ~pi01401 & w14911;
assign w14913 = ~w14882 & ~w14885;
assign w14914 = ~w14887 & ~w14890;
assign w14915 = ~w14892 & ~w14894;
assign w14916 = ~w14897 & ~w14900;
assign w14917 = ~w14902 & ~w14904;
assign w14918 = ~w14906 & ~w14908;
assign w14919 = ~w14910 & ~w14912;
assign w14920 = w14918 & w14919;
assign w14921 = w14916 & w14917;
assign w14922 = w14914 & w14915;
assign w14923 = w14913 & w14922;
assign w14924 = w14920 & w14921;
assign w14925 = w14923 & w14924;
assign w14926 = w12993 & ~w14925;
assign w14927 = ~w14875 & ~w14880;
assign w14928 = ~w14926 & w14927;
assign w14929 = (~pi02668 & w14874) | (~pi02668 & w57333) | (w14874 & w57333);
assign w14930 = w14878 & w57334;
assign w14931 = ~pi01226 & w14886;
assign w14932 = ~pi10323 & w14901;
assign w14933 = ~pi10217 & w14889;
assign w14934 = ~pi01370 & w14905;
assign w14935 = ~pi10070 & w14891;
assign w14936 = ~pi10003 & w14907;
assign w14937 = ~pi10279 & w14884;
assign w14938 = ~pi02689 & w14909;
assign w14939 = ~pi10131 & w14903;
assign w14940 = ~pi10116 & w14911;
assign w14941 = ~pi10184 & w14899;
assign w14942 = ~pi01416 & w14881;
assign w14943 = ~pi10081 & w14896;
assign w14944 = ~pi02694 & w14893;
assign w14945 = ~w14931 & ~w14932;
assign w14946 = ~w14933 & ~w14934;
assign w14947 = ~w14935 & ~w14936;
assign w14948 = ~w14937 & ~w14938;
assign w14949 = ~w14939 & ~w14940;
assign w14950 = ~w14941 & ~w14942;
assign w14951 = ~w14943 & ~w14944;
assign w14952 = w14950 & w14951;
assign w14953 = w14948 & w14949;
assign w14954 = w14946 & w14947;
assign w14955 = w14945 & w14954;
assign w14956 = w14952 & w14953;
assign w14957 = w14955 & w14956;
assign w14958 = w12993 & ~w14957;
assign w14959 = ~w14929 & ~w14930;
assign w14960 = ~w14958 & w14959;
assign w14961 = (~pi01336 & w14874) | (~pi01336 & w57335) | (w14874 & w57335);
assign w14962 = w14878 & w57336;
assign w14963 = ~pi10039 & w14889;
assign w14964 = ~pi01225 & w14886;
assign w14965 = ~pi10337 & w14891;
assign w14966 = ~pi02217 & w14909;
assign w14967 = ~pi10326 & w14896;
assign w14968 = ~pi01323 & w14884;
assign w14969 = ~pi10055 & w14907;
assign w14970 = ~pi01371 & w14905;
assign w14971 = ~pi10117 & w14911;
assign w14972 = ~pi01448 & w14893;
assign w14973 = ~pi01298 & w14899;
assign w14974 = ~pi10302 & w14903;
assign w14975 = ~pi10283 & w14881;
assign w14976 = ~pi01360 & w14901;
assign w14977 = ~w14963 & ~w14964;
assign w14978 = ~w14965 & ~w14966;
assign w14979 = ~w14967 & ~w14968;
assign w14980 = ~w14969 & ~w14970;
assign w14981 = ~w14971 & ~w14972;
assign w14982 = ~w14973 & ~w14974;
assign w14983 = ~w14975 & ~w14976;
assign w14984 = w14982 & w14983;
assign w14985 = w14980 & w14981;
assign w14986 = w14978 & w14979;
assign w14987 = w14977 & w14986;
assign w14988 = w14984 & w14985;
assign w14989 = w14987 & w14988;
assign w14990 = w12993 & ~w14989;
assign w14991 = ~w14961 & ~w14962;
assign w14992 = ~w14990 & w14991;
assign w14993 = (~pi02669 & w14874) | (~pi02669 & w57337) | (w14874 & w57337);
assign w14994 = w14878 & w57338;
assign w14995 = ~pi01372 & w14905;
assign w14996 = ~pi10172 & w14884;
assign w14997 = ~pi01329 & w14889;
assign w14998 = ~pi01440 & w14893;
assign w14999 = ~pi10048 & w14907;
assign w15000 = ~pi10094 & w14901;
assign w15001 = ~pi01386 & w14909;
assign w15002 = ~pi01220 & w14896;
assign w15003 = ~pi10132 & w14903;
assign w15004 = ~pi01417 & w14881;
assign w15005 = ~pi01236 & w14899;
assign w15006 = ~pi10118 & w14911;
assign w15007 = ~pi10071 & w14891;
assign w15008 = ~pi10294 & w14886;
assign w15009 = ~w14995 & ~w14996;
assign w15010 = ~w14997 & ~w14998;
assign w15011 = ~w14999 & ~w15000;
assign w15012 = ~w15001 & ~w15002;
assign w15013 = ~w15003 & ~w15004;
assign w15014 = ~w15005 & ~w15006;
assign w15015 = ~w15007 & ~w15008;
assign w15016 = w15014 & w15015;
assign w15017 = w15012 & w15013;
assign w15018 = w15010 & w15011;
assign w15019 = w15009 & w15018;
assign w15020 = w15016 & w15017;
assign w15021 = w15019 & w15020;
assign w15022 = w12993 & ~w15021;
assign w15023 = ~w14993 & ~w14994;
assign w15024 = ~w15022 & w15023;
assign w15025 = (~pi01337 & w14874) | (~pi01337 & w57339) | (w14874 & w57339);
assign w15026 = w14878 & w57340;
assign w15027 = ~pi10133 & w14903;
assign w15028 = ~pi01373 & w14905;
assign w15029 = ~pi01227 & w14886;
assign w15030 = ~pi01295 & w14889;
assign w15031 = ~pi10321 & w14901;
assign w15032 = ~pi10272 & w14907;
assign w15033 = ~pi01387 & w14909;
assign w15034 = ~pi10082 & w14896;
assign w15035 = ~pi01402 & w14911;
assign w15036 = ~pi10161 & w14881;
assign w15037 = ~pi10269 & w14899;
assign w15038 = ~pi01348 & w14891;
assign w15039 = ~pi10278 & w14884;
assign w15040 = ~pi10205 & w14893;
assign w15041 = ~w15027 & ~w15028;
assign w15042 = ~w15029 & ~w15030;
assign w15043 = ~w15031 & ~w15032;
assign w15044 = ~w15033 & ~w15034;
assign w15045 = ~w15035 & ~w15036;
assign w15046 = ~w15037 & ~w15038;
assign w15047 = ~w15039 & ~w15040;
assign w15048 = w15046 & w15047;
assign w15049 = w15044 & w15045;
assign w15050 = w15042 & w15043;
assign w15051 = w15041 & w15050;
assign w15052 = w15048 & w15049;
assign w15053 = w15051 & w15052;
assign w15054 = w12993 & ~w15053;
assign w15055 = ~w15025 & ~w15026;
assign w15056 = ~w15054 & w15055;
assign w15057 = (~pi01338 & w14874) | (~pi01338 & w57341) | (w14874 & w57341);
assign w15058 = w14878 & w57342;
assign w15059 = ~pi01441 & w14893;
assign w15060 = ~pi10309 & w14911;
assign w15061 = ~pi01330 & w14889;
assign w15062 = ~pi01388 & w14909;
assign w15063 = ~pi10173 & w14884;
assign w15064 = ~pi01349 & w14891;
assign w15065 = ~pi10134 & w14903;
assign w15066 = ~pi01237 & w14899;
assign w15067 = ~pi01221 & w14896;
assign w15068 = ~pi01361 & w14901;
assign w15069 = ~pi10285 & w14881;
assign w15070 = ~pi01313 & w14907;
assign w15071 = ~pi10147 & w14886;
assign w15072 = ~pi02685 & w14905;
assign w15073 = ~w15059 & ~w15060;
assign w15074 = ~w15061 & ~w15062;
assign w15075 = ~w15063 & ~w15064;
assign w15076 = ~w15065 & ~w15066;
assign w15077 = ~w15067 & ~w15068;
assign w15078 = ~w15069 & ~w15070;
assign w15079 = ~w15071 & ~w15072;
assign w15080 = w15078 & w15079;
assign w15081 = w15076 & w15077;
assign w15082 = w15074 & w15075;
assign w15083 = w15073 & w15082;
assign w15084 = w15080 & w15081;
assign w15085 = w15083 & w15084;
assign w15086 = w12993 & ~w15085;
assign w15087 = ~w15057 & ~w15058;
assign w15088 = ~w15086 & w15087;
assign w15089 = (~pi02671 & w14874) | (~pi02671 & w57343) | (w14874 & w57343);
assign w15090 = w14878 & w57344;
assign w15091 = ~pi10083 & w14896;
assign w15092 = ~pi10174 & w14884;
assign w15093 = ~pi01350 & w14891;
assign w15094 = ~pi10218 & w14889;
assign w15095 = ~pi01362 & w14901;
assign w15096 = ~pi10162 & w14881;
assign w15097 = ~pi01389 & w14909;
assign w15098 = ~pi01374 & w14905;
assign w15099 = ~pi10148 & w14886;
assign w15100 = ~pi10341 & w14907;
assign w15101 = ~pi10185 & w14899;
assign w15102 = ~pi10053 & w14893;
assign w15103 = ~pi10119 & w14911;
assign w15104 = ~pi01412 & w14903;
assign w15105 = ~w15091 & ~w15092;
assign w15106 = ~w15093 & ~w15094;
assign w15107 = ~w15095 & ~w15096;
assign w15108 = ~w15097 & ~w15098;
assign w15109 = ~w15099 & ~w15100;
assign w15110 = ~w15101 & ~w15102;
assign w15111 = ~w15103 & ~w15104;
assign w15112 = w15110 & w15111;
assign w15113 = w15108 & w15109;
assign w15114 = w15106 & w15107;
assign w15115 = w15105 & w15114;
assign w15116 = w15112 & w15113;
assign w15117 = w15115 & w15116;
assign w15118 = w12993 & ~w15117;
assign w15119 = ~w15089 & ~w15090;
assign w15120 = ~w15118 & w15119;
assign w15121 = (~pi01339 & w14874) | (~pi01339 & w57345) | (w14874 & w57345);
assign w15122 = w14878 & w57346;
assign w15123 = ~pi10175 & w14884;
assign w15124 = ~pi01442 & w14893;
assign w15125 = ~pi10084 & w14896;
assign w15126 = ~pi01395 & w14909;
assign w15127 = ~pi02228 & w14905;
assign w15128 = ~pi10120 & w14911;
assign w15129 = ~pi01351 & w14891;
assign w15130 = ~pi01410 & w14903;
assign w15131 = ~pi01238 & w14899;
assign w15132 = ~pi10056 & w14907;
assign w15133 = ~pi10095 & w14901;
assign w15134 = ~pi10032 & w14889;
assign w15135 = ~pi10149 & w14886;
assign w15136 = ~pi01418 & w14881;
assign w15137 = ~w15123 & ~w15124;
assign w15138 = ~w15125 & ~w15126;
assign w15139 = ~w15127 & ~w15128;
assign w15140 = ~w15129 & ~w15130;
assign w15141 = ~w15131 & ~w15132;
assign w15142 = ~w15133 & ~w15134;
assign w15143 = ~w15135 & ~w15136;
assign w15144 = w15142 & w15143;
assign w15145 = w15140 & w15141;
assign w15146 = w15138 & w15139;
assign w15147 = w15137 & w15146;
assign w15148 = w15144 & w15145;
assign w15149 = w15147 & w15148;
assign w15150 = w12993 & ~w15149;
assign w15151 = ~w15121 & ~w15122;
assign w15152 = ~w15150 & w15151;
assign w15153 = (~pi01340 & w14874) | (~pi01340 & w57347) | (w14874 & w57347);
assign w15154 = w14878 & w57348;
assign w15155 = ~pi01285 & w14911;
assign w15156 = ~pi01352 & w14891;
assign w15157 = ~pi10273 & w14884;
assign w15158 = ~pi10332 & w14896;
assign w15159 = ~pi10106 & w14905;
assign w15160 = ~pi10268 & w14899;
assign w15161 = ~pi01411 & w14903;
assign w15162 = ~pi10057 & w14907;
assign w15163 = ~pi01443 & w14893;
assign w15164 = ~pi10322 & w14901;
assign w15165 = ~pi10295 & w14886;
assign w15166 = ~pi01419 & w14881;
assign w15167 = ~pi01390 & w14909;
assign w15168 = ~pi10219 & w14889;
assign w15169 = ~w15155 & ~w15156;
assign w15170 = ~w15157 & ~w15158;
assign w15171 = ~w15159 & ~w15160;
assign w15172 = ~w15161 & ~w15162;
assign w15173 = ~w15163 & ~w15164;
assign w15174 = ~w15165 & ~w15166;
assign w15175 = ~w15167 & ~w15168;
assign w15176 = w15174 & w15175;
assign w15177 = w15172 & w15173;
assign w15178 = w15170 & w15171;
assign w15179 = w15169 & w15178;
assign w15180 = w15176 & w15177;
assign w15181 = w15179 & w15180;
assign w15182 = w12993 & ~w15181;
assign w15183 = ~w15153 & ~w15154;
assign w15184 = ~w15182 & w15183;
assign w15185 = (~pi02256 & w14874) | (~pi02256 & w57349) | (w14874 & w57349);
assign w15186 = w14878 & w57350;
assign w15187 = ~pi02216 & w14909;
assign w15188 = ~pi01228 & w14886;
assign w15189 = ~pi01420 & w14881;
assign w15190 = ~pi10317 & w14905;
assign w15191 = ~pi01322 & w14884;
assign w15192 = ~pi10096 & w14901;
assign w15193 = ~pi01279 & w14891;
assign w15194 = ~pi01296 & w14899;
assign w15195 = ~pi01314 & w14907;
assign w15196 = ~pi10121 & w14911;
assign w15197 = ~pi01222 & w14896;
assign w15198 = ~pi10206 & w14893;
assign w15199 = ~pi10038 & w14889;
assign w15200 = ~pi10303 & w14903;
assign w15201 = ~w15187 & ~w15188;
assign w15202 = ~w15189 & ~w15190;
assign w15203 = ~w15191 & ~w15192;
assign w15204 = ~w15193 & ~w15194;
assign w15205 = ~w15195 & ~w15196;
assign w15206 = ~w15197 & ~w15198;
assign w15207 = ~w15199 & ~w15200;
assign w15208 = w15206 & w15207;
assign w15209 = w15204 & w15205;
assign w15210 = w15202 & w15203;
assign w15211 = w15201 & w15210;
assign w15212 = w15208 & w15209;
assign w15213 = w15211 & w15212;
assign w15214 = w12993 & ~w15213;
assign w15215 = ~w15185 & ~w15186;
assign w15216 = ~w15214 & w15215;
assign w15217 = (~pi02673 & w14874) | (~pi02673 & w57351) | (w14874 & w57351);
assign w15218 = w14878 & w57352;
assign w15219 = ~pi01421 & w14881;
assign w15220 = ~pi10135 & w14903;
assign w15221 = ~pi10058 & w14907;
assign w15222 = ~pi10308 & w14911;
assign w15223 = ~pi01232 & w14884;
assign w15224 = ~pi10085 & w14896;
assign w15225 = ~pi10186 & w14899;
assign w15226 = ~pi10220 & w14889;
assign w15227 = ~pi10107 & w14905;
assign w15228 = ~pi01444 & w14893;
assign w15229 = ~pi10097 & w14901;
assign w15230 = ~pi01320 & w14886;
assign w15231 = ~pi01391 & w14909;
assign w15232 = ~pi01353 & w14891;
assign w15233 = ~w15219 & ~w15220;
assign w15234 = ~w15221 & ~w15222;
assign w15235 = ~w15223 & ~w15224;
assign w15236 = ~w15225 & ~w15226;
assign w15237 = ~w15227 & ~w15228;
assign w15238 = ~w15229 & ~w15230;
assign w15239 = ~w15231 & ~w15232;
assign w15240 = w15238 & w15239;
assign w15241 = w15236 & w15237;
assign w15242 = w15234 & w15235;
assign w15243 = w15233 & w15242;
assign w15244 = w15240 & w15241;
assign w15245 = w15243 & w15244;
assign w15246 = w12993 & ~w15245;
assign w15247 = ~w15217 & ~w15218;
assign w15248 = ~w15246 & w15247;
assign w15249 = (~pi02672 & w14874) | (~pi02672 & w57353) | (w14874 & w57353);
assign w15250 = w14878 & w57354;
assign w15251 = ~pi10122 & w14911;
assign w15252 = ~pi10221 & w14889;
assign w15253 = ~pi01422 & w14881;
assign w15254 = ~pi10346 & w14907;
assign w15255 = ~pi01375 & w14905;
assign w15256 = ~pi10300 & w14903;
assign w15257 = ~pi01239 & w14899;
assign w15258 = ~pi10098 & w14901;
assign w15259 = ~pi10072 & w14891;
assign w15260 = ~pi10150 & w14886;
assign w15261 = ~pi01300 & w14884;
assign w15262 = ~pi01280 & w14893;
assign w15263 = ~pi01392 & w14909;
assign w15264 = ~pi10329 & w14896;
assign w15265 = ~w15251 & ~w15252;
assign w15266 = ~w15253 & ~w15254;
assign w15267 = ~w15255 & ~w15256;
assign w15268 = ~w15257 & ~w15258;
assign w15269 = ~w15259 & ~w15260;
assign w15270 = ~w15261 & ~w15262;
assign w15271 = ~w15263 & ~w15264;
assign w15272 = w15270 & w15271;
assign w15273 = w15268 & w15269;
assign w15274 = w15266 & w15267;
assign w15275 = w15265 & w15274;
assign w15276 = w15272 & w15273;
assign w15277 = w15275 & w15276;
assign w15278 = w12993 & ~w15277;
assign w15279 = ~w15249 & ~w15250;
assign w15280 = ~w15278 & w15279;
assign w15281 = (~pi02253 & w14874) | (~pi02253 & w57355) | (w14874 & w57355);
assign w15282 = w14878 & w57356;
assign w15283 = ~pi10108 & w14905;
assign w15284 = ~pi10176 & w14884;
assign w15285 = ~pi01282 & w14881;
assign w15286 = ~pi02683 & w14891;
assign w15287 = ~pi10151 & w14886;
assign w15288 = ~pi10207 & w14893;
assign w15289 = ~pi10136 & w14903;
assign w15290 = ~pi10331 & w14896;
assign w15291 = ~pi10123 & w14911;
assign w15292 = ~pi01363 & w14901;
assign w15293 = ~pi01240 & w14899;
assign w15294 = ~pi01331 & w14889;
assign w15295 = ~pi01393 & w14909;
assign w15296 = ~pi10059 & w14907;
assign w15297 = ~w15283 & ~w15284;
assign w15298 = ~w15285 & ~w15286;
assign w15299 = ~w15287 & ~w15288;
assign w15300 = ~w15289 & ~w15290;
assign w15301 = ~w15291 & ~w15292;
assign w15302 = ~w15293 & ~w15294;
assign w15303 = ~w15295 & ~w15296;
assign w15304 = w15302 & w15303;
assign w15305 = w15300 & w15301;
assign w15306 = w15298 & w15299;
assign w15307 = w15297 & w15306;
assign w15308 = w15304 & w15305;
assign w15309 = w15307 & w15308;
assign w15310 = w12993 & ~w15309;
assign w15311 = ~w15281 & ~w15282;
assign w15312 = ~w15310 & w15311;
assign w15313 = (~pi01341 & w14874) | (~pi01341 & w57357) | (w14874 & w57357);
assign w15314 = w14878 & w57358;
assign w15315 = ~pi10124 & w14911;
assign w15316 = ~pi10330 & w14896;
assign w15317 = ~pi01394 & w14909;
assign w15318 = ~pi10284 & w14881;
assign w15319 = ~pi10152 & w14886;
assign w15320 = ~pi10222 & w14889;
assign w15321 = ~pi01292 & w14901;
assign w15322 = ~pi10276 & w14884;
assign w15323 = ~pi10073 & w14891;
assign w15324 = ~pi10267 & w14899;
assign w15325 = ~pi10060 & w14907;
assign w15326 = ~pi10301 & w14903;
assign w15327 = ~pi01376 & w14905;
assign w15328 = ~pi10208 & w14893;
assign w15329 = ~w15315 & ~w15316;
assign w15330 = ~w15317 & ~w15318;
assign w15331 = ~w15319 & ~w15320;
assign w15332 = ~w15321 & ~w15322;
assign w15333 = ~w15323 & ~w15324;
assign w15334 = ~w15325 & ~w15326;
assign w15335 = ~w15327 & ~w15328;
assign w15336 = w15334 & w15335;
assign w15337 = w15332 & w15333;
assign w15338 = w15330 & w15331;
assign w15339 = w15329 & w15338;
assign w15340 = w15336 & w15337;
assign w15341 = w15339 & w15340;
assign w15342 = w12993 & ~w15341;
assign w15343 = ~w15313 & ~w15314;
assign w15344 = ~w15342 & w15343;
assign w15345 = (~pi01342 & w14874) | (~pi01342 & w57359) | (w14874 & w57359);
assign w15346 = w14878 & w57360;
assign w15347 = ~pi01283 & w14903;
assign w15348 = ~pi10111 & w14909;
assign w15349 = ~pi10291 & w14886;
assign w15350 = ~pi02235 & w14891;
assign w15351 = ~pi10109 & w14905;
assign w15352 = ~pi10320 & w14901;
assign w15353 = ~pi10187 & w14899;
assign w15354 = ~pi10036 & w14889;
assign w15355 = ~pi10043 & w14893;
assign w15356 = ~pi01423 & w14881;
assign w15357 = ~pi10061 & w14907;
assign w15358 = ~pi10274 & w14884;
assign w15359 = ~pi10305 & w14911;
assign w15360 = ~pi01316 & w14896;
assign w15361 = ~w15347 & ~w15348;
assign w15362 = ~w15349 & ~w15350;
assign w15363 = ~w15351 & ~w15352;
assign w15364 = ~w15353 & ~w15354;
assign w15365 = ~w15355 & ~w15356;
assign w15366 = ~w15357 & ~w15358;
assign w15367 = ~w15359 & ~w15360;
assign w15368 = w15366 & w15367;
assign w15369 = w15364 & w15365;
assign w15370 = w15362 & w15363;
assign w15371 = w15361 & w15370;
assign w15372 = w15368 & w15369;
assign w15373 = w15371 & w15372;
assign w15374 = w12993 & ~w15373;
assign w15375 = ~w15345 & ~w15346;
assign w15376 = ~w15374 & w15375;
assign w15377 = (~pi02674 & w14874) | (~pi02674 & w57361) | (w14874 & w57361);
assign w15378 = w14878 & w57362;
assign w15379 = ~pi01377 & w14905;
assign w15380 = ~pi01364 & w14901;
assign w15381 = ~pi10223 & w14889;
assign w15382 = ~pi10154 & w14886;
assign w15383 = ~pi10163 & w14881;
assign w15384 = ~pi01241 & w14899;
assign w15385 = ~pi01413 & w14903;
assign w15386 = ~pi10316 & w14909;
assign w15387 = ~pi01354 & w14891;
assign w15388 = ~pi10342 & w14907;
assign w15389 = ~pi01325 & w14884;
assign w15390 = ~pi10209 & w14893;
assign w15391 = ~pi10125 & w14911;
assign w15392 = ~pi10086 & w14896;
assign w15393 = ~w15379 & ~w15380;
assign w15394 = ~w15381 & ~w15382;
assign w15395 = ~w15383 & ~w15384;
assign w15396 = ~w15385 & ~w15386;
assign w15397 = ~w15387 & ~w15388;
assign w15398 = ~w15389 & ~w15390;
assign w15399 = ~w15391 & ~w15392;
assign w15400 = w15398 & w15399;
assign w15401 = w15396 & w15397;
assign w15402 = w15394 & w15395;
assign w15403 = w15393 & w15402;
assign w15404 = w15400 & w15401;
assign w15405 = w15403 & w15404;
assign w15406 = w12993 & ~w15405;
assign w15407 = ~w15377 & ~w15378;
assign w15408 = ~w15406 & w15407;
assign w15409 = (~pi01343 & w14874) | (~pi01343 & w57363) | (w14874 & w57363);
assign w15410 = w14878 & w57364;
assign w15411 = ~pi10099 & w14901;
assign w15412 = ~pi10087 & w14896;
assign w15413 = ~pi01233 & w14884;
assign w15414 = ~pi10164 & w14881;
assign w15415 = ~pi10062 & w14907;
assign w15416 = ~pi10307 & w14911;
assign w15417 = ~pi10314 & w14905;
assign w15418 = ~pi10137 & w14903;
assign w15419 = ~pi01447 & w14893;
assign w15420 = ~pi10112 & w14909;
assign w15421 = ~pi10188 & w14899;
assign w15422 = ~pi10224 & w14889;
assign w15423 = ~pi10336 & w14891;
assign w15424 = ~pi10292 & w14886;
assign w15425 = ~w15411 & ~w15412;
assign w15426 = ~w15413 & ~w15414;
assign w15427 = ~w15415 & ~w15416;
assign w15428 = ~w15417 & ~w15418;
assign w15429 = ~w15419 & ~w15420;
assign w15430 = ~w15421 & ~w15422;
assign w15431 = ~w15423 & ~w15424;
assign w15432 = w15430 & w15431;
assign w15433 = w15428 & w15429;
assign w15434 = w15426 & w15427;
assign w15435 = w15425 & w15434;
assign w15436 = w15432 & w15433;
assign w15437 = w15435 & w15436;
assign w15438 = w12993 & ~w15437;
assign w15439 = ~w15409 & ~w15410;
assign w15440 = ~w15438 & w15439;
assign w15441 = (~pi02675 & w14874) | (~pi02675 & w57365) | (w14874 & w57365);
assign w15442 = w14878 & w57366;
assign w15443 = ~pi01223 & w14896;
assign w15444 = ~pi01301 & w14886;
assign w15445 = ~pi10044 & w14893;
assign w15446 = ~pi10100 & w14901;
assign w15447 = ~pi10113 & w14909;
assign w15448 = ~pi01324 & w14884;
assign w15449 = ~pi01169 & w14899;
assign w15450 = ~pi10074 & w14891;
assign w15451 = ~pi01414 & w14903;
assign w15452 = ~pi10165 & w14881;
assign w15453 = ~pi10344 & w14907;
assign w15454 = ~pi01333 & w14889;
assign w15455 = ~pi01403 & w14911;
assign w15456 = ~pi01378 & w14905;
assign w15457 = ~w15443 & ~w15444;
assign w15458 = ~w15445 & ~w15446;
assign w15459 = ~w15447 & ~w15448;
assign w15460 = ~w15449 & ~w15450;
assign w15461 = ~w15451 & ~w15452;
assign w15462 = ~w15453 & ~w15454;
assign w15463 = ~w15455 & ~w15456;
assign w15464 = w15462 & w15463;
assign w15465 = w15460 & w15461;
assign w15466 = w15458 & w15459;
assign w15467 = w15457 & w15466;
assign w15468 = w15464 & w15465;
assign w15469 = w15467 & w15468;
assign w15470 = w12993 & ~w15469;
assign w15471 = ~w15441 & ~w15442;
assign w15472 = ~w15470 & w15471;
assign w15473 = (~pi01344 & w14874) | (~pi01344 & w57367) | (w14874 & w57367);
assign w15474 = w14878 & w57368;
assign w15475 = ~pi10282 & w14881;
assign w15476 = ~pi10101 & w14901;
assign w15477 = ~pi01290 & w14905;
assign w15478 = ~pi01234 & w14884;
assign w15479 = ~pi10114 & w14909;
assign w15480 = ~pi10045 & w14893;
assign w15481 = ~pi01404 & w14911;
assign w15482 = ~pi10138 & w14903;
assign w15483 = ~pi10155 & w14886;
assign w15484 = ~pi10334 & w14891;
assign w15485 = ~pi10189 & w14899;
assign w15486 = ~pi10088 & w14896;
assign w15487 = ~pi01332 & w14889;
assign w15488 = ~pi10063 & w14907;
assign w15489 = ~w15475 & ~w15476;
assign w15490 = ~w15477 & ~w15478;
assign w15491 = ~w15479 & ~w15480;
assign w15492 = ~w15481 & ~w15482;
assign w15493 = ~w15483 & ~w15484;
assign w15494 = ~w15485 & ~w15486;
assign w15495 = ~w15487 & ~w15488;
assign w15496 = w15494 & w15495;
assign w15497 = w15492 & w15493;
assign w15498 = w15490 & w15491;
assign w15499 = w15489 & w15498;
assign w15500 = w15496 & w15497;
assign w15501 = w15499 & w15500;
assign w15502 = w12993 & ~w15501;
assign w15503 = ~w15473 & ~w15474;
assign w15504 = ~w15502 & w15503;
assign w15505 = (~pi01345 & w14874) | (~pi01345 & w57369) | (w14874 & w57369);
assign w15506 = w14878 & w57370;
assign w15507 = ~pi02686 & w14905;
assign w15508 = ~pi10126 & w14911;
assign w15509 = ~pi10275 & w14884;
assign w15510 = ~pi10046 & w14893;
assign w15511 = ~pi10225 & w14889;
assign w15512 = ~pi01218 & w14907;
assign w15513 = ~pi01317 & w14896;
assign w15514 = ~pi02684 & w14891;
assign w15515 = ~pi10289 & w14886;
assign w15516 = ~pi02691 & w14881;
assign w15517 = ~pi01242 & w14899;
assign w15518 = ~pi02690 & w14909;
assign w15519 = ~pi10139 & w14903;
assign w15520 = ~pi01365 & w14901;
assign w15521 = ~w15507 & ~w15508;
assign w15522 = ~w15509 & ~w15510;
assign w15523 = ~w15511 & ~w15512;
assign w15524 = ~w15513 & ~w15514;
assign w15525 = ~w15515 & ~w15516;
assign w15526 = ~w15517 & ~w15518;
assign w15527 = ~w15519 & ~w15520;
assign w15528 = w15526 & w15527;
assign w15529 = w15524 & w15525;
assign w15530 = w15522 & w15523;
assign w15531 = w15521 & w15530;
assign w15532 = w15528 & w15529;
assign w15533 = w15531 & w15532;
assign w15534 = w12993 & ~w15533;
assign w15535 = ~w15505 & ~w15506;
assign w15536 = ~w15534 & w15535;
assign w15537 = (~pi02676 & w14874) | (~pi02676 & w57371) | (w14874 & w57371);
assign w15538 = w14878 & w57372;
assign w15539 = ~pi01405 & w14911;
assign w15540 = ~pi01327 & w14884;
assign w15541 = ~pi10075 & w14891;
assign w15542 = ~pi10210 & w14893;
assign w15543 = ~pi10299 & w14903;
assign w15544 = ~pi01379 & w14905;
assign w15545 = ~pi01243 & w14899;
assign w15546 = ~pi10312 & w14909;
assign w15547 = ~pi10037 & w14889;
assign w15548 = ~pi10166 & w14881;
assign w15549 = ~pi01318 & w14896;
assign w15550 = ~pi10156 & w14886;
assign w15551 = ~pi10343 & w14907;
assign w15552 = ~pi10319 & w14901;
assign w15553 = ~w15539 & ~w15540;
assign w15554 = ~w15541 & ~w15542;
assign w15555 = ~w15543 & ~w15544;
assign w15556 = ~w15545 & ~w15546;
assign w15557 = ~w15547 & ~w15548;
assign w15558 = ~w15549 & ~w15550;
assign w15559 = ~w15551 & ~w15552;
assign w15560 = w15558 & w15559;
assign w15561 = w15556 & w15557;
assign w15562 = w15554 & w15555;
assign w15563 = w15553 & w15562;
assign w15564 = w15560 & w15561;
assign w15565 = w15563 & w15564;
assign w15566 = w12993 & ~w15565;
assign w15567 = ~w15537 & ~w15538;
assign w15568 = ~w15566 & w15567;
assign w15569 = (~pi02250 & w14874) | (~pi02250 & w57373) | (w14874 & w57373);
assign w15570 = w14878 & w57374;
assign w15571 = ~pi10226 & w14889;
assign w15572 = ~pi10281 & w14881;
assign w15573 = ~pi10211 & w14893;
assign w15574 = ~pi10306 & w14911;
assign w15575 = ~pi10328 & w14896;
assign w15576 = ~pi10177 & w14884;
assign w15577 = ~pi01219 & w14907;
assign w15578 = ~pi10140 & w14903;
assign w15579 = ~pi10190 & w14899;
assign w15580 = ~pi01396 & w14909;
assign w15581 = ~pi01380 & w14905;
assign w15582 = ~pi10335 & w14891;
assign w15583 = ~pi01366 & w14901;
assign w15584 = ~pi01299 & w14886;
assign w15585 = ~w15571 & ~w15572;
assign w15586 = ~w15573 & ~w15574;
assign w15587 = ~w15575 & ~w15576;
assign w15588 = ~w15577 & ~w15578;
assign w15589 = ~w15579 & ~w15580;
assign w15590 = ~w15581 & ~w15582;
assign w15591 = ~w15583 & ~w15584;
assign w15592 = w15590 & w15591;
assign w15593 = w15588 & w15589;
assign w15594 = w15586 & w15587;
assign w15595 = w15585 & w15594;
assign w15596 = w15592 & w15593;
assign w15597 = w15595 & w15596;
assign w15598 = w12993 & ~w15597;
assign w15599 = ~w15569 & ~w15570;
assign w15600 = ~w15598 & w15599;
assign w15601 = (~pi02677 & w14874) | (~pi02677 & w57375) | (w14874 & w57375);
assign w15602 = w14878 & w57376;
assign w15603 = ~pi10127 & w14911;
assign w15604 = ~pi10167 & w14881;
assign w15605 = ~pi10290 & w14886;
assign w15606 = ~pi02201 & w14903;
assign w15607 = ~pi01287 & w14909;
assign w15608 = ~pi01291 & w14901;
assign w15609 = ~pi01288 & w14905;
assign w15610 = ~pi10064 & w14907;
assign w15611 = ~pi10191 & w14899;
assign w15612 = ~pi10178 & w14884;
assign w15613 = ~pi01355 & w14891;
assign w15614 = ~pi10212 & w14893;
assign w15615 = ~pi10089 & w14896;
assign w15616 = ~pi10227 & w14889;
assign w15617 = ~w15603 & ~w15604;
assign w15618 = ~w15605 & ~w15606;
assign w15619 = ~w15607 & ~w15608;
assign w15620 = ~w15609 & ~w15610;
assign w15621 = ~w15611 & ~w15612;
assign w15622 = ~w15613 & ~w15614;
assign w15623 = ~w15615 & ~w15616;
assign w15624 = w15622 & w15623;
assign w15625 = w15620 & w15621;
assign w15626 = w15618 & w15619;
assign w15627 = w15617 & w15626;
assign w15628 = w15624 & w15625;
assign w15629 = w15627 & w15628;
assign w15630 = w12993 & ~w15629;
assign w15631 = ~w15601 & ~w15602;
assign w15632 = ~w15630 & w15631;
assign w15633 = (~pi02678 & w14874) | (~pi02678 & w57377) | (w14874 & w57377);
assign w15634 = w14878 & w57378;
assign w15635 = ~pi10115 & w14909;
assign w15636 = ~pi10042 & w14893;
assign w15637 = ~pi01302 & w14896;
assign w15638 = ~pi10327 & w14907;
assign w15639 = ~pi01294 & w14889;
assign w15640 = ~pi10076 & w14891;
assign w15641 = ~pi10102 & w14901;
assign w15642 = ~pi10141 & w14903;
assign w15643 = ~pi10157 & w14886;
assign w15644 = ~pi10128 & w14911;
assign w15645 = ~pi02194 & w14881;
assign w15646 = ~pi10179 & w14884;
assign w15647 = ~pi01244 & w14899;
assign w15648 = ~pi01381 & w14905;
assign w15649 = ~w15635 & ~w15636;
assign w15650 = ~w15637 & ~w15638;
assign w15651 = ~w15639 & ~w15640;
assign w15652 = ~w15641 & ~w15642;
assign w15653 = ~w15643 & ~w15644;
assign w15654 = ~w15645 & ~w15646;
assign w15655 = ~w15647 & ~w15648;
assign w15656 = w15654 & w15655;
assign w15657 = w15652 & w15653;
assign w15658 = w15650 & w15651;
assign w15659 = w15649 & w15658;
assign w15660 = w15656 & w15657;
assign w15661 = w15659 & w15660;
assign w15662 = w12993 & ~w15661;
assign w15663 = ~w15633 & ~w15634;
assign w15664 = ~w15662 & w15663;
assign w15665 = (~pi02246 & w14874) | (~pi02246 & w57379) | (w14874 & w57379);
assign w15666 = w14878 & w57380;
assign w15667 = ~pi01229 & w14886;
assign w15668 = ~pi10280 & w14881;
assign w15669 = ~pi01397 & w14909;
assign w15670 = ~pi10129 & w14911;
assign w15671 = ~pi01356 & w14891;
assign w15672 = ~pi10262 & w14884;
assign w15673 = ~pi10228 & w14889;
assign w15674 = ~pi10192 & w14899;
assign w15675 = ~pi10103 & w14901;
assign w15676 = ~pi10213 & w14893;
assign w15677 = ~pi10090 & w14896;
assign w15678 = ~pi01382 & w14905;
assign w15679 = ~pi10065 & w14907;
assign w15680 = ~pi10142 & w14903;
assign w15681 = ~w15667 & ~w15668;
assign w15682 = ~w15669 & ~w15670;
assign w15683 = ~w15671 & ~w15672;
assign w15684 = ~w15673 & ~w15674;
assign w15685 = ~w15675 & ~w15676;
assign w15686 = ~w15677 & ~w15678;
assign w15687 = ~w15679 & ~w15680;
assign w15688 = w15686 & w15687;
assign w15689 = w15684 & w15685;
assign w15690 = w15682 & w15683;
assign w15691 = w15681 & w15690;
assign w15692 = w15688 & w15689;
assign w15693 = w15691 & w15692;
assign w15694 = w12993 & ~w15693;
assign w15695 = ~w15665 & ~w15666;
assign w15696 = ~w15694 & w15695;
assign w15697 = (~pi01346 & w14874) | (~pi01346 & w57381) | (w14874 & w57381);
assign w15698 = w14878 & w57382;
assign w15699 = ~pi10214 & w14893;
assign w15700 = ~pi01367 & w14901;
assign w15701 = ~pi01315 & w14907;
assign w15702 = ~pi10033 & w14889;
assign w15703 = ~pi01224 & w14896;
assign w15704 = ~pi01326 & w14884;
assign w15705 = ~pi01247 & w14899;
assign w15706 = ~pi10297 & w14903;
assign w15707 = ~pi01293 & w14891;
assign w15708 = ~pi10287 & w14886;
assign w15709 = ~pi01424 & w14881;
assign w15710 = ~pi10304 & w14909;
assign w15711 = ~pi01406 & w14911;
assign w15712 = ~pi01383 & w14905;
assign w15713 = ~w15699 & ~w15700;
assign w15714 = ~w15701 & ~w15702;
assign w15715 = ~w15703 & ~w15704;
assign w15716 = ~w15705 & ~w15706;
assign w15717 = ~w15707 & ~w15708;
assign w15718 = ~w15709 & ~w15710;
assign w15719 = ~w15711 & ~w15712;
assign w15720 = w15718 & w15719;
assign w15721 = w15716 & w15717;
assign w15722 = w15714 & w15715;
assign w15723 = w15713 & w15722;
assign w15724 = w15720 & w15721;
assign w15725 = w15723 & w15724;
assign w15726 = w12993 & ~w15725;
assign w15727 = ~w15697 & ~w15698;
assign w15728 = ~w15726 & w15727;
assign w15729 = (~pi02680 & w14874) | (~pi02680 & w57383) | (w14874 & w57383);
assign w15730 = w14878 & w57384;
assign w15731 = ~pi01445 & w14893;
assign w15732 = ~pi10077 & w14891;
assign w15733 = ~pi10180 & w14884;
assign w15734 = ~pi01398 & w14909;
assign w15735 = ~pi01407 & w14911;
assign w15736 = ~pi10091 & w14896;
assign w15737 = ~pi01328 & w14899;
assign w15738 = ~pi10168 & w14881;
assign w15739 = ~pi10143 & w14903;
assign w15740 = ~pi10340 & w14907;
assign w15741 = ~pi01321 & w14886;
assign w15742 = ~pi02688 & w14905;
assign w15743 = ~pi10229 & w14889;
assign w15744 = ~pi01368 & w14901;
assign w15745 = ~w15731 & ~w15732;
assign w15746 = ~w15733 & ~w15734;
assign w15747 = ~w15735 & ~w15736;
assign w15748 = ~w15737 & ~w15738;
assign w15749 = ~w15739 & ~w15740;
assign w15750 = ~w15741 & ~w15742;
assign w15751 = ~w15743 & ~w15744;
assign w15752 = w15750 & w15751;
assign w15753 = w15748 & w15749;
assign w15754 = w15746 & w15747;
assign w15755 = w15745 & w15754;
assign w15756 = w15752 & w15753;
assign w15757 = w15755 & w15756;
assign w15758 = w12993 & ~w15757;
assign w15759 = ~w15729 & ~w15730;
assign w15760 = ~w15758 & w15759;
assign w15761 = (~pi02679 & w14874) | (~pi02679 & w57385) | (w14874 & w57385);
assign w15762 = w14878 & w57386;
assign w15763 = ~pi01230 & w14886;
assign w15764 = ~pi10169 & w14881;
assign w15765 = ~pi01399 & w14909;
assign w15766 = ~pi10066 & w14907;
assign w15767 = ~pi10078 & w14891;
assign w15768 = ~pi10144 & w14903;
assign w15769 = ~pi10181 & w14884;
assign w15770 = ~pi10104 & w14901;
assign w15771 = ~pi10215 & w14893;
assign w15772 = ~pi01385 & w14905;
assign w15773 = ~pi01245 & w14899;
assign w15774 = ~pi01408 & w14911;
assign w15775 = ~pi01334 & w14889;
assign w15776 = ~pi10324 & w14896;
assign w15777 = ~w15763 & ~w15764;
assign w15778 = ~w15765 & ~w15766;
assign w15779 = ~w15767 & ~w15768;
assign w15780 = ~w15769 & ~w15770;
assign w15781 = ~w15771 & ~w15772;
assign w15782 = ~w15773 & ~w15774;
assign w15783 = ~w15775 & ~w15776;
assign w15784 = w15782 & w15783;
assign w15785 = w15780 & w15781;
assign w15786 = w15778 & w15779;
assign w15787 = w15777 & w15786;
assign w15788 = w15784 & w15785;
assign w15789 = w15787 & w15788;
assign w15790 = w12993 & ~w15789;
assign w15791 = ~w15761 & ~w15762;
assign w15792 = ~w15790 & w15791;
assign w15793 = (~pi01347 & w14874) | (~pi01347 & w57387) | (w14874 & w57387);
assign w15794 = w14878 & w57388;
assign w15795 = ~pi10182 & w14884;
assign w15796 = ~pi10145 & w14903;
assign w15797 = ~pi10158 & w14886;
assign w15798 = ~pi10067 & w14907;
assign w15799 = ~pi01319 & w14896;
assign w15800 = ~pi10286 & w14911;
assign w15801 = ~pi01425 & w14881;
assign w15802 = ~pi01286 & w14909;
assign w15803 = ~pi02687 & w14905;
assign w15804 = ~pi10333 & w14891;
assign w15805 = ~pi01246 & w14899;
assign w15806 = ~pi10035 & w14889;
assign w15807 = ~pi01369 & w14901;
assign w15808 = ~pi02695 & w14893;
assign w15809 = ~w15795 & ~w15796;
assign w15810 = ~w15797 & ~w15798;
assign w15811 = ~w15799 & ~w15800;
assign w15812 = ~w15801 & ~w15802;
assign w15813 = ~w15803 & ~w15804;
assign w15814 = ~w15805 & ~w15806;
assign w15815 = ~w15807 & ~w15808;
assign w15816 = w15814 & w15815;
assign w15817 = w15812 & w15813;
assign w15818 = w15810 & w15811;
assign w15819 = w15809 & w15818;
assign w15820 = w15816 & w15817;
assign w15821 = w15819 & w15820;
assign w15822 = w12993 & ~w15821;
assign w15823 = ~w15793 & ~w15794;
assign w15824 = ~w15822 & w15823;
assign w15825 = (~pi02238 & w14874) | (~pi02238 & w57389) | (w14874 & w57389);
assign w15826 = w14878 & w57390;
assign w15827 = ~pi01409 & w14911;
assign w15828 = ~pi10040 & w14893;
assign w15829 = ~pi10230 & w14889;
assign w15830 = ~pi01384 & w14905;
assign w15831 = ~pi10068 & w14907;
assign w15832 = ~pi10296 & w14903;
assign w15833 = ~pi01297 & w14899;
assign w15834 = ~pi10270 & w14884;
assign w15835 = ~pi01357 & w14891;
assign w15836 = ~pi10318 & w14901;
assign w15837 = ~pi10170 & w14881;
assign w15838 = ~pi10092 & w14896;
assign w15839 = ~pi10159 & w14886;
assign w15840 = ~pi10311 & w14909;
assign w15841 = ~w15827 & ~w15828;
assign w15842 = ~w15829 & ~w15830;
assign w15843 = ~w15831 & ~w15832;
assign w15844 = ~w15833 & ~w15834;
assign w15845 = ~w15835 & ~w15836;
assign w15846 = ~w15837 & ~w15838;
assign w15847 = ~w15839 & ~w15840;
assign w15848 = w15846 & w15847;
assign w15849 = w15844 & w15845;
assign w15850 = w15842 & w15843;
assign w15851 = w15841 & w15850;
assign w15852 = w15848 & w15849;
assign w15853 = w15851 & w15852;
assign w15854 = w12993 & ~w15853;
assign w15855 = ~w15825 & ~w15826;
assign w15856 = ~w15854 & w15855;
assign w15857 = (~pi02682 & w14874) | (~pi02682 & w57391) | (w14874 & w57391);
assign w15858 = w14878 & w57392;
assign w15859 = ~pi10216 & w14893;
assign w15860 = ~pi10325 & w14896;
assign w15861 = ~pi10110 & w14905;
assign w15862 = ~pi10310 & w14909;
assign w15863 = ~pi01231 & w14886;
assign w15864 = ~pi01235 & w14884;
assign w15865 = ~pi10105 & w14901;
assign w15866 = ~pi01335 & w14889;
assign w15867 = ~pi10146 & w14903;
assign w15868 = ~pi01248 & w14899;
assign w15869 = ~pi01426 & w14881;
assign w15870 = ~pi01284 & w14911;
assign w15871 = ~pi10339 & w14907;
assign w15872 = ~pi10079 & w14891;
assign w15873 = ~w15859 & ~w15860;
assign w15874 = ~w15861 & ~w15862;
assign w15875 = ~w15863 & ~w15864;
assign w15876 = ~w15865 & ~w15866;
assign w15877 = ~w15867 & ~w15868;
assign w15878 = ~w15869 & ~w15870;
assign w15879 = ~w15871 & ~w15872;
assign w15880 = w15878 & w15879;
assign w15881 = w15876 & w15877;
assign w15882 = w15874 & w15875;
assign w15883 = w15873 & w15882;
assign w15884 = w15880 & w15881;
assign w15885 = w15883 & w15884;
assign w15886 = w12993 & ~w15885;
assign w15887 = ~w15857 & ~w15858;
assign w15888 = ~w15886 & w15887;
assign w15889 = (~pi02681 & w14874) | (~pi02681 & w57393) | (w14874 & w57393);
assign w15890 = ~pi10203 & w14879;
assign w15891 = ~pi02226 & w14901;
assign w15892 = ~pi01358 & w14891;
assign w15893 = ~pi10160 & w14886;
assign w15894 = ~pi10093 & w14896;
assign w15895 = ~pi10183 & w14884;
assign w15896 = ~pi10130 & w14911;
assign w15897 = ~pi01446 & w14893;
assign w15898 = ~pi10193 & w14899;
assign w15899 = ~pi10034 & w14889;
assign w15900 = ~pi10288 & w14903;
assign w15901 = ~pi10069 & w14907;
assign w15902 = ~pi01400 & w14909;
assign w15903 = ~pi10315 & w14905;
assign w15904 = ~pi10277 & w14881;
assign w15905 = ~w15891 & ~w15892;
assign w15906 = ~w15893 & ~w15894;
assign w15907 = ~w15895 & ~w15896;
assign w15908 = ~w15897 & ~w15898;
assign w15909 = ~w15899 & ~w15900;
assign w15910 = ~w15901 & ~w15902;
assign w15911 = ~w15903 & ~w15904;
assign w15912 = w15910 & w15911;
assign w15913 = w15908 & w15909;
assign w15914 = w15906 & w15907;
assign w15915 = w15905 & w15914;
assign w15916 = w15912 & w15913;
assign w15917 = w15915 & w15916;
assign w15918 = w12993 & ~w15917;
assign w15919 = ~w15889 & ~w15890;
assign w15920 = ~w15918 & w15919;
assign w15921 = w538 & ~w574;
assign w15922 = pi01204 & ~w11337;
assign w15923 = ~w11338 & ~w15922;
assign w15924 = (pi09862 & ~w14191) | (pi09862 & w57394) | (~w14191 & w57394);
assign w15925 = w11341 & ~w14195;
assign w15926 = ~w15924 & w15925;
assign w15927 = ~w15923 & ~w15926;
assign w15928 = pi01205 & ~w11340;
assign w15929 = (pi01206 & ~w11335) | (pi01206 & w57395) | (~w11335 & w57395);
assign w15930 = ~w11337 & ~w15929;
assign w15931 = (pi09861 & ~w14191) | (pi09861 & w57396) | (~w14191 & w57396);
assign w15932 = w11341 & ~w14194;
assign w15933 = ~w15931 & w15932;
assign w15934 = ~w15930 & ~w15933;
assign w15935 = ~w12878 & w57397;
assign w15936 = ~pi01207 & w12884;
assign w15937 = ~w12879 & ~w12884;
assign w15938 = pi01207 & w15937;
assign w15939 = ~w15935 & ~w15936;
assign w15940 = ~w15938 & w15939;
assign w15941 = pi00869 & ~w1494;
assign w15942 = ~pi00869 & pi01208;
assign w15943 = ~w15941 & ~w15942;
assign w15944 = pi00870 & pi01463;
assign w15945 = w11149 & w15944;
assign w15946 = ~w12989 & w57398;
assign w15947 = w12984 & ~w12987;
assign w15948 = ~w12990 & ~w15946;
assign w15949 = (pi01209 & w12987) | (pi01209 & w57399) | (w12987 & w57399);
assign w15950 = ~w15948 & w15949;
assign w15951 = (w12993 & w15946) | (w12993 & w57400) | (w15946 & w57400);
assign w15952 = ~w15950 & w15951;
assign w15953 = (~pi01210 & ~w11340) | (~pi01210 & w57401) | (~w11340 & w57401);
assign w15954 = w14136 & w57402;
assign w15955 = ~pi00957 & w15954;
assign w15956 = ~w15953 & ~w15955;
assign w15957 = (~pi01211 & ~w11340) | (~pi01211 & w57403) | (~w11340 & w57403);
assign w15958 = w11340 & w57404;
assign w15959 = pi01213 & pi01275;
assign w15960 = w11340 & w57405;
assign w15961 = pi01308 & w15960;
assign w15962 = ~pi00957 & pi01305;
assign w15963 = pi01309 & w15962;
assign w15964 = w11356 & w15963;
assign w15965 = w15960 & w57406;
assign w15966 = ~w15957 & ~w15965;
assign w15967 = pi00869 & ~w1424;
assign w15968 = ~pi00869 & pi01212;
assign w15969 = ~w15967 & ~w15968;
assign w15970 = (~pi01213 & ~w11340) | (~pi01213 & w57407) | (~w11340 & w57407);
assign w15971 = w11340 & w57408;
assign w15972 = ~w15970 & ~w15971;
assign w15973 = (pi01214 & ~w11337) | (pi01214 & w57409) | (~w11337 & w57409);
assign w15974 = ~w11339 & ~w15973;
assign w15975 = pi09808 & ~w14195;
assign w15976 = w11341 & ~w14196;
assign w15977 = ~w15975 & w15976;
assign w15978 = ~w15974 & ~w15977;
assign w15979 = ~w12878 & w57410;
assign w15980 = (pi01215 & w12878) | (pi01215 & w57411) | (w12878 & w57411);
assign w15981 = ~w12886 & ~w15980;
assign w15982 = ~w12887 & ~w15981;
assign w15983 = ~w15979 & ~w15982;
assign w15984 = pi01216 & ~w11706;
assign w15985 = w1192 & ~w11709;
assign w15986 = ~w1192 & w11709;
assign w15987 = ~w15985 & ~w15986;
assign w15988 = w15984 & w15987;
assign w15989 = ~w15984 & ~w15987;
assign w15990 = ~w15988 & ~w15989;
assign w15991 = ~w12989 & w57412;
assign w15992 = w12989 & w57413;
assign w15993 = ~w15991 & ~w15992;
assign w15994 = ~w15993 & w57414;
assign w15995 = (~pi01217 & w15948) | (~pi01217 & w57415) | (w15948 & w57415);
assign w15996 = ~w15994 & w15995;
assign w15997 = ~w12989 & w15945;
assign w15998 = w12986 & w15947;
assign w15999 = ~w15997 & ~w15998;
assign w16000 = ~w12992 & ~w15999;
assign w16001 = w12993 & ~w16000;
assign w16002 = ~w15996 & w16001;
assign w16003 = pi09825 & ~pi09856;
assign w16004 = pi09855 & w12993;
assign w16005 = w14864 & w57416;
assign w16006 = w16003 & w16005;
assign w16007 = (pi01218 & ~w16005) | (pi01218 & w57417) | (~w16005 & w57417);
assign w16008 = w16005 & w57418;
assign w16009 = ~w16007 & ~w16008;
assign w16010 = (pi01219 & ~w16005) | (pi01219 & w57419) | (~w16005 & w57419);
assign w16011 = w16005 & w57420;
assign w16012 = ~w16010 & ~w16011;
assign w16013 = ~pi09825 & pi09856;
assign w16014 = w16005 & w16013;
assign w16015 = (pi01220 & ~w16005) | (pi01220 & w57421) | (~w16005 & w57421);
assign w16016 = w16005 & w57422;
assign w16017 = ~w16015 & ~w16016;
assign w16018 = (pi01221 & ~w16005) | (pi01221 & w57423) | (~w16005 & w57423);
assign w16019 = w16005 & w57424;
assign w16020 = ~w16018 & ~w16019;
assign w16021 = (pi01222 & ~w16005) | (pi01222 & w57425) | (~w16005 & w57425);
assign w16022 = w16005 & w57426;
assign w16023 = ~w16021 & ~w16022;
assign w16024 = (pi01223 & ~w16005) | (pi01223 & w57427) | (~w16005 & w57427);
assign w16025 = w16005 & w57428;
assign w16026 = ~w16024 & ~w16025;
assign w16027 = (pi01224 & ~w16005) | (pi01224 & w57429) | (~w16005 & w57429);
assign w16028 = w16005 & w57430;
assign w16029 = ~w16027 & ~w16028;
assign w16030 = pi01451 & w14864;
assign w16031 = w14864 & w57431;
assign w16032 = w16003 & w16031;
assign w16033 = (pi01225 & ~w16031) | (pi01225 & w57432) | (~w16031 & w57432);
assign w16034 = w16031 & w57433;
assign w16035 = ~w16033 & ~w16034;
assign w16036 = (pi01226 & ~w16031) | (pi01226 & w57434) | (~w16031 & w57434);
assign w16037 = w16031 & w57435;
assign w16038 = ~w16036 & ~w16037;
assign w16039 = (pi01227 & ~w16031) | (pi01227 & w57436) | (~w16031 & w57436);
assign w16040 = w16031 & w57437;
assign w16041 = ~w16039 & ~w16040;
assign w16042 = (pi01228 & ~w16031) | (pi01228 & w57438) | (~w16031 & w57438);
assign w16043 = w16031 & w57439;
assign w16044 = ~w16042 & ~w16043;
assign w16045 = (pi01229 & ~w16031) | (pi01229 & w57440) | (~w16031 & w57440);
assign w16046 = w16031 & w57441;
assign w16047 = ~w16045 & ~w16046;
assign w16048 = (pi01230 & ~w16031) | (pi01230 & w57442) | (~w16031 & w57442);
assign w16049 = w16031 & w57443;
assign w16050 = ~w16048 & ~w16049;
assign w16051 = (pi01231 & ~w16031) | (pi01231 & w57444) | (~w16031 & w57444);
assign w16052 = w16031 & w57445;
assign w16053 = ~w16051 & ~w16052;
assign w16054 = w16013 & w16031;
assign w16055 = (pi01232 & ~w16031) | (pi01232 & w57446) | (~w16031 & w57446);
assign w16056 = w16031 & w57447;
assign w16057 = ~w16055 & ~w16056;
assign w16058 = (pi01233 & ~w16031) | (pi01233 & w57448) | (~w16031 & w57448);
assign w16059 = w16031 & w57449;
assign w16060 = ~w16058 & ~w16059;
assign w16061 = (pi01234 & ~w16031) | (pi01234 & w57450) | (~w16031 & w57450);
assign w16062 = w16031 & w57451;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = (pi01235 & ~w16031) | (pi01235 & w57452) | (~w16031 & w57452);
assign w16065 = w16031 & w57453;
assign w16066 = ~w16064 & ~w16065;
assign w16067 = (pi01236 & ~w14865) | (pi01236 & w57454) | (~w14865 & w57454);
assign w16068 = w14865 & w57455;
assign w16069 = ~w16067 & ~w16068;
assign w16070 = (pi01237 & ~w14865) | (pi01237 & w57456) | (~w14865 & w57456);
assign w16071 = w14865 & w57457;
assign w16072 = ~w16070 & ~w16071;
assign w16073 = (pi01238 & ~w14865) | (pi01238 & w57458) | (~w14865 & w57458);
assign w16074 = w14865 & w57459;
assign w16075 = ~w16073 & ~w16074;
assign w16076 = (pi01239 & ~w14865) | (pi01239 & w57460) | (~w14865 & w57460);
assign w16077 = w14865 & w57461;
assign w16078 = ~w16076 & ~w16077;
assign w16079 = (pi01240 & ~w14865) | (pi01240 & w57462) | (~w14865 & w57462);
assign w16080 = w14865 & w57463;
assign w16081 = ~w16079 & ~w16080;
assign w16082 = (pi01241 & ~w14865) | (pi01241 & w57464) | (~w14865 & w57464);
assign w16083 = w14865 & w57465;
assign w16084 = ~w16082 & ~w16083;
assign w16085 = (pi01242 & ~w14865) | (pi01242 & w57466) | (~w14865 & w57466);
assign w16086 = w14865 & w57467;
assign w16087 = ~w16085 & ~w16086;
assign w16088 = (pi01243 & ~w14865) | (pi01243 & w57468) | (~w14865 & w57468);
assign w16089 = w14865 & w57469;
assign w16090 = ~w16088 & ~w16089;
assign w16091 = (pi01244 & ~w14865) | (pi01244 & w57470) | (~w14865 & w57470);
assign w16092 = w14865 & w57471;
assign w16093 = ~w16091 & ~w16092;
assign w16094 = (pi01245 & ~w14865) | (pi01245 & w57472) | (~w14865 & w57472);
assign w16095 = w14865 & w57473;
assign w16096 = ~w16094 & ~w16095;
assign w16097 = (pi01246 & ~w14865) | (pi01246 & w57474) | (~w14865 & w57474);
assign w16098 = w14865 & w57475;
assign w16099 = ~w16097 & ~w16098;
assign w16100 = (pi01247 & ~w14865) | (pi01247 & w57476) | (~w14865 & w57476);
assign w16101 = w14865 & w57477;
assign w16102 = ~w16100 & ~w16101;
assign w16103 = (pi01248 & ~w14865) | (pi01248 & w57478) | (~w14865 & w57478);
assign w16104 = w14865 & w57479;
assign w16105 = ~w16103 & ~w16104;
assign w16106 = (~pi01249 & ~w11340) | (~pi01249 & w57480) | (~w11340 & w57480);
assign w16107 = ~pi01306 & ~pi01309;
assign w16108 = w11368 & w16107;
assign w16109 = ~w16106 & ~w16108;
assign w16110 = pi00869 & ~w1417;
assign w16111 = ~pi00869 & pi01250;
assign w16112 = ~w16110 & ~w16111;
assign w16113 = (pi01251 & ~w11485) | (pi01251 & w57481) | (~w11485 & w57481);
assign w16114 = w11485 & w57482;
assign w16115 = ~w16113 & ~w16114;
assign w16116 = (pi01252 & ~w11485) | (pi01252 & w57483) | (~w11485 & w57483);
assign w16117 = w11485 & w57484;
assign w16118 = ~w16116 & ~w16117;
assign w16119 = (pi01253 & ~w11485) | (pi01253 & w57485) | (~w11485 & w57485);
assign w16120 = w11485 & w57486;
assign w16121 = ~w16119 & ~w16120;
assign w16122 = (pi01254 & ~w11485) | (pi01254 & w57487) | (~w11485 & w57487);
assign w16123 = w11485 & w57488;
assign w16124 = ~w16122 & ~w16123;
assign w16125 = (pi01255 & ~w11485) | (pi01255 & w57489) | (~w11485 & w57489);
assign w16126 = w11485 & w57490;
assign w16127 = ~w16125 & ~w16126;
assign w16128 = (pi01256 & ~w11485) | (pi01256 & w57491) | (~w11485 & w57491);
assign w16129 = w11485 & w57492;
assign w16130 = ~w16128 & ~w16129;
assign w16131 = (pi01257 & ~w11485) | (pi01257 & w57493) | (~w11485 & w57493);
assign w16132 = w11485 & w57494;
assign w16133 = ~w16131 & ~w16132;
assign w16134 = (pi01258 & ~w11485) | (pi01258 & w57495) | (~w11485 & w57495);
assign w16135 = w11485 & w57496;
assign w16136 = ~w16134 & ~w16135;
assign w16137 = (pi01259 & ~w11485) | (pi01259 & w57497) | (~w11485 & w57497);
assign w16138 = w11485 & w57498;
assign w16139 = ~w16137 & ~w16138;
assign w16140 = (pi01260 & ~w11485) | (pi01260 & w57499) | (~w11485 & w57499);
assign w16141 = w11485 & w57500;
assign w16142 = ~w16140 & ~w16141;
assign w16143 = w1209 & w57501;
assign w16144 = (~pi01261 & ~w16143) | (~pi01261 & w57502) | (~w16143 & w57502);
assign w16145 = w16143 & w57503;
assign w16146 = ~pi10351 & ~w16144;
assign w16147 = ~w16145 & w16146;
assign w16148 = ~pi01262 & w15993;
assign w16149 = (w12993 & w15993) | (w12993 & w57504) | (w15993 & w57504);
assign w16150 = ~w16148 & w16149;
assign w16151 = (pi01263 & ~w11485) | (pi01263 & w57505) | (~w11485 & w57505);
assign w16152 = w11485 & w57506;
assign w16153 = ~w16151 & ~w16152;
assign w16154 = (pi01264 & ~w11485) | (pi01264 & w57507) | (~w11485 & w57507);
assign w16155 = w11485 & w57508;
assign w16156 = ~w16154 & ~w16155;
assign w16157 = (pi01265 & ~w11485) | (pi01265 & w57509) | (~w11485 & w57509);
assign w16158 = w11485 & w57510;
assign w16159 = ~w16157 & ~w16158;
assign w16160 = (pi01266 & ~w11485) | (pi01266 & w57511) | (~w11485 & w57511);
assign w16161 = w11485 & w57512;
assign w16162 = ~w16160 & ~w16161;
assign w16163 = (pi01267 & ~w11485) | (pi01267 & w57513) | (~w11485 & w57513);
assign w16164 = w11485 & w57514;
assign w16165 = ~w16163 & ~w16164;
assign w16166 = (pi01268 & ~w11485) | (pi01268 & w57515) | (~w11485 & w57515);
assign w16167 = w11485 & w57516;
assign w16168 = ~w16166 & ~w16167;
assign w16169 = (pi01269 & ~w11485) | (pi01269 & w57517) | (~w11485 & w57517);
assign w16170 = w11485 & w57518;
assign w16171 = ~w16169 & ~w16170;
assign w16172 = ~pi10366 & pi10518;
assign w16173 = pi00845 & ~w11126;
assign w16174 = ~w11126 & w57519;
assign w16175 = (pi01270 & w11126) | (pi01270 & w57520) | (w11126 & w57520);
assign w16176 = ~w11180 & ~w16174;
assign w16177 = ~w16175 & w16176;
assign w16178 = ~w11193 & w16172;
assign w16179 = ~w16177 & w16178;
assign w16180 = (pi01271 & w11126) | (pi01271 & w57521) | (w11126 & w57521);
assign w16181 = ~w11176 & ~w11182;
assign w16182 = w16173 & w16181;
assign w16183 = ~w11193 & ~w16180;
assign w16184 = ~w16182 & w16183;
assign w16185 = (w16172 & ~w11193) | (w16172 & w57522) | (~w11193 & w57522);
assign w16186 = ~w16184 & w16185;
assign w16187 = pi01273 & ~w11160;
assign w16188 = pi00034 & pi00036;
assign w16189 = pi10375 & ~w16188;
assign w16190 = w13021 & w16189;
assign w16191 = ~w16187 & ~w16190;
assign w16192 = pi01216 & pi01450;
assign w16193 = (~w16192 & w11709) | (~w16192 & w57523) | (w11709 & w57523);
assign w16194 = (~w10686 & ~w11709) | (~w10686 & w57524) | (~w11709 & w57524);
assign w16195 = ~w16193 & ~w16194;
assign w16196 = (~w15985 & ~w16195) | (~w15985 & w57525) | (~w16195 & w57525);
assign w16197 = pi01312 & ~w1192;
assign w16198 = ~w10688 & ~w16197;
assign w16199 = (~pi01274 & w16196) | (~pi01274 & w57526) | (w16196 & w57526);
assign w16200 = ~w16196 & w57527;
assign w16201 = ~w11706 & ~w16199;
assign w16202 = ~w16200 & w16201;
assign w16203 = (pi01275 & ~w11340) | (pi01275 & w57528) | (~w11340 & w57528);
assign w16204 = ~w11346 & ~w15959;
assign w16205 = w11340 & w57529;
assign w16206 = ~w16203 & ~w16205;
assign w16207 = w671 & ~w805;
assign w16208 = (w12833 & ~w141) | (w12833 & w57530) | (~w141 & w57530);
assign w16209 = w2432 & ~w16208;
assign w16210 = (pi01278 & ~w11485) | (pi01278 & w57531) | (~w11485 & w57531);
assign w16211 = w11485 & w57532;
assign w16212 = ~w16210 & ~w16211;
assign w16213 = w14864 & w57533;
assign w16214 = w16003 & w16213;
assign w16215 = (pi01279 & ~w16213) | (pi01279 & w57534) | (~w16213 & w57534);
assign w16216 = w16213 & w57439;
assign w16217 = ~w16215 & ~w16216;
assign w16218 = ~pi09825 & ~pi09856;
assign w16219 = w16005 & w16218;
assign w16220 = (pi01280 & ~w16005) | (pi01280 & w57535) | (~w16005 & w57535);
assign w16221 = w16005 & w57536;
assign w16222 = ~w16220 & ~w16221;
assign w16223 = w14864 & w57537;
assign w16224 = w14864 & w57538;
assign w16225 = w14864 & w57539;
assign w16226 = pi01281 & ~w16225;
assign w16227 = ~pi10633 & w16225;
assign w16228 = ~w16226 & ~w16227;
assign w16229 = w14865 & w16013;
assign w16230 = (pi01282 & ~w14865) | (pi01282 & w57540) | (~w14865 & w57540);
assign w16231 = w14865 & w57541;
assign w16232 = ~w16230 & ~w16231;
assign w16233 = w14865 & w16003;
assign w16234 = (pi01283 & ~w14865) | (pi01283 & w57542) | (~w14865 & w57542);
assign w16235 = w14865 & w57543;
assign w16236 = ~w16234 & ~w16235;
assign w16237 = w16031 & w16218;
assign w16238 = (pi01284 & ~w16031) | (pi01284 & w57544) | (~w16031 & w57544);
assign w16239 = w16031 & w57545;
assign w16240 = ~w16238 & ~w16239;
assign w16241 = (pi01285 & ~w16031) | (pi01285 & w57546) | (~w16031 & w57546);
assign w16242 = w16031 & w57547;
assign w16243 = ~w16241 & ~w16242;
assign w16244 = w14861 & w16213;
assign w16245 = (pi01286 & ~w16213) | (pi01286 & w57548) | (~w16213 & w57548);
assign w16246 = w16213 & w57475;
assign w16247 = ~w16245 & ~w16246;
assign w16248 = (pi01287 & ~w16213) | (pi01287 & w57549) | (~w16213 & w57549);
assign w16249 = w16213 & w57550;
assign w16250 = ~w16248 & ~w16249;
assign w16251 = w14861 & w16005;
assign w16252 = (pi01288 & ~w16005) | (pi01288 & w57551) | (~w16005 & w57551);
assign w16253 = w16005 & w57550;
assign w16254 = ~w16252 & ~w16253;
assign w16255 = (pi01289 & ~w16213) | (pi01289 & w57552) | (~w16213 & w57552);
assign w16256 = w16213 & w57553;
assign w16257 = ~w16255 & ~w16256;
assign w16258 = (pi01290 & ~w16005) | (pi01290 & w57554) | (~w16005 & w57554);
assign w16259 = w16005 & w57555;
assign w16260 = ~w16258 & ~w16259;
assign w16261 = w16013 & w16213;
assign w16262 = (pi01291 & ~w16213) | (pi01291 & w57556) | (~w16213 & w57556);
assign w16263 = w16213 & w57557;
assign w16264 = ~w16262 & ~w16263;
assign w16265 = (pi01292 & ~w16213) | (pi01292 & w57558) | (~w16213 & w57558);
assign w16266 = w16213 & w57559;
assign w16267 = ~w16265 & ~w16266;
assign w16268 = (pi01293 & ~w16213) | (pi01293 & w57560) | (~w16213 & w57560);
assign w16269 = w16213 & w57561;
assign w16270 = ~w16268 & ~w16269;
assign w16271 = w16213 & w16218;
assign w16272 = (pi01294 & ~w16213) | (pi01294 & w57562) | (~w16213 & w57562);
assign w16273 = w16213 & w57563;
assign w16274 = ~w16272 & ~w16273;
assign w16275 = (pi01295 & ~w16213) | (pi01295 & w57564) | (~w16213 & w57564);
assign w16276 = w16213 & w57565;
assign w16277 = ~w16275 & ~w16276;
assign w16278 = (pi01296 & ~w14865) | (pi01296 & w57566) | (~w14865 & w57566);
assign w16279 = w14865 & w57567;
assign w16280 = ~w16278 & ~w16279;
assign w16281 = (pi01297 & ~w14865) | (pi01297 & w57568) | (~w14865 & w57568);
assign w16282 = w14865 & w57569;
assign w16283 = ~w16281 & ~w16282;
assign w16284 = (pi01298 & ~w14865) | (pi01298 & w57570) | (~w14865 & w57570);
assign w16285 = w14865 & w57571;
assign w16286 = ~w16284 & ~w16285;
assign w16287 = (pi01299 & ~w16031) | (pi01299 & w57572) | (~w16031 & w57572);
assign w16288 = w16031 & w57420;
assign w16289 = ~w16287 & ~w16288;
assign w16290 = (pi01300 & ~w16031) | (pi01300 & w57573) | (~w16031 & w57573);
assign w16291 = w16031 & w57574;
assign w16292 = ~w16290 & ~w16291;
assign w16293 = (pi01301 & ~w16031) | (pi01301 & w57575) | (~w16031 & w57575);
assign w16294 = w16031 & w57576;
assign w16295 = ~w16293 & ~w16294;
assign w16296 = (pi01302 & ~w16005) | (pi01302 & w57577) | (~w16005 & w57577);
assign w16297 = w16005 & w57578;
assign w16298 = ~w16296 & ~w16297;
assign w16299 = pi10423 & w12844;
assign w16300 = (pi01303 & ~w523) | (pi01303 & w57579) | (~w523 & w57579);
assign w16301 = pi01252 & pi10376;
assign w16302 = w523 & w57580;
assign w16303 = ~w16300 & ~w16302;
assign w16304 = ~w12878 & w57581;
assign w16305 = (~pi01304 & ~w12881) | (~pi01304 & w57582) | (~w12881 & w57582);
assign w16306 = w15937 & ~w16305;
assign w16307 = ~w16304 & ~w16306;
assign w16308 = ~w14137 & ~w15961;
assign w16309 = (pi01307 & w15961) | (pi01307 & w57583) | (w15961 & w57583);
assign w16310 = (~pi01305 & ~w16309) | (~pi01305 & w57584) | (~w16309 & w57584);
assign w16311 = ~w14137 & ~w14149;
assign w16312 = ~w16310 & w16311;
assign w16313 = (pi01306 & ~w11340) | (pi01306 & w57585) | (~w11340 & w57585);
assign w16314 = ~w14150 & w16313;
assign w16315 = ~w15954 & ~w16314;
assign w16316 = (~pi01307 & ~w15960) | (~pi01307 & w57586) | (~w15960 & w57586);
assign w16317 = ~w16309 & ~w16316;
assign w16318 = ~pi01308 & ~w15960;
assign w16319 = w16308 & ~w16318;
assign w16320 = w11355 & w57587;
assign w16321 = ~w14148 & ~w16320;
assign w16322 = w15958 & ~w16321;
assign w16323 = ~pi01309 & ~w16322;
assign w16324 = (pi01309 & w14149) | (pi01309 & w57588) | (w14149 & w57588);
assign w16325 = ~w16323 & ~w16324;
assign w16326 = (pi01310 & ~w11340) | (pi01310 & w57589) | (~w11340 & w57589);
assign w16327 = ~w15958 & ~w16326;
assign w16328 = ~w12878 & w57590;
assign w16329 = (pi01311 & w12878) | (pi01311 & w57591) | (w12878 & w57591);
assign w16330 = ~w12885 & ~w16329;
assign w16331 = ~w12886 & ~w16330;
assign w16332 = ~w16328 & ~w16331;
assign w16333 = w1192 & ~w10687;
assign w16334 = (~pi01312 & w16196) | (~pi01312 & w57592) | (w16196 & w57592);
assign w16335 = ~w16196 & w57593;
assign w16336 = ~w11706 & ~w16334;
assign w16337 = ~w16335 & w16336;
assign w16338 = (pi01313 & ~w16005) | (pi01313 & w57594) | (~w16005 & w57594);
assign w16339 = w16005 & w57595;
assign w16340 = ~w16338 & ~w16339;
assign w16341 = (pi01314 & ~w16005) | (pi01314 & w57596) | (~w16005 & w57596);
assign w16342 = w16005 & w57439;
assign w16343 = ~w16341 & ~w16342;
assign w16344 = (pi01315 & ~w16005) | (pi01315 & w57597) | (~w16005 & w57597);
assign w16345 = w16005 & w57561;
assign w16346 = ~w16344 & ~w16345;
assign w16347 = (pi01316 & ~w16005) | (pi01316 & w57598) | (~w16005 & w57598);
assign w16348 = w16005 & w57599;
assign w16349 = ~w16347 & ~w16348;
assign w16350 = (pi01317 & ~w16005) | (pi01317 & w57600) | (~w16005 & w57600);
assign w16351 = w16005 & w57601;
assign w16352 = ~w16350 & ~w16351;
assign w16353 = (pi01318 & ~w16005) | (pi01318 & w57602) | (~w16005 & w57602);
assign w16354 = w16005 & w57603;
assign w16355 = ~w16353 & ~w16354;
assign w16356 = (pi01319 & ~w16005) | (pi01319 & w57604) | (~w16005 & w57604);
assign w16357 = w16005 & w57605;
assign w16358 = ~w16356 & ~w16357;
assign w16359 = (pi01320 & ~w16031) | (pi01320 & w57606) | (~w16031 & w57606);
assign w16360 = w16031 & w57607;
assign w16361 = ~w16359 & ~w16360;
assign w16362 = (pi01321 & ~w16031) | (pi01321 & w57608) | (~w16031 & w57608);
assign w16363 = w16031 & w57609;
assign w16364 = ~w16362 & ~w16363;
assign w16365 = (pi01322 & ~w16031) | (pi01322 & w57610) | (~w16031 & w57610);
assign w16366 = w16031 & w57426;
assign w16367 = ~w16365 & ~w16366;
assign w16368 = (pi01323 & ~w16031) | (pi01323 & w57611) | (~w16031 & w57611);
assign w16369 = w16031 & w57612;
assign w16370 = ~w16368 & ~w16369;
assign w16371 = (pi01324 & ~w16031) | (pi01324 & w57613) | (~w16031 & w57613);
assign w16372 = w16031 & w57428;
assign w16373 = ~w16371 & ~w16372;
assign w16374 = (pi01325 & ~w16031) | (pi01325 & w57614) | (~w16031 & w57614);
assign w16375 = w16031 & w57615;
assign w16376 = ~w16374 & ~w16375;
assign w16377 = (pi01326 & ~w16031) | (pi01326 & w57616) | (~w16031 & w57616);
assign w16378 = w16031 & w57430;
assign w16379 = ~w16377 & ~w16378;
assign w16380 = (pi01327 & ~w16031) | (pi01327 & w57617) | (~w16031 & w57617);
assign w16381 = w16031 & w57603;
assign w16382 = ~w16380 & ~w16381;
assign w16383 = (pi01328 & ~w14865) | (pi01328 & w57618) | (~w14865 & w57618);
assign w16384 = w14865 & w57619;
assign w16385 = ~w16383 & ~w16384;
assign w16386 = (pi01329 & ~w16213) | (pi01329 & w57620) | (~w16213 & w57620);
assign w16387 = w16213 & w57621;
assign w16388 = ~w16386 & ~w16387;
assign w16389 = (pi01330 & ~w16213) | (pi01330 & w57622) | (~w16213 & w57622);
assign w16390 = w16213 & w57623;
assign w16391 = ~w16389 & ~w16390;
assign w16392 = (pi01331 & ~w16213) | (pi01331 & w57624) | (~w16213 & w57624);
assign w16393 = w16213 & w57625;
assign w16394 = ~w16392 & ~w16393;
assign w16395 = (pi01332 & ~w16213) | (pi01332 & w57626) | (~w16213 & w57626);
assign w16396 = w16213 & w57627;
assign w16397 = ~w16395 & ~w16396;
assign w16398 = (pi01333 & ~w16213) | (pi01333 & w57628) | (~w16213 & w57628);
assign w16399 = w16213 & w57629;
assign w16400 = ~w16398 & ~w16399;
assign w16401 = (pi01334 & ~w16213) | (pi01334 & w57630) | (~w16213 & w57630);
assign w16402 = w16213 & w57631;
assign w16403 = ~w16401 & ~w16402;
assign w16404 = (pi01335 & ~w16213) | (pi01335 & w57632) | (~w16213 & w57632);
assign w16405 = w16213 & w57545;
assign w16406 = ~w16404 & ~w16405;
assign w16407 = w1789 & ~w12993;
assign w16408 = (~w16407 & ~w14865) | (~w16407 & w57633) | (~w14865 & w57633);
assign w16409 = pi10633 & ~w16408;
assign w16410 = (~w14865 & w57634) | (~w14865 & w57635) | (w57634 & w57635);
assign w16411 = ~w16409 & ~w16410;
assign w16412 = (w14865 & w57636) | (w14865 & w57637) | (w57636 & w57637);
assign w16413 = (~w14865 & w57638) | (~w14865 & w57639) | (w57638 & w57639);
assign w16414 = ~w16412 & ~w16413;
assign w16415 = (w14865 & w57640) | (w14865 & w57641) | (w57640 & w57641);
assign w16416 = (~w14865 & w57642) | (~w14865 & w57643) | (w57642 & w57643);
assign w16417 = ~w16415 & ~w16416;
assign w16418 = (w14865 & w57644) | (w14865 & w57645) | (w57644 & w57645);
assign w16419 = (~w14865 & w57646) | (~w14865 & w57647) | (w57646 & w57647);
assign w16420 = ~w16418 & ~w16419;
assign w16421 = (w14865 & w57648) | (w14865 & w57649) | (w57648 & w57649);
assign w16422 = (~w14865 & w57650) | (~w14865 & w57651) | (w57650 & w57651);
assign w16423 = ~w16421 & ~w16422;
assign w16424 = (w14865 & w57652) | (w14865 & w57653) | (w57652 & w57653);
assign w16425 = (~w14865 & w57654) | (~w14865 & w57655) | (w57654 & w57655);
assign w16426 = ~w16424 & ~w16425;
assign w16427 = (w14865 & w57656) | (w14865 & w57657) | (w57656 & w57657);
assign w16428 = (~w14865 & w57658) | (~w14865 & w57659) | (w57658 & w57659);
assign w16429 = ~w16427 & ~w16428;
assign w16430 = (w14865 & w57660) | (w14865 & w57661) | (w57660 & w57661);
assign w16431 = (~w14865 & w57662) | (~w14865 & w57663) | (w57662 & w57663);
assign w16432 = ~w16430 & ~w16431;
assign w16433 = (w14865 & w57664) | (w14865 & w57665) | (w57664 & w57665);
assign w16434 = (~w14865 & w57666) | (~w14865 & w57667) | (w57666 & w57667);
assign w16435 = ~w16433 & ~w16434;
assign w16436 = (w14865 & w57668) | (w14865 & w57669) | (w57668 & w57669);
assign w16437 = (~w14865 & w57670) | (~w14865 & w57671) | (w57670 & w57671);
assign w16438 = ~w16436 & ~w16437;
assign w16439 = (w14865 & w57672) | (w14865 & w57673) | (w57672 & w57673);
assign w16440 = (~w14865 & w57674) | (~w14865 & w57675) | (w57674 & w57675);
assign w16441 = ~w16439 & ~w16440;
assign w16442 = (w14865 & w57676) | (w14865 & w57677) | (w57676 & w57677);
assign w16443 = (~w14865 & w57678) | (~w14865 & w57679) | (w57678 & w57679);
assign w16444 = ~w16442 & ~w16443;
assign w16445 = (pi01348 & ~w16213) | (pi01348 & w57680) | (~w16213 & w57680);
assign w16446 = w16213 & w57437;
assign w16447 = ~w16445 & ~w16446;
assign w16448 = (pi01349 & ~w16213) | (pi01349 & w57681) | (~w16213 & w57681);
assign w16449 = w16213 & w57595;
assign w16450 = ~w16448 & ~w16449;
assign w16451 = (pi01350 & ~w16213) | (pi01350 & w57682) | (~w16213 & w57682);
assign w16452 = w16213 & w57683;
assign w16453 = ~w16451 & ~w16452;
assign w16454 = (pi01351 & ~w16213) | (pi01351 & w57684) | (~w16213 & w57684);
assign w16455 = w16213 & w57685;
assign w16456 = ~w16454 & ~w16455;
assign w16457 = (pi01352 & ~w16213) | (pi01352 & w57686) | (~w16213 & w57686);
assign w16458 = w16213 & w57687;
assign w16459 = ~w16457 & ~w16458;
assign w16460 = (pi01353 & ~w16213) | (pi01353 & w57688) | (~w16213 & w57688);
assign w16461 = w16213 & w57607;
assign w16462 = ~w16460 & ~w16461;
assign w16463 = (pi01354 & ~w16213) | (pi01354 & w57689) | (~w16213 & w57689);
assign w16464 = w16213 & w57690;
assign w16465 = ~w16463 & ~w16464;
assign w16466 = (pi01355 & ~w16213) | (pi01355 & w57691) | (~w16213 & w57691);
assign w16467 = w16213 & w57692;
assign w16468 = ~w16466 & ~w16467;
assign w16469 = (pi01356 & ~w16213) | (pi01356 & w57693) | (~w16213 & w57693);
assign w16470 = w16213 & w57441;
assign w16471 = ~w16469 & ~w16470;
assign w16472 = (pi01357 & ~w16213) | (pi01357 & w57694) | (~w16213 & w57694);
assign w16473 = w16213 & w57695;
assign w16474 = ~w16472 & ~w16473;
assign w16475 = (pi01358 & ~w16213) | (pi01358 & w57696) | (~w16213 & w57696);
assign w16476 = w16213 & w57697;
assign w16477 = ~w16475 & ~w16476;
assign w16478 = (pi01359 & ~w16213) | (pi01359 & w57698) | (~w16213 & w57698);
assign w16479 = w16213 & w57699;
assign w16480 = ~w16478 & ~w16479;
assign w16481 = (pi01360 & ~w16213) | (pi01360 & w57700) | (~w16213 & w57700);
assign w16482 = w16213 & w57612;
assign w16483 = ~w16481 & ~w16482;
assign w16484 = (pi01361 & ~w16213) | (pi01361 & w57701) | (~w16213 & w57701);
assign w16485 = w16213 & w57424;
assign w16486 = ~w16484 & ~w16485;
assign w16487 = (pi01362 & ~w16213) | (pi01362 & w57702) | (~w16213 & w57702);
assign w16488 = w16213 & w57703;
assign w16489 = ~w16487 & ~w16488;
assign w16490 = (pi01363 & ~w16213) | (pi01363 & w57704) | (~w16213 & w57704);
assign w16491 = w16213 & w57541;
assign w16492 = ~w16490 & ~w16491;
assign w16493 = (pi01364 & ~w16213) | (pi01364 & w57705) | (~w16213 & w57705);
assign w16494 = w16213 & w57615;
assign w16495 = ~w16493 & ~w16494;
assign w16496 = (pi01365 & ~w16213) | (pi01365 & w57706) | (~w16213 & w57706);
assign w16497 = w16213 & w57601;
assign w16498 = ~w16496 & ~w16497;
assign w16499 = (pi01366 & ~w16213) | (pi01366 & w57707) | (~w16213 & w57707);
assign w16500 = w16213 & w57708;
assign w16501 = ~w16499 & ~w16500;
assign w16502 = (pi01367 & ~w16213) | (pi01367 & w57709) | (~w16213 & w57709);
assign w16503 = w16213 & w57430;
assign w16504 = ~w16502 & ~w16503;
assign w16505 = (pi01368 & ~w16213) | (pi01368 & w57710) | (~w16213 & w57710);
assign w16506 = w16213 & w57711;
assign w16507 = ~w16505 & ~w16506;
assign w16508 = (pi01369 & ~w16213) | (pi01369 & w57712) | (~w16213 & w57712);
assign w16509 = w16213 & w57605;
assign w16510 = ~w16508 & ~w16509;
assign w16511 = (pi01370 & ~w16005) | (pi01370 & w57713) | (~w16005 & w57713);
assign w16512 = w16005 & w57714;
assign w16513 = ~w16511 & ~w16512;
assign w16514 = (pi01371 & ~w16005) | (pi01371 & w57715) | (~w16005 & w57715);
assign w16515 = w16005 & w57571;
assign w16516 = ~w16514 & ~w16515;
assign w16517 = (pi01372 & ~w16005) | (pi01372 & w57716) | (~w16005 & w57716);
assign w16518 = w16005 & w57455;
assign w16519 = ~w16517 & ~w16518;
assign w16520 = (pi01373 & ~w16005) | (pi01373 & w57717) | (~w16005 & w57717);
assign w16521 = w16005 & w57718;
assign w16522 = ~w16520 & ~w16521;
assign w16523 = (pi01374 & ~w16005) | (pi01374 & w57719) | (~w16005 & w57719);
assign w16524 = w16005 & w57720;
assign w16525 = ~w16523 & ~w16524;
assign w16526 = (pi01375 & ~w16005) | (pi01375 & w57721) | (~w16005 & w57721);
assign w16527 = w16005 & w57461;
assign w16528 = ~w16526 & ~w16527;
assign w16529 = (pi01376 & ~w16005) | (pi01376 & w57722) | (~w16005 & w57722);
assign w16530 = w16005 & w57723;
assign w16531 = ~w16529 & ~w16530;
assign w16532 = (pi01377 & ~w16005) | (pi01377 & w57724) | (~w16005 & w57724);
assign w16533 = w16005 & w57465;
assign w16534 = ~w16532 & ~w16533;
assign w16535 = (pi01378 & ~w16005) | (pi01378 & w57725) | (~w16005 & w57725);
assign w16536 = w16005 & w57329;
assign w16537 = ~w16535 & ~w16536;
assign w16538 = (pi01379 & ~w16005) | (pi01379 & w57726) | (~w16005 & w57726);
assign w16539 = w16005 & w57469;
assign w16540 = ~w16538 & ~w16539;
assign w16541 = (pi01380 & ~w16005) | (pi01380 & w57727) | (~w16005 & w57727);
assign w16542 = w16005 & w57728;
assign w16543 = ~w16541 & ~w16542;
assign w16544 = (pi01381 & ~w16005) | (pi01381 & w57729) | (~w16005 & w57729);
assign w16545 = w16005 & w57471;
assign w16546 = ~w16544 & ~w16545;
assign w16547 = (pi01382 & ~w16005) | (pi01382 & w57730) | (~w16005 & w57730);
assign w16548 = w16005 & w57731;
assign w16549 = ~w16547 & ~w16548;
assign w16550 = (pi01383 & ~w16005) | (pi01383 & w57732) | (~w16005 & w57732);
assign w16551 = w16005 & w57477;
assign w16552 = ~w16550 & ~w16551;
assign w16553 = (pi01384 & ~w16005) | (pi01384 & w57733) | (~w16005 & w57733);
assign w16554 = w16005 & w57569;
assign w16555 = ~w16553 & ~w16554;
assign w16556 = (pi01385 & ~w16005) | (pi01385 & w57734) | (~w16005 & w57734);
assign w16557 = w16005 & w57473;
assign w16558 = ~w16556 & ~w16557;
assign w16559 = (pi01386 & ~w16213) | (pi01386 & w57735) | (~w16213 & w57735);
assign w16560 = w16213 & w57455;
assign w16561 = ~w16559 & ~w16560;
assign w16562 = (pi01387 & ~w16213) | (pi01387 & w57736) | (~w16213 & w57736);
assign w16563 = w16213 & w57718;
assign w16564 = ~w16562 & ~w16563;
assign w16565 = (pi01388 & ~w16213) | (pi01388 & w57737) | (~w16213 & w57737);
assign w16566 = w16213 & w57457;
assign w16567 = ~w16565 & ~w16566;
assign w16568 = (pi01389 & ~w16213) | (pi01389 & w57738) | (~w16213 & w57738);
assign w16569 = w16213 & w57720;
assign w16570 = ~w16568 & ~w16569;
assign w16571 = (pi01390 & ~w16213) | (pi01390 & w57739) | (~w16213 & w57739);
assign w16572 = w16213 & w57740;
assign w16573 = ~w16571 & ~w16572;
assign w16574 = (pi01391 & ~w16213) | (pi01391 & w57741) | (~w16213 & w57741);
assign w16575 = w16213 & w57742;
assign w16576 = ~w16574 & ~w16575;
assign w16577 = (pi01392 & ~w16213) | (pi01392 & w57743) | (~w16213 & w57743);
assign w16578 = w16213 & w57461;
assign w16579 = ~w16577 & ~w16578;
assign w16580 = (pi01393 & ~w16213) | (pi01393 & w57744) | (~w16213 & w57744);
assign w16581 = w16213 & w57463;
assign w16582 = ~w16580 & ~w16581;
assign w16583 = (pi01394 & ~w16213) | (pi01394 & w57745) | (~w16213 & w57745);
assign w16584 = w16213 & w57723;
assign w16585 = ~w16583 & ~w16584;
assign w16586 = (pi01395 & ~w16213) | (pi01395 & w57746) | (~w16213 & w57746);
assign w16587 = w16213 & w57459;
assign w16588 = ~w16586 & ~w16587;
assign w16589 = (pi01396 & ~w16213) | (pi01396 & w57747) | (~w16213 & w57747);
assign w16590 = w16213 & w57728;
assign w16591 = ~w16589 & ~w16590;
assign w16592 = (pi01397 & ~w16213) | (pi01397 & w57748) | (~w16213 & w57748);
assign w16593 = w16213 & w57731;
assign w16594 = ~w16592 & ~w16593;
assign w16595 = (pi01398 & ~w16213) | (pi01398 & w57749) | (~w16213 & w57749);
assign w16596 = w16213 & w57619;
assign w16597 = ~w16595 & ~w16596;
assign w16598 = (pi01399 & ~w16213) | (pi01399 & w57750) | (~w16213 & w57750);
assign w16599 = w16213 & w57473;
assign w16600 = ~w16598 & ~w16599;
assign w16601 = (pi01400 & ~w16213) | (pi01400 & w57751) | (~w16213 & w57751);
assign w16602 = w16213 & w57752;
assign w16603 = ~w16601 & ~w16602;
assign w16604 = (pi01401 & ~w16031) | (pi01401 & w57753) | (~w16031 & w57753);
assign w16605 = w16031 & w57754;
assign w16606 = ~w16604 & ~w16605;
assign w16607 = (pi01402 & ~w16031) | (pi01402 & w57755) | (~w16031 & w57755);
assign w16608 = w16031 & w57565;
assign w16609 = ~w16607 & ~w16608;
assign w16610 = (pi01403 & ~w16031) | (pi01403 & w57756) | (~w16031 & w57756);
assign w16611 = w16031 & w57629;
assign w16612 = ~w16610 & ~w16611;
assign w16613 = (pi01404 & ~w16031) | (pi01404 & w57757) | (~w16031 & w57757);
assign w16614 = w16031 & w57627;
assign w16615 = ~w16613 & ~w16614;
assign w16616 = (pi01405 & ~w16031) | (pi01405 & w57758) | (~w16031 & w57758);
assign w16617 = w16031 & w57759;
assign w16618 = ~w16616 & ~w16617;
assign w16619 = (pi01406 & ~w16031) | (pi01406 & w57760) | (~w16031 & w57760);
assign w16620 = w16031 & w57761;
assign w16621 = ~w16619 & ~w16620;
assign w16622 = (pi01407 & ~w16031) | (pi01407 & w57762) | (~w16031 & w57762);
assign w16623 = w16031 & w57763;
assign w16624 = ~w16622 & ~w16623;
assign w16625 = (pi01408 & ~w16031) | (pi01408 & w57764) | (~w16031 & w57764);
assign w16626 = w16031 & w57631;
assign w16627 = ~w16625 & ~w16626;
assign w16628 = (pi01409 & ~w16031) | (pi01409 & w57765) | (~w16031 & w57765);
assign w16629 = w16031 & w57766;
assign w16630 = ~w16628 & ~w16629;
assign w16631 = (pi01410 & ~w14865) | (pi01410 & w57767) | (~w14865 & w57767);
assign w16632 = w14865 & w57685;
assign w16633 = ~w16631 & ~w16632;
assign w16634 = (pi01411 & ~w14865) | (pi01411 & w57768) | (~w14865 & w57768);
assign w16635 = w14865 & w57687;
assign w16636 = ~w16634 & ~w16635;
assign w16637 = (pi01412 & ~w14865) | (pi01412 & w57769) | (~w14865 & w57769);
assign w16638 = w14865 & w57683;
assign w16639 = ~w16637 & ~w16638;
assign w16640 = (pi01413 & ~w14865) | (pi01413 & w57770) | (~w14865 & w57770);
assign w16641 = w14865 & w57690;
assign w16642 = ~w16640 & ~w16641;
assign w16643 = (pi01414 & ~w14865) | (pi01414 & w57771) | (~w14865 & w57771);
assign w16644 = w14865 & w57576;
assign w16645 = ~w16643 & ~w16644;
assign w16646 = (pi01415 & ~w14865) | (pi01415 & w57772) | (~w14865 & w57772);
assign w16647 = w14865 & w57699;
assign w16648 = ~w16646 & ~w16647;
assign w16649 = (pi01416 & ~w14865) | (pi01416 & w57773) | (~w14865 & w57773);
assign w16650 = w14865 & w57774;
assign w16651 = ~w16649 & ~w16650;
assign w16652 = (pi01417 & ~w14865) | (pi01417 & w57775) | (~w14865 & w57775);
assign w16653 = w14865 & w57422;
assign w16654 = ~w16652 & ~w16653;
assign w16655 = (pi01418 & ~w14865) | (pi01418 & w57776) | (~w14865 & w57776);
assign w16656 = w14865 & w57777;
assign w16657 = ~w16655 & ~w16656;
assign w16658 = (pi01419 & ~w14865) | (pi01419 & w57778) | (~w14865 & w57778);
assign w16659 = w14865 & w57779;
assign w16660 = ~w16658 & ~w16659;
assign w16661 = (pi01420 & ~w14865) | (pi01420 & w57780) | (~w14865 & w57780);
assign w16662 = w14865 & w57426;
assign w16663 = ~w16661 & ~w16662;
assign w16664 = (pi01421 & ~w14865) | (pi01421 & w57781) | (~w14865 & w57781);
assign w16665 = w14865 & w57447;
assign w16666 = ~w16664 & ~w16665;
assign w16667 = (pi01422 & ~w14865) | (pi01422 & w57782) | (~w14865 & w57782);
assign w16668 = w14865 & w57574;
assign w16669 = ~w16667 & ~w16668;
assign w16670 = (pi01423 & ~w14865) | (pi01423 & w57783) | (~w14865 & w57783);
assign w16671 = w14865 & w57599;
assign w16672 = ~w16670 & ~w16671;
assign w16673 = (pi01424 & ~w14865) | (pi01424 & w57784) | (~w14865 & w57784);
assign w16674 = w14865 & w57430;
assign w16675 = ~w16673 & ~w16674;
assign w16676 = (pi01425 & ~w14865) | (pi01425 & w57785) | (~w14865 & w57785);
assign w16677 = w14865 & w57605;
assign w16678 = ~w16676 & ~w16677;
assign w16679 = (pi01426 & ~w14865) | (pi01426 & w57786) | (~w14865 & w57786);
assign w16680 = w14865 & w57453;
assign w16681 = ~w16679 & ~w16680;
assign w16682 = pi01427 & ~w16225;
assign w16683 = ~pi10622 & w16225;
assign w16684 = ~w16682 & ~w16683;
assign w16685 = pi01428 & ~w16225;
assign w16686 = ~pi10635 & w16225;
assign w16687 = ~w16685 & ~w16686;
assign w16688 = pi01429 & ~w16225;
assign w16689 = ~pi10634 & w16225;
assign w16690 = ~w16688 & ~w16689;
assign w16691 = pi01430 & ~w16225;
assign w16692 = ~pi10637 & w16225;
assign w16693 = ~w16691 & ~w16692;
assign w16694 = pi01431 & ~w16225;
assign w16695 = ~pi10639 & w16225;
assign w16696 = ~w16694 & ~w16695;
assign w16697 = pi01432 & ~w16225;
assign w16698 = ~pi10640 & w16225;
assign w16699 = ~w16697 & ~w16698;
assign w16700 = pi01433 & ~w16225;
assign w16701 = ~pi10623 & w16225;
assign w16702 = ~w16700 & ~w16701;
assign w16703 = pi01434 & ~w16225;
assign w16704 = ~pi10641 & w16225;
assign w16705 = ~w16703 & ~w16704;
assign w16706 = pi01435 & ~w16225;
assign w16707 = ~pi10624 & w16225;
assign w16708 = ~w16706 & ~w16707;
assign w16709 = pi01436 & ~w16225;
assign w16710 = ~pi10652 & w16225;
assign w16711 = ~w16709 & ~w16710;
assign w16712 = pi01437 & ~w16225;
assign w16713 = ~pi10653 & w16225;
assign w16714 = ~w16712 & ~w16713;
assign w16715 = pi01438 & ~w16225;
assign w16716 = ~pi10627 & w16225;
assign w16717 = ~w16715 & ~w16716;
assign w16718 = pi01439 & ~w16225;
assign w16719 = ~pi10630 & w16225;
assign w16720 = ~w16718 & ~w16719;
assign w16721 = (pi01440 & ~w16005) | (pi01440 & w57787) | (~w16005 & w57787);
assign w16722 = w16005 & w57621;
assign w16723 = ~w16721 & ~w16722;
assign w16724 = (pi01441 & ~w16005) | (pi01441 & w57788) | (~w16005 & w57788);
assign w16725 = w16005 & w57623;
assign w16726 = ~w16724 & ~w16725;
assign w16727 = (pi01442 & ~w16005) | (pi01442 & w57789) | (~w16005 & w57789);
assign w16728 = w16005 & w57790;
assign w16729 = ~w16727 & ~w16728;
assign w16730 = (pi01443 & ~w16005) | (pi01443 & w57791) | (~w16005 & w57791);
assign w16731 = w16005 & w57547;
assign w16732 = ~w16730 & ~w16731;
assign w16733 = (pi01444 & ~w16005) | (pi01444 & w57792) | (~w16005 & w57792);
assign w16734 = w16005 & w57793;
assign w16735 = ~w16733 & ~w16734;
assign w16736 = (pi01445 & ~w16005) | (pi01445 & w57794) | (~w16005 & w57794);
assign w16737 = w16005 & w57763;
assign w16738 = ~w16736 & ~w16737;
assign w16739 = (pi01446 & ~w16005) | (pi01446 & w57795) | (~w16005 & w57795);
assign w16740 = w16005 & w57796;
assign w16741 = ~w16739 & ~w16740;
assign w16742 = (pi01447 & ~w16005) | (pi01447 & w57797) | (~w16005 & w57797);
assign w16743 = w16005 & w57798;
assign w16744 = ~w16742 & ~w16743;
assign w16745 = (pi01448 & ~w16005) | (pi01448 & w57799) | (~w16005 & w57799);
assign w16746 = w16005 & w57800;
assign w16747 = ~w16745 & ~w16746;
assign w16748 = w12853 & w57801;
assign w16749 = pi02800 & w12910;
assign w16750 = pi02791 & w12897;
assign w16751 = pi01471 & w12915;
assign w16752 = pi00857 & pi01449;
assign w16753 = pi09899 & w12902;
assign w16754 = pi09941 & w12908;
assign w16755 = pi09880 & w12906;
assign w16756 = w12853 & w57802;
assign w16757 = (~w16752 & ~w12901) | (~w16752 & w57803) | (~w12901 & w57803);
assign w16758 = ~w16749 & w16757;
assign w16759 = ~w16753 & ~w16754;
assign w16760 = ~w16755 & w16759;
assign w16761 = w16758 & w57804;
assign w16762 = w16760 & w57805;
assign w16763 = w16761 & w16762;
assign w16764 = ~w10686 & ~w16192;
assign w16765 = ~w11709 & w57806;
assign w16766 = w11709 & w57807;
assign w16767 = pi01450 & w15987;
assign w16768 = ~w16765 & ~w16766;
assign w16769 = ~w16767 & w16768;
assign w16770 = ~w11706 & ~w16769;
assign w16771 = ~pi01451 & ~w14864;
assign w16772 = (w12993 & ~w14864) | (w12993 & w57808) | (~w14864 & w57808);
assign w16773 = ~w16771 & w16772;
assign w16774 = ~w16407 & ~w16773;
assign w16775 = ~pi01168 & ~w14858;
assign w16776 = ~pi00477 & ~pi00478;
assign w16777 = ~pi00479 & ~pi00480;
assign w16778 = ~pi00481 & ~pi00482;
assign w16779 = ~pi00483 & ~pi00484;
assign w16780 = w16778 & w16779;
assign w16781 = w16776 & w16777;
assign w16782 = w16780 & w16781;
assign w16783 = pi09804 & ~w16782;
assign w16784 = ~w16782 & w57809;
assign w16785 = ~w16775 & ~w16784;
assign w16786 = (pi00139 & w16782) | (pi00139 & w57810) | (w16782 & w57810);
assign w16787 = pi02796 & ~pi09802;
assign w16788 = pi09867 & ~w16787;
assign w16789 = pi01455 & pi02796;
assign w16790 = w16788 & w16789;
assign w16791 = pi01452 & pi09866;
assign w16792 = w16788 & w57811;
assign w16793 = w16786 & ~w16792;
assign w16794 = ~w16785 & ~w16793;
assign w16795 = w16786 & ~w16790;
assign w16796 = ~w16785 & ~w16795;
assign w16797 = pi09866 & w16796;
assign w16798 = (~pi01452 & ~w16796) | (~pi01452 & w57812) | (~w16796 & w57812);
assign w16799 = ~w16794 & ~w16798;
assign w16800 = w16775 & w16786;
assign w16801 = (pi01453 & ~w16800) | (pi01453 & w57813) | (~w16800 & w57813);
assign w16802 = ~pi01453 & w16794;
assign w16803 = ~w16801 & ~w16802;
assign w16804 = ~pi01454 & ~w16195;
assign w16805 = (~w11706 & ~w16195) | (~w11706 & w57814) | (~w16195 & w57814);
assign w16806 = ~w16804 & w16805;
assign w16807 = pi02796 & w16800;
assign w16808 = w16800 & w57815;
assign w16809 = (~pi01455 & ~w16800) | (~pi01455 & w57816) | (~w16800 & w57816);
assign w16810 = ~w16796 & ~w16809;
assign w16811 = (pi01456 & ~w11485) | (pi01456 & w57817) | (~w11485 & w57817);
assign w16812 = w11485 & w57818;
assign w16813 = ~w16811 & ~w16812;
assign w16814 = (pi01457 & ~w11485) | (pi01457 & w57819) | (~w11485 & w57819);
assign w16815 = w11485 & w57820;
assign w16816 = ~w16814 & ~w16815;
assign w16817 = (pi01458 & ~w11485) | (pi01458 & w57821) | (~w11485 & w57821);
assign w16818 = w11485 & w57822;
assign w16819 = ~w16817 & ~w16818;
assign w16820 = (pi01459 & ~w11485) | (pi01459 & w57823) | (~w11485 & w57823);
assign w16821 = w11485 & w57824;
assign w16822 = ~w16820 & ~w16821;
assign w16823 = (pi01460 & ~w11485) | (pi01460 & w57825) | (~w11485 & w57825);
assign w16824 = w11485 & w57826;
assign w16825 = ~w16823 & ~w16824;
assign w16826 = (pi01461 & ~w11485) | (pi01461 & w57827) | (~w11485 & w57827);
assign w16827 = w11485 & w57828;
assign w16828 = ~w16826 & ~w16827;
assign w16829 = (pi01462 & ~w11485) | (pi01462 & w57829) | (~w11485 & w57829);
assign w16830 = w11485 & w57830;
assign w16831 = ~w16829 & ~w16830;
assign w16832 = pi01463 & w12992;
assign w16833 = ~w12985 & ~w15944;
assign w16834 = w12989 & w57831;
assign w16835 = ~w12989 & w57832;
assign w16836 = ~w16834 & ~w16835;
assign w16837 = ~w16832 & w16836;
assign w16838 = w12993 & ~w16837;
assign w16839 = (pi01464 & ~w11485) | (pi01464 & w57833) | (~w11485 & w57833);
assign w16840 = w11485 & w57834;
assign w16841 = ~w16839 & ~w16840;
assign w16842 = (pi01465 & ~w11485) | (pi01465 & w57835) | (~w11485 & w57835);
assign w16843 = w11485 & w57836;
assign w16844 = ~w16842 & ~w16843;
assign w16845 = (pi01466 & ~w11485) | (pi01466 & w57837) | (~w11485 & w57837);
assign w16846 = w11485 & w57838;
assign w16847 = ~w16845 & ~w16846;
assign w16848 = (pi01467 & ~w11485) | (pi01467 & w57839) | (~w11485 & w57839);
assign w16849 = w11485 & w57840;
assign w16850 = ~w16848 & ~w16849;
assign w16851 = (pi01468 & ~w11485) | (pi01468 & w57841) | (~w11485 & w57841);
assign w16852 = w11485 & w57842;
assign w16853 = ~w16851 & ~w16852;
assign w16854 = (pi01469 & ~w11485) | (pi01469 & w57843) | (~w11485 & w57843);
assign w16855 = w11485 & w57844;
assign w16856 = ~w16854 & ~w16855;
assign w16857 = (pi01470 & ~w11485) | (pi01470 & w57845) | (~w11485 & w57845);
assign w16858 = w11485 & w57846;
assign w16859 = ~w16857 & ~w16858;
assign w16860 = (pi01471 & ~w11485) | (pi01471 & w57847) | (~w11485 & w57847);
assign w16861 = w11485 & w57848;
assign w16862 = ~w16860 & ~w16861;
assign w16863 = (pi01472 & ~w11485) | (pi01472 & w57849) | (~w11485 & w57849);
assign w16864 = w11485 & w57850;
assign w16865 = ~w16863 & ~w16864;
assign w16866 = (pi01473 & ~w11485) | (pi01473 & w57851) | (~w11485 & w57851);
assign w16867 = w11485 & w57852;
assign w16868 = ~w16866 & ~w16867;
assign w16869 = (pi01474 & ~w11485) | (pi01474 & w57853) | (~w11485 & w57853);
assign w16870 = w11485 & w57854;
assign w16871 = ~w16869 & ~w16870;
assign w16872 = (pi01475 & ~w11485) | (pi01475 & w57855) | (~w11485 & w57855);
assign w16873 = w11485 & w57856;
assign w16874 = ~w16872 & ~w16873;
assign w16875 = (pi01476 & ~w11485) | (pi01476 & w57857) | (~w11485 & w57857);
assign w16876 = w11485 & w57858;
assign w16877 = ~w16875 & ~w16876;
assign w16878 = w13057 & w14844;
assign w16879 = w14844 & w57859;
assign w16880 = (~w11706 & ~w14844) | (~w11706 & w57860) | (~w14844 & w57860);
assign w16881 = (w14844 & w57861) | (w14844 & w57862) | (w57861 & w57862);
assign w16882 = pi01477 & ~w16881;
assign w16883 = ~w16878 & ~w16882;
assign w16884 = (pi01478 & ~w11485) | (pi01478 & w57863) | (~w11485 & w57863);
assign w16885 = w11485 & w57864;
assign w16886 = ~w16884 & ~w16885;
assign w16887 = pi00869 & ~w1413;
assign w16888 = ~pi00869 & pi01479;
assign w16889 = ~w16887 & ~w16888;
assign w16890 = (~w12877 & w14858) | (~w12877 & w57865) | (w14858 & w57865);
assign w16891 = pi10029 & w3878;
assign w16892 = w16890 & ~w16891;
assign w16893 = ~pi02699 & ~pi02700;
assign w16894 = pi02180 & ~pi02696;
assign w16895 = w16893 & w16894;
assign w16896 = pi02697 & pi02701;
assign w16897 = pi02698 & ~pi02702;
assign w16898 = w16896 & w16897;
assign w16899 = w16895 & w16898;
assign w16900 = (w16899 & ~w16890) | (w16899 & w57866) | (~w16890 & w57866);
assign w16901 = pi01482 & ~w16900;
assign w16902 = ~pi02705 & w16900;
assign w16903 = ~w16901 & ~w16902;
assign w16904 = pi09998 & w3878;
assign w16905 = w16890 & ~w16904;
assign w16906 = ~pi02697 & pi02702;
assign w16907 = pi02698 & ~pi02701;
assign w16908 = w16906 & w16907;
assign w16909 = ~pi02180 & pi02699;
assign w16910 = pi02696 & pi02700;
assign w16911 = w16909 & w16910;
assign w16912 = w16908 & w16911;
assign w16913 = (w16912 & ~w16890) | (w16912 & w57867) | (~w16890 & w57867);
assign w16914 = pi01483 & ~w16913;
assign w16915 = ~pi02711 & w16913;
assign w16916 = ~w16914 & ~w16915;
assign w16917 = pi02180 & pi02699;
assign w16918 = ~pi02696 & pi02700;
assign w16919 = w16917 & w16918;
assign w16920 = pi02697 & ~pi02701;
assign w16921 = w16897 & w16920;
assign w16922 = w16919 & w16921;
assign w16923 = (w16922 & ~w16890) | (w16922 & w57868) | (~w16890 & w57868);
assign w16924 = pi01484 & ~w16923;
assign w16925 = ~pi02710 & w16923;
assign w16926 = ~w16924 & ~w16925;
assign w16927 = pi10028 & w3878;
assign w16928 = w16890 & ~w16927;
assign w16929 = pi02698 & pi02702;
assign w16930 = w16896 & w16929;
assign w16931 = w16919 & w16930;
assign w16932 = (w16931 & ~w16890) | (w16931 & w57869) | (~w16890 & w57869);
assign w16933 = pi01485 & ~w16932;
assign w16934 = ~pi09812 & w16932;
assign w16935 = ~w16933 & ~w16934;
assign w16936 = ~pi02699 & pi02700;
assign w16937 = pi02180 & pi02696;
assign w16938 = w16936 & w16937;
assign w16939 = ~pi02698 & ~pi02702;
assign w16940 = w16896 & w16939;
assign w16941 = w16938 & w16940;
assign w16942 = (w16941 & ~w16890) | (w16941 & w57870) | (~w16890 & w57870);
assign w16943 = pi01486 & ~w16942;
assign w16944 = ~pi02711 & w16942;
assign w16945 = ~w16943 & ~w16944;
assign w16946 = ~pi02696 & ~pi02700;
assign w16947 = w16917 & w16946;
assign w16948 = w16940 & w16947;
assign w16949 = (w16948 & ~w16890) | (w16948 & w57871) | (~w16890 & w57871);
assign w16950 = pi01487 & ~w16949;
assign w16951 = ~pi02705 & w16949;
assign w16952 = ~w16950 & ~w16951;
assign w16953 = w16894 & w16936;
assign w16954 = w16908 & w16953;
assign w16955 = (w16954 & ~w16890) | (w16954 & w57872) | (~w16890 & w57872);
assign w16956 = pi01488 & ~w16955;
assign w16957 = ~pi09848 & w16955;
assign w16958 = ~w16956 & ~w16957;
assign w16959 = pi02696 & ~pi02700;
assign w16960 = w16909 & w16959;
assign w16961 = w16930 & w16960;
assign w16962 = (w16961 & ~w16890) | (w16961 & w57873) | (~w16890 & w57873);
assign w16963 = pi01489 & ~w16962;
assign w16964 = ~pi02709 & w16962;
assign w16965 = ~w16963 & ~w16964;
assign w16966 = ~pi02698 & ~pi02701;
assign w16967 = w16906 & w16966;
assign w16968 = ~pi02180 & pi02696;
assign w16969 = w16936 & w16968;
assign w16970 = w16967 & w16969;
assign w16971 = (w16970 & ~w16890) | (w16970 & w57874) | (~w16890 & w57874);
assign w16972 = pi01490 & ~w16971;
assign w16973 = (~pi02717 & ~w16890) | (~pi02717 & w57875) | (~w16890 & w57875);
assign w16974 = (~w16890 & w57876) | (~w16890 & w57877) | (w57876 & w57877);
assign w16975 = ~w16972 & ~w16974;
assign w16976 = ~pi02698 & pi02702;
assign w16977 = w16920 & w16976;
assign w16978 = w16911 & w16977;
assign w16979 = (w16978 & ~w16890) | (w16978 & w57878) | (~w16890 & w57878);
assign w16980 = pi01491 & ~w16979;
assign w16981 = ~pi02711 & w16979;
assign w16982 = ~w16980 & ~w16981;
assign w16983 = w16893 & w16968;
assign w16984 = ~pi02697 & ~pi02702;
assign w16985 = w16966 & w16984;
assign w16986 = w16983 & w16985;
assign w16987 = (w16986 & ~w16890) | (w16986 & w57879) | (~w16890 & w57879);
assign w16988 = pi01492 & ~w16987;
assign w16989 = ~pi02714 & w16987;
assign w16990 = ~w16988 & ~w16989;
assign w16991 = pi10232 & w3878;
assign w16992 = w16890 & ~w16991;
assign w16993 = w16917 & w16959;
assign w16994 = w16967 & w16993;
assign w16995 = (w16994 & ~w16890) | (w16994 & w57880) | (~w16890 & w57880);
assign w16996 = pi01493 & ~w16995;
assign w16997 = ~pi02722 & w16995;
assign w16998 = ~w16996 & ~w16997;
assign w16999 = w16953 & w16985;
assign w17000 = (w16999 & ~w16890) | (w16999 & w57881) | (~w16890 & w57881);
assign w17001 = pi01494 & ~w17000;
assign w17002 = ~pi09848 & w17000;
assign w17003 = ~w17001 & ~w17002;
assign w17004 = ~pi02180 & ~pi02696;
assign w17005 = w16893 & w17004;
assign w17006 = w16967 & w17005;
assign w17007 = (w17006 & ~w16890) | (w17006 & w57882) | (~w16890 & w57882);
assign w17008 = pi01495 & ~w17007;
assign w17009 = ~pi02711 & w17007;
assign w17010 = ~w17008 & ~w17009;
assign w17011 = w16940 & w17005;
assign w17012 = (w17011 & ~w16890) | (w17011 & w57883) | (~w16890 & w57883);
assign w17013 = pi01496 & ~w17012;
assign w17014 = ~pi02169 & w17012;
assign w17015 = ~w17013 & ~w17014;
assign w17016 = w16893 & w16937;
assign w17017 = w16908 & w17016;
assign w17018 = (w17017 & ~w16890) | (w17017 & w57884) | (~w16890 & w57884);
assign w17019 = pi01497 & ~w17018;
assign w17020 = (~pi02712 & ~w16890) | (~pi02712 & w57885) | (~w16890 & w57885);
assign w17021 = (~w16890 & w57886) | (~w16890 & w57887) | (w57886 & w57887);
assign w17022 = ~w17019 & ~w17021;
assign w17023 = w16985 & w17016;
assign w17024 = (w17023 & ~w16890) | (w17023 & w57888) | (~w16890 & w57888);
assign w17025 = pi01498 & ~w17024;
assign w17026 = ~pi09812 & w17024;
assign w17027 = ~w17025 & ~w17026;
assign w17028 = w16898 & w16919;
assign w17029 = (w17028 & ~w16890) | (w17028 & w57889) | (~w16890 & w57889);
assign w17030 = pi01499 & ~w17029;
assign w17031 = ~pi02714 & w17029;
assign w17032 = ~w17030 & ~w17031;
assign w17033 = pi01500 & ~w16979;
assign w17034 = ~pi02715 & w16979;
assign w17035 = ~w17033 & ~w17034;
assign w17036 = pi02698 & pi02701;
assign w17037 = w16984 & w17036;
assign w17038 = w16909 & w16946;
assign w17039 = w17037 & w17038;
assign w17040 = (w17039 & ~w16890) | (w17039 & w57890) | (~w16890 & w57890);
assign w17041 = pi01501 & ~w17040;
assign w17042 = ~pi02160 & w17040;
assign w17043 = ~w17041 & ~w17042;
assign w17044 = pi01502 & ~w16979;
assign w17045 = ~pi02717 & w16979;
assign w17046 = ~w17044 & ~w17045;
assign w17047 = w16895 & w16921;
assign w17048 = (w17047 & ~w16890) | (w17047 & w57891) | (~w16890 & w57891);
assign w17049 = pi01503 & ~w17048;
assign w17050 = ~pi09812 & w17048;
assign w17051 = ~w17049 & ~w17050;
assign w17052 = w16910 & w16917;
assign w17053 = w16898 & w17052;
assign w17054 = (w17053 & ~w16890) | (w17053 & w57892) | (~w16890 & w57892);
assign w17055 = pi01504 & ~w17054;
assign w17056 = ~pi02711 & w17054;
assign w17057 = ~w17055 & ~w17056;
assign w17058 = ~pi02698 & pi02701;
assign w17059 = w16984 & w17058;
assign w17060 = w16938 & w17059;
assign w17061 = (w17060 & ~w16890) | (w17060 & w57893) | (~w16890 & w57893);
assign w17062 = pi01505 & ~w17061;
assign w17063 = ~pi02705 & w17061;
assign w17064 = ~w17062 & ~w17063;
assign w17065 = pi09963 & pi09969;
assign w17066 = pi09926 & w17065;
assign w17067 = w11114 & w17066;
assign w17068 = w25 & w57894;
assign w17069 = ~w17067 & ~w17068;
assign w17070 = pi00250 & ~w17069;
assign w17071 = (w16994 & ~w16890) | (w16994 & w57895) | (~w16890 & w57895);
assign w17072 = pi01507 & ~w17071;
assign w17073 = ~pi02711 & w17071;
assign w17074 = ~w17072 & ~w17073;
assign w17075 = pi01508 & ~w16923;
assign w17076 = ~pi02723 & w16923;
assign w17077 = ~w17075 & ~w17076;
assign w17078 = w16967 & w17052;
assign w17079 = (w17078 & ~w16890) | (w17078 & w57896) | (~w16890 & w57896);
assign w17080 = pi01509 & ~w17079;
assign w17081 = ~pi09954 & w17079;
assign w17082 = ~w17080 & ~w17081;
assign w17083 = w16936 & w17004;
assign w17084 = w16967 & w17083;
assign w17085 = (w17084 & ~w16890) | (w17084 & w57897) | (~w16890 & w57897);
assign w17086 = pi01510 & ~w17085;
assign w17087 = ~pi02704 & w17085;
assign w17088 = ~w17086 & ~w17087;
assign w17089 = pi01511 & ~w16995;
assign w17090 = ~pi02721 & w16995;
assign w17091 = ~w17089 & ~w17090;
assign w17092 = pi01512 & ~w16923;
assign w17093 = ~pi02705 & w16923;
assign w17094 = ~w17092 & ~w17093;
assign w17095 = pi01513 & ~w17079;
assign w17096 = ~pi09848 & w17079;
assign w17097 = ~w17095 & ~w17096;
assign w17098 = w17005 & w17037;
assign w17099 = (w17098 & ~w16890) | (w17098 & w57898) | (~w16890 & w57898);
assign w17100 = pi01514 & ~w17099;
assign w17101 = ~pi02705 & w17099;
assign w17102 = ~w17100 & ~w17101;
assign w17103 = w16919 & w16967;
assign w17104 = (w17103 & ~w16890) | (w17103 & w57899) | (~w16890 & w57899);
assign w17105 = pi01515 & ~w17104;
assign w17106 = ~pi09954 & w17104;
assign w17107 = ~w17105 & ~w17106;
assign w17108 = w16940 & w16983;
assign w17109 = (w17108 & ~w16890) | (w17108 & w57900) | (~w16890 & w57900);
assign w17110 = pi01516 & ~w17109;
assign w17111 = ~pi02164 & w17109;
assign w17112 = ~w17110 & ~w17111;
assign w17113 = w16907 & w16984;
assign w17114 = w17016 & w17113;
assign w17115 = (w17114 & ~w16890) | (w17114 & w57901) | (~w16890 & w57901);
assign w17116 = pi01517 & ~w17115;
assign w17117 = ~pi02719 & w17115;
assign w17118 = ~w17116 & ~w17117;
assign w17119 = w16985 & w17038;
assign w17120 = (w17119 & ~w16890) | (w17119 & w57902) | (~w16890 & w57902);
assign w17121 = pi01518 & ~w17120;
assign w17122 = ~pi09961 & w17120;
assign w17123 = ~w17121 & ~w17122;
assign w17124 = w16909 & w16918;
assign w17125 = w17059 & w17124;
assign w17126 = (w17125 & ~w16890) | (w17125 & w57903) | (~w16890 & w57903);
assign w17127 = pi01519 & ~w17126;
assign w17128 = (~pi02720 & ~w16890) | (~pi02720 & w57904) | (~w16890 & w57904);
assign w17129 = (~w16890 & w57905) | (~w16890 & w57906) | (w57905 & w57906);
assign w17130 = ~w17127 & ~w17129;
assign w17131 = w16947 & w17037;
assign w17132 = (w17131 & ~w16890) | (w17131 & w57907) | (~w16890 & w57907);
assign w17133 = pi01520 & ~w17132;
assign w17134 = ~pi02723 & w17132;
assign w17135 = ~w17133 & ~w17134;
assign w17136 = w16920 & w16929;
assign w17137 = w16895 & w17136;
assign w17138 = (w17137 & ~w16890) | (w17137 & w57908) | (~w16890 & w57908);
assign w17139 = pi01521 & ~w17138;
assign w17140 = ~pi02712 & w17138;
assign w17141 = ~w17139 & ~w17140;
assign w17142 = pi01522 & ~w17018;
assign w17143 = ~pi02715 & w17018;
assign w17144 = ~w17142 & ~w17143;
assign w17145 = pi01523 & ~w16949;
assign w17146 = ~pi02723 & w16949;
assign w17147 = ~w17145 & ~w17146;
assign w17148 = w16908 & w16993;
assign w17149 = (w17148 & ~w16890) | (w17148 & w57909) | (~w16890 & w57909);
assign w17150 = pi01524 & ~w17149;
assign w17151 = ~pi02720 & w17149;
assign w17152 = ~w17150 & ~w17151;
assign w17153 = w16908 & w16938;
assign w17154 = (w17153 & ~w16890) | (w17153 & w57910) | (~w16890 & w57910);
assign w17155 = pi01525 & ~w17154;
assign w17156 = ~pi02720 & w17154;
assign w17157 = ~w17155 & ~w17156;
assign w17158 = (w16912 & ~w16890) | (w16912 & w57911) | (~w16890 & w57911);
assign w17159 = pi01526 & ~w17158;
assign w17160 = ~pi09962 & w17158;
assign w17161 = ~w17159 & ~w17160;
assign w17162 = w16967 & w17016;
assign w17163 = (w17162 & ~w16890) | (w17162 & w57912) | (~w16890 & w57912);
assign w17164 = pi01527 & ~w17163;
assign w17165 = ~pi09812 & w17163;
assign w17166 = ~w17164 & ~w17165;
assign w17167 = w16983 & w17113;
assign w17168 = (w17167 & ~w16890) | (w17167 & w57913) | (~w16890 & w57913);
assign w17169 = pi01528 & ~w17168;
assign w17170 = ~pi09812 & w17168;
assign w17171 = ~w17169 & ~w17170;
assign w17172 = w16895 & w16985;
assign w17173 = (w17172 & ~w16890) | (w17172 & w57914) | (~w16890 & w57914);
assign w17174 = pi01529 & ~w17173;
assign w17175 = ~pi02720 & w17173;
assign w17176 = ~w17174 & ~w17175;
assign w17177 = w16911 & w17136;
assign w17178 = (w17177 & ~w16890) | (w17177 & w57915) | (~w16890 & w57915);
assign w17179 = pi01530 & ~w17178;
assign w17180 = ~pi09962 & w17178;
assign w17181 = ~w17179 & ~w17180;
assign w17182 = w16920 & w16939;
assign w17183 = w17038 & w17182;
assign w17184 = (w17183 & ~w16890) | (w17183 & w57916) | (~w16890 & w57916);
assign w17185 = pi01531 & ~w17184;
assign w17186 = (~pi09848 & ~w16890) | (~pi09848 & w57917) | (~w16890 & w57917);
assign w17187 = (~w16890 & w57918) | (~w16890 & w57919) | (w57918 & w57919);
assign w17188 = ~w17185 & ~w17187;
assign w17189 = w16906 & w17036;
assign w17190 = w16969 & w17189;
assign w17191 = (w17190 & ~w16890) | (w17190 & w57920) | (~w16890 & w57920);
assign w17192 = pi01532 & ~w17191;
assign w17193 = (~pi09812 & ~w16890) | (~pi09812 & w57921) | (~w16890 & w57921);
assign w17194 = (~w16890 & w57922) | (~w16890 & w57923) | (w57922 & w57923);
assign w17195 = ~w17192 & ~w17194;
assign w17196 = (w17047 & ~w16890) | (w17047 & w57924) | (~w16890 & w57924);
assign w17197 = pi01533 & ~w17196;
assign w17198 = ~pi02718 & w17196;
assign w17199 = ~w17197 & ~w17198;
assign w17200 = w16898 & w16911;
assign w17201 = (w17200 & ~w16890) | (w17200 & w57925) | (~w16890 & w57925);
assign w17202 = pi01534 & ~w17201;
assign w17203 = (~w16890 & w57926) | (~w16890 & w57927) | (w57926 & w57927);
assign w17204 = ~w17202 & ~w17203;
assign w17205 = w16911 & w17037;
assign w17206 = (w17205 & ~w16890) | (w17205 & w57928) | (~w16890 & w57928);
assign w17207 = pi01535 & ~w17206;
assign w17208 = ~pi02718 & w17206;
assign w17209 = ~w17207 & ~w17208;
assign w17210 = w16953 & w17059;
assign w17211 = (w17210 & ~w16890) | (w17210 & w57929) | (~w16890 & w57929);
assign w17212 = pi01536 & ~w17211;
assign w17213 = ~pi09962 & w17211;
assign w17214 = ~w17212 & ~w17213;
assign w17215 = pi01537 & ~w17178;
assign w17216 = ~pi02704 & w17178;
assign w17217 = ~w17215 & ~w17216;
assign w17218 = w16993 & w17059;
assign w17219 = (w17218 & ~w16890) | (w17218 & w57930) | (~w16890 & w57930);
assign w17220 = pi01538 & ~w17219;
assign w17221 = ~pi02723 & w17219;
assign w17222 = ~w17220 & ~w17221;
assign w17223 = pi01539 & ~w17211;
assign w17224 = ~pi02704 & w17211;
assign w17225 = ~w17223 & ~w17224;
assign w17226 = w16921 & w17052;
assign w17227 = (w17226 & ~w16890) | (w17226 & w57931) | (~w16890 & w57931);
assign w17228 = pi01540 & ~w17227;
assign w17229 = ~pi09962 & w17227;
assign w17230 = ~w17228 & ~w17229;
assign w17231 = w16993 & w17037;
assign w17232 = (w17231 & ~w16890) | (w17231 & w57932) | (~w16890 & w57932);
assign w17233 = pi01541 & ~w17232;
assign w17234 = ~pi09954 & w17232;
assign w17235 = ~w17233 & ~w17234;
assign w17236 = pi01542 & ~w16955;
assign w17237 = ~pi09954 & w16955;
assign w17238 = ~w17236 & ~w17237;
assign w17239 = w16911 & w16940;
assign w17240 = (w17239 & ~w16890) | (w17239 & w57933) | (~w16890 & w57933);
assign w17241 = pi01543 & ~w17240;
assign w17242 = ~pi09812 & w17240;
assign w17243 = ~w17241 & ~w17242;
assign w17244 = w16895 & w16977;
assign w17245 = (w17244 & ~w16890) | (w17244 & w57934) | (~w16890 & w57934);
assign w17246 = pi01544 & ~w17245;
assign w17247 = (~w16890 & w57935) | (~w16890 & w57936) | (w57935 & w57936);
assign w17248 = ~w17246 & ~w17247;
assign w17249 = w16921 & w17005;
assign w17250 = (w17249 & ~w16890) | (w17249 & w57937) | (~w16890 & w57937);
assign w17251 = pi01545 & ~w17250;
assign w17252 = ~pi02719 & w17250;
assign w17253 = ~w17251 & ~w17252;
assign w17254 = w16977 & w17052;
assign w17255 = (w17254 & ~w16890) | (w17254 & w57938) | (~w16890 & w57938);
assign w17256 = pi01546 & ~w17255;
assign w17257 = ~pi09812 & w17255;
assign w17258 = ~w17256 & ~w17257;
assign w17259 = w16895 & w17059;
assign w17260 = (w17259 & ~w16890) | (w17259 & w57939) | (~w16890 & w57939);
assign w17261 = pi01547 & ~w17260;
assign w17262 = ~pi09962 & w17260;
assign w17263 = ~w17261 & ~w17262;
assign w17264 = w16969 & w17113;
assign w17265 = (w17264 & ~w16890) | (w17264 & w57940) | (~w16890 & w57940);
assign w17266 = pi01548 & ~w17265;
assign w17267 = (~w16890 & w57941) | (~w16890 & w57942) | (w57941 & w57942);
assign w17268 = ~w17266 & ~w17267;
assign w17269 = (w17205 & ~w16890) | (w17205 & w57943) | (~w16890 & w57943);
assign w17270 = pi01549 & ~w17269;
assign w17271 = ~pi02716 & w17269;
assign w17272 = ~w17270 & ~w17271;
assign w17273 = pi01550 & ~w17255;
assign w17274 = (~w16890 & w57944) | (~w16890 & w57945) | (w57944 & w57945);
assign w17275 = ~w17273 & ~w17274;
assign w17276 = pi01551 & ~w16900;
assign w17277 = ~pi02723 & w16900;
assign w17278 = ~w17276 & ~w17277;
assign w17279 = w16908 & w16983;
assign w17280 = (w17279 & ~w16890) | (w17279 & w57946) | (~w16890 & w57946);
assign w17281 = pi01552 & ~w17280;
assign w17282 = ~pi09962 & w17280;
assign w17283 = ~w17281 & ~w17282;
assign w17284 = w17124 & w17136;
assign w17285 = (w17284 & ~w16890) | (w17284 & w57947) | (~w16890 & w57947);
assign w17286 = pi01553 & ~w17285;
assign w17287 = ~pi02704 & w17285;
assign w17288 = ~w17286 & ~w17287;
assign w17289 = w17005 & w17059;
assign w17290 = (w17289 & ~w16890) | (w17289 & w57948) | (~w16890 & w57948);
assign w17291 = pi01554 & ~w17290;
assign w17292 = ~pi02716 & w17290;
assign w17293 = ~w17291 & ~w17292;
assign w17294 = pi01555 & ~w17163;
assign w17295 = ~pi02720 & w17163;
assign w17296 = ~w17294 & ~w17295;
assign w17297 = pi01556 & ~w17109;
assign w17298 = ~pi02721 & w17109;
assign w17299 = ~w17297 & ~w17298;
assign w17300 = w16919 & w16977;
assign w17301 = (w17300 & ~w16890) | (w17300 & w57949) | (~w16890 & w57949);
assign w17302 = pi01557 & ~w17301;
assign w17303 = ~pi09812 & w17301;
assign w17304 = ~w17302 & ~w17303;
assign w17305 = w16930 & w16947;
assign w17306 = (w17305 & ~w16890) | (w17305 & w57950) | (~w16890 & w57950);
assign w17307 = pi01558 & ~w17306;
assign w17308 = ~pi02720 & w17306;
assign w17309 = ~w17307 & ~w17308;
assign w17310 = pi01559 & ~w17158;
assign w17311 = (~pi02704 & ~w16890) | (~pi02704 & w57951) | (~w16890 & w57951);
assign w17312 = (~w16890 & w57952) | (~w16890 & w57953) | (w57952 & w57953);
assign w17313 = ~w17310 & ~w17312;
assign w17314 = w16898 & w16969;
assign w17315 = (w17314 & ~w16890) | (w17314 & w57954) | (~w16890 & w57954);
assign w17316 = pi01560 & ~w17315;
assign w17317 = (~pi02716 & ~w16890) | (~pi02716 & w57955) | (~w16890 & w57955);
assign w17318 = (~w16890 & w57956) | (~w16890 & w57957) | (w57956 & w57957);
assign w17319 = ~w17316 & ~w17318;
assign w17320 = w16911 & w16930;
assign w17321 = (w17320 & ~w16890) | (w17320 & w57958) | (~w16890 & w57958);
assign w17322 = pi01561 & ~w17321;
assign w17323 = ~pi02720 & w17321;
assign w17324 = ~w17322 & ~w17323;
assign w17325 = w17083 & w17182;
assign w17326 = ~w16928 & w17325;
assign w17327 = pi01562 & ~w17326;
assign w17328 = ~pi09812 & w17326;
assign w17329 = ~w17327 & ~w17328;
assign w17330 = ~w16928 & w17314;
assign w17331 = pi01563 & ~w17330;
assign w17332 = ~pi09812 & w17330;
assign w17333 = ~w17331 & ~w17332;
assign w17334 = w16985 & w17124;
assign w17335 = ~w16928 & w17334;
assign w17336 = pi01564 & ~w17335;
assign w17337 = w17193 & w17334;
assign w17338 = ~w17336 & ~w17337;
assign w17339 = w16938 & w17136;
assign w17340 = ~w16892 & w17339;
assign w17341 = pi01565 & ~w17340;
assign w17342 = ~pi02708 & w17340;
assign w17343 = ~w17341 & ~w17342;
assign w17344 = w16895 & w16967;
assign w17345 = ~w16928 & w17344;
assign w17346 = pi01566 & ~w17345;
assign w17347 = ~pi09812 & w17345;
assign w17348 = ~w17346 & ~w17347;
assign w17349 = w16898 & w16993;
assign w17350 = ~w16928 & w17349;
assign w17351 = pi01567 & ~w17350;
assign w17352 = ~pi09848 & w17350;
assign w17353 = ~w17351 & ~w17352;
assign w17354 = ~w16928 & w16978;
assign w17355 = pi01568 & ~w17354;
assign w17356 = w16978 & w17311;
assign w17357 = ~w17355 & ~w17356;
assign w17358 = pi01569 & ~w17115;
assign w17359 = ~pi02718 & w17115;
assign w17360 = ~w17358 & ~w17359;
assign w17361 = w16960 & w16985;
assign w17362 = ~w16905 & w17361;
assign w17363 = pi01570 & ~w17362;
assign w17364 = ~pi02714 & w17362;
assign w17365 = ~w17363 & ~w17364;
assign w17366 = w16898 & w17124;
assign w17367 = ~w16928 & w17366;
assign w17368 = pi01571 & ~w17367;
assign w17369 = ~pi02720 & w17367;
assign w17370 = ~w17368 & ~w17369;
assign w17371 = pi01572 & ~w17260;
assign w17372 = ~pi02704 & w17260;
assign w17373 = ~w17371 & ~w17372;
assign w17374 = w16906 & w17058;
assign w17375 = w16911 & w17374;
assign w17376 = ~w16905 & w17375;
assign w17377 = pi01573 & ~w17376;
assign w17378 = ~pi02713 & w17376;
assign w17379 = ~w17377 & ~w17378;
assign w17380 = w17016 & w17037;
assign w17381 = ~w16892 & w17380;
assign w17382 = pi01574 & ~w17381;
assign w17383 = ~pi02723 & w17381;
assign w17384 = ~w17382 & ~w17383;
assign w17385 = w16898 & w16947;
assign w17386 = ~w16928 & w17385;
assign w17387 = pi01575 & ~w17386;
assign w17388 = ~pi09954 & w17386;
assign w17389 = ~w17387 & ~w17388;
assign w17390 = w16908 & w17083;
assign w17391 = ~w16992 & w17390;
assign w17392 = pi01576 & ~w17391;
assign w17393 = ~pi02721 & w17391;
assign w17394 = ~w17392 & ~w17393;
assign w17395 = pi01577 & ~w17029;
assign w17396 = ~pi02711 & w17029;
assign w17397 = ~w17395 & ~w17396;
assign w17398 = w16895 & w17113;
assign w17399 = ~w16992 & w17398;
assign w17400 = pi01578 & ~w17399;
assign w17401 = ~pi02722 & w17399;
assign w17402 = ~w17400 & ~w17401;
assign w17403 = pi01579 & ~w17306;
assign w17404 = ~pi09812 & w17306;
assign w17405 = ~w17403 & ~w17404;
assign w17406 = w17038 & w17113;
assign w17407 = ~w16992 & w17406;
assign w17408 = pi01580 & ~w17407;
assign w17409 = ~pi02167 & w17407;
assign w17410 = ~w17408 & ~w17409;
assign w17411 = w16993 & w17189;
assign w17412 = ~w16928 & w17411;
assign w17413 = pi01581 & ~w17412;
assign w17414 = ~pi09812 & w17412;
assign w17415 = ~w17413 & ~w17414;
assign w17416 = w17037 & w17083;
assign w17417 = ~w16928 & w17416;
assign w17418 = pi01582 & ~w17417;
assign w17419 = ~pi09812 & w17417;
assign w17420 = ~w17418 & ~w17419;
assign w17421 = ~w16928 & w17339;
assign w17422 = pi01583 & ~w17421;
assign w17423 = ~pi02720 & w17421;
assign w17424 = ~w17422 & ~w17423;
assign w17425 = pi01584 & ~w17321;
assign w17426 = ~pi09812 & w17321;
assign w17427 = ~w17425 & ~w17426;
assign w17428 = w16911 & w16921;
assign w17429 = ~w16905 & w17428;
assign w17430 = pi01585 & ~w17429;
assign w17431 = ~pi02716 & w17429;
assign w17432 = ~w17430 & ~w17431;
assign w17433 = pi01586 & ~w17421;
assign w17434 = ~pi09812 & w17421;
assign w17435 = ~w17433 & ~w17434;
assign w17436 = w16967 & w17124;
assign w17437 = ~w16928 & w17436;
assign w17438 = pi01587 & ~w17437;
assign w17439 = ~pi09962 & ~w16928;
assign w17440 = w17436 & w17439;
assign w17441 = ~w17438 & ~w17440;
assign w17442 = pi01588 & ~w17386;
assign w17443 = ~pi09848 & w17386;
assign w17444 = ~w17442 & ~w17443;
assign w17445 = w16977 & w17016;
assign w17446 = ~w16905 & w17445;
assign w17447 = pi01589 & ~w17446;
assign w17448 = ~pi02712 & w17446;
assign w17449 = ~w17447 & ~w17448;
assign w17450 = w16969 & w17136;
assign w17451 = ~w16928 & w17450;
assign w17452 = pi01590 & ~w17451;
assign w17453 = ~pi02704 & w17451;
assign w17454 = ~w17452 & ~w17453;
assign w17455 = pi01591 & ~w17437;
assign w17456 = ~pi02704 & w17437;
assign w17457 = ~w17455 & ~w17456;
assign w17458 = pi01592 & ~w17367;
assign w17459 = ~pi09812 & w17367;
assign w17460 = ~w17458 & ~w17459;
assign w17461 = w16921 & w16938;
assign w17462 = ~w16928 & w17461;
assign w17463 = pi01593 & ~w17462;
assign w17464 = ~pi02178 & w17462;
assign w17465 = ~w17463 & ~w17464;
assign w17466 = w16953 & w17136;
assign w17467 = ~w16928 & w17466;
assign w17468 = pi01594 & ~w17467;
assign w17469 = ~pi09812 & w17467;
assign w17470 = ~w17468 & ~w17469;
assign w17471 = pi01595 & ~w17362;
assign w17472 = ~pi02712 & w17362;
assign w17473 = ~w17471 & ~w17472;
assign w17474 = w16930 & w17124;
assign w17475 = ~w16928 & w17474;
assign w17476 = pi01596 & ~w17475;
assign w17477 = ~pi09812 & w17475;
assign w17478 = ~w17476 & ~w17477;
assign w17479 = w17016 & w17182;
assign w17480 = ~w16992 & w17479;
assign w17481 = pi01597 & ~w17480;
assign w17482 = ~pi02718 & w17480;
assign w17483 = ~w17481 & ~w17482;
assign w17484 = pi01598 & ~w17326;
assign w17485 = ~pi02720 & w17326;
assign w17486 = ~w17484 & ~w17485;
assign w17487 = pi01599 & ~w17480;
assign w17488 = ~pi02719 & w17480;
assign w17489 = ~w17487 & ~w17488;
assign w17490 = w16947 & w16985;
assign w17491 = ~w16905 & w17490;
assign w17492 = pi01600 & ~w17491;
assign w17493 = ~pi02713 & w17491;
assign w17494 = ~w17492 & ~w17493;
assign w17495 = w16921 & w17038;
assign w17496 = ~w16928 & w17495;
assign w17497 = pi01601 & ~w17496;
assign w17498 = ~pi02720 & w17496;
assign w17499 = ~w17497 & ~w17498;
assign w17500 = w16947 & w17113;
assign w17501 = ~w16928 & w17500;
assign w17502 = pi01602 & ~w17501;
assign w17503 = ~pi09848 & w17501;
assign w17504 = ~w17502 & ~w17503;
assign w17505 = w17083 & w17113;
assign w17506 = ~w16928 & w17505;
assign w17507 = pi01603 & ~w17506;
assign w17508 = ~pi09954 & w17506;
assign w17509 = ~w17507 & ~w17508;
assign w17510 = w16960 & w17374;
assign w17511 = ~w16928 & w17510;
assign w17512 = pi01604 & ~w17511;
assign w17513 = ~pi09954 & ~w16928;
assign w17514 = w17510 & w17513;
assign w17515 = ~w17512 & ~w17514;
assign w17516 = w16983 & w17189;
assign w17517 = ~w16905 & w17516;
assign w17518 = pi01605 & ~w17517;
assign w17519 = ~pi02716 & w17517;
assign w17520 = ~w17518 & ~w17519;
assign w17521 = w16911 & w17189;
assign w17522 = ~w16928 & w17521;
assign w17523 = pi01607 & ~w17522;
assign w17524 = ~pi09812 & w17522;
assign w17525 = ~w17523 & ~w17524;
assign w17526 = w16953 & w17189;
assign w17527 = ~w16892 & w17526;
assign w17528 = pi01608 & ~w17527;
assign w17529 = ~pi02709 & w17527;
assign w17530 = ~w17528 & ~w17529;
assign w17531 = pi01609 & ~w17480;
assign w17532 = ~pi02703 & ~w16992;
assign w17533 = w17479 & w17532;
assign w17534 = ~w17531 & ~w17533;
assign w17535 = w16895 & w16940;
assign w17536 = ~w16905 & w17535;
assign w17537 = pi01610 & ~w17536;
assign w17538 = ~pi02714 & w17536;
assign w17539 = ~w17537 & ~w17538;
assign w17540 = w16930 & w17016;
assign w17541 = ~w16992 & w17540;
assign w17542 = pi01611 & ~w17541;
assign w17543 = ~pi02722 & w17541;
assign w17544 = ~w17542 & ~w17543;
assign w17545 = pi01612 & ~w17541;
assign w17546 = ~pi02703 & w17541;
assign w17547 = ~w17545 & ~w17546;
assign w17548 = ~w16905 & w17249;
assign w17549 = pi01613 & ~w17548;
assign w17550 = ~pi02712 & w17548;
assign w17551 = ~w17549 & ~w17550;
assign w17552 = ~w16992 & w17289;
assign w17553 = pi01614 & ~w17552;
assign w17554 = ~pi02721 & w17552;
assign w17555 = ~w17553 & ~w17554;
assign w17556 = w16953 & w17182;
assign w17557 = ~w16892 & w17556;
assign w17558 = pi01615 & ~w17557;
assign w17559 = ~pi02710 & w17557;
assign w17560 = ~w17558 & ~w17559;
assign w17561 = ~w16905 & w17047;
assign w17562 = pi01616 & ~w17561;
assign w17563 = ~pi02712 & w17561;
assign w17564 = ~w17562 & ~w17563;
assign w17565 = w16983 & w17374;
assign w17566 = ~w16992 & w17565;
assign w17567 = pi01617 & ~w17566;
assign w17568 = ~pi02169 & w17566;
assign w17569 = ~w17567 & ~w17568;
assign w17570 = pi01618 & ~w17536;
assign w17571 = w17020 & w17535;
assign w17572 = ~w17570 & ~w17571;
assign w17573 = w17037 & w17052;
assign w17574 = ~w16905 & w17573;
assign w17575 = pi01619 & ~w17574;
assign w17576 = ~pi02711 & w17574;
assign w17577 = ~w17575 & ~w17576;
assign w17578 = ~w16992 & w17137;
assign w17579 = pi01620 & ~w17578;
assign w17580 = ~pi02721 & w17578;
assign w17581 = ~w17579 & ~w17580;
assign w17582 = w16896 & w16976;
assign w17583 = w17052 & w17582;
assign w17584 = ~w16992 & w17583;
assign w17585 = pi01621 & ~w17584;
assign w17586 = ~pi02718 & ~w16992;
assign w17587 = w17583 & w17586;
assign w17588 = ~w17585 & ~w17587;
assign w17589 = pi01622 & ~w17578;
assign w17590 = ~pi02164 & w17578;
assign w17591 = ~w17589 & ~w17590;
assign w17592 = ~w16992 & w17023;
assign w17593 = pi01623 & ~w17592;
assign w17594 = ~pi02719 & ~w16992;
assign w17595 = w17023 & w17594;
assign w17596 = ~w17593 & ~w17595;
assign w17597 = pi01624 & ~w16962;
assign w17598 = ~pi02707 & w16962;
assign w17599 = ~w17597 & ~w17598;
assign w17600 = w16930 & w16969;
assign w17601 = ~w16905 & w17600;
assign w17602 = pi01625 & ~w17601;
assign w17603 = ~pi02711 & ~w16905;
assign w17604 = w17600 & w17603;
assign w17605 = ~w17602 & ~w17604;
assign w17606 = pi01626 & ~w17407;
assign w17607 = ~pi02703 & w17407;
assign w17608 = ~w17606 & ~w17607;
assign w17609 = w16921 & w17083;
assign w17610 = ~w16992 & w17609;
assign w17611 = pi01627 & ~w17610;
assign w17612 = ~pi02169 & w17610;
assign w17613 = ~w17611 & ~w17612;
assign w17614 = w16938 & w17582;
assign w17615 = ~w16992 & w17614;
assign w17616 = pi01628 & ~w17615;
assign w17617 = ~pi02167 & w17615;
assign w17618 = ~w17616 & ~w17617;
assign w17619 = pi01629 & ~w17584;
assign w17620 = ~pi02164 & ~w16992;
assign w17621 = w17583 & w17620;
assign w17622 = ~w17619 & ~w17621;
assign w17623 = pi01630 & ~w17429;
assign w17624 = ~pi02712 & w17429;
assign w17625 = ~w17623 & ~w17624;
assign w17626 = w16938 & w16967;
assign w17627 = ~w16928 & w17626;
assign w17628 = pi01631 & ~w17627;
assign w17629 = ~pi09954 & w17627;
assign w17630 = ~w17628 & ~w17629;
assign w17631 = w16940 & w17083;
assign w17632 = ~w16928 & w17631;
assign w17633 = pi01632 & ~w17632;
assign w17634 = ~pi09812 & w17632;
assign w17635 = ~w17633 & ~w17634;
assign w17636 = w16960 & w17189;
assign w17637 = ~w16892 & w17636;
assign w17638 = pi01633 & ~w17637;
assign w17639 = ~pi02709 & w17637;
assign w17640 = ~w17638 & ~w17639;
assign w17641 = w16930 & w16953;
assign w17642 = ~w16892 & w17641;
assign w17643 = pi01634 & ~w17642;
assign w17644 = ~pi02723 & w17642;
assign w17645 = ~w17643 & ~w17644;
assign w17646 = ~w16992 & w17505;
assign w17647 = pi01635 & ~w17646;
assign w17648 = ~pi02722 & w17646;
assign w17649 = ~w17647 & ~w17648;
assign w17650 = w16969 & w17582;
assign w17651 = ~w16992 & w17650;
assign w17652 = pi01636 & ~w17651;
assign w17653 = ~pi02164 & w17651;
assign w17654 = ~w17652 & ~w17653;
assign w17655 = pi01637 & ~w17315;
assign w17656 = ~pi02712 & w17315;
assign w17657 = ~w17655 & ~w17656;
assign w17658 = w17052 & w17136;
assign w17659 = ~w16905 & w17658;
assign w17660 = pi01638 & ~w17659;
assign w17661 = ~pi02716 & w17659;
assign w17662 = ~w17660 & ~w17661;
assign w17663 = w16908 & w16919;
assign w17664 = ~w16992 & w17663;
assign w17665 = pi01639 & ~w17664;
assign w17666 = w17532 & w17663;
assign w17667 = ~w17665 & ~w17666;
assign w17668 = w16960 & w17582;
assign w17669 = ~w16892 & w17668;
assign w17670 = pi01640 & ~w17669;
assign w17671 = ~pi02723 & ~w16892;
assign w17672 = w17668 & w17671;
assign w17673 = ~w17670 & ~w17672;
assign w17674 = ~w16905 & w17416;
assign w17675 = pi01641 & ~w17674;
assign w17676 = ~pi02716 & w17674;
assign w17677 = ~w17675 & ~w17676;
assign w17678 = pi01642 & ~w17610;
assign w17679 = ~pi02722 & w17610;
assign w17680 = ~w17678 & ~w17679;
assign w17681 = w16908 & w17052;
assign w17682 = ~w16905 & w17681;
assign w17683 = pi01643 & ~w17682;
assign w17684 = ~pi02170 & w17682;
assign w17685 = ~w17683 & ~w17684;
assign w17686 = w16953 & w17582;
assign w17687 = ~w16905 & w17686;
assign w17688 = pi01644 & ~w17687;
assign w17689 = ~pi02711 & w17687;
assign w17690 = ~w17688 & ~w17689;
assign w17691 = pi01645 & ~w17376;
assign w17692 = ~pi02712 & w17376;
assign w17693 = ~w17691 & ~w17692;
assign w17694 = w16947 & w16967;
assign w17695 = ~w16992 & w17694;
assign w17696 = pi01646 & ~w17695;
assign w17697 = ~pi02164 & w17695;
assign w17698 = ~w17696 & ~w17697;
assign w17699 = pi01647 & ~w17642;
assign w17700 = ~pi02706 & w17642;
assign w17701 = ~w17699 & ~w17700;
assign w17702 = ~w16992 & w17162;
assign w17703 = pi01648 & ~w17702;
assign w17704 = ~pi02719 & w17702;
assign w17705 = ~w17703 & ~w17704;
assign w17706 = ~w16892 & w17119;
assign w17707 = pi01649 & ~w17706;
assign w17708 = ~pi02723 & w17706;
assign w17709 = ~w17707 & ~w17708;
assign w17710 = w17059 & w17083;
assign w17711 = ~w16928 & w17710;
assign w17712 = pi01650 & ~w17711;
assign w17713 = ~pi09812 & w17711;
assign w17714 = ~w17712 & ~w17713;
assign w17715 = pi01651 & ~w17669;
assign w17716 = ~pi02707 & w17669;
assign w17717 = ~w17715 & ~w17716;
assign w17718 = w17005 & w17113;
assign w17719 = ~w16928 & w17718;
assign w17720 = pi01652 & ~w17719;
assign w17721 = ~pi02720 & w17719;
assign w17722 = ~w17720 & ~w17721;
assign w17723 = pi01653 & ~w17651;
assign w17724 = ~pi02703 & w17651;
assign w17725 = ~w17723 & ~w17724;
assign w17726 = ~w16992 & w17385;
assign w17727 = pi01654 & ~w17726;
assign w17728 = ~pi02721 & w17726;
assign w17729 = ~w17727 & ~w17728;
assign w17730 = ~w16992 & w17017;
assign w17731 = pi01655 & ~w17730;
assign w17732 = ~pi02721 & w17730;
assign w17733 = ~w17731 & ~w17732;
assign w17734 = w16967 & w16983;
assign w17735 = ~w16992 & w17734;
assign w17736 = pi01656 & ~w17735;
assign w17737 = ~pi02169 & w17735;
assign w17738 = ~w17736 & ~w17737;
assign w17739 = w16969 & w17182;
assign w17740 = ~w16905 & w17739;
assign w17741 = pi01657 & ~w17740;
assign w17742 = ~pi02714 & ~w16905;
assign w17743 = w17739 & w17742;
assign w17744 = ~w17741 & ~w17743;
assign w17745 = ~w16905 & w17436;
assign w17746 = pi01658 & ~w17745;
assign w17747 = ~pi02711 & w17745;
assign w17748 = ~w17746 & ~w17747;
assign w17749 = w16919 & w17136;
assign w17750 = ~w16905 & w17749;
assign w17751 = pi01659 & ~w17750;
assign w17752 = ~pi02716 & w17750;
assign w17753 = ~w17751 & ~w17752;
assign w17754 = w17005 & w17182;
assign w17755 = ~w16905 & w17754;
assign w17756 = pi01660 & ~w17755;
assign w17757 = ~pi02170 & w17755;
assign w17758 = ~w17756 & ~w17757;
assign w17759 = pi01661 & ~w17592;
assign w17760 = w17023 & w17586;
assign w17761 = ~w17759 & ~w17760;
assign w17762 = w17016 & w17059;
assign w17763 = ~w16905 & w17762;
assign w17764 = pi01662 & ~w17763;
assign w17765 = ~pi02712 & w17763;
assign w17766 = ~w17764 & ~w17765;
assign w17767 = w16938 & w17374;
assign w17768 = ~w16905 & w17767;
assign w17769 = pi01663 & ~w17768;
assign w17770 = ~pi02715 & w17768;
assign w17771 = ~w17769 & ~w17770;
assign w17772 = pi01664 & ~w17706;
assign w17773 = ~pi02705 & w17706;
assign w17774 = ~w17772 & ~w17773;
assign w17775 = w16919 & w17037;
assign w17776 = ~w16905 & w17775;
assign w17777 = pi01665 & ~w17776;
assign w17778 = ~pi02714 & w17776;
assign w17779 = ~w17777 & ~w17778;
assign w17780 = ~w16892 & w17416;
assign w17781 = pi01666 & ~w17780;
assign w17782 = w17416 & w17671;
assign w17783 = ~w17781 & ~w17782;
assign w17784 = pi01667 & ~w17776;
assign w17785 = w17603 & w17775;
assign w17786 = ~w17784 & ~w17785;
assign w17787 = pi01668 & ~w17627;
assign w17788 = ~pi09848 & w17627;
assign w17789 = ~w17787 & ~w17788;
assign w17790 = ~w16992 & w17200;
assign w17791 = pi01669 & ~w17790;
assign w17792 = ~pi02719 & w17790;
assign w17793 = ~w17791 & ~w17792;
assign w17794 = ~w16992 & w17686;
assign w17795 = pi01670 & ~w17794;
assign w17796 = ~pi02167 & w17794;
assign w17797 = ~w17795 & ~w17796;
assign w17798 = ~w16905 & w17450;
assign w17799 = pi01671 & ~w17798;
assign w17800 = ~pi02714 & w17798;
assign w17801 = ~w17799 & ~w17800;
assign w17802 = pi01672 & ~w17232;
assign w17803 = ~pi02178 & w17232;
assign w17804 = ~w17802 & ~w17803;
assign w17805 = pi01673 & ~w17674;
assign w17806 = ~pi02714 & w17674;
assign w17807 = ~w17805 & ~w17806;
assign w17808 = w16977 & w17083;
assign w17809 = ~w16992 & w17808;
assign w17810 = pi01674 & ~w17809;
assign w17811 = ~pi02721 & ~w16992;
assign w17812 = w17808 & w17811;
assign w17813 = ~w17810 & ~w17812;
assign w17814 = w16919 & w16940;
assign w17815 = ~w16905 & w17814;
assign w17816 = pi01675 & ~w17815;
assign w17817 = ~pi02711 & w17815;
assign w17818 = ~w17816 & ~w17817;
assign w17819 = pi01676 & ~w17809;
assign w17820 = ~pi02703 & w17809;
assign w17821 = ~w17819 & ~w17820;
assign w17822 = w16940 & w17052;
assign w17823 = ~w16905 & w17822;
assign w17824 = pi01677 & ~w17823;
assign w17825 = w17603 & w17822;
assign w17826 = ~w17824 & ~w17825;
assign w17827 = ~w16892 & w17461;
assign w17828 = pi01678 & ~w17827;
assign w17829 = ~pi02706 & w17827;
assign w17830 = ~w17828 & ~w17829;
assign w17831 = pi01679 & ~w17232;
assign w17832 = ~pi09961 & w17232;
assign w17833 = ~w17831 & ~w17832;
assign w17834 = pi01680 & ~w17815;
assign w17835 = ~pi02714 & w17815;
assign w17836 = ~w17834 & ~w17835;
assign w17837 = w16898 & w16938;
assign w17838 = ~w16905 & w17837;
assign w17839 = pi01681 & ~w17838;
assign w17840 = ~pi02715 & w17838;
assign w17841 = ~w17839 & ~w17840;
assign w17842 = pi01682 & ~w17750;
assign w17843 = ~pi02170 & w17750;
assign w17844 = ~w17842 & ~w17843;
assign w17845 = pi01683 & ~w17566;
assign w17846 = ~pi02719 & w17566;
assign w17847 = ~w17845 & ~w17846;
assign w17848 = w16970 & ~w16992;
assign w17849 = pi01684 & ~w17848;
assign w17850 = ~pi02703 & w17848;
assign w17851 = ~w17849 & ~w17850;
assign w17852 = pi01685 & ~w17711;
assign w17853 = ~pi02720 & w17711;
assign w17854 = ~w17852 & ~w17853;
assign w17855 = w16953 & w17113;
assign w17856 = ~w16892 & w17855;
assign w17857 = pi01686 & ~w17856;
assign w17858 = ~pi02709 & w17856;
assign w17859 = ~w17857 & ~w17858;
assign w17860 = pi01687 & ~w17695;
assign w17861 = ~pi02721 & w17695;
assign w17862 = ~w17860 & ~w17861;
assign w17863 = pi01688 & ~w17566;
assign w17864 = ~pi02164 & w17566;
assign w17865 = ~w17863 & ~w17864;
assign w17866 = ~w16992 & w17681;
assign w17867 = pi01689 & ~w17866;
assign w17868 = w17586 & w17681;
assign w17869 = ~w17867 & ~w17868;
assign w17870 = pi01690 & ~w17735;
assign w17871 = ~pi02703 & w17735;
assign w17872 = ~w17870 & ~w17871;
assign w17873 = ~w16992 & w17172;
assign w17874 = pi01691 & ~w17873;
assign w17875 = w17172 & w17594;
assign w17876 = ~w17874 & ~w17875;
assign w17877 = pi01692 & ~w17682;
assign w17878 = w16973 & w17681;
assign w17879 = ~w17877 & ~w17878;
assign w17880 = pi01693 & ~w17856;
assign w17881 = ~pi02160 & w17856;
assign w17882 = ~w17880 & ~w17881;
assign w17883 = pi01694 & ~w17496;
assign w17884 = ~pi02704 & w17496;
assign w17885 = ~w17883 & ~w17884;
assign w17886 = pi01695 & ~w17763;
assign w17887 = ~pi02716 & w17763;
assign w17888 = ~w17886 & ~w17887;
assign w17889 = ~w16992 & w17445;
assign w17890 = pi01696 & ~w17889;
assign w17891 = ~pi02164 & w17889;
assign w17892 = ~w17890 & ~w17891;
assign w17893 = pi01697 & ~w17798;
assign w17894 = ~pi02711 & w17798;
assign w17895 = ~w17893 & ~w17894;
assign w17896 = ~w16928 & w17390;
assign w17897 = pi01698 & ~w17896;
assign w17898 = w17311 & w17390;
assign w17899 = ~w17897 & ~w17898;
assign w17900 = ~w16992 & w17084;
assign w17901 = pi01699 & ~w17900;
assign w17902 = ~pi02703 & w17900;
assign w17903 = ~w17901 & ~w17902;
assign w17904 = pi01700 & ~w17889;
assign w17905 = ~pi02721 & w17889;
assign w17906 = ~w17904 & ~w17905;
assign w17907 = w17113 & w17124;
assign w17908 = ~w16905 & w17907;
assign w17909 = pi01701 & ~w17908;
assign w17910 = w17020 & w17907;
assign w17911 = ~w17909 & ~w17910;
assign w17912 = w16908 & w16947;
assign w17913 = ~w16928 & w17912;
assign w17914 = pi01702 & ~w17913;
assign w17915 = w17513 & w17912;
assign w17916 = ~w17914 & ~w17915;
assign w17917 = w16985 & w17083;
assign w17918 = ~w16892 & w17917;
assign w17919 = pi01703 & ~w17918;
assign w17920 = ~pi02709 & w17918;
assign w17921 = ~w17919 & ~w17920;
assign w17922 = w16938 & w17189;
assign w17923 = ~w16892 & w17922;
assign w17924 = pi01704 & ~w17923;
assign w17925 = ~pi02706 & ~w16892;
assign w17926 = w17922 & w17925;
assign w17927 = ~w17924 & ~w17926;
assign w17928 = pi01705 & ~w17561;
assign w17929 = ~pi02713 & ~w16905;
assign w17930 = w17047 & w17929;
assign w17931 = ~w17928 & ~w17930;
assign w17932 = pi01706 & ~w17664;
assign w17933 = ~pi02164 & w17664;
assign w17934 = ~w17932 & ~w17933;
assign w17935 = pi01707 & ~w17601;
assign w17936 = ~pi02713 & w17601;
assign w17937 = ~w17935 & ~w17936;
assign w17938 = w16983 & w17059;
assign w17939 = ~w16928 & w17938;
assign w17940 = pi01708 & ~w17939;
assign w17941 = ~pi09812 & w17939;
assign w17942 = ~w17940 & ~w17941;
assign w17943 = pi01709 & ~w17154;
assign w17944 = ~pi09812 & w17154;
assign w17945 = ~w17943 & ~w17944;
assign w17946 = ~w16905 & w17259;
assign w17947 = pi01710 & ~w17946;
assign w17948 = w17259 & w17742;
assign w17949 = ~w17947 & ~w17948;
assign w17950 = ~w16992 & w17767;
assign w17951 = pi01711 & ~w17950;
assign w17952 = ~pi02167 & w17950;
assign w17953 = ~w17951 & ~w17952;
assign w17954 = ~w16905 & w17411;
assign w17955 = pi01712 & ~w17954;
assign w17956 = ~pi02715 & w17954;
assign w17957 = ~w17955 & ~w17956;
assign w17958 = pi01713 & ~w17664;
assign w17959 = ~pi02721 & w17664;
assign w17960 = ~w17958 & ~w17959;
assign w17961 = ~w16905 & w17663;
assign w17962 = pi01714 & ~w17961;
assign w17963 = ~pi02717 & w17961;
assign w17964 = ~w17962 & ~w17963;
assign w17965 = w16947 & w16977;
assign w17966 = ~w16928 & w17965;
assign w17967 = pi01715 & ~w17966;
assign w17968 = ~pi09954 & w17966;
assign w17969 = ~w17967 & ~w17968;
assign w17970 = pi01716 & ~w17961;
assign w17971 = ~pi02714 & w17961;
assign w17972 = ~w17970 & ~w17971;
assign w17973 = ~w16892 & w17631;
assign w17974 = pi01717 & ~w17973;
assign w17975 = ~pi02706 & w17973;
assign w17976 = ~w17974 & ~w17975;
assign w17977 = w16898 & w17016;
assign w17978 = ~w16928 & w17977;
assign w17979 = pi01718 & ~w17978;
assign w17980 = ~pi09962 & w17978;
assign w17981 = ~w17979 & ~w17980;
assign w17982 = pi01719 & ~w17552;
assign w17983 = ~pi02722 & w17552;
assign w17984 = ~w17982 & ~w17983;
assign w17985 = pi01720 & ~w17790;
assign w17986 = w17200 & w17586;
assign w17987 = ~w17985 & ~w17986;
assign w17988 = ~w16928 & w17808;
assign w17989 = pi01721 & ~w17988;
assign w17990 = ~pi09962 & w17988;
assign w17991 = ~w17989 & ~w17990;
assign w17992 = ~w16992 & w17366;
assign w17993 = pi01722 & ~w17992;
assign w17994 = w17366 & w17594;
assign w17995 = ~w17993 & ~w17994;
assign w17996 = w16940 & w16993;
assign w17997 = ~w16992 & w17996;
assign w17998 = pi01723 & ~w17997;
assign w17999 = w17811 & w17996;
assign w18000 = ~w17998 & ~w17999;
assign w18001 = w16898 & w16953;
assign w18002 = ~w16905 & w18001;
assign w18003 = pi01724 & ~w18002;
assign w18004 = ~pi02713 & w18002;
assign w18005 = ~w18003 & ~w18004;
assign w18006 = pi01725 & ~w17417;
assign w18007 = ~pi02720 & w17417;
assign w18008 = ~w18006 & ~w18007;
assign w18009 = w17083 & w17374;
assign w18010 = ~w16992 & w18009;
assign w18011 = pi01726 & ~w18010;
assign w18012 = ~pi02167 & w18010;
assign w18013 = ~w18011 & ~w18012;
assign w18014 = ~w16892 & w17450;
assign w18015 = pi01727 & ~w18014;
assign w18016 = ~pi02706 & w18014;
assign w18017 = ~w18015 & ~w18016;
assign w18018 = ~w16928 & w16994;
assign w18019 = pi01728 & ~w18018;
assign w18020 = ~pi09954 & w18018;
assign w18021 = ~w18019 & ~w18020;
assign w18022 = w16930 & w16993;
assign w18023 = ~w16905 & w18022;
assign w18024 = pi01729 & ~w18023;
assign w18025 = w17603 & w18022;
assign w18026 = ~w18024 & ~w18025;
assign w18027 = w16947 & w17059;
assign w18028 = ~w16928 & w18027;
assign w18029 = pi01730 & ~w18028;
assign w18030 = ~pi09962 & w18028;
assign w18031 = ~w18029 & ~w18030;
assign w18032 = w17016 & w17189;
assign w18033 = ~w16992 & w18032;
assign w18034 = pi01731 & ~w18033;
assign w18035 = w17620 & w18032;
assign w18036 = ~w18034 & ~w18035;
assign w18037 = pi01732 & ~w17548;
assign w18038 = ~pi02716 & w17548;
assign w18039 = ~w18037 & ~w18038;
assign w18040 = w17038 & w17374;
assign w18041 = ~w16892 & w18040;
assign w18042 = pi01733 & ~w18041;
assign w18043 = ~pi02709 & w18041;
assign w18044 = ~w18042 & ~w18043;
assign w18045 = pi01734 & ~w18028;
assign w18046 = ~pi02178 & w18028;
assign w18047 = ~w18045 & ~w18046;
assign w18048 = pi01735 & ~w17988;
assign w18049 = ~pi02704 & w17988;
assign w18050 = ~w18048 & ~w18049;
assign w18051 = w17124 & w17374;
assign w18052 = ~w16905 & w18051;
assign w18053 = pi01736 & ~w18052;
assign w18054 = w17020 & w18051;
assign w18055 = ~w18053 & ~w18054;
assign w18056 = w16930 & w17083;
assign w18057 = ~w16905 & w18056;
assign w18058 = pi01737 & ~w18057;
assign w18059 = ~pi02715 & ~w16905;
assign w18060 = w18056 & w18059;
assign w18061 = ~w18058 & ~w18060;
assign w18062 = ~w16928 & w17098;
assign w18063 = pi01738 & ~w18062;
assign w18064 = ~pi09812 & w18062;
assign w18065 = ~w18063 & ~w18064;
assign w18066 = pi01739 & ~w18041;
assign w18067 = ~pi02707 & ~w16892;
assign w18068 = w18040 & w18067;
assign w18069 = ~w18066 & ~w18068;
assign w18070 = w17083 & w17189;
assign w18071 = ~w16905 & w18070;
assign w18072 = pi01740 & ~w18071;
assign w18073 = ~pi02712 & w18071;
assign w18074 = ~w18072 & ~w18073;
assign w18075 = ~w16905 & w17305;
assign w18076 = pi01741 & ~w18075;
assign w18077 = ~pi02715 & w18075;
assign w18078 = ~w18076 & ~w18077;
assign w18079 = ~w16905 & w17264;
assign w18080 = pi01742 & ~w18079;
assign w18081 = ~pi02716 & w18079;
assign w18082 = ~w18080 & ~w18081;
assign w18083 = pi01743 & ~w17695;
assign w18084 = ~pi02703 & w17695;
assign w18085 = ~w18083 & ~w18084;
assign w18086 = ~w16992 & w17739;
assign w18087 = pi01744 & ~w18086;
assign w18088 = ~pi02719 & w18086;
assign w18089 = ~w18087 & ~w18088;
assign w18090 = ~w16892 & w17500;
assign w18091 = pi01745 & ~w18090;
assign w18092 = ~pi02709 & ~w16892;
assign w18093 = w17500 & w18092;
assign w18094 = ~w18091 & ~w18093;
assign w18095 = pi01746 & ~w18057;
assign w18096 = ~pi02712 & w18057;
assign w18097 = ~w18095 & ~w18096;
assign w18098 = pi01747 & ~w17973;
assign w18099 = ~pi02723 & w17973;
assign w18100 = ~w18098 & ~w18099;
assign w18101 = ~w16905 & w17495;
assign w18102 = pi01748 & ~w18101;
assign w18103 = ~pi02711 & w18101;
assign w18104 = ~w18102 & ~w18103;
assign w18105 = ~w16928 & w17039;
assign w18106 = pi01749 & ~w18105;
assign w18107 = ~pi09812 & w18105;
assign w18108 = ~w18106 & ~w18107;
assign w18109 = pi01750 & ~w17966;
assign w18110 = w17186 & w17965;
assign w18111 = ~w18109 & ~w18110;
assign w18112 = ~w16892 & w17565;
assign w18113 = pi01751 & ~w18112;
assign w18114 = ~pi02710 & w18112;
assign w18115 = ~w18113 & ~w18114;
assign w18116 = w17083 & w17582;
assign w18117 = ~w16905 & w18116;
assign w18118 = pi01752 & ~w18117;
assign w18119 = ~pi02712 & w18117;
assign w18120 = ~w18118 & ~w18119;
assign w18121 = pi01753 & ~w18117;
assign w18122 = w18059 & w18116;
assign w18123 = ~w18121 & ~w18122;
assign w18124 = pi01754 & ~w18033;
assign w18125 = ~pi02169 & w18033;
assign w18126 = ~w18124 & ~w18125;
assign w18127 = ~w16905 & w17190;
assign w18128 = pi01755 & ~w18127;
assign w18129 = w17190 & w17742;
assign w18130 = ~w18128 & ~w18129;
assign w18131 = pi01756 & ~w17557;
assign w18132 = ~pi02160 & w17557;
assign w18133 = ~w18131 & ~w18132;
assign w18134 = ~w16992 & w17183;
assign w18135 = pi01757 & ~w18134;
assign w18136 = ~pi02167 & w18134;
assign w18137 = ~w18135 & ~w18136;
assign w18138 = ~w16928 & w17445;
assign w18139 = pi01758 & ~w18138;
assign w18140 = w17186 & w17445;
assign w18141 = ~w18139 & ~w18140;
assign w18142 = ~w16892 & w17177;
assign w18143 = pi01759 & ~w18142;
assign w18144 = ~pi02710 & w18142;
assign w18145 = ~w18143 & ~w18144;
assign w18146 = w16969 & w17374;
assign w18147 = ~w16905 & w18146;
assign w18148 = pi01760 & ~w18147;
assign w18149 = w17020 & w18146;
assign w18150 = ~w18148 & ~w18149;
assign w18151 = ~w16992 & w17053;
assign w18152 = pi01761 & ~w18151;
assign w18153 = ~pi02167 & w18151;
assign w18154 = ~w18152 & ~w18153;
assign w18155 = w16930 & w17038;
assign w18156 = ~w16905 & w18155;
assign w18157 = pi01762 & ~w18156;
assign w18158 = w18059 & w18155;
assign w18159 = ~w18157 & ~w18158;
assign w18160 = ~w16928 & w17137;
assign w18161 = pi01763 & ~w18160;
assign w18162 = ~pi09954 & w18160;
assign w18163 = ~w18161 & ~w18162;
assign w18164 = ~w16892 & w17718;
assign w18165 = pi01764 & ~w18164;
assign w18166 = ~pi02710 & w18164;
assign w18167 = ~w18165 & ~w18166;
assign w18168 = pi01765 & ~w17950;
assign w18169 = ~pi02169 & w17950;
assign w18170 = ~w18168 & ~w18169;
assign w18171 = pi01766 & ~w18160;
assign w18172 = ~pi09848 & w18160;
assign w18173 = ~w18171 & ~w18172;
assign w18174 = pi01767 & ~w18156;
assign w18175 = w17020 & w18155;
assign w18176 = ~w18174 & ~w18175;
assign w18177 = w17005 & w17374;
assign w18178 = ~w16892 & w18177;
assign w18179 = pi01768 & ~w18178;
assign w18180 = ~pi02710 & w18178;
assign w18181 = ~w18179 & ~w18180;
assign w18182 = ~w16992 & w17231;
assign w18183 = pi01769 & ~w18182;
assign w18184 = ~pi02719 & w18182;
assign w18185 = ~w18183 & ~w18184;
assign w18186 = w16960 & w17136;
assign w18187 = ~w16992 & w18186;
assign w18188 = pi01770 & ~w18187;
assign w18189 = ~pi02703 & w18187;
assign w18190 = ~w18188 & ~w18189;
assign w18191 = pi01771 & ~w18002;
assign w18192 = ~pi02711 & w18002;
assign w18193 = ~w18191 & ~w18192;
assign w18194 = ~w16928 & w17017;
assign w18195 = pi01772 & ~w18194;
assign w18196 = ~pi09954 & w18194;
assign w18197 = ~w18195 & ~w18196;
assign w18198 = pi01773 & ~w17719;
assign w18199 = ~pi09812 & w17719;
assign w18200 = ~w18198 & ~w18199;
assign w18201 = pi01774 & ~w18010;
assign w18202 = ~pi02703 & w18010;
assign w18203 = ~w18201 & ~w18202;
assign w18204 = pi01775 & ~w18079;
assign w18205 = ~pi02170 & w18079;
assign w18206 = ~w18204 & ~w18205;
assign w18207 = pi01776 & ~w18134;
assign w18208 = ~pi02721 & w18134;
assign w18209 = ~w18207 & ~w18208;
assign w18210 = ~w16928 & w17028;
assign w18211 = pi01777 & ~w18210;
assign w18212 = ~pi02178 & w18210;
assign w18213 = ~w18211 & ~w18212;
assign w18214 = pi01778 & ~w18010;
assign w18215 = ~pi02718 & w18010;
assign w18216 = ~w18214 & ~w18215;
assign w18217 = w17016 & w17136;
assign w18218 = ~w16905 & w18217;
assign w18219 = pi01779 & ~w18218;
assign w18220 = ~pi02712 & w18218;
assign w18221 = ~w18219 & ~w18220;
assign w18222 = ~w16892 & w16999;
assign w18223 = pi01780 & ~w18222;
assign w18224 = ~pi02723 & w18222;
assign w18225 = ~w18223 & ~w18224;
assign w18226 = pi01781 & ~w18164;
assign w18227 = ~pi02706 & w18164;
assign w18228 = ~w18226 & ~w18227;
assign w18229 = ~w16905 & w17254;
assign w18230 = pi01782 & ~w18229;
assign w18231 = ~pi02716 & w18229;
assign w18232 = ~w18230 & ~w18231;
assign w18233 = pi01783 & ~w18178;
assign w18234 = ~pi02160 & ~w16892;
assign w18235 = w18177 & w18234;
assign w18236 = ~w18233 & ~w18235;
assign w18237 = pi01784 & ~w18151;
assign w18238 = w17053 & w17620;
assign w18239 = ~w18237 & ~w18238;
assign w18240 = pi01785 & ~w18138;
assign w18241 = ~pi09954 & w18138;
assign w18242 = ~w18240 & ~w18241;
assign w18243 = ~w16892 & w17614;
assign w18244 = pi01786 & ~w18243;
assign w18245 = w17614 & w17671;
assign w18246 = ~w18244 & ~w18245;
assign w18247 = w16930 & w16983;
assign w18248 = ~w16905 & w18247;
assign w18249 = pi01787 & ~w18248;
assign w18250 = ~pi02715 & w18248;
assign w18251 = ~w18249 & ~w18250;
assign w18252 = ~w16928 & w18051;
assign w18253 = pi01788 & ~w18252;
assign w18254 = ~pi09954 & w18252;
assign w18255 = ~w18253 & ~w18254;
assign w18256 = w16961 & ~w16992;
assign w18257 = pi01789 & ~w18256;
assign w18258 = ~pi02718 & w18256;
assign w18259 = ~w18257 & ~w18258;
assign w18260 = pi01790 & ~w18222;
assign w18261 = ~pi02705 & w18222;
assign w18262 = ~w18260 & ~w18261;
assign w18263 = w17038 & w17189;
assign w18264 = ~w16905 & w18263;
assign w18265 = pi01791 & ~w18264;
assign w18266 = ~pi02712 & w18264;
assign w18267 = ~w18265 & ~w18266;
assign w18268 = pi01792 & ~w18256;
assign w18269 = ~pi02167 & w18256;
assign w18270 = ~w18268 & ~w18269;
assign w18271 = ~w16892 & w17686;
assign w18272 = pi01793 & ~w18271;
assign w18273 = ~pi02706 & w18271;
assign w18274 = ~w18272 & ~w18273;
assign w18275 = pi01794 & ~w17040;
assign w18276 = ~pi02709 & w17040;
assign w18277 = ~w18275 & ~w18276;
assign w18278 = w16938 & w17037;
assign w18279 = ~w16905 & w18278;
assign w18280 = pi01795 & ~w18279;
assign w18281 = ~pi02711 & w18279;
assign w18282 = ~w18280 & ~w18281;
assign w18283 = ~w16992 & w17344;
assign w18284 = pi01796 & ~w18283;
assign w18285 = ~pi02703 & w18283;
assign w18286 = ~w18284 & ~w18285;
assign w18287 = ~w16892 & w17284;
assign w18288 = pi01797 & ~w18287;
assign w18289 = ~pi02710 & w18287;
assign w18290 = ~w18288 & ~w18289;
assign w18291 = w16947 & w17189;
assign w18292 = ~w16928 & w18291;
assign w18293 = pi01798 & ~w18292;
assign w18294 = ~pi02720 & w18292;
assign w18295 = ~w18293 & ~w18294;
assign w18296 = ~w16928 & w18056;
assign w18297 = pi01799 & ~w18296;
assign w18298 = ~pi09954 & w18296;
assign w18299 = ~w18297 & ~w18298;
assign w18300 = w17124 & w17182;
assign w18301 = ~w16905 & w18300;
assign w18302 = pi01800 & ~w18301;
assign w18303 = w17020 & w18300;
assign w18304 = ~w18302 & ~w18303;
assign w18305 = pi01801 & ~w18151;
assign w18306 = ~pi02721 & w18151;
assign w18307 = ~w18305 & ~w18306;
assign w18308 = w17038 & w17582;
assign w18309 = ~w16905 & w18308;
assign w18310 = pi01802 & ~w18309;
assign w18311 = ~pi02715 & w18309;
assign w18312 = ~w18310 & ~w18311;
assign w18313 = pi01803 & ~w18296;
assign w18314 = ~pi09848 & w18296;
assign w18315 = ~w18313 & ~w18314;
assign w18316 = pi01804 & ~w18271;
assign w18317 = ~pi02723 & w18271;
assign w18318 = ~w18316 & ~w18317;
assign w18319 = ~w16905 & w17510;
assign w18320 = pi01805 & ~w18319;
assign w18321 = ~pi02712 & w18319;
assign w18322 = ~w18320 & ~w18321;
assign w18323 = pi01806 & ~w18287;
assign w18324 = ~pi02160 & w18287;
assign w18325 = ~w18323 & ~w18324;
assign w18326 = ~w16928 & w18146;
assign w18327 = pi01807 & ~w18326;
assign w18328 = ~pi09954 & w18326;
assign w18329 = ~w18327 & ~w18328;
assign w18330 = ~w16992 & w18177;
assign w18331 = pi01808 & ~w18330;
assign w18332 = ~pi02164 & w18330;
assign w18333 = ~w18331 & ~w18332;
assign w18334 = pi01809 & ~w18075;
assign w18335 = ~pi02713 & w18075;
assign w18336 = ~w18334 & ~w18335;
assign w18337 = ~w16928 & w18116;
assign w18338 = pi01810 & ~w18337;
assign w18339 = ~pi09954 & w18337;
assign w18340 = ~w18338 & ~w18339;
assign w18341 = pi01811 & ~w18309;
assign w18342 = ~pi02712 & w18309;
assign w18343 = ~w18341 & ~w18342;
assign w18344 = ~w16928 & w18070;
assign w18345 = pi01812 & ~w18344;
assign w18346 = ~pi09954 & w18344;
assign w18347 = ~w18345 & ~w18346;
assign w18348 = w17124 & w17189;
assign w18349 = ~w16928 & w18348;
assign w18350 = pi01813 & ~w18349;
assign w18351 = ~pi02720 & w18349;
assign w18352 = ~w18350 & ~w18351;
assign w18353 = pi01814 & ~w18151;
assign w18354 = ~pi02703 & w18151;
assign w18355 = ~w18353 & ~w18354;
assign w18356 = pi01815 & ~w17085;
assign w18357 = ~pi09962 & w17085;
assign w18358 = ~w18356 & ~w18357;
assign w18359 = pi01816 & ~w18182;
assign w18360 = ~pi02169 & w18182;
assign w18361 = ~w18359 & ~w18360;
assign w18362 = ~w16892 & w16912;
assign w18363 = pi01817 & ~w18362;
assign w18364 = ~pi02710 & ~w16892;
assign w18365 = w16912 & w18364;
assign w18366 = ~w18363 & ~w18365;
assign w18367 = pi01818 & ~w17206;
assign w18368 = ~pi02719 & w17206;
assign w18369 = ~w18367 & ~w18368;
assign w18370 = w16921 & w16983;
assign w18371 = ~w16892 & w18370;
assign w18372 = pi01819 & ~w18371;
assign w18373 = ~pi02705 & w18371;
assign w18374 = ~w18372 & ~w18373;
assign w18375 = pi01820 & ~w18362;
assign w18376 = ~pi02705 & w18362;
assign w18377 = ~w18375 & ~w18376;
assign w18378 = ~w16892 & w17710;
assign w18379 = pi01821 & ~w18378;
assign w18380 = ~pi02706 & w18378;
assign w18381 = ~w18379 & ~w18380;
assign w18382 = ~w16905 & w17631;
assign w18383 = pi01822 & ~w18382;
assign w18384 = w17631 & w17929;
assign w18385 = ~w18383 & ~w18384;
assign w18386 = pi01823 & ~w18337;
assign w18387 = ~pi09848 & w18337;
assign w18388 = ~w18386 & ~w18387;
assign w18389 = ~w16892 & w16978;
assign w18390 = pi01824 & ~w18389;
assign w18391 = ~pi02723 & w18389;
assign w18392 = ~w18390 & ~w18391;
assign w18393 = ~w16892 & w17767;
assign w18394 = pi01825 & ~w18393;
assign w18395 = w17767 & w17925;
assign w18396 = ~w18394 & ~w18395;
assign w18397 = pi01826 & ~w18330;
assign w18398 = ~pi02703 & w18330;
assign w18399 = ~w18397 & ~w18398;
assign w18400 = ~w16992 & w17028;
assign w18401 = pi01827 & ~w18400;
assign w18402 = ~pi02167 & w18400;
assign w18403 = ~w18401 & ~w18402;
assign w18404 = ~w16928 & w18308;
assign w18405 = pi01828 & ~w18404;
assign w18406 = ~pi09848 & w18404;
assign w18407 = ~w18405 & ~w18406;
assign w18408 = pi01829 & ~w17552;
assign w18409 = ~pi02718 & w17552;
assign w18410 = ~w18408 & ~w18409;
assign w18411 = ~w16892 & w18022;
assign w18412 = pi01830 & ~w18411;
assign w18413 = ~pi02710 & w18411;
assign w18414 = ~w18412 & ~w18413;
assign w18415 = pi01831 & ~w18127;
assign w18416 = ~pi02712 & w18127;
assign w18417 = ~w18415 & ~w18416;
assign w18418 = ~w16905 & w17300;
assign w18419 = pi01832 & ~w18418;
assign w18420 = ~pi02717 & w18418;
assign w18421 = ~w18419 & ~w18420;
assign w18422 = w16921 & w16993;
assign w18423 = ~w16892 & w18422;
assign w18424 = pi01833 & ~w18423;
assign w18425 = ~pi02723 & w18423;
assign w18426 = ~w18424 & ~w18425;
assign w18427 = ~w16928 & w16970;
assign w18428 = pi01834 & ~w18427;
assign w18429 = ~pi02704 & w18427;
assign w18430 = ~w18428 & ~w18429;
assign w18431 = w16930 & w17005;
assign w18432 = ~w16905 & w18431;
assign w18433 = pi01835 & ~w18432;
assign w18434 = ~pi02712 & w18432;
assign w18435 = ~w18433 & ~w18434;
assign w18436 = pi01836 & ~w18389;
assign w18437 = ~pi02705 & w18389;
assign w18438 = ~w18436 & ~w18437;
assign w18439 = ~w16928 & w18155;
assign w18440 = pi01837 & ~w18439;
assign w18441 = ~pi09954 & w18439;
assign w18442 = ~w18440 & ~w18441;
assign w18443 = pi01838 & ~w18105;
assign w18444 = ~pi09954 & w18105;
assign w18445 = ~w18443 & ~w18444;
assign w18446 = pi01839 & ~w18423;
assign w18447 = ~pi02705 & w18423;
assign w18448 = ~w18446 & ~w18447;
assign w18449 = w16938 & w16977;
assign w18450 = ~w16928 & w18449;
assign w18451 = pi01840 & ~w18450;
assign w18452 = ~pi09812 & w18450;
assign w18453 = ~w18451 & ~w18452;
assign w18454 = w16898 & w16960;
assign w18455 = ~w16892 & w18454;
assign w18456 = pi01841 & ~w18455;
assign w18457 = w17925 & w18454;
assign w18458 = ~w18456 & ~w18457;
assign w18459 = pi01842 & ~w18439;
assign w18460 = ~pi09848 & w18439;
assign w18461 = ~w18459 & ~w18460;
assign w18462 = pi01843 & ~w18411;
assign w18463 = ~pi02723 & w18411;
assign w18464 = ~w18462 & ~w18463;
assign w18465 = pi01844 & ~w18292;
assign w18466 = ~pi09812 & w18292;
assign w18467 = ~w18465 & ~w18466;
assign w18468 = w16969 & w17059;
assign w18469 = ~w16928 & w18468;
assign w18470 = pi01845 & ~w18469;
assign w18471 = ~pi09812 & w18469;
assign w18472 = ~w18470 & ~w18471;
assign w18473 = pi01846 & ~w18349;
assign w18474 = ~pi09812 & w18349;
assign w18475 = ~w18473 & ~w18474;
assign w18476 = pi01847 & ~w18014;
assign w18477 = ~pi02708 & w18014;
assign w18478 = ~w18476 & ~w18477;
assign w18479 = pi01848 & ~w18248;
assign w18480 = w17020 & w18247;
assign w18481 = ~w18479 & ~w18480;
assign w18482 = ~w16928 & w18263;
assign w18483 = pi01849 & ~w18482;
assign w18484 = ~pi09954 & w18482;
assign w18485 = ~w18483 & ~w18484;
assign w18486 = pi01850 & ~w18400;
assign w18487 = ~pi02703 & w18400;
assign w18488 = ~w18486 & ~w18487;
assign w18489 = pi01851 & ~w17997;
assign w18490 = ~pi02169 & w17997;
assign w18491 = ~w18489 & ~w18490;
assign w18492 = w16986 & ~w16992;
assign w18493 = pi01852 & ~w18492;
assign w18494 = ~pi02718 & w18492;
assign w18495 = ~w18493 & ~w18494;
assign w18496 = ~w16892 & w17436;
assign w18497 = pi01853 & ~w18496;
assign w18498 = ~pi02706 & w18496;
assign w18499 = ~w18497 & ~w18498;
assign w18500 = pi01854 & ~w18404;
assign w18501 = w17513 & w18308;
assign w18502 = ~w18500 & ~w18501;
assign w18503 = ~w16992 & w18051;
assign w18504 = pi01855 & ~w18503;
assign w18505 = ~pi02164 & w18503;
assign w18506 = ~w18504 & ~w18505;
assign w18507 = ~w16905 & w17668;
assign w18508 = pi01856 & ~w18507;
assign w18509 = ~pi02716 & w18507;
assign w18510 = ~w18508 & ~w18509;
assign w18511 = pi01857 & ~w17506;
assign w18512 = w17193 & w17505;
assign w18513 = ~w18511 & ~w18512;
assign w18514 = ~w16928 & w17540;
assign w18515 = pi01858 & ~w18514;
assign w18516 = ~pi02720 & w18514;
assign w18517 = ~w18515 & ~w18516;
assign w18518 = ~w16992 & w17636;
assign w18519 = pi01859 & ~w18518;
assign w18520 = ~pi02722 & w18518;
assign w18521 = ~w18519 & ~w18520;
assign w18522 = ~w16905 & w17650;
assign w18523 = pi01860 & ~w18522;
assign w18524 = w17317 & w17650;
assign w18525 = ~w18523 & ~w18524;
assign w18526 = w16993 & w17582;
assign w18527 = ~w16905 & w18526;
assign w18528 = pi01861 & ~w18527;
assign w18529 = w17603 & w18526;
assign w18530 = ~w18528 & ~w18529;
assign w18531 = ~w16892 & w17775;
assign w18532 = pi01862 & ~w18531;
assign w18533 = ~pi02723 & w18531;
assign w18534 = ~w18532 & ~w18533;
assign w18535 = ~w16892 & w17047;
assign w18536 = pi01863 & ~w18535;
assign w18537 = ~pi02709 & w18535;
assign w18538 = ~w18536 & ~w18537;
assign w18539 = pi01864 & ~w16971;
assign w18540 = ~pi02711 & w16971;
assign w18541 = ~w18539 & ~w18540;
assign w18542 = w16983 & w17182;
assign w18543 = ~w16892 & w18542;
assign w18544 = pi01865 & ~w18543;
assign w18545 = ~pi02160 & w18543;
assign w18546 = ~w18544 & ~w18545;
assign w18547 = ~w16892 & w17305;
assign w18548 = pi01866 & ~w18547;
assign w18549 = ~pi02706 & w18547;
assign w18550 = ~w18548 & ~w18549;
assign w18551 = pi01867 & ~w18090;
assign w18552 = w17500 & w18234;
assign w18553 = ~w18551 & ~w18552;
assign w18554 = w16940 & w17038;
assign w18555 = ~w16928 & w18554;
assign w18556 = pi01868 & ~w18555;
assign w18557 = w17193 & w18554;
assign w18558 = ~w18556 & ~w18557;
assign w18559 = ~w16992 & w17775;
assign w18560 = pi01869 & ~w18559;
assign w18561 = w17594 & w17775;
assign w18562 = ~w18560 & ~w18561;
assign w18563 = w16947 & w17136;
assign w18564 = ~w16928 & w18563;
assign w18565 = pi01870 & ~w18564;
assign w18566 = ~pi09812 & w18564;
assign w18567 = ~w18565 & ~w18566;
assign w18568 = ~w16992 & w17320;
assign w18569 = pi01871 & ~w18568;
assign w18570 = ~pi02167 & w18568;
assign w18571 = ~w18569 & ~w18570;
assign w18572 = w16960 & w17113;
assign w18573 = ~w16992 & w18572;
assign w18574 = pi01872 & ~w18573;
assign w18575 = ~pi02721 & w18573;
assign w18576 = ~w18574 & ~w18575;
assign w18577 = pi01873 & ~w18090;
assign w18578 = ~pi02705 & ~w16892;
assign w18579 = w17500 & w18578;
assign w18580 = ~w18577 & ~w18579;
assign w18581 = ~w16992 & w17177;
assign w18582 = pi01874 & ~w18581;
assign w18583 = ~pi02167 & w18581;
assign w18584 = ~w18582 & ~w18583;
assign w18585 = w16947 & w17582;
assign w18586 = ~w16892 & w18585;
assign w18587 = pi01875 & ~w18586;
assign w18588 = ~pi02706 & w18586;
assign w18589 = ~w18587 & ~w18588;
assign w18590 = ~w16992 & w17822;
assign w18591 = pi01876 & ~w18590;
assign w18592 = ~pi02719 & w18590;
assign w18593 = ~w18591 & ~w18592;
assign w18594 = pi01877 & ~w16971;
assign w18595 = ~pi02714 & w16971;
assign w18596 = ~w18594 & ~w18595;
assign w18597 = ~w16905 & w17210;
assign w18598 = pi01878 & ~w18597;
assign w18599 = ~pi02715 & w18597;
assign w18600 = ~w18598 & ~w18599;
assign w18601 = ~w16892 & w18554;
assign w18602 = pi01879 & ~w18601;
assign w18603 = w18364 & w18554;
assign w18604 = ~w18602 & ~w18603;
assign w18605 = ~w16892 & w17411;
assign w18606 = pi01880 & ~w18605;
assign w18607 = w17411 & w17925;
assign w18608 = ~w18606 & ~w18607;
assign w18609 = pi01881 & ~w18601;
assign w18610 = ~pi02160 & w18601;
assign w18611 = ~w18609 & ~w18610;
assign w18612 = w17005 & w17189;
assign w18613 = ~w16905 & w18612;
assign w18614 = pi01882 & ~w18613;
assign w18615 = ~pi02716 & w18613;
assign w18616 = ~w18614 & ~w18615;
assign w18617 = w16960 & w17059;
assign w18618 = ~w16892 & w18617;
assign w18619 = pi01883 & ~w18618;
assign w18620 = ~pi02705 & w18618;
assign w18621 = ~w18619 & ~w18620;
assign w18622 = w16969 & w16985;
assign w18623 = ~w16905 & w18622;
assign w18624 = pi01884 & ~w18623;
assign w18625 = ~pi02712 & w18623;
assign w18626 = ~w18624 & ~w18625;
assign w18627 = ~w16928 & w18572;
assign w18628 = pi01885 & ~w18627;
assign w18629 = ~pi02704 & w18627;
assign w18630 = ~w18628 & ~w18629;
assign w18631 = w17052 & w17374;
assign w18632 = ~w16928 & w18631;
assign w18633 = pi01886 & ~w18632;
assign w18634 = ~pi09812 & w18632;
assign w18635 = ~w18633 & ~w18634;
assign w18636 = w16977 & w17038;
assign w18637 = ~w16992 & w18636;
assign w18638 = pi01887 & ~w18637;
assign w18639 = ~pi02718 & w18637;
assign w18640 = ~w18638 & ~w18639;
assign w18641 = ~w16892 & w18291;
assign w18642 = pi01888 & ~w18641;
assign w18643 = ~pi02708 & w18641;
assign w18644 = ~w18642 & ~w18643;
assign w18645 = w16947 & w17182;
assign w18646 = ~w16892 & w18645;
assign w18647 = pi01889 & ~w18646;
assign w18648 = w18234 & w18645;
assign w18649 = ~w18647 & ~w18648;
assign w18650 = pi01890 & ~w18646;
assign w18651 = ~pi02705 & w18646;
assign w18652 = ~w18650 & ~w18651;
assign w18653 = pi01891 & ~w18597;
assign w18654 = w17210 & w17603;
assign w18655 = ~w18653 & ~w18654;
assign w18656 = pi01892 & ~w18641;
assign w18657 = ~pi02706 & w18641;
assign w18658 = ~w18656 & ~w18657;
assign w18659 = pi01893 & ~w18618;
assign w18660 = ~pi02160 & w18618;
assign w18661 = ~w18659 & ~w18660;
assign w18662 = w17038 & w17059;
assign w18663 = ~w16892 & w18662;
assign w18664 = pi01894 & ~w18663;
assign w18665 = w18092 & w18662;
assign w18666 = ~w18664 & ~w18665;
assign w18667 = ~w16905 & w17084;
assign w18668 = pi01895 & ~w18667;
assign w18669 = w17084 & w17603;
assign w18670 = ~w18668 & ~w18669;
assign w18671 = ~w16905 & w17349;
assign w18672 = pi01896 & ~w18671;
assign w18673 = ~pi02715 & w18671;
assign w18674 = ~w18672 & ~w18673;
assign w18675 = ~w16992 & w17284;
assign w18676 = pi01897 & ~w18675;
assign w18677 = ~pi02164 & w18675;
assign w18678 = ~w18676 & ~w18677;
assign w18679 = ~w16892 & w18526;
assign w18680 = pi01898 & ~w18679;
assign w18681 = ~pi02706 & w18679;
assign w18682 = ~w18680 & ~w18681;
assign w18683 = w16911 & w17582;
assign w18684 = ~w16928 & w18683;
assign w18685 = pi01899 & ~w18684;
assign w18686 = ~pi09812 & w18684;
assign w18687 = ~w18685 & ~w18686;
assign w18688 = pi01900 & ~w18586;
assign w18689 = ~pi02708 & ~w16892;
assign w18690 = w18585 & w18689;
assign w18691 = ~w18688 & ~w18690;
assign w18692 = ~w16892 & w17490;
assign w18693 = pi01901 & ~w18692;
assign w18694 = ~pi02706 & w18692;
assign w18695 = ~w18693 & ~w18694;
assign w18696 = ~w16905 & w18186;
assign w18697 = pi01902 & ~w18696;
assign w18698 = ~pi02715 & w18696;
assign w18699 = ~w18697 & ~w18698;
assign w18700 = pi01903 & ~w18543;
assign w18701 = ~pi02709 & w18543;
assign w18702 = ~w18700 & ~w18701;
assign w18703 = ~w16992 & w17814;
assign w18704 = pi01904 & ~w18703;
assign w18705 = w17594 & w17814;
assign w18706 = ~w18704 & ~w18705;
assign w18707 = pi01905 & ~w18613;
assign w18708 = ~pi02713 & w18613;
assign w18709 = ~w18707 & ~w18708;
assign w18710 = ~w16928 & w18247;
assign w18711 = pi01906 & ~w18710;
assign w18712 = ~pi09954 & w18710;
assign w18713 = ~w18711 & ~w18712;
assign w18714 = ~w16892 & w17495;
assign w18715 = pi01907 & ~w18714;
assign w18716 = ~pi02706 & w18714;
assign w18717 = ~w18715 & ~w18716;
assign w18718 = ~w16928 & w18186;
assign w18719 = pi01908 & ~w18718;
assign w18720 = ~pi02704 & w18718;
assign w18721 = ~w18719 & ~w18720;
assign w18722 = ~w16928 & w18585;
assign w18723 = pi01909 & ~w18722;
assign w18724 = ~pi02720 & w18722;
assign w18725 = ~w18723 & ~w18724;
assign w18726 = w16960 & w16967;
assign w18727 = ~w16928 & w18726;
assign w18728 = pi01910 & ~w18727;
assign w18729 = ~pi02720 & w18727;
assign w18730 = ~w18728 & ~w18729;
assign w18731 = w17124 & w17582;
assign w18732 = ~w16928 & w18731;
assign w18733 = pi01911 & ~w18732;
assign w18734 = ~pi02720 & w18732;
assign w18735 = ~w18733 & ~w18734;
assign w18736 = ~w16928 & w18526;
assign w18737 = pi01912 & ~w18736;
assign w18738 = ~pi09812 & w18736;
assign w18739 = ~w18737 & ~w18738;
assign w18740 = w16895 & w17182;
assign w18741 = ~w16905 & w18740;
assign w18742 = pi01913 & ~w18741;
assign w18743 = ~pi02716 & w18741;
assign w18744 = ~w18742 & ~w18743;
assign w18745 = w16895 & w17037;
assign w18746 = ~w16928 & w18745;
assign w18747 = pi01914 & ~w18746;
assign w18748 = ~pi09962 & w18746;
assign w18749 = ~w18747 & ~w18748;
assign w18750 = pi01915 & ~w18732;
assign w18751 = ~pi09812 & w18732;
assign w18752 = ~w18750 & ~w18751;
assign w18753 = ~w16928 & w18662;
assign w18754 = pi01916 & ~w18753;
assign w18755 = ~pi09812 & w18753;
assign w18756 = ~w18754 & ~w18755;
assign w18757 = ~w16905 & w17114;
assign w18758 = pi01917 & ~w18757;
assign w18759 = w17114 & w17742;
assign w18760 = ~w18758 & ~w18759;
assign w18761 = ~w16905 & w17718;
assign w18762 = pi01918 & ~w18761;
assign w18763 = ~pi02711 & w18761;
assign w18764 = ~w18762 & ~w18763;
assign w18765 = ~w16928 & w17375;
assign w18766 = pi01919 & ~w18765;
assign w18767 = ~pi09812 & w18765;
assign w18768 = ~w18766 & ~w18767;
assign w18769 = pi01920 & ~w18503;
assign w18770 = w17532 & w18051;
assign w18771 = ~w18769 & ~w18770;
assign w18772 = w16930 & w17052;
assign w18773 = ~w16905 & w18772;
assign w18774 = pi01921 & ~w18773;
assign w18775 = ~pi02716 & w18773;
assign w18776 = ~w18774 & ~w18775;
assign w18777 = ~w16928 & w17600;
assign w18778 = pi01922 & ~w18777;
assign w18779 = ~pi02704 & w18777;
assign w18780 = ~w18778 & ~w18779;
assign w18781 = w16953 & w16967;
assign w18782 = ~w16928 & w18781;
assign w18783 = pi01923 & ~w18782;
assign w18784 = ~pi09812 & w18782;
assign w18785 = ~w18783 & ~w18784;
assign w18786 = ~w16992 & w18056;
assign w18787 = pi01924 & ~w18786;
assign w18788 = w17811 & w18056;
assign w18789 = ~w18787 & ~w18788;
assign w18790 = ~w16928 & w18431;
assign w18791 = pi01925 & ~w18790;
assign w18792 = ~pi09954 & w18790;
assign w18793 = ~w18791 & ~w18792;
assign w18794 = ~w16892 & w18186;
assign w18795 = pi01926 & ~w18794;
assign w18796 = ~pi02710 & w18794;
assign w18797 = ~w18795 & ~w18796;
assign w18798 = pi01927 & ~w18710;
assign w18799 = ~pi09848 & w18710;
assign w18800 = ~w18798 & ~w18799;
assign w18801 = pi01928 & ~w18722;
assign w18802 = ~pi09812 & w18722;
assign w18803 = ~w18801 & ~w18802;
assign w18804 = ~w16905 & w17226;
assign w18805 = pi01929 & ~w18804;
assign w18806 = w17020 & w17226;
assign w18807 = ~w18805 & ~w18806;
assign w18808 = w16908 & w17038;
assign w18809 = ~w16928 & w18808;
assign w18810 = pi01930 & ~w18809;
assign w18811 = w17439 & w18808;
assign w18812 = ~w18810 & ~w18811;
assign w18813 = w16993 & w17136;
assign w18814 = ~w16928 & w18813;
assign w18815 = pi01931 & ~w18814;
assign w18816 = ~pi02720 & w18814;
assign w18817 = ~w18815 & ~w18816;
assign w18818 = ~w16928 & w17516;
assign w18819 = pi01932 & ~w18818;
assign w18820 = ~pi09954 & w18818;
assign w18821 = ~w18819 & ~w18820;
assign w18822 = w16983 & w17582;
assign w18823 = ~w16905 & w18822;
assign w18824 = pi01933 & ~w18823;
assign w18825 = ~pi02712 & w18823;
assign w18826 = ~w18824 & ~w18825;
assign w18827 = ~w16892 & w17390;
assign w18828 = pi01934 & ~w18827;
assign w18829 = ~pi02708 & w18827;
assign w18830 = ~w18828 & ~w18829;
assign w18831 = w17005 & w17582;
assign w18832 = ~w16905 & w18831;
assign w18833 = pi01935 & ~w18832;
assign w18834 = ~pi02715 & w18832;
assign w18835 = ~w18833 & ~w18834;
assign w18836 = pi01936 & ~w18832;
assign w18837 = ~pi02712 & w18832;
assign w18838 = ~w18836 & ~w18837;
assign w18839 = pi01937 & ~w18827;
assign w18840 = ~pi02706 & w18827;
assign w18841 = ~w18839 & ~w18840;
assign w18842 = pi01938 & ~w18818;
assign w18843 = w17186 & w17516;
assign w18844 = ~w18842 & ~w18843;
assign w18845 = pi01939 & ~w18761;
assign w18846 = ~pi02714 & w18761;
assign w18847 = ~w18845 & ~w18846;
assign w18848 = ~w16928 & w18636;
assign w18849 = pi01940 & ~w18848;
assign w18850 = ~pi02178 & w18848;
assign w18851 = ~w18849 & ~w18850;
assign w18852 = ~w16928 & w18612;
assign w18853 = pi01941 & ~w18852;
assign w18854 = w17513 & w18612;
assign w18855 = ~w18853 & ~w18854;
assign w18856 = ~w16928 & w18822;
assign w18857 = pi01942 & ~w18856;
assign w18858 = ~pi09954 & w18856;
assign w18859 = ~w18857 & ~w18858;
assign w18860 = pi01943 & ~w18809;
assign w18861 = ~pi02178 & ~w16928;
assign w18862 = w18808 & w18861;
assign w18863 = ~w18860 & ~w18862;
assign w18864 = ~w16992 & w18146;
assign w18865 = pi01944 & ~w18864;
assign w18866 = ~pi02721 & w18864;
assign w18867 = ~w18865 & ~w18866;
assign w18868 = pi01945 & ~w18814;
assign w18869 = ~pi09812 & w18814;
assign w18870 = ~w18868 & ~w18869;
assign w18871 = w16921 & w16960;
assign w18872 = ~w16905 & w18871;
assign w18873 = pi01946 & ~w18872;
assign w18874 = ~pi02712 & w18872;
assign w18875 = ~w18873 & ~w18874;
assign w18876 = pi01947 & ~w18872;
assign w18877 = ~pi02715 & w18872;
assign w18878 = ~w18876 & ~w18877;
assign w18879 = ~w16892 & w17808;
assign w18880 = pi01948 & ~w18879;
assign w18881 = ~pi02160 & w18879;
assign w18882 = ~w18880 & ~w18881;
assign w18883 = pi01949 & ~w18632;
assign w18884 = ~pi02720 & w18632;
assign w18885 = ~w18883 & ~w18884;
assign w18886 = pi01950 & ~w18856;
assign w18887 = ~pi09848 & w18856;
assign w18888 = ~w18886 & ~w18887;
assign w18889 = ~w16928 & w18831;
assign w18890 = pi01951 & ~w18889;
assign w18891 = ~pi09954 & w18889;
assign w18892 = ~w18890 & ~w18891;
assign w18893 = ~w16892 & w16970;
assign w18894 = pi01952 & ~w18893;
assign w18895 = ~pi02160 & w18893;
assign w18896 = ~w18894 & ~w18895;
assign w18897 = w16908 & w17124;
assign w18898 = ~w16905 & w18897;
assign w18899 = pi01953 & ~w18898;
assign w18900 = ~pi02715 & w18898;
assign w18901 = ~w18899 & ~w18900;
assign w18902 = pi01954 & ~w18893;
assign w18903 = w16970 & w18364;
assign w18904 = ~w18902 & ~w18903;
assign w18905 = ~w16928 & w18871;
assign w18906 = pi01955 & ~w18905;
assign w18907 = ~pi09954 & w18905;
assign w18908 = ~w18906 & ~w18907;
assign w18909 = ~w16992 & w18070;
assign w18910 = pi01956 & ~w18909;
assign w18911 = ~pi02721 & w18909;
assign w18912 = ~w18910 & ~w18911;
assign w18913 = w16977 & w17124;
assign w18914 = ~w16928 & w18913;
assign w18915 = pi01957 & ~w18914;
assign w18916 = ~pi09954 & w18914;
assign w18917 = ~w18915 & ~w18916;
assign w18918 = ~w16905 & w17385;
assign w18919 = pi01958 & ~w18918;
assign w18920 = w17385 & w18059;
assign w18921 = ~w18919 & ~w18920;
assign w18922 = pi01959 & ~w18777;
assign w18923 = w17439 & w17600;
assign w18924 = ~w18922 & ~w18923;
assign w18925 = w17083 & w17136;
assign w18926 = ~w16928 & w18925;
assign w18927 = pi01960 & ~w18926;
assign w18928 = w17186 & w18925;
assign w18929 = ~w18927 & ~w18928;
assign w18930 = pi01961 & ~w18898;
assign w18931 = w17020 & w18897;
assign w18932 = ~w18930 & ~w18931;
assign w18933 = pi01962 & ~w18905;
assign w18934 = ~pi09848 & w18905;
assign w18935 = ~w18933 & ~w18934;
assign w18936 = ~w16928 & w18897;
assign w18937 = pi01963 & ~w18936;
assign w18938 = ~pi09954 & w18936;
assign w18939 = ~w18937 & ~w18938;
assign w18940 = ~w16905 & w18913;
assign w18941 = pi01964 & ~w18940;
assign w18942 = ~pi02712 & w18940;
assign w18943 = ~w18941 & ~w18942;
assign w18944 = w16911 & w16967;
assign w18945 = ~w16905 & w18944;
assign w18946 = pi01965 & ~w18945;
assign w18947 = ~pi02715 & w18945;
assign w18948 = ~w18946 & ~w18947;
assign w18949 = w16993 & w17374;
assign w18950 = ~w16928 & w18949;
assign w18951 = pi01966 & ~w18950;
assign w18952 = ~pi09812 & w18950;
assign w18953 = ~w18951 & ~w18952;
assign w18954 = ~w16928 & w18944;
assign w18955 = pi01967 & ~w18954;
assign w18956 = ~pi09954 & w18954;
assign w18957 = ~w18955 & ~w18956;
assign w18958 = pi01968 & ~w18945;
assign w18959 = ~pi02712 & w18945;
assign w18960 = ~w18958 & ~w18959;
assign w18961 = pi01969 & ~w18914;
assign w18962 = ~pi09848 & w18914;
assign w18963 = ~w18961 & ~w18962;
assign w18964 = pi01970 & ~w18864;
assign w18965 = ~pi02719 & w18864;
assign w18966 = ~w18964 & ~w18965;
assign w18967 = ~w16992 & w18116;
assign w18968 = pi01971 & ~w18967;
assign w18969 = ~pi02721 & w18967;
assign w18970 = ~w18968 & ~w18969;
assign w18971 = ~w16892 & w17084;
assign w18972 = pi01972 & ~w18971;
assign w18973 = w17084 & w18234;
assign w18974 = ~w18972 & ~w18973;
assign w18975 = pi01973 & ~w18926;
assign w18976 = ~pi09954 & w18926;
assign w18977 = ~w18975 & ~w18976;
assign w18978 = ~w16905 & w18925;
assign w18979 = pi01974 & ~w18978;
assign w18980 = ~pi02713 & w18978;
assign w18981 = ~w18979 & ~w18980;
assign w18982 = ~w16892 & w18949;
assign w18983 = pi01975 & ~w18982;
assign w18984 = ~pi02160 & w18982;
assign w18985 = ~w18983 & ~w18984;
assign w18986 = w16908 & w16969;
assign w18987 = ~w16905 & w18986;
assign w18988 = pi01976 & ~w18987;
assign w18989 = ~pi02715 & w18987;
assign w18990 = ~w18988 & ~w18989;
assign w18991 = ~w16992 & w18155;
assign w18992 = pi01977 & ~w18991;
assign w18993 = ~pi02721 & w18991;
assign w18994 = ~w18992 & ~w18993;
assign w18995 = w16908 & w16960;
assign w18996 = ~w16928 & w18995;
assign w18997 = pi01978 & ~w18996;
assign w18998 = ~pi09848 & w18996;
assign w18999 = ~w18997 & ~w18998;
assign w19000 = ~w16892 & w18726;
assign w19001 = pi01979 & ~w19000;
assign w19002 = w17671 & w18726;
assign w19003 = ~w19001 & ~w19002;
assign w19004 = ~w16992 & w18263;
assign w19005 = pi01980 & ~w19004;
assign w19006 = ~pi02721 & w19004;
assign w19007 = ~w19005 & ~w19006;
assign w19008 = ~w16928 & w17131;
assign w19009 = pi01981 & ~w19008;
assign w19010 = ~pi09848 & w19008;
assign w19011 = ~w19009 & ~w19010;
assign w19012 = w17052 & w17182;
assign w19013 = ~w16992 & w19012;
assign w19014 = pi01982 & ~w19013;
assign w19015 = ~pi02164 & w19013;
assign w19016 = ~w19014 & ~w19015;
assign w19017 = ~w16992 & w18247;
assign w19018 = pi01983 & ~w19017;
assign w19019 = ~pi02721 & w19017;
assign w19020 = ~w19018 & ~w19019;
assign w19021 = pi01984 & ~w17646;
assign w19022 = ~pi02167 & w17646;
assign w19023 = ~w19021 & ~w19022;
assign w19024 = pi01985 & ~w18703;
assign w19025 = w17532 & w17814;
assign w19026 = ~w19024 & ~w19025;
assign w19027 = ~w16928 & w18986;
assign w19028 = pi01986 & ~w19027;
assign w19029 = ~pi09954 & w19027;
assign w19030 = ~w19028 & ~w19029;
assign w19031 = pi01987 & ~w18987;
assign w19032 = ~pi02712 & w18987;
assign w19033 = ~w19031 & ~w19032;
assign w19034 = w16969 & w16977;
assign w19035 = ~w16905 & w19034;
assign w19036 = pi01988 & ~w19035;
assign w19037 = ~pi02712 & w19035;
assign w19038 = ~w19036 & ~w19037;
assign w19039 = ~w16992 & w18027;
assign w19040 = pi01989 & ~w19039;
assign w19041 = w17532 & w18027;
assign w19042 = ~w19040 & ~w19041;
assign w19043 = ~w16928 & w19034;
assign w19044 = pi01990 & ~w19043;
assign w19045 = ~pi09954 & w19043;
assign w19046 = ~w19044 & ~w19045;
assign w19047 = pi01991 & ~w18991;
assign w19048 = ~pi02164 & w18991;
assign w19049 = ~w19047 & ~w19048;
assign w19050 = pi01992 & ~w18794;
assign w19051 = ~pi02160 & w18794;
assign w19052 = ~w19050 & ~w19051;
assign w19053 = w17038 & w17136;
assign w19054 = ~w16928 & w19053;
assign w19055 = pi01993 & ~w19054;
assign w19056 = ~pi09954 & w19054;
assign w19057 = ~w19055 & ~w19056;
assign w19058 = pi01994 & ~w19043;
assign w19059 = ~pi09848 & w19043;
assign w19060 = ~w19058 & ~w19059;
assign w19061 = ~w16905 & w19053;
assign w19062 = pi01995 & ~w19061;
assign w19063 = ~pi02712 & w19061;
assign w19064 = ~w19062 & ~w19063;
assign w19065 = ~w16905 & w18995;
assign w19066 = pi01996 & ~w19065;
assign w19067 = ~pi02715 & w19065;
assign w19068 = ~w19066 & ~w19067;
assign w19069 = pi01997 & ~w19004;
assign w19070 = ~pi02719 & w19004;
assign w19071 = ~w19069 & ~w19070;
assign w19072 = pi01998 & ~w18996;
assign w19073 = ~pi09954 & w18996;
assign w19074 = ~w19072 & ~w19073;
assign w19075 = w16960 & w16977;
assign w19076 = ~w16905 & w19075;
assign w19077 = pi01999 & ~w19076;
assign w19078 = ~pi02715 & w19076;
assign w19079 = ~w19077 & ~w19078;
assign w19080 = ~w16928 & w19075;
assign w19081 = pi02000 & ~w19080;
assign w19082 = ~pi09954 & w19080;
assign w19083 = ~w19081 & ~w19082;
assign w19084 = pi02001 & ~w19076;
assign w19085 = ~pi02712 & w19076;
assign w19086 = ~w19084 & ~w19085;
assign w19087 = w16983 & w17136;
assign w19088 = ~w16928 & w19087;
assign w19089 = pi02002 & ~w19088;
assign w19090 = ~pi02178 & w19088;
assign w19091 = ~w19089 & ~w19090;
assign w19092 = ~w16905 & w19087;
assign w19093 = pi02003 & ~w19092;
assign w19094 = ~pi02712 & w19092;
assign w19095 = ~w19093 & ~w19094;
assign w19096 = ~w16992 & w18308;
assign w19097 = pi02004 & ~w19096;
assign w19098 = w17811 & w18308;
assign w19099 = ~w19097 & ~w19098;
assign w19100 = pi02005 & ~w17462;
assign w19101 = ~pi09961 & w17462;
assign w19102 = ~w19100 & ~w19101;
assign w19103 = pi02006 & ~w19092;
assign w19104 = ~pi02715 & w19092;
assign w19105 = ~w19103 & ~w19104;
assign w19106 = w16940 & w16953;
assign w19107 = ~w16928 & w19106;
assign w19108 = pi02007 & ~w19107;
assign w19109 = w17513 & w19106;
assign w19110 = ~w19108 & ~w19109;
assign w19111 = ~w16892 & w18808;
assign w19112 = pi02008 & ~w19111;
assign w19113 = ~pi02160 & w19111;
assign w19114 = ~w19112 & ~w19113;
assign w19115 = w17005 & w17136;
assign w19116 = ~w16928 & w19115;
assign w19117 = pi02009 & ~w19116;
assign w19118 = ~pi02178 & w19116;
assign w19119 = ~w19117 & ~w19118;
assign w19120 = ~w16992 & w17510;
assign w19121 = pi02010 & ~w19120;
assign w19122 = ~pi02164 & w19120;
assign w19123 = ~w19121 & ~w19122;
assign w19124 = pi02011 & ~w19111;
assign w19125 = ~pi02705 & w19111;
assign w19126 = ~w19124 & ~w19125;
assign w19127 = pi02012 & ~w19120;
assign w19128 = ~pi02719 & w19120;
assign w19129 = ~w19127 & ~w19128;
assign w19130 = w17052 & w17059;
assign w19131 = ~w16928 & w19130;
assign w19132 = pi02013 & ~w19131;
assign w19133 = ~pi02178 & w19131;
assign w19134 = ~w19132 & ~w19133;
assign w19135 = pi02014 & ~w19131;
assign w19136 = ~pi09961 & w19131;
assign w19137 = ~w19135 & ~w19136;
assign w19138 = ~w16892 & w18572;
assign w19139 = pi02015 & ~w19138;
assign w19140 = ~pi02723 & w19138;
assign w19141 = ~w19139 & ~w19140;
assign w19142 = pi02016 & ~w19120;
assign w19143 = ~pi02721 & w19120;
assign w19144 = ~w19142 & ~w19143;
assign w19145 = ~w16992 & w17361;
assign w19146 = pi02017 & ~w19145;
assign w19147 = ~pi02719 & w19145;
assign w19148 = ~w19146 & ~w19147;
assign w19149 = w16953 & w17037;
assign w19150 = ~w16928 & w19149;
assign w19151 = pi02018 & ~w19150;
assign w19152 = ~pi09961 & w19150;
assign w19153 = ~w19151 & ~w19152;
assign w19154 = ~w16992 & w17325;
assign w19155 = pi02019 & ~w19154;
assign w19156 = ~pi02167 & w19154;
assign w19157 = ~w19155 & ~w19156;
assign w19158 = ~w16992 & w18431;
assign w19159 = pi02020 & ~w19158;
assign w19160 = ~pi02164 & w19158;
assign w19161 = ~w19159 & ~w19160;
assign w19162 = ~w16992 & w18612;
assign w19163 = pi02021 & ~w19162;
assign w19164 = w17620 & w18612;
assign w19165 = ~w19163 & ~w19164;
assign w19166 = w16919 & w17059;
assign w19167 = ~w16928 & w19166;
assign w19168 = pi02022 & ~w19167;
assign w19169 = ~pi09954 & w19167;
assign w19170 = ~w19168 & ~w19169;
assign w19171 = ~w16992 & w17254;
assign w19172 = pi02023 & ~w19171;
assign w19173 = ~pi02719 & w19171;
assign w19174 = ~w19172 & ~w19173;
assign w19175 = pi02024 & ~w19158;
assign w19176 = ~pi02721 & w19158;
assign w19177 = ~w19175 & ~w19176;
assign w19178 = pi02025 & ~w19171;
assign w19179 = ~pi02718 & w19171;
assign w19180 = ~w19178 & ~w19179;
assign w19181 = ~w16992 & w17516;
assign w19182 = pi02026 & ~w19181;
assign w19183 = w17516 & w17811;
assign w19184 = ~w19182 & ~w19183;
assign w19185 = pi02027 & ~w19162;
assign w19186 = ~pi02721 & w19162;
assign w19187 = ~w19185 & ~w19186;
assign w19188 = ~w16992 & w18822;
assign w19189 = pi02028 & ~w19188;
assign w19190 = ~pi02169 & w19188;
assign w19191 = ~w19189 & ~w19190;
assign w19192 = ~w16905 & w19166;
assign w19193 = pi02029 & ~w19192;
assign w19194 = ~pi02714 & w19192;
assign w19195 = ~w19193 & ~w19194;
assign w19196 = pi02030 & ~w19188;
assign w19197 = ~pi02721 & w19188;
assign w19198 = ~w19196 & ~w19197;
assign w19199 = pi02031 & ~w19150;
assign w19200 = ~pi02178 & w19150;
assign w19201 = ~w19199 & ~w19200;
assign w19202 = ~w16992 & w17167;
assign w19203 = pi02032 & ~w19202;
assign w19204 = ~pi02719 & w19202;
assign w19205 = ~w19203 & ~w19204;
assign w19206 = ~w16905 & w19130;
assign w19207 = pi02033 & ~w19206;
assign w19208 = ~pi02712 & w19206;
assign w19209 = ~w19207 & ~w19208;
assign w19210 = ~w16892 & w18636;
assign w19211 = pi02034 & ~w19210;
assign w19212 = ~pi02723 & w19210;
assign w19213 = ~w19211 & ~w19212;
assign w19214 = pi02035 & ~w19192;
assign w19215 = ~pi02712 & w19192;
assign w19216 = ~w19214 & ~w19215;
assign w19217 = ~w16992 & w18831;
assign w19218 = pi02036 & ~w19217;
assign w19219 = ~pi02721 & w19217;
assign w19220 = ~w19218 & ~w19219;
assign w19221 = pi02037 & ~w19107;
assign w19222 = ~pi02704 & w19107;
assign w19223 = ~w19221 & ~w19222;
assign w19224 = ~w16905 & w19149;
assign w19225 = pi02038 & ~w19224;
assign w19226 = ~pi02712 & w19224;
assign w19227 = ~w19225 & ~w19226;
assign w19228 = ~w16992 & w18871;
assign w19229 = pi02039 & ~w19228;
assign w19230 = ~pi02164 & w19228;
assign w19231 = ~w19229 & ~w19230;
assign w19232 = pi02040 & ~w19228;
assign w19233 = ~pi02718 & w19228;
assign w19234 = ~w19232 & ~w19233;
assign w19235 = pi02041 & ~w18918;
assign w19236 = ~pi02170 & w18918;
assign w19237 = ~w19235 & ~w19236;
assign w19238 = ~w16905 & w19106;
assign w19239 = pi02042 & ~w19238;
assign w19240 = ~pi02712 & w19238;
assign w19241 = ~w19239 & ~w19240;
assign w19242 = ~w16905 & w17060;
assign w19243 = pi02043 & ~w19242;
assign w19244 = w17060 & w18059;
assign w19245 = ~w19243 & ~w19244;
assign w19246 = pi02044 & ~w19242;
assign w19247 = ~pi02712 & w19242;
assign w19248 = ~w19246 & ~w19247;
assign w19249 = ~w16928 & w17060;
assign w19250 = pi02045 & ~w19249;
assign w19251 = ~pi09848 & w19249;
assign w19252 = ~w19250 & ~w19251;
assign w19253 = ~w16905 & w17131;
assign w19254 = pi02046 & ~w19253;
assign w19255 = ~pi02713 & w19253;
assign w19256 = ~w19254 & ~w19255;
assign w19257 = pi02047 & ~w19008;
assign w19258 = w17131 & w17513;
assign w19259 = ~w19257 & ~w19258;
assign w19260 = pi02048 & ~w19210;
assign w19261 = ~pi02705 & w19210;
assign w19262 = ~w19260 & ~w19261;
assign w19263 = pi02049 & ~w18746;
assign w19264 = ~pi02178 & w18746;
assign w19265 = ~w19263 & ~w19264;
assign w19266 = pi10665 & w11484;
assign w19267 = w1240 & w19266;
assign w19268 = pi02050 & ~w19267;
assign w19269 = pi10604 & w19267;
assign w19270 = ~w19268 & ~w19269;
assign w19271 = ~w16992 & w18897;
assign w19272 = pi02051 & ~w19271;
assign w19273 = ~pi02167 & ~w16992;
assign w19274 = w18897 & w19273;
assign w19275 = ~w19272 & ~w19274;
assign w19276 = pi02052 & ~w19271;
assign w19277 = ~pi02721 & w19271;
assign w19278 = ~w19276 & ~w19277;
assign w19279 = pi02053 & ~w19267;
assign w19280 = pi10600 & w19267;
assign w19281 = ~w19279 & ~w19280;
assign w19282 = w16967 & w17038;
assign w19283 = ~w16892 & w19282;
assign w19284 = pi02054 & ~w19283;
assign w19285 = ~pi02723 & w19283;
assign w19286 = ~w19284 & ~w19285;
assign w19287 = ~w16905 & w17218;
assign w19288 = pi02055 & ~w19287;
assign w19289 = w17218 & w18059;
assign w19290 = ~w19288 & ~w19289;
assign w19291 = ~w16905 & w16948;
assign w19292 = pi02056 & ~w19291;
assign w19293 = ~pi02712 & w19291;
assign w19294 = ~w19292 & ~w19293;
assign w19295 = pi02057 & ~w19287;
assign w19296 = ~pi02712 & w19287;
assign w19297 = ~w19295 & ~w19296;
assign w19298 = ~w16992 & w18944;
assign w19299 = pi02058 & ~w19298;
assign w19300 = ~pi02169 & w19298;
assign w19301 = ~w19299 & ~w19300;
assign w19302 = ~w16992 & w18913;
assign w19303 = pi02059 & ~w19302;
assign w19304 = w17811 & w18913;
assign w19305 = ~w19303 & ~w19304;
assign w19306 = w16895 & w16908;
assign w19307 = ~w16905 & w19306;
assign w19308 = pi02060 & ~w19307;
assign w19309 = ~pi02712 & w19307;
assign w19310 = ~w19308 & ~w19309;
assign w19311 = pi02061 & ~w19298;
assign w19312 = ~pi02722 & ~w16992;
assign w19313 = w18944 & w19312;
assign w19314 = ~w19311 & ~w19313;
assign w19315 = w16899 & ~w16905;
assign w19316 = pi02062 & ~w19315;
assign w19317 = ~pi02715 & w19315;
assign w19318 = ~w19316 & ~w19317;
assign w19319 = ~w16905 & w17380;
assign w19320 = pi02063 & ~w19319;
assign w19321 = ~pi02715 & w19319;
assign w19322 = ~w19320 & ~w19321;
assign w19323 = ~w16928 & w16948;
assign w19324 = pi02064 & ~w19323;
assign w19325 = ~pi09848 & w19323;
assign w19326 = ~w19324 & ~w19325;
assign w19327 = w16985 & w17052;
assign w19328 = ~w16892 & w19327;
assign w19329 = pi02065 & ~w19328;
assign w19330 = ~pi02706 & w19328;
assign w19331 = ~w19329 & ~w19330;
assign w19332 = pi02066 & ~w19319;
assign w19333 = w17380 & w17603;
assign w19334 = ~w19332 & ~w19333;
assign w19335 = ~w16928 & w17218;
assign w19336 = pi02067 & ~w19335;
assign w19337 = ~pi09954 & w19335;
assign w19338 = ~w19336 & ~w19337;
assign w19339 = ~w16992 & w18925;
assign w19340 = pi02068 & ~w19339;
assign w19341 = ~pi02164 & w19339;
assign w19342 = ~w19340 & ~w19341;
assign w19343 = w16940 & w17016;
assign w19344 = ~w16892 & w19343;
assign w19345 = pi02069 & ~w19344;
assign w19346 = ~pi02706 & w19344;
assign w19347 = ~w19345 & ~w19346;
assign w19348 = w17052 & w17113;
assign w19349 = ~w16892 & w19348;
assign w19350 = pi02070 & ~w19349;
assign w19351 = w18067 & w19348;
assign w19352 = ~w19350 & ~w19351;
assign w19353 = pi02071 & ~w19335;
assign w19354 = ~pi09961 & w19335;
assign w19355 = ~w19353 & ~w19354;
assign w19356 = pi02072 & ~w19339;
assign w19357 = ~pi02721 & w19339;
assign w19358 = ~w19356 & ~w19357;
assign w19359 = ~w16992 & w18986;
assign w19360 = pi02073 & ~w19359;
assign w19361 = ~pi02167 & w19359;
assign w19362 = ~w19360 & ~w19361;
assign w19363 = ~w16928 & w17380;
assign w19364 = pi02074 & ~w19363;
assign w19365 = ~pi09961 & ~w16928;
assign w19366 = w17380 & w19365;
assign w19367 = ~w19364 & ~w19366;
assign w19368 = pi02075 & ~w19349;
assign w19369 = w18578 & w19348;
assign w19370 = ~w19368 & ~w19369;
assign w19371 = pi02076 & ~w18522;
assign w19372 = w17020 & w17650;
assign w19373 = ~w19371 & ~w19372;
assign w19374 = w16919 & w17113;
assign w19375 = ~w16892 & w19374;
assign w19376 = pi02077 & ~w19375;
assign w19377 = ~pi02706 & w19375;
assign w19378 = ~w19376 & ~w19377;
assign w19379 = w16985 & w17005;
assign w19380 = ~w16928 & w19379;
assign w19381 = pi02078 & ~w19380;
assign w19382 = w17439 & w19379;
assign w19383 = ~w19381 & ~w19382;
assign w19384 = ~w16892 & w19012;
assign w19385 = pi02079 & ~w19384;
assign w19386 = ~pi02708 & w19384;
assign w19387 = ~w19385 & ~w19386;
assign w19388 = ~w16992 & w19034;
assign w19389 = pi02080 & ~w19388;
assign w19390 = ~pi02164 & w19388;
assign w19391 = ~w19389 & ~w19390;
assign w19392 = pi02081 & ~w19384;
assign w19393 = ~pi02706 & w19384;
assign w19394 = ~w19392 & ~w19393;
assign w19395 = w16899 & ~w16928;
assign w19396 = pi02082 & ~w19395;
assign w19397 = ~pi09848 & w19395;
assign w19398 = ~w19396 & ~w19397;
assign w19399 = pi02083 & ~w19388;
assign w19400 = ~pi02719 & w19388;
assign w19401 = ~w19399 & ~w19400;
assign w19402 = ~w16905 & w18808;
assign w19403 = pi02084 & ~w19402;
assign w19404 = ~pi02714 & w19402;
assign w19405 = ~w19403 & ~w19404;
assign w19406 = ~w16905 & w16922;
assign w19407 = pi02085 & ~w19406;
assign w19408 = ~pi02714 & w19406;
assign w19409 = ~w19407 & ~w19408;
assign w19410 = pi02086 & ~w19363;
assign w19411 = w17380 & w17513;
assign w19412 = ~w19410 & ~w19411;
assign w19413 = pi02087 & ~w19328;
assign w19414 = ~pi02710 & w19328;
assign w19415 = ~w19413 & ~w19414;
assign w19416 = ~w16992 & w19053;
assign w19417 = pi02088 & ~w19416;
assign w19418 = ~pi02719 & w19416;
assign w19419 = ~w19417 & ~w19418;
assign w19420 = w16921 & w16953;
assign w19421 = ~w16892 & w19420;
assign w19422 = pi02089 & ~w19421;
assign w19423 = ~pi02706 & w19421;
assign w19424 = ~w19422 & ~w19423;
assign w19425 = pi02090 & ~w19406;
assign w19426 = ~pi02712 & w19406;
assign w19427 = ~w19425 & ~w19426;
assign w19428 = ~w16992 & w19343;
assign w19429 = pi02091 & ~w19428;
assign w19430 = ~pi02721 & w19428;
assign w19431 = ~w19429 & ~w19430;
assign w19432 = pi02092 & ~w19283;
assign w19433 = ~pi02705 & w19283;
assign w19434 = ~w19432 & ~w19433;
assign w19435 = w16993 & w17182;
assign w19436 = ~w16892 & w19435;
assign w19437 = pi02093 & ~w19436;
assign w19438 = ~pi02706 & w19436;
assign w19439 = ~w19437 & ~w19438;
assign w19440 = ~w16992 & w19348;
assign w19441 = pi02094 & ~w19440;
assign w19442 = ~pi02164 & w19440;
assign w19443 = ~w19441 & ~w19442;
assign w19444 = w16919 & w16985;
assign w19445 = ~w16892 & w19444;
assign w19446 = pi02095 & ~w19445;
assign w19447 = ~pi02708 & w19445;
assign w19448 = ~w19446 & ~w19447;
assign w19449 = pi02096 & ~w17954;
assign w19450 = ~pi02711 & w17954;
assign w19451 = ~w19449 & ~w19450;
assign w19452 = pi02097 & ~w19445;
assign w19453 = ~pi02706 & w19445;
assign w19454 = ~w19452 & ~w19453;
assign w19455 = ~w16992 & w17474;
assign w19456 = pi02098 & ~w19455;
assign w19457 = ~pi02703 & w19455;
assign w19458 = ~w19456 & ~w19457;
assign w19459 = w16938 & w17113;
assign w19460 = ~w16892 & w19459;
assign w19461 = pi02099 & ~w19460;
assign w19462 = ~pi02706 & w19460;
assign w19463 = ~w19461 & ~w19462;
assign w19464 = pi02100 & ~w19460;
assign w19465 = w18689 & w19459;
assign w19466 = ~w19464 & ~w19465;
assign w19467 = pi02101 & ~w18518;
assign w19468 = ~pi02703 & w18518;
assign w19469 = ~w19467 & ~w19468;
assign w19470 = pi02102 & ~w19455;
assign w19471 = ~pi02167 & w19455;
assign w19472 = ~w19470 & ~w19471;
assign w19473 = pi02103 & ~w19307;
assign w19474 = ~pi02714 & w19307;
assign w19475 = ~w19473 & ~w19474;
assign w19476 = ~w16992 & w17239;
assign w19477 = pi02104 & ~w19476;
assign w19478 = ~pi02719 & w19476;
assign w19479 = ~w19477 & ~w19478;
assign w19480 = w16938 & w17182;
assign w19481 = ~w16892 & w19480;
assign w19482 = pi02105 & ~w19481;
assign w19483 = w17925 & w19480;
assign w19484 = ~w19482 & ~w19483;
assign w19485 = ~w16905 & w17339;
assign w19486 = pi02106 & ~w19485;
assign w19487 = w16973 & w17339;
assign w19488 = ~w19486 & ~w19487;
assign w19489 = pi02107 & ~w19485;
assign w19490 = ~pi02713 & w19485;
assign w19491 = ~w19489 & ~w19490;
assign w19492 = w16938 & w16985;
assign w19493 = ~w16892 & w19492;
assign w19494 = pi02108 & ~w19493;
assign w19495 = ~pi02708 & w19493;
assign w19496 = ~w19494 & ~w19495;
assign w19497 = ~w16928 & w18370;
assign w19498 = pi02109 & ~w19497;
assign w19499 = w17513 & w18370;
assign w19500 = ~w19498 & ~w19499;
assign w19501 = ~w16992 & w18995;
assign w19502 = pi02110 & ~w19501;
assign w19503 = ~pi02164 & w19501;
assign w19504 = ~w19502 & ~w19503;
assign w19505 = pi02111 & ~w19416;
assign w19506 = ~pi02721 & w19416;
assign w19507 = ~w19505 & ~w19506;
assign w19508 = ~w16992 & w19374;
assign w19509 = pi02112 & ~w19508;
assign w19510 = ~pi02721 & w19508;
assign w19511 = ~w19509 & ~w19510;
assign w19512 = pi02113 & ~w19501;
assign w19513 = ~pi02169 & w19501;
assign w19514 = ~w19512 & ~w19513;
assign w19515 = pi02114 & ~w19039;
assign w19516 = ~pi02167 & w19039;
assign w19517 = ~w19515 & ~w19516;
assign w19518 = w16921 & w16947;
assign w19519 = ~w16892 & w19518;
assign w19520 = pi02115 & ~w19519;
assign w19521 = w18578 & w19518;
assign w19522 = ~w19520 & ~w19521;
assign w19523 = ~w16892 & w17279;
assign w19524 = pi02116 & ~w19523;
assign w19525 = w17279 & w17671;
assign w19526 = ~w19524 & ~w19525;
assign w19527 = pi02117 & ~w19440;
assign w19528 = ~pi02721 & w19440;
assign w19529 = ~w19527 & ~w19528;
assign w19530 = w16993 & w17113;
assign w19531 = ~w16892 & w19530;
assign w19532 = pi02118 & ~w19531;
assign w19533 = ~pi02708 & w19531;
assign w19534 = ~w19532 & ~w19533;
assign w19535 = pi02119 & ~w19531;
assign w19536 = ~pi02706 & w19531;
assign w19537 = ~w19535 & ~w19536;
assign w19538 = pi02120 & ~w19013;
assign w19539 = ~pi02721 & w19013;
assign w19540 = ~w19538 & ~w19539;
assign w19541 = ~w16905 & w17153;
assign w19542 = pi02121 & ~w19541;
assign w19543 = ~pi02717 & w19541;
assign w19544 = ~w19542 & ~w19543;
assign w19545 = ~w16992 & w17428;
assign w19546 = pi02122 & ~w19545;
assign w19547 = ~pi02721 & w19545;
assign w19548 = ~w19546 & ~w19547;
assign w19549 = pi02123 & ~w14136;
assign w19550 = ~pi01210 & w14136;
assign w19551 = ~w19549 & ~w19550;
assign w19552 = w16985 & w16993;
assign w19553 = ~w16892 & w19552;
assign w19554 = pi02124 & ~w19553;
assign w19555 = ~pi02709 & w19553;
assign w19556 = ~w19554 & ~w19555;
assign w19557 = ~w16992 & w19075;
assign w19558 = pi02125 & ~w19557;
assign w19559 = ~pi02164 & w19557;
assign w19560 = ~w19558 & ~w19559;
assign w19561 = w16921 & w17016;
assign w19562 = ~w16892 & w19561;
assign w19563 = pi02126 & ~w19562;
assign w19564 = ~pi02706 & w19562;
assign w19565 = ~w19563 & ~w19564;
assign w19566 = pi02127 & ~w19557;
assign w19567 = ~pi02721 & w19557;
assign w19568 = ~w19566 & ~w19567;
assign w19569 = pi02128 & ~w19557;
assign w19570 = ~pi02703 & w19557;
assign w19571 = ~w19569 & ~w19570;
assign w19572 = ~w16992 & w19087;
assign w19573 = pi02129 & ~w19572;
assign w19574 = ~pi02721 & w19572;
assign w19575 = ~w19573 & ~w19574;
assign w19576 = w16898 & w17083;
assign w19577 = ~w16892 & w19576;
assign w19578 = pi02130 & ~w19577;
assign w19579 = ~pi02709 & w19577;
assign w19580 = ~w19578 & ~w19579;
assign w19581 = pi02131 & ~w19476;
assign w19582 = ~pi02718 & w19476;
assign w19583 = ~w19581 & ~w19582;
assign w19584 = ~w16992 & w19115;
assign w19585 = pi02132 & ~w19584;
assign w19586 = ~pi02721 & w19584;
assign w19587 = ~w19585 & ~w19586;
assign w19588 = pi02133 & ~w19584;
assign w19589 = ~pi02164 & w19584;
assign w19590 = ~w19588 & ~w19589;
assign w19591 = w16919 & w17182;
assign w19592 = ~w16992 & w19591;
assign w19593 = pi02134 & ~w19592;
assign w19594 = w17811 & w19591;
assign w19595 = ~w19593 & ~w19594;
assign w19596 = w16908 & w17005;
assign w19597 = ~w16892 & w19596;
assign w19598 = pi02135 & ~w19597;
assign w19599 = ~pi02723 & w19597;
assign w19600 = ~w19598 & ~w19599;
assign w19601 = w17037 & w17124;
assign w19602 = ~w16892 & w19601;
assign w19603 = pi02136 & ~w19602;
assign w19604 = ~pi02706 & w19602;
assign w19605 = ~w19603 & ~w19604;
assign w19606 = w16940 & w17124;
assign w19607 = ~w16892 & w19606;
assign w19608 = pi02137 & ~w19607;
assign w19609 = ~pi02708 & w19607;
assign w19610 = ~w19608 & ~w19609;
assign w19611 = ~w16992 & w19327;
assign w19612 = pi02138 & ~w19611;
assign w19613 = w17620 & w19327;
assign w19614 = ~w19612 & ~w19613;
assign w19615 = pi02139 & ~w19607;
assign w19616 = ~pi02706 & w19607;
assign w19617 = ~w19615 & ~w19616;
assign w19618 = pi02140 & ~w19611;
assign w19619 = ~pi02721 & w19611;
assign w19620 = ~w19618 & ~w19619;
assign w19621 = pi02141 & ~w19597;
assign w19622 = w18578 & w19596;
assign w19623 = ~w19621 & ~w19622;
assign w19624 = w16911 & w17059;
assign w19625 = ~w16892 & w19624;
assign w19626 = pi02142 & ~w19625;
assign w19627 = ~pi02706 & w19625;
assign w19628 = ~w19626 & ~w19627;
assign w19629 = w16977 & w17005;
assign w19630 = ~w16892 & w19629;
assign w19631 = pi02143 & ~w19630;
assign w19632 = ~pi02723 & w19630;
assign w19633 = ~w19631 & ~w19632;
assign w19634 = ~w16992 & w17259;
assign w19635 = pi02144 & ~w19634;
assign w19636 = w17259 & w17594;
assign w19637 = ~w19635 & ~w19636;
assign w19638 = ~w16992 & w19420;
assign w19639 = pi02145 & ~w19638;
assign w19640 = ~pi02721 & w19638;
assign w19641 = ~w19639 & ~w19640;
assign w19642 = pi02146 & ~w19577;
assign w19643 = ~pi02707 & w19577;
assign w19644 = ~w19642 & ~w19643;
assign w19645 = w16969 & w17037;
assign w19646 = ~w16892 & w19645;
assign w19647 = pi02147 & ~w19646;
assign w19648 = ~pi02707 & w19646;
assign w19649 = ~w19647 & ~w19648;
assign w19650 = w16940 & w16969;
assign w19651 = ~w16892 & w19650;
assign w19652 = pi02148 & ~w19651;
assign w19653 = ~pi02709 & w19651;
assign w19654 = ~w19652 & ~w19653;
assign w19655 = w16977 & w16983;
assign w19656 = ~w16892 & w19655;
assign w19657 = pi02149 & ~w19656;
assign w19658 = ~pi02723 & w19656;
assign w19659 = ~w19657 & ~w19658;
assign w19660 = w16960 & w17037;
assign w19661 = ~w16892 & w19660;
assign w19662 = pi02150 & ~w19661;
assign w19663 = w18092 & w19660;
assign w19664 = ~w19662 & ~w19663;
assign w19665 = ~w16992 & w17416;
assign w19666 = pi02151 & ~w19665;
assign w19667 = w17416 & w17532;
assign w19668 = ~w19666 & ~w19667;
assign w19669 = pi02152 & ~w19485;
assign w19670 = ~pi02711 & w19485;
assign w19671 = ~w19669 & ~w19670;
assign w19672 = pi02153 & ~w19651;
assign w19673 = ~pi02707 & w19651;
assign w19674 = ~w19672 & ~w19673;
assign w19675 = ~w16992 & w19444;
assign w19676 = pi02154 & ~w19675;
assign w19677 = w17811 & w19444;
assign w19678 = ~w19676 & ~w19677;
assign w19679 = w16898 & w17038;
assign w19680 = ~w16892 & w19679;
assign w19681 = pi02155 & ~w19680;
assign w19682 = ~pi02707 & w19680;
assign w19683 = ~w19681 & ~w19682;
assign w19684 = pi02156 & ~w19638;
assign w19685 = ~pi02164 & w19638;
assign w19686 = ~w19684 & ~w19685;
assign w19687 = pi00468 & w14250;
assign w19688 = pi02157 & ~w14250;
assign w19689 = ~w19687 & ~w19688;
assign w19690 = ~w16992 & w19480;
assign w19691 = pi02158 & ~w19690;
assign w19692 = ~pi02721 & w19690;
assign w19693 = ~w19691 & ~w19692;
assign w19694 = ~w16992 & w17762;
assign w19695 = pi02159 & ~w19694;
assign w19696 = ~pi02718 & w19694;
assign w19697 = ~w19695 & ~w19696;
assign w19698 = pi10480 & pi10539;
assign w19699 = ~pi10480 & ~pi10539;
assign w19700 = pi10393 & w19699;
assign w19701 = pi10408 & ~pi10539;
assign w19702 = ~pi10540 & ~w19698;
assign w19703 = ~w19701 & w19702;
assign w19704 = ~w19700 & w19703;
assign w19705 = pi10609 & w19704;
assign w19706 = pi10480 & ~pi10540;
assign w19707 = pi10540 & w19699;
assign w19708 = ~pi10393 & w19707;
assign w19709 = ~w19706 & ~w19708;
assign w19710 = w19701 & ~w19709;
assign w19711 = ~w19704 & ~w19710;
assign w19712 = pi10393 & w19707;
assign w19713 = w19711 & ~w19712;
assign w19714 = ~pi02160 & w19713;
assign w19715 = pi10369 & w19712;
assign w19716 = ~pi00258 & w19710;
assign w19717 = ~w19705 & ~w19715;
assign w19718 = ~w19716 & w19717;
assign w19719 = ~w19714 & w19718;
assign w19720 = pi02161 & ~w19661;
assign w19721 = w18067 & w19660;
assign w19722 = ~w19720 & ~w19721;
assign w19723 = w16940 & w16960;
assign w19724 = ~w16892 & w19723;
assign w19725 = pi02162 & ~w19724;
assign w19726 = ~pi02707 & w19724;
assign w19727 = ~w19725 & ~w19726;
assign w19728 = w16898 & w16983;
assign w19729 = ~w16892 & w19728;
assign w19730 = pi02163 & ~w19729;
assign w19731 = ~pi02709 & w19729;
assign w19732 = ~w19730 & ~w19731;
assign w19733 = pi10595 & w19704;
assign w19734 = ~pi02164 & w19713;
assign w19735 = pi10477 & w19712;
assign w19736 = pi00048 & w19710;
assign w19737 = ~w19733 & ~w19735;
assign w19738 = ~w19736 & w19737;
assign w19739 = ~w19734 & w19738;
assign w19740 = w16898 & w17005;
assign w19741 = ~w16892 & w19740;
assign w19742 = pi02165 & ~w19741;
assign w19743 = ~pi02723 & w19741;
assign w19744 = ~w19742 & ~w19743;
assign w19745 = pi02166 & ~w19729;
assign w19746 = ~pi02707 & w19729;
assign w19747 = ~w19745 & ~w19746;
assign w19748 = pi10594 & w19704;
assign w19749 = ~pi02167 & w19713;
assign w19750 = pi10537 & w19712;
assign w19751 = pi00047 & w19710;
assign w19752 = ~w19748 & ~w19750;
assign w19753 = ~w19751 & w19752;
assign w19754 = ~w19749 & w19753;
assign w19755 = ~w16992 & w19459;
assign w19756 = pi02168 & ~w19755;
assign w19757 = ~pi02703 & w19755;
assign w19758 = ~w19756 & ~w19757;
assign w19759 = pi10592 & w19704;
assign w19760 = ~pi02169 & w19713;
assign w19761 = pi10524 & w19712;
assign w19762 = pi00046 & w19710;
assign w19763 = ~w19759 & ~w19761;
assign w19764 = ~w19762 & w19763;
assign w19765 = ~w19760 & w19764;
assign w19766 = pi10616 & w19704;
assign w19767 = ~pi02170 & w19713;
assign w19768 = ~pi00960 & w19712;
assign w19769 = ~pi00193 & w19710;
assign w19770 = ~w19766 & ~w19768;
assign w19771 = ~w19769 & w19770;
assign w19772 = ~w19767 & w19771;
assign w19773 = ~w16992 & w19130;
assign w19774 = pi02171 & ~w19773;
assign w19775 = ~pi02169 & w19773;
assign w19776 = ~w19774 & ~w19775;
assign w19777 = pi02172 & ~w19741;
assign w19778 = ~pi02707 & w19741;
assign w19779 = ~w19777 & ~w19778;
assign w19780 = pi02173 & ~w19690;
assign w19781 = w17620 & w19480;
assign w19782 = ~w19780 & ~w19781;
assign w19783 = ~w16992 & w19435;
assign w19784 = pi02174 & ~w19783;
assign w19785 = ~pi02721 & w19783;
assign w19786 = ~w19784 & ~w19785;
assign w19787 = ~w16892 & w17734;
assign w19788 = pi02175 & ~w19787;
assign w19789 = ~pi02723 & w19787;
assign w19790 = ~w19788 & ~w19789;
assign w19791 = ~w16992 & w17125;
assign w19792 = pi02176 & ~w19791;
assign w19793 = ~pi02719 & w19791;
assign w19794 = ~w19792 & ~w19793;
assign w19795 = ~w16992 & w19492;
assign w19796 = pi02177 & ~w19795;
assign w19797 = ~pi02169 & ~w16992;
assign w19798 = w19492 & w19797;
assign w19799 = ~w19796 & ~w19798;
assign w19800 = pi10604 & w19704;
assign w19801 = ~pi02178 & w19713;
assign w19802 = ~pi00133 & w19712;
assign w19803 = ~pi00140 & w19710;
assign w19804 = ~w19800 & ~w19802;
assign w19805 = ~w19803 & w19804;
assign w19806 = ~w19801 & w19805;
assign w19807 = ~w16992 & w19166;
assign w19808 = pi02179 & ~w19807;
assign w19809 = ~pi02169 & w19807;
assign w19810 = ~w19808 & ~w19809;
assign w19811 = pi10660 & w19704;
assign w19812 = pi02180 & w19713;
assign w19813 = pi01215 & w19712;
assign w19814 = pi01452 & w19710;
assign w19815 = ~w19811 & ~w19813;
assign w19816 = ~w19814 & w19815;
assign w19817 = ~w19812 & w19816;
assign w19818 = w16921 & w17124;
assign w19819 = ~w16892 & w19818;
assign w19820 = pi02181 & ~w19819;
assign w19821 = w18092 & w19818;
assign w19822 = ~w19820 & ~w19821;
assign w19823 = pi02182 & ~w19819;
assign w19824 = ~pi02707 & w19819;
assign w19825 = ~w19823 & ~w19824;
assign w19826 = w16911 & w17113;
assign w19827 = ~w16892 & w19826;
assign w19828 = pi02183 & ~w19827;
assign w19829 = ~pi02707 & w19827;
assign w19830 = ~w19828 & ~w19829;
assign w19831 = ~w16992 & w19518;
assign w19832 = pi02184 & ~w19831;
assign w19833 = ~pi02164 & w19831;
assign w19834 = ~w19832 & ~w19833;
assign w19835 = pi02185 & ~w19831;
assign w19836 = ~pi02721 & w19831;
assign w19837 = ~w19835 & ~w19836;
assign w19838 = w16911 & w17182;
assign w19839 = ~w16892 & w19838;
assign w19840 = pi02186 & ~w19839;
assign w19841 = ~pi02709 & w19839;
assign w19842 = ~w19840 & ~w19841;
assign w19843 = pi02187 & ~w19630;
assign w19844 = ~pi02705 & w19630;
assign w19845 = ~w19843 & ~w19844;
assign w19846 = pi02188 & ~w19839;
assign w19847 = ~pi02160 & w19839;
assign w19848 = ~w19846 & ~w19847;
assign w19849 = pi02189 & ~w16225;
assign w19850 = ~pi10628 & w16225;
assign w19851 = ~w19849 & ~w19850;
assign w19852 = w16911 & w16985;
assign w19853 = ~w16892 & w19852;
assign w19854 = pi02190 & ~w19853;
assign w19855 = w18092 & w19852;
assign w19856 = ~w19854 & ~w19855;
assign w19857 = pi02191 & ~w16225;
assign w19858 = ~pi10625 & w16225;
assign w19859 = ~w19857 & ~w19858;
assign w19860 = ~w16992 & w19149;
assign w19861 = pi02192 & ~w19860;
assign w19862 = ~pi02169 & w19860;
assign w19863 = ~w19861 & ~w19862;
assign w19864 = pi02193 & ~w16225;
assign w19865 = ~pi10647 & w16225;
assign w19866 = ~w19864 & ~w19865;
assign w19867 = pi02194 & ~w16229;
assign w19868 = ~pi10652 & w16229;
assign w19869 = ~w19867 & ~w19868;
assign w19870 = pi02195 & ~w19853;
assign w19871 = w18067 & w19852;
assign w19872 = ~w19870 & ~w19871;
assign w19873 = pi02196 & ~w19145;
assign w19874 = w17361 & w17586;
assign w19875 = ~w19873 & ~w19874;
assign w19876 = ~w16892 & w17406;
assign w19877 = pi02197 & ~w19876;
assign w19878 = ~pi02723 & w19876;
assign w19879 = ~w19877 & ~w19878;
assign w19880 = ~w16905 & w18291;
assign w19881 = pi02198 & ~w19880;
assign w19882 = ~pi02711 & w19880;
assign w19883 = ~w19881 & ~w19882;
assign w19884 = ~w16992 & w19106;
assign w19885 = pi02199 & ~w19884;
assign w19886 = ~pi02169 & w19884;
assign w19887 = ~w19885 & ~w19886;
assign w19888 = ~w16992 & w19530;
assign w19889 = pi02200 & ~w19888;
assign w19890 = ~pi02721 & w19888;
assign w19891 = ~w19889 & ~w19890;
assign w19892 = pi02201 & ~w16233;
assign w19893 = ~pi10624 & w16233;
assign w19894 = ~w19892 & ~w19893;
assign w19895 = ~w16992 & w17060;
assign w19896 = pi02202 & ~w19895;
assign w19897 = ~pi02722 & w19895;
assign w19898 = ~w19896 & ~w19897;
assign w19899 = ~w16992 & w17131;
assign w19900 = pi02203 & ~w19899;
assign w19901 = ~pi02164 & w19899;
assign w19902 = ~w19900 & ~w19901;
assign w19903 = pi02204 & ~w19895;
assign w19904 = w17060 & w19797;
assign w19905 = ~w19903 & ~w19904;
assign w19906 = pi02205 & ~w19783;
assign w19907 = w17620 & w19435;
assign w19908 = ~w19906 & ~w19907;
assign w19909 = w16953 & w17374;
assign w19910 = ~w16892 & w19909;
assign w19911 = pi02206 & ~w19910;
assign w19912 = ~pi02706 & w19910;
assign w19913 = ~w19911 & ~w19912;
assign w19914 = ~w16992 & w17380;
assign w19915 = pi02207 & ~w19914;
assign w19916 = w17380 & w19797;
assign w19917 = ~w19915 & ~w19916;
assign w19918 = w16948 & ~w16992;
assign w19919 = pi02208 & ~w19918;
assign w19920 = ~pi02722 & w19918;
assign w19921 = ~w19919 & ~w19920;
assign w19922 = ~w16992 & w19561;
assign w19923 = pi02209 & ~w19922;
assign w19924 = w17811 & w19561;
assign w19925 = ~w19923 & ~w19924;
assign w19926 = ~w16892 & w17006;
assign w19927 = pi02210 & ~w19926;
assign w19928 = ~pi02723 & w19926;
assign w19929 = ~w19927 & ~w19928;
assign w19930 = w16921 & w16969;
assign w19931 = ~w16892 & w19930;
assign w19932 = pi02211 & ~w19931;
assign w19933 = ~pi02710 & w19931;
assign w19934 = ~w19932 & ~w19933;
assign w19935 = pi02212 & ~w19497;
assign w19936 = ~pi09848 & w19497;
assign w19937 = ~w19935 & ~w19936;
assign w19938 = pi02213 & ~w19931;
assign w19939 = ~pi02706 & w19931;
assign w19940 = ~w19938 & ~w19939;
assign w19941 = w16947 & w17374;
assign w19942 = ~w16892 & w19941;
assign w19943 = pi02214 & ~w19942;
assign w19944 = ~pi02709 & w19942;
assign w19945 = ~w19943 & ~w19944;
assign w19946 = ~w16992 & w19552;
assign w19947 = pi02215 & ~w19946;
assign w19948 = ~pi02721 & w19946;
assign w19949 = ~w19947 & ~w19948;
assign w19950 = pi02216 & ~w16244;
assign w19951 = ~pi10640 & w16244;
assign w19952 = ~w19950 & ~w19951;
assign w19953 = pi02217 & ~w16244;
assign w19954 = ~pi10633 & w16244;
assign w19955 = ~w19953 & ~w19954;
assign w19956 = pi02218 & ~w19918;
assign w19957 = ~pi02169 & w19918;
assign w19958 = ~w19956 & ~w19957;
assign w19959 = ~w16992 & w17218;
assign w19960 = pi02219 & ~w19959;
assign w19961 = w17218 & w19797;
assign w19962 = ~w19960 & ~w19961;
assign w19963 = ~w16905 & w18009;
assign w19964 = pi02220 & ~w19963;
assign w19965 = ~pi02712 & w19963;
assign w19966 = ~w19964 & ~w19965;
assign w19967 = ~w16905 & w18468;
assign w19968 = pi02221 & ~w19967;
assign w19969 = ~pi02714 & w19967;
assign w19970 = ~w19968 & ~w19969;
assign w19971 = pi02222 & ~w19922;
assign w19972 = w17620 & w19561;
assign w19973 = ~w19971 & ~w19972;
assign w19974 = ~w16992 & w17977;
assign w19975 = pi02223 & ~w19974;
assign w19976 = ~pi02722 & w19974;
assign w19977 = ~w19975 & ~w19976;
assign w19978 = ~w16992 & w19601;
assign w19979 = pi02224 & ~w19978;
assign w19980 = ~pi02721 & w19978;
assign w19981 = ~w19979 & ~w19980;
assign w19982 = pi02225 & ~w19942;
assign w19983 = w18067 & w19941;
assign w19984 = ~w19982 & ~w19983;
assign w19985 = pi02226 & ~w16261;
assign w19986 = ~pi10631 & w16261;
assign w19987 = ~w19985 & ~w19986;
assign w19988 = w16895 & w16930;
assign w19989 = ~w16892 & w19988;
assign w19990 = pi02227 & ~w19989;
assign w19991 = ~pi02707 & w19989;
assign w19992 = ~w19990 & ~w19991;
assign w19993 = pi02228 & ~w16251;
assign w19994 = ~pi10638 & w16251;
assign w19995 = ~w19993 & ~w19994;
assign w19996 = w16899 & ~w16992;
assign w19997 = pi02229 & ~w19996;
assign w19998 = ~pi02722 & w19996;
assign w19999 = ~w19997 & ~w19998;
assign w20000 = ~w16992 & w17754;
assign w20001 = pi02230 & ~w20000;
assign w20002 = w17754 & w19797;
assign w20003 = ~w20001 & ~w20002;
assign w20004 = pi02231 & ~w19996;
assign w20005 = ~pi02169 & w19996;
assign w20006 = ~w20004 & ~w20005;
assign w20007 = ~w16992 & w19606;
assign w20008 = pi02232 & ~w20007;
assign w20009 = ~pi02721 & w20007;
assign w20010 = ~w20008 & ~w20009;
assign w20011 = pi02233 & ~w19787;
assign w20012 = ~pi02705 & w19787;
assign w20013 = ~w20011 & ~w20012;
assign w20014 = w16895 & w17189;
assign w20015 = ~w16892 & w20014;
assign w20016 = pi02234 & ~w20015;
assign w20017 = ~pi02160 & w20015;
assign w20018 = ~w20016 & ~w20017;
assign w20019 = pi02235 & ~w16214;
assign w20020 = ~pi10644 & w16214;
assign w20021 = ~w20019 & ~w20020;
assign w20022 = pi02236 & ~w20007;
assign w20023 = ~pi02164 & w20007;
assign w20024 = ~w20022 & ~w20023;
assign w20025 = pi02237 & ~w19914;
assign w20026 = ~pi02164 & w19914;
assign w20027 = ~w20025 & ~w20026;
assign w20028 = pi10629 & ~w16408;
assign w20029 = ~pi02238 & w16408;
assign w20030 = ~w20028 & ~w20029;
assign w20031 = pi02239 & ~w19974;
assign w20032 = ~pi02721 & w19974;
assign w20033 = ~w20031 & ~w20032;
assign w20034 = ~w16892 & w17912;
assign w20035 = pi02240 & ~w20034;
assign w20036 = ~pi02709 & w20034;
assign w20037 = ~w20035 & ~w20036;
assign w20038 = ~w16992 & w19660;
assign w20039 = pi02241 & ~w20038;
assign w20040 = ~pi02721 & w20038;
assign w20041 = ~w20039 & ~w20040;
assign w20042 = pi02242 & ~w20038;
assign w20043 = ~pi02164 & w20038;
assign w20044 = ~w20042 & ~w20043;
assign w20045 = ~w16992 & w19645;
assign w20046 = pi02243 & ~w20045;
assign w20047 = ~pi02721 & w20045;
assign w20048 = ~w20046 & ~w20047;
assign w20049 = pi02244 & ~w18848;
assign w20050 = ~pi02720 & w18848;
assign w20051 = ~w20049 & ~w20050;
assign w20052 = ~w16992 & w19576;
assign w20053 = pi02245 & ~w20052;
assign w20054 = ~pi02164 & w20052;
assign w20055 = ~w20053 & ~w20054;
assign w20056 = pi10653 & ~w16408;
assign w20057 = ~pi02246 & w16408;
assign w20058 = ~w20056 & ~w20057;
assign w20059 = w16895 & w17582;
assign w20060 = ~w16892 & w20059;
assign w20061 = pi02247 & ~w20060;
assign w20062 = ~pi02707 & w20060;
assign w20063 = ~w20061 & ~w20062;
assign w20064 = ~w16992 & w19624;
assign w20065 = pi02248 & ~w20064;
assign w20066 = ~pi02721 & w20064;
assign w20067 = ~w20065 & ~w20066;
assign w20068 = ~w16905 & w17183;
assign w20069 = pi02249 & ~w20068;
assign w20070 = ~pi02717 & w20068;
assign w20071 = ~w20069 & ~w20070;
assign w20072 = pi10651 & ~w16408;
assign w20073 = ~pi02250 & w16408;
assign w20074 = ~w20072 & ~w20073;
assign w20075 = w17016 & w17374;
assign w20076 = ~w16892 & w20075;
assign w20077 = pi02251 & ~w20076;
assign w20078 = ~pi02709 & w20076;
assign w20079 = ~w20077 & ~w20078;
assign w20080 = ~w16892 & w17078;
assign w20081 = pi02252 & ~w20080;
assign w20082 = w17078 & w18067;
assign w20083 = ~w20081 & ~w20082;
assign w20084 = pi10642 & ~w16408;
assign w20085 = ~pi02253 & w16408;
assign w20086 = ~w20084 & ~w20085;
assign w20087 = pi02254 & ~w20076;
assign w20088 = ~pi02707 & w20076;
assign w20089 = ~w20087 & ~w20088;
assign w20090 = ~w16928 & w16941;
assign w20091 = pi02255 & ~w20090;
assign w20092 = ~pi02720 & w20090;
assign w20093 = ~w20091 & ~w20092;
assign w20094 = pi10640 & ~w16408;
assign w20095 = ~pi02256 & w16408;
assign w20096 = ~w20094 & ~w20095;
assign w20097 = ~w16892 & w17103;
assign w20098 = pi02257 & ~w20097;
assign w20099 = ~pi02709 & w20097;
assign w20100 = ~w20098 & ~w20099;
assign w20101 = pi02258 & ~w20097;
assign w20102 = ~pi02707 & w20097;
assign w20103 = ~w20101 & ~w20102;
assign w20104 = ~w16992 & w19650;
assign w20105 = pi02259 & ~w20104;
assign w20106 = ~pi02164 & w20104;
assign w20107 = ~w20105 & ~w20106;
assign w20108 = pi02260 & ~w19402;
assign w20109 = ~pi02711 & w19402;
assign w20110 = ~w20108 & ~w20109;
assign w20111 = ~w16892 & w17053;
assign w20112 = pi02261 & ~w20111;
assign w20113 = ~pi02705 & w20111;
assign w20114 = ~w20112 & ~w20113;
assign w20115 = ~w16892 & w16954;
assign w20116 = pi02262 & ~w20115;
assign w20117 = ~pi02707 & w20115;
assign w20118 = ~w20116 & ~w20117;
assign w20119 = w16953 & w16977;
assign w20120 = ~w16892 & w20119;
assign w20121 = pi02263 & ~w20120;
assign w20122 = ~pi02709 & w20120;
assign w20123 = ~w20121 & ~w20122;
assign w20124 = pi02264 & ~w20111;
assign w20125 = ~pi02723 & w20111;
assign w20126 = ~w20124 & ~w20125;
assign w20127 = pi02265 & ~w20120;
assign w20128 = ~pi02707 & w20120;
assign w20129 = ~w20127 & ~w20128;
assign w20130 = pi02266 & ~w20104;
assign w20131 = w17811 & w19650;
assign w20132 = ~w20130 & ~w20131;
assign w20133 = pi02267 & ~w19974;
assign w20134 = ~pi02167 & w19974;
assign w20135 = ~w20133 & ~w20134;
assign w20136 = ~w16892 & w17626;
assign w20137 = pi02268 & ~w20136;
assign w20138 = ~pi02707 & w20136;
assign w20139 = ~w20137 & ~w20138;
assign w20140 = ~w16992 & w19679;
assign w20141 = pi02269 & ~w20140;
assign w20142 = ~pi02721 & w20140;
assign w20143 = ~w20141 & ~w20142;
assign w20144 = pi02270 & ~w20034;
assign w20145 = ~pi02707 & w20034;
assign w20146 = ~w20144 & ~w20145;
assign w20147 = ~w16892 & w17028;
assign w20148 = pi02271 & ~w20147;
assign w20149 = w17028 & w17671;
assign w20150 = ~w20148 & ~w20149;
assign w20151 = ~w16905 & w16961;
assign w20152 = pi02272 & ~w20151;
assign w20153 = ~pi02716 & w20151;
assign w20154 = ~w20152 & ~w20153;
assign w20155 = ~w16905 & w17461;
assign w20156 = pi02273 & ~w20155;
assign w20157 = ~pi02713 & w20155;
assign w20158 = ~w20156 & ~w20157;
assign w20159 = pi02274 & ~w20000;
assign w20160 = w17754 & w17811;
assign w20161 = ~w20159 & ~w20160;
assign w20162 = ~w16992 & w17314;
assign w20163 = pi02275 & ~w20162;
assign w20164 = ~pi02719 & w20162;
assign w20165 = ~w20163 & ~w20164;
assign w20166 = ~w16992 & w17535;
assign w20167 = pi02276 & ~w20166;
assign w20168 = w17535 & w17594;
assign w20169 = ~w20167 & ~w20168;
assign w20170 = w17052 & w17189;
assign w20171 = ~w16905 & w20170;
assign w20172 = pi02277 & ~w20171;
assign w20173 = ~pi02717 & w20171;
assign w20174 = ~w20172 & ~w20173;
assign w20175 = pi02278 & ~w19694;
assign w20176 = w17594 & w17762;
assign w20177 = ~w20175 & ~w20176;
assign w20178 = pi02279 & ~w20162;
assign w20179 = ~pi02718 & w20162;
assign w20180 = ~w20178 & ~w20179;
assign w20181 = ~w16905 & w17710;
assign w20182 = pi02280 & ~w20181;
assign w20183 = ~pi02711 & w20181;
assign w20184 = ~w20182 & ~w20183;
assign w20185 = ~w16905 & w16931;
assign w20186 = pi02281 & ~w20185;
assign w20187 = ~pi02716 & w20185;
assign w20188 = ~w20186 & ~w20187;
assign w20189 = ~w16905 & w17119;
assign w20190 = pi02282 & ~w20189;
assign w20191 = w17020 & w17119;
assign w20192 = ~w20190 & ~w20191;
assign w20193 = ~w16905 & w17398;
assign w20194 = pi02283 & ~w20193;
assign w20195 = ~pi02716 & w20193;
assign w20196 = ~w20194 & ~w20195;
assign w20197 = pi02284 & ~w20181;
assign w20198 = ~pi02714 & w20181;
assign w20199 = ~w20197 & ~w20198;
assign w20200 = ~w16992 & w18217;
assign w20201 = pi02285 & ~w20200;
assign w20202 = ~pi02719 & w20200;
assign w20203 = ~w20201 & ~w20202;
assign w20204 = ~w16992 & w17334;
assign w20205 = pi02286 & ~w20204;
assign w20206 = ~pi02718 & w20204;
assign w20207 = ~w20205 & ~w20206;
assign w20208 = pi02287 & ~w20185;
assign w20209 = ~pi02170 & ~w16905;
assign w20210 = w16931 & w20209;
assign w20211 = ~w20208 & ~w20210;
assign w20212 = pi02288 & ~w20193;
assign w20213 = ~pi02712 & w20193;
assign w20214 = ~w20212 & ~w20213;
assign w20215 = ~w16928 & w17011;
assign w20216 = pi02289 & ~w20215;
assign w20217 = w17011 & w17128;
assign w20218 = ~w20216 & ~w20217;
assign w20219 = pi02290 & ~w18527;
assign w20220 = w18059 & w18526;
assign w20221 = ~w20219 & ~w20220;
assign w20222 = ~w16905 & w17466;
assign w20223 = pi02291 & ~w20222;
assign w20224 = ~pi02170 & w20222;
assign w20225 = ~w20223 & ~w20224;
assign w20226 = ~w16992 & w17907;
assign w20227 = pi02292 & ~w20226;
assign w20228 = ~pi02167 & w20226;
assign w20229 = ~w20227 & ~w20228;
assign w20230 = ~w16905 & w17231;
assign w20231 = pi02293 & ~w20230;
assign w20232 = w17231 & w18059;
assign w20233 = ~w20231 & ~w20232;
assign w20234 = pi02294 & ~w20171;
assign w20235 = ~pi02712 & w20171;
assign w20236 = ~w20234 & ~w20235;
assign w20237 = ~w16892 & w18032;
assign w20238 = pi02295 & ~w20237;
assign w20239 = ~pi02708 & w20237;
assign w20240 = ~w20238 & ~w20239;
assign w20241 = pi02296 & ~w18535;
assign w20242 = w17047 & w18578;
assign w20243 = ~w20241 & ~w20242;
assign w20244 = w16983 & w17037;
assign w20245 = ~w16892 & w20244;
assign w20246 = pi02297 & ~w20245;
assign w20247 = w17671 & w20244;
assign w20248 = ~w20246 & ~w20247;
assign w20249 = ~w16992 & w19282;
assign w20250 = pi02298 & ~w20249;
assign w20251 = ~pi02164 & w20249;
assign w20252 = ~w20250 & ~w20251;
assign w20253 = ~w16992 & w19723;
assign w20254 = pi02299 & ~w20253;
assign w20255 = ~pi02721 & w20253;
assign w20256 = ~w20254 & ~w20255;
assign w20257 = w16912 & ~w16992;
assign w20258 = pi02300 & ~w20257;
assign w20259 = ~pi02164 & w20257;
assign w20260 = ~w20258 & ~w20259;
assign w20261 = ~w16905 & w17344;
assign w20262 = pi02301 & ~w20261;
assign w20263 = w17344 & w17929;
assign w20264 = ~w20262 & ~w20263;
assign w20265 = ~w16992 & w17521;
assign w20266 = pi02302 & ~w20265;
assign w20267 = ~pi02167 & w20265;
assign w20268 = ~w20266 & ~w20267;
assign w20269 = ~w16905 & w17479;
assign w20270 = pi02303 & ~w20269;
assign w20271 = ~pi02714 & w20269;
assign w20272 = ~w20270 & ~w20271;
assign w20273 = ~w16892 & w17249;
assign w20274 = pi02304 & ~w20273;
assign w20275 = w17249 & w18689;
assign w20276 = ~w20274 & ~w20275;
assign w20277 = ~w16892 & w16994;
assign w20278 = pi02305 & ~w20277;
assign w20279 = ~pi02709 & w20277;
assign w20280 = ~w20278 & ~w20279;
assign w20281 = ~w16928 & w18454;
assign w20282 = pi02306 & ~w20281;
assign w20283 = ~pi09812 & w20281;
assign w20284 = ~w20282 & ~w20283;
assign w20285 = ~w16905 & w18572;
assign w20286 = pi02307 & ~w20285;
assign w20287 = ~pi02170 & w20285;
assign w20288 = ~w20286 & ~w20287;
assign w20289 = pi02308 & ~w20265;
assign w20290 = ~pi02719 & w20265;
assign w20291 = ~w20289 & ~w20290;
assign w20292 = ~w16992 & w17668;
assign w20293 = pi02309 & ~w20292;
assign w20294 = w17668 & w19273;
assign w20295 = ~w20293 & ~w20294;
assign w20296 = pi02310 & ~w20200;
assign w20297 = ~pi02718 & w20200;
assign w20298 = ~w20296 & ~w20297;
assign w20299 = ~w16992 & w18726;
assign w20300 = pi02311 & ~w20299;
assign w20301 = ~pi02164 & w20299;
assign w20302 = ~w20300 & ~w20301;
assign w20303 = pi02312 & ~w20068;
assign w20304 = ~pi02711 & w20068;
assign w20305 = ~w20303 & ~w20304;
assign w20306 = ~w16905 & w17996;
assign w20307 = pi02313 & ~w20306;
assign w20308 = ~pi02711 & w20306;
assign w20309 = ~w20307 & ~w20308;
assign w20310 = ~w16905 & w18636;
assign w20311 = pi02314 & ~w20310;
assign w20312 = ~pi02711 & w20310;
assign w20313 = ~w20311 & ~w20312;
assign w20314 = ~w16905 & w17636;
assign w20315 = pi02315 & ~w20314;
assign w20316 = ~pi02716 & w20314;
assign w20317 = ~w20315 & ~w20316;
assign w20318 = ~w16892 & w17114;
assign w20319 = pi02316 & ~w20318;
assign w20320 = ~pi02709 & w20318;
assign w20321 = ~w20319 & ~w20320;
assign w20322 = ~w16905 & w18726;
assign w20323 = pi02317 & ~w20322;
assign w20324 = w17603 & w18726;
assign w20325 = ~w20323 & ~w20324;
assign w20326 = ~w16992 & w18348;
assign w20327 = pi02318 & ~w20326;
assign w20328 = ~pi02167 & w20326;
assign w20329 = ~w20327 & ~w20328;
assign w20330 = ~w16905 & w17244;
assign w20331 = pi02319 & ~w20330;
assign w20332 = ~pi02712 & w20330;
assign w20333 = ~w20331 & ~w20332;
assign w20334 = pi02320 & ~w20310;
assign w20335 = ~pi02717 & w20310;
assign w20336 = ~w20334 & ~w20335;
assign w20337 = ~w16905 & w17162;
assign w20338 = pi02321 & ~w20337;
assign w20339 = ~pi02716 & w20337;
assign w20340 = ~w20338 & ~w20339;
assign w20341 = pi02322 & ~w20257;
assign w20342 = ~pi02703 & w20257;
assign w20343 = ~w20341 & ~w20342;
assign w20344 = pi02323 & ~w20318;
assign w20345 = ~pi02160 & w20318;
assign w20346 = ~w20344 & ~w20345;
assign w20347 = pi02324 & ~w20322;
assign w20348 = ~pi02714 & w20322;
assign w20349 = ~w20347 & ~w20348;
assign w20350 = pi02325 & ~w20306;
assign w20351 = w17742 & w17996;
assign w20352 = ~w20350 & ~w20351;
assign w20353 = ~w16892 & w17965;
assign w20354 = pi02326 & ~w20353;
assign w20355 = ~pi02707 & w20353;
assign w20356 = ~w20354 & ~w20355;
assign w20357 = pi02327 & ~w20261;
assign w20358 = ~pi02717 & w20261;
assign w20359 = ~w20357 & ~w20358;
assign w20360 = pi02328 & ~w20318;
assign w20361 = ~pi02705 & w20318;
assign w20362 = ~w20360 & ~w20361;
assign w20363 = pi02329 & ~w20314;
assign w20364 = ~pi02712 & w20314;
assign w20365 = ~w20363 & ~w20364;
assign w20366 = ~w16928 & w18542;
assign w20367 = pi02330 & ~w20366;
assign w20368 = ~pi09812 & w20366;
assign w20369 = ~w20367 & ~w20368;
assign w20370 = ~w16928 & w18617;
assign w20371 = pi02331 & ~w20370;
assign w20372 = ~pi02720 & w20370;
assign w20373 = ~w20371 & ~w20372;
assign w20374 = pi02332 & ~w20366;
assign w20375 = ~pi02720 & w20366;
assign w20376 = ~w20374 & ~w20375;
assign w20377 = pi02333 & ~w20269;
assign w20378 = ~pi02712 & w20269;
assign w20379 = ~w20377 & ~w20378;
assign w20380 = pi02334 & ~w20226;
assign w20381 = ~pi02721 & w20226;
assign w20382 = ~w20380 & ~w20381;
assign w20383 = pi02335 & ~w18062;
assign w20384 = ~pi02720 & w18062;
assign w20385 = ~w20383 & ~w20384;
assign w20386 = ~w16892 & w17573;
assign w20387 = pi02336 & ~w20386;
assign w20388 = ~pi02705 & w20386;
assign w20389 = ~w20387 & ~w20388;
assign w20390 = ~w16892 & w17609;
assign w20391 = pi02337 & ~w20390;
assign w20392 = ~pi02706 & w20390;
assign w20393 = ~w20391 & ~w20392;
assign w20394 = ~w16905 & w18454;
assign w20395 = pi02338 & ~w20394;
assign w20396 = ~pi02715 & w20394;
assign w20397 = ~w20395 & ~w20396;
assign w20398 = pi02339 & ~w20386;
assign w20399 = w17573 & w17671;
assign w20400 = ~w20398 & ~w20399;
assign w20401 = pi02340 & ~w20245;
assign w20402 = ~pi02705 & w20245;
assign w20403 = ~w20401 & ~w20402;
assign w20404 = pi02341 & ~w14136;
assign w20405 = pi10357 & w14136;
assign w20406 = ~w20404 & ~w20405;
assign w20407 = ~w16892 & w18070;
assign w20408 = pi02342 & ~w20407;
assign w20409 = ~pi02707 & w20407;
assign w20410 = ~w20408 & ~w20409;
assign w20411 = ~w16892 & w17017;
assign w20412 = pi02343 & ~w20411;
assign w20413 = ~pi02709 & w20411;
assign w20414 = ~w20412 & ~w20413;
assign w20415 = ~w16892 & w17822;
assign w20416 = pi02344 & ~w20415;
assign w20417 = w17822 & w18578;
assign w20418 = ~w20416 & ~w20417;
assign w20419 = pi02345 & ~w20237;
assign w20420 = ~pi02706 & w20237;
assign w20421 = ~w20419 & ~w20420;
assign w20422 = pi02346 & ~w18741;
assign w20423 = ~pi02712 & w18741;
assign w20424 = ~w20422 & ~w20423;
assign w20425 = ~w16992 & w17279;
assign w20426 = pi02347 & ~w20425;
assign w20427 = ~pi02164 & w20425;
assign w20428 = ~w20426 & ~w20427;
assign w20429 = ~pi00880 & pi02348;
assign w20430 = ~w12984 & w20429;
assign w20431 = w12993 & w20430;
assign w20432 = ~pi00209 & w11150;
assign w20433 = w2040 & w20432;
assign w20434 = ~w15945 & ~w20433;
assign w20435 = pi09927 & ~pi10030;
assign w20436 = w10683 & w20435;
assign w20437 = ~w20434 & w20436;
assign w20438 = ~w20431 & ~w20437;
assign w20439 = pi02349 & ~w20415;
assign w20440 = ~pi02723 & w20415;
assign w20441 = ~w20439 & ~w20440;
assign w20442 = ~w16905 & w17320;
assign w20443 = pi02350 & ~w20442;
assign w20444 = ~pi02717 & w20442;
assign w20445 = ~w20443 & ~w20444;
assign w20446 = ~w16892 & w17108;
assign w20447 = pi02351 & ~w20446;
assign w20448 = ~pi02723 & w20446;
assign w20449 = ~w20447 & ~w20448;
assign w20450 = ~w16892 & w17231;
assign w20451 = pi02352 & ~w20450;
assign w20452 = w17231 & w18092;
assign w20453 = ~w20451 & ~w20452;
assign w20454 = pi02353 & ~w20277;
assign w20455 = ~pi02707 & w20277;
assign w20456 = ~w20454 & ~w20455;
assign w20457 = ~w16892 & w17814;
assign w20458 = pi02354 & ~w20457;
assign w20459 = ~pi02723 & w20457;
assign w20460 = ~w20458 & ~w20459;
assign w20461 = ~w16992 & w17631;
assign w20462 = pi02355 & ~w20461;
assign w20463 = w17631 & w19273;
assign w20464 = ~w20462 & ~w20463;
assign w20465 = w16960 & w17182;
assign w20466 = ~w16892 & w20465;
assign w20467 = pi02356 & ~w20466;
assign w20468 = ~pi02723 & w20466;
assign w20469 = ~w20467 & ~w20468;
assign w20470 = w17016 & w17582;
assign w20471 = ~w16892 & w20470;
assign w20472 = pi02357 & ~w20471;
assign w20473 = ~pi02706 & w20471;
assign w20474 = ~w20472 & ~w20473;
assign w20475 = pi02358 & ~w20446;
assign w20476 = ~pi02705 & w20446;
assign w20477 = ~w20475 & ~w20476;
assign w20478 = ~w16892 & w17837;
assign w20479 = pi02359 & ~w20478;
assign w20480 = w17837 & w18689;
assign w20481 = ~w20479 & ~w20480;
assign w20482 = pi02360 & ~w20466;
assign w20483 = ~pi02705 & w20466;
assign w20484 = ~w20482 & ~w20483;
assign w20485 = ~w16992 & w18745;
assign w20486 = pi02361 & ~w20485;
assign w20487 = ~pi02722 & w20485;
assign w20488 = ~w20486 & ~w20487;
assign w20489 = ~w16892 & w17011;
assign w20490 = pi02362 & ~w20489;
assign w20491 = ~pi02707 & w20489;
assign w20492 = ~w20490 & ~w20491;
assign w20493 = ~w16905 & w18027;
assign w20494 = pi02363 & ~w20493;
assign w20495 = ~pi02711 & w20493;
assign w20496 = ~w20494 & ~w20495;
assign w20497 = ~w16992 & w19728;
assign w20498 = pi02364 & ~w20497;
assign w20499 = ~pi02164 & w20497;
assign w20500 = ~w20498 & ~w20499;
assign w20501 = ~w16905 & w17366;
assign w20502 = pi02365 & ~w20501;
assign w20503 = ~pi02712 & w20501;
assign w20504 = ~w20502 & ~w20503;
assign w20505 = ~w16928 & w20075;
assign w20506 = pi02366 & ~w20505;
assign w20507 = ~pi09954 & w20505;
assign w20508 = ~w20506 & ~w20507;
assign w20509 = pi02367 & ~w20485;
assign w20510 = ~pi02721 & w20485;
assign w20511 = ~w20509 & ~w20510;
assign w20512 = ~w16992 & w18022;
assign w20513 = pi02368 & ~w20512;
assign w20514 = w17620 & w18022;
assign w20515 = ~w20513 & ~w20514;
assign w20516 = pi02369 & ~w20489;
assign w20517 = ~pi02705 & w20489;
assign w20518 = ~w20516 & ~w20517;
assign w20519 = ~w16892 & w17658;
assign w20520 = pi02370 & ~w20519;
assign w20521 = ~pi02723 & w20519;
assign w20522 = ~w20520 & ~w20521;
assign w20523 = ~w16892 & w17479;
assign w20524 = pi02371 & ~w20523;
assign w20525 = ~pi02708 & w20523;
assign w20526 = ~w20524 & ~w20525;
assign w20527 = ~w16892 & w17398;
assign w20528 = pi02372 & ~w20527;
assign w20529 = ~pi02705 & w20527;
assign w20530 = ~w20528 & ~w20529;
assign w20531 = ~w16992 & w17917;
assign w20532 = pi02373 & ~w20531;
assign w20533 = w17917 & w19312;
assign w20534 = ~w20532 & ~w20533;
assign w20535 = pi02374 & ~w20512;
assign w20536 = w17532 & w18022;
assign w20537 = ~w20535 & ~w20536;
assign w20538 = ~w16892 & w18001;
assign w20539 = pi02375 & ~w20538;
assign w20540 = ~pi02708 & w20538;
assign w20541 = ~w20539 & ~w20540;
assign w20542 = pi02376 & ~w20497;
assign w20543 = ~pi02721 & w20497;
assign w20544 = ~w20542 & ~w20543;
assign w20545 = ~w16892 & w18278;
assign w20546 = pi02377 & ~w20545;
assign w20547 = ~pi02708 & w20545;
assign w20548 = ~w20546 & ~w20547;
assign w20549 = ~w16892 & w17137;
assign w20550 = pi02378 & ~w20549;
assign w20551 = ~pi02707 & w20549;
assign w20552 = ~w20550 & ~w20551;
assign w20553 = ~w16992 & w17305;
assign w20554 = pi02379 & ~w20553;
assign w20555 = ~pi02722 & w20553;
assign w20556 = ~w20554 & ~w20555;
assign w20557 = ~w16992 & w19740;
assign w20558 = pi02380 & ~w20557;
assign w20559 = ~pi02721 & w20557;
assign w20560 = ~w20558 & ~w20559;
assign w20561 = w16895 & w17374;
assign w20562 = ~w16892 & w20561;
assign w20563 = pi02381 & ~w20562;
assign w20564 = ~pi02707 & w20562;
assign w20565 = ~w20563 & ~w20564;
assign w20566 = w16919 & w17189;
assign w20567 = ~w16905 & w20566;
assign w20568 = pi02382 & ~w20567;
assign w20569 = ~pi02715 & w20567;
assign w20570 = ~w20568 & ~w20569;
assign w20571 = pi02383 & ~w20538;
assign w20572 = ~pi02706 & w20538;
assign w20573 = ~w20571 & ~w20572;
assign w20574 = ~w16892 & w17938;
assign w20575 = pi02384 & ~w20574;
assign w20576 = w17938 & w18689;
assign w20577 = ~w20575 & ~w20576;
assign w20578 = pi02385 & ~w20519;
assign w20579 = ~pi02710 & w20519;
assign w20580 = ~w20578 & ~w20579;
assign w20581 = ~w16892 & w18056;
assign w20582 = pi02386 & ~w20581;
assign w20583 = ~pi02707 & w20581;
assign w20584 = ~w20582 & ~w20583;
assign w20585 = pi02387 & ~w20574;
assign w20586 = w17938 & w18578;
assign w20587 = ~w20585 & ~w20586;
assign w20588 = ~w16892 & w16941;
assign w20589 = pi02388 & ~w20588;
assign w20590 = ~pi02708 & w20588;
assign w20591 = ~w20589 & ~w20590;
assign w20592 = ~w16905 & w19343;
assign w20593 = pi02389 & ~w20592;
assign w20594 = ~pi02716 & w20592;
assign w20595 = ~w20593 & ~w20594;
assign w20596 = ~w16892 & w17428;
assign w20597 = pi02390 & ~w20596;
assign w20598 = w17428 & w18067;
assign w20599 = ~w20597 & ~w20598;
assign w20600 = ~w16892 & w17289;
assign w20601 = pi02391 & ~w20600;
assign w20602 = ~pi02707 & w20600;
assign w20603 = ~w20601 & ~w20602;
assign w20604 = ~w16905 & w19374;
assign w20605 = pi02392 & ~w20604;
assign w20606 = ~pi02714 & w20604;
assign w20607 = ~w20605 & ~w20606;
assign w20608 = pi02393 & ~w20592;
assign w20609 = ~pi02712 & w20592;
assign w20610 = ~w20608 & ~w20609;
assign w20611 = pi02394 & ~w20411;
assign w20612 = ~pi02707 & w20411;
assign w20613 = ~w20611 & ~w20612;
assign w20614 = pi02395 & ~w20493;
assign w20615 = ~pi02717 & w20493;
assign w20616 = ~w20614 & ~w20615;
assign w20617 = ~w16892 & w17445;
assign w20618 = pi02396 & ~w20617;
assign w20619 = ~pi02707 & w20617;
assign w20620 = ~w20618 & ~w20619;
assign w20621 = ~w16928 & w17490;
assign w20622 = pi02397 & ~w20621;
assign w20623 = ~pi09954 & w20621;
assign w20624 = ~w20622 & ~w20623;
assign w20625 = ~w16892 & w18740;
assign w20626 = pi02398 & ~w20625;
assign w20627 = ~pi02723 & w20625;
assign w20628 = ~w20626 & ~w20627;
assign w20629 = ~w16892 & w17210;
assign w20630 = pi02399 & ~w20629;
assign w20631 = ~pi02709 & w20629;
assign w20632 = ~w20630 & ~w20631;
assign w20633 = ~w16905 & w19348;
assign w20634 = pi02400 & ~w20633;
assign w20635 = w17020 & w19348;
assign w20636 = ~w20634 & ~w20635;
assign w20637 = ~w16892 & w18051;
assign w20638 = pi02401 & ~w20637;
assign w20639 = ~pi02709 & w20637;
assign w20640 = ~w20638 & ~w20639;
assign w20641 = pi02402 & ~w20523;
assign w20642 = ~pi02705 & w20523;
assign w20643 = ~w20641 & ~w20642;
assign w20644 = pi02403 & ~w20588;
assign w20645 = ~pi02706 & w20588;
assign w20646 = ~w20644 & ~w20645;
assign w20647 = ~w16892 & w17749;
assign w20648 = pi02404 & ~w20647;
assign w20649 = w17671 & w17749;
assign w20650 = ~w20648 & ~w20649;
assign w20651 = pi02405 & ~w20600;
assign w20652 = ~pi02708 & w20600;
assign w20653 = ~w20651 & ~w20652;
assign w20654 = pi02406 & ~w20647;
assign w20655 = ~pi02710 & w20647;
assign w20656 = ~w20654 & ~w20655;
assign w20657 = pi02407 & ~w20637;
assign w20658 = ~pi02707 & w20637;
assign w20659 = ~w20657 & ~w20658;
assign w20660 = ~w16892 & w17349;
assign w20661 = pi02408 & ~w20660;
assign w20662 = ~pi02709 & w20660;
assign w20663 = ~w20661 & ~w20662;
assign w20664 = ~w16892 & w17681;
assign w20665 = pi02409 & ~w20664;
assign w20666 = ~pi02706 & w20664;
assign w20667 = ~w20665 & ~w20666;
assign w20668 = pi02410 & ~w19541;
assign w20669 = ~pi02715 & w19541;
assign w20670 = ~w20668 & ~w20669;
assign w20671 = pi02411 & ~w20660;
assign w20672 = w17349 & w18067;
assign w20673 = ~w20671 & ~w20672;
assign w20674 = pi02412 & ~w20604;
assign w20675 = ~pi02716 & w20604;
assign w20676 = ~w20674 & ~w20675;
assign w20677 = pi02413 & ~w20647;
assign w20678 = ~pi02706 & w20647;
assign w20679 = ~w20677 & ~w20678;
assign w20680 = ~w16905 & w17855;
assign w20681 = pi02414 & ~w20680;
assign w20682 = ~pi02712 & w20680;
assign w20683 = ~w20681 & ~w20682;
assign w20684 = ~w16892 & w17385;
assign w20685 = pi02415 & ~w20684;
assign w20686 = ~pi02709 & w20684;
assign w20687 = ~w20685 & ~w20686;
assign w20688 = pi02416 & ~w20625;
assign w20689 = w18578 & w18740;
assign w20690 = ~w20688 & ~w20689;
assign w20691 = pi02417 & ~w20493;
assign w20692 = ~pi02714 & w20493;
assign w20693 = ~w20691 & ~w20692;
assign w20694 = ~w16928 & w18645;
assign w20695 = pi02418 & ~w20694;
assign w20696 = ~pi09848 & w20694;
assign w20697 = ~w20695 & ~w20696;
assign w20698 = ~w16992 & w17837;
assign w20699 = pi02419 & ~w20698;
assign w20700 = w17586 & w17837;
assign w20701 = ~w20699 & ~w20700;
assign w20702 = ~w16892 & w17183;
assign w20703 = pi02420 & ~w20702;
assign w20704 = ~pi02709 & w20702;
assign w20705 = ~w20703 & ~w20704;
assign w20706 = ~w16928 & w20244;
assign w20707 = pi02421 & ~w20706;
assign w20708 = w17193 & w20244;
assign w20709 = ~w20707 & ~w20708;
assign w20710 = pi02422 & ~w17501;
assign w20711 = ~pi09954 & w17501;
assign w20712 = ~w20710 & ~w20711;
assign w20713 = ~w16992 & w17749;
assign w20714 = pi02423 & ~w20713;
assign w20715 = ~pi02703 & w20713;
assign w20716 = ~w20714 & ~w20715;
assign w20717 = pi02424 & ~w20567;
assign w20718 = ~pi02713 & w20567;
assign w20719 = ~w20717 & ~w20718;
assign w20720 = w16919 & w17374;
assign w20721 = ~w16992 & w20720;
assign w20722 = pi02425 & ~w20721;
assign w20723 = ~pi02718 & w20721;
assign w20724 = ~w20722 & ~w20723;
assign w20725 = pi02426 & ~w20461;
assign w20726 = ~pi02703 & w20461;
assign w20727 = ~w20725 & ~w20726;
assign w20728 = pi02427 & ~w17149;
assign w20729 = ~pi09812 & w17149;
assign w20730 = ~w20728 & ~w20729;
assign w20731 = ~w16892 & w17663;
assign w20732 = pi02428 & ~w20731;
assign w20733 = ~pi02706 & w20731;
assign w20734 = ~w20732 & ~w20733;
assign w20735 = ~w16928 & w17535;
assign w20736 = pi02429 & ~w20735;
assign w20737 = ~pi02704 & w20735;
assign w20738 = ~w20736 & ~w20737;
assign w20739 = ~w16928 & w19282;
assign w20740 = pi02430 & ~w20739;
assign w20741 = ~pi09848 & w20739;
assign w20742 = ~w20740 & ~w20741;
assign w20743 = ~w16905 & w17023;
assign w20744 = pi02431 & ~w20743;
assign w20745 = ~pi02715 & w20743;
assign w20746 = ~w20744 & ~w20745;
assign w20747 = ~w16992 & w20470;
assign w20748 = pi02432 & ~w20747;
assign w20749 = ~pi02703 & w20747;
assign w20750 = ~w20748 & ~w20749;
assign w20751 = ~w16905 & w17039;
assign w20752 = pi02433 & ~w20751;
assign w20753 = ~pi02712 & w20751;
assign w20754 = ~w20752 & ~w20753;
assign w20755 = pi02434 & ~w20702;
assign w20756 = ~pi02707 & w20702;
assign w20757 = ~w20755 & ~w20756;
assign w20758 = ~w16905 & w18585;
assign w20759 = pi02435 & ~w20758;
assign w20760 = ~pi02715 & w20758;
assign w20761 = ~w20759 & ~w20760;
assign w20762 = pi02436 & ~w20553;
assign w20763 = ~pi02703 & w20553;
assign w20764 = ~w20762 & ~w20763;
assign w20765 = pi02437 & ~w20721;
assign w20766 = w17594 & w20720;
assign w20767 = ~w20765 & ~w20766;
assign w20768 = pi02438 & ~w20739;
assign w20769 = ~pi09954 & w20739;
assign w20770 = ~w20768 & ~w20769;
assign w20771 = ~w16992 & w17226;
assign w20772 = pi02439 & ~w20771;
assign w20773 = ~pi02719 & w20771;
assign w20774 = ~w20772 & ~w20773;
assign w20775 = w16919 & w17582;
assign w20776 = ~w16905 & w20775;
assign w20777 = pi02440 & ~w20776;
assign w20778 = w17317 & w20775;
assign w20779 = ~w20777 & ~w20778;
assign w20780 = ~w16992 & w17718;
assign w20781 = pi02441 & ~w20780;
assign w20782 = ~pi02703 & w20780;
assign w20783 = ~w20781 & ~w20782;
assign w20784 = pi02442 & ~w20735;
assign w20785 = ~pi09962 & w20735;
assign w20786 = ~w20784 & ~w20785;
assign w20787 = ~w16905 & w17172;
assign w20788 = pi02443 & ~w20787;
assign w20789 = ~pi02716 & w20787;
assign w20790 = ~w20788 & ~w20789;
assign w20791 = ~w16992 & w17411;
assign w20792 = pi02444 & ~w20791;
assign w20793 = ~pi02722 & w20791;
assign w20794 = ~w20792 & ~w20793;
assign w20795 = ~w16992 & w18300;
assign w20796 = pi02445 & ~w20795;
assign w20797 = ~pi02164 & w20795;
assign w20798 = ~w20796 & ~w20797;
assign w20799 = ~w16928 & w18622;
assign w20800 = pi02446 & ~w20799;
assign w20801 = w17128 & w18622;
assign w20802 = ~w20800 & ~w20801;
assign w20803 = pi02447 & ~w20758;
assign w20804 = ~pi02170 & w20758;
assign w20805 = ~w20803 & ~w20804;
assign w20806 = ~w16892 & w17172;
assign w20807 = pi02448 & ~w20806;
assign w20808 = ~pi02723 & w20806;
assign w20809 = ~w20807 & ~w20808;
assign w20810 = ~w16905 & w17583;
assign w20811 = pi02449 & ~w20810;
assign w20812 = ~pi02170 & w20810;
assign w20813 = ~w20811 & ~w20812;
assign w20814 = pi02450 & ~w20771;
assign w20815 = ~pi02718 & w20771;
assign w20816 = ~w20814 & ~w20815;
assign w20817 = ~w16905 & w17556;
assign w20818 = pi02451 & ~w20817;
assign w20819 = ~pi02716 & w20817;
assign w20820 = ~w20818 & ~w20819;
assign w20821 = ~w16928 & w17479;
assign w20822 = pi02452 & ~w20821;
assign w20823 = w17193 & w17479;
assign w20824 = ~w20822 & ~w20823;
assign w20825 = ~w16992 & w17461;
assign w20826 = pi02453 & ~w20825;
assign w20827 = ~pi02719 & w20825;
assign w20828 = ~w20826 & ~w20827;
assign w20829 = pi02454 & ~w20731;
assign w20830 = ~pi02708 & w20731;
assign w20831 = ~w20829 & ~w20830;
assign w20832 = pi02455 & ~w20596;
assign w20833 = ~pi02705 & w20596;
assign w20834 = ~w20832 & ~w20833;
assign w20835 = ~w16992 & w17119;
assign w20836 = pi02456 & ~w20835;
assign w20837 = ~pi02719 & w20835;
assign w20838 = ~w20836 & ~w20837;
assign w20839 = ~w16992 & w18468;
assign w20840 = pi02457 & ~w20839;
assign w20841 = ~pi02703 & w20839;
assign w20842 = ~w20840 & ~w20841;
assign w20843 = w16922 & ~w16992;
assign w20844 = pi02458 & ~w20843;
assign w20845 = w16922 & w17594;
assign w20846 = ~w20844 & ~w20845;
assign w20847 = pi02459 & ~w20839;
assign w20848 = ~pi02167 & w20839;
assign w20849 = ~w20847 & ~w20848;
assign w20850 = pi02460 & ~w20835;
assign w20851 = ~pi02718 & w20835;
assign w20852 = ~w20850 & ~w20851;
assign w20853 = pi02461 & ~w20407;
assign w20854 = ~pi02709 & w20407;
assign w20855 = ~w20853 & ~w20854;
assign w20856 = ~w16992 & w17710;
assign w20857 = pi02462 & ~w20856;
assign w20858 = ~pi02703 & w20856;
assign w20859 = ~w20857 & ~w20858;
assign w20860 = ~w16892 & w17023;
assign w20861 = pi02463 & ~w20860;
assign w20862 = ~pi02705 & w20860;
assign w20863 = ~w20861 & ~w20862;
assign w20864 = pi02464 & ~w20531;
assign w20865 = w17532 & w17917;
assign w20866 = ~w20864 & ~w20865;
assign w20867 = ~w16992 & w17855;
assign w20868 = pi02465 & ~w20867;
assign w20869 = ~pi02719 & w20867;
assign w20870 = ~w20868 & ~w20869;
assign w20871 = ~w16905 & w17977;
assign w20872 = pi02466 & ~w20871;
assign w20873 = ~pi02711 & w20871;
assign w20874 = ~w20872 & ~w20873;
assign w20875 = ~w16928 & w17249;
assign w20876 = pi02467 & ~w20875;
assign w20877 = ~pi09812 & w20875;
assign w20878 = ~w20876 & ~w20877;
assign w20879 = ~w16905 & w19327;
assign w20880 = pi02468 & ~w20879;
assign w20881 = ~pi02714 & w20879;
assign w20882 = ~w20880 & ~w20881;
assign w20883 = ~w16905 & w18554;
assign w20884 = pi02469 & ~w20883;
assign w20885 = w17603 & w18554;
assign w20886 = ~w20884 & ~w20885;
assign w20887 = ~w16928 & w18009;
assign w20888 = pi02470 & ~w20887;
assign w20889 = ~pi02720 & w20887;
assign w20890 = ~w20888 & ~w20889;
assign w20891 = ~w16905 & w19012;
assign w20892 = pi02471 & ~w20891;
assign w20893 = ~pi02716 & w20891;
assign w20894 = ~w20892 & ~w20893;
assign w20895 = ~w16905 & w18745;
assign w20896 = pi02472 & ~w20895;
assign w20897 = w18745 & w20209;
assign w20898 = ~w20896 & ~w20897;
assign w20899 = pi02473 & ~w20817;
assign w20900 = w17020 & w17556;
assign w20901 = ~w20899 & ~w20900;
assign w20902 = ~w16928 & w17636;
assign w20903 = pi02474 & ~w20902;
assign w20904 = ~pi02720 & w20902;
assign w20905 = ~w20903 & ~w20904;
assign w20906 = ~w16992 & w18454;
assign w20907 = pi02475 & ~w20906;
assign w20908 = ~pi02167 & w20906;
assign w20909 = ~w20907 & ~w20908;
assign w20910 = pi02476 & ~w20531;
assign w20911 = w17917 & w19273;
assign w20912 = ~w20910 & ~w20911;
assign w20913 = pi02477 & ~w17280;
assign w20914 = w17279 & w17311;
assign w20915 = ~w20913 & ~w20914;
assign w20916 = pi02478 & ~w20806;
assign w20917 = ~pi02705 & w20806;
assign w20918 = ~w20916 & ~w20917;
assign w20919 = ~w16928 & w18740;
assign w20920 = pi02479 & ~w20919;
assign w20921 = ~pi02720 & w20919;
assign w20922 = ~w20920 & ~w20921;
assign w20923 = w16977 & w16993;
assign w20924 = ~w16928 & w20923;
assign w20925 = pi02480 & ~w20924;
assign w20926 = ~pi09812 & w20924;
assign w20927 = ~w20925 & ~w20926;
assign w20928 = ~w16905 & w17334;
assign w20929 = pi02481 & ~w20928;
assign w20930 = ~pi02716 & w20928;
assign w20931 = ~w20929 & ~w20930;
assign w20932 = ~w16928 & w17754;
assign w20933 = pi02482 & ~w20932;
assign w20934 = ~pi02704 & w20932;
assign w20935 = ~w20933 & ~w20934;
assign w20936 = pi02483 & ~w18514;
assign w20937 = ~pi09812 & w18514;
assign w20938 = ~w20936 & ~w20937;
assign w20939 = ~w16905 & w18617;
assign w20940 = pi02484 & ~w20939;
assign w20941 = ~pi02713 & w20939;
assign w20942 = ~w20940 & ~w20941;
assign w20943 = pi02485 & ~w16932;
assign w20944 = ~pi02720 & w16932;
assign w20945 = ~w20943 & ~w20944;
assign w20946 = ~w16905 & w18949;
assign w20947 = pi02486 & ~w20946;
assign w20948 = w18059 & w18949;
assign w20949 = ~w20947 & ~w20948;
assign w20950 = pi02487 & ~w20799;
assign w20951 = w17193 & w18622;
assign w20952 = ~w20950 & ~w20951;
assign w20953 = ~w16992 & w18001;
assign w20954 = pi02488 & ~w20953;
assign w20955 = w17586 & w18001;
assign w20956 = ~w20954 & ~w20955;
assign w20957 = pi02489 & ~w20787;
assign w20958 = w17020 & w17172;
assign w20959 = ~w20957 & ~w20958;
assign w20960 = pi02490 & ~w20370;
assign w20961 = w17193 & w18617;
assign w20962 = ~w20960 & ~w20961;
assign w20963 = pi02491 & ~w20939;
assign w20964 = ~pi02716 & w20939;
assign w20965 = ~w20963 & ~w20964;
assign w20966 = ~w16992 & w18291;
assign w20967 = pi02492 & ~w20966;
assign w20968 = ~pi02722 & w20966;
assign w20969 = ~w20967 & ~w20968;
assign w20970 = ~w16928 & w20720;
assign w20971 = pi02493 & ~w20970;
assign w20972 = ~pi09812 & w20970;
assign w20973 = ~w20971 & ~w20972;
assign w20974 = ~w16928 & w19596;
assign w20975 = pi02494 & ~w20974;
assign w20976 = w18861 & w19596;
assign w20977 = ~w20975 & ~w20976;
assign w20978 = pi02495 & ~w20928;
assign w20979 = ~pi02170 & w20928;
assign w20980 = ~w20978 & ~w20979;
assign w20981 = ~w16905 & w18631;
assign w20982 = pi02496 & ~w20981;
assign w20983 = ~pi02716 & w20981;
assign w20984 = ~w20982 & ~w20983;
assign w20985 = pi02497 & ~w20895;
assign w20986 = w18059 & w18745;
assign w20987 = ~w20985 & ~w20986;
assign w20988 = ~w16928 & w17855;
assign w20989 = pi02498 & ~w20988;
assign w20990 = w17186 & w17855;
assign w20991 = ~w20989 & ~w20990;
assign w20992 = ~w16905 & w18662;
assign w20993 = pi02499 & ~w20992;
assign w20994 = ~pi02170 & w20992;
assign w20995 = ~w20993 & ~w20994;
assign w20996 = ~w16928 & w17609;
assign w20997 = pi02500 & ~w20996;
assign w20998 = ~pi09812 & w20996;
assign w20999 = ~w20997 & ~w20998;
assign w21000 = ~w16928 & w19655;
assign w21001 = pi02501 & ~w21000;
assign w21002 = ~pi02720 & w21000;
assign w21003 = ~w21001 & ~w21002;
assign w21004 = ~w16928 & w17650;
assign w21005 = pi02502 & ~w21004;
assign w21006 = ~pi09812 & w21004;
assign w21007 = ~w21005 & ~w21006;
assign w21008 = pi02503 & ~w20992;
assign w21009 = ~pi02711 & w20992;
assign w21010 = ~w21008 & ~w21009;
assign w21011 = ~w16892 & w17264;
assign w21012 = pi02504 & ~w21011;
assign w21013 = w17264 & w17925;
assign w21014 = ~w21012 & ~w21013;
assign w21015 = pi02505 & ~w20891;
assign w21016 = ~pi02712 & w20891;
assign w21017 = ~w21015 & ~w21016;
assign w21018 = ~w16892 & w18116;
assign w21019 = pi02506 & ~w21018;
assign w21020 = ~pi02707 & w21018;
assign w21021 = ~w21019 & ~w21020;
assign w21022 = ~w16905 & w17200;
assign w21023 = pi02507 & ~w21022;
assign w21024 = ~pi02713 & w21022;
assign w21025 = ~w21023 & ~w21024;
assign w21026 = ~w16992 & w19818;
assign w21027 = pi02508 & ~w21026;
assign w21028 = ~pi02721 & w21026;
assign w21029 = ~w21027 & ~w21028;
assign w21030 = ~w16892 & w17754;
assign w21031 = pi02509 & ~w21030;
assign w21032 = ~pi02707 & w21030;
assign w21033 = ~w21031 & ~w21032;
assign w21034 = pi02510 & ~w20875;
assign w21035 = ~pi02720 & w20875;
assign w21036 = ~w21034 & ~w21035;
assign w21037 = ~w16905 & w20720;
assign w21038 = pi02511 & ~w21037;
assign w21039 = ~pi02713 & w21037;
assign w21040 = ~w21038 & ~w21039;
assign w21041 = ~w16992 & w18813;
assign w21042 = pi02512 & ~w21041;
assign w21043 = ~pi02719 & w21041;
assign w21044 = ~w21042 & ~w21043;
assign w21045 = ~w16892 & w17200;
assign w21046 = pi02513 & ~w21045;
assign w21047 = ~pi02705 & w21045;
assign w21048 = ~w21046 & ~w21047;
assign w21049 = pi02514 & ~w20946;
assign w21050 = ~pi02170 & w20946;
assign w21051 = ~w21049 & ~w21050;
assign w21052 = ~w16905 & w16999;
assign w21053 = pi02515 & ~w21052;
assign w21054 = ~pi02715 & w21052;
assign w21055 = ~w21053 & ~w21054;
assign w21056 = ~w16892 & w17254;
assign w21057 = pi02516 & ~w21056;
assign w21058 = ~pi02706 & w21056;
assign w21059 = ~w21057 & ~w21058;
assign w21060 = ~w16892 & w17996;
assign w21061 = pi02517 & ~w21060;
assign w21062 = ~pi02709 & w21060;
assign w21063 = ~w21061 & ~w21062;
assign w21064 = pi02518 & ~w20425;
assign w21065 = ~pi02719 & w20425;
assign w21066 = ~w21064 & ~w21065;
assign w21067 = pi02519 & ~w20953;
assign w21068 = ~pi02703 & w20953;
assign w21069 = ~w21067 & ~w21068;
assign w21070 = ~w16992 & w18585;
assign w21071 = pi02520 & ~w21070;
assign w21072 = w17620 & w18585;
assign w21073 = ~w21071 & ~w21072;
assign w21074 = pi02521 & ~w21022;
assign w21075 = ~pi02712 & w21022;
assign w21076 = ~w21074 & ~w21075;
assign w21077 = pi02522 & ~w21056;
assign w21078 = w17254 & w18689;
assign w21079 = ~w21077 & ~w21078;
assign w21080 = ~w16905 & w17474;
assign w21081 = pi02523 & ~w21080;
assign w21082 = ~pi02717 & w21080;
assign w21083 = ~w21081 & ~w21082;
assign w21084 = ~w16905 & w19591;
assign w21085 = pi02524 & ~w21084;
assign w21086 = ~pi02712 & w21084;
assign w21087 = ~w21085 & ~w21086;
assign w21088 = ~w16905 & w18542;
assign w21089 = pi02525 & ~w21088;
assign w21090 = ~pi02713 & w21088;
assign w21091 = ~w21089 & ~w21090;
assign w21092 = pi02526 & ~w20906;
assign w21093 = ~pi02703 & w20906;
assign w21094 = ~w21092 & ~w21093;
assign w21095 = ~w16892 & w18146;
assign w21096 = pi02527 & ~w21095;
assign w21097 = ~pi02709 & w21095;
assign w21098 = ~w21096 & ~w21097;
assign w21099 = pi02528 & ~w21000;
assign w21100 = w17193 & w19655;
assign w21101 = ~w21099 & ~w21100;
assign w21102 = pi02529 & ~w21060;
assign w21103 = ~pi02707 & w21060;
assign w21104 = ~w21102 & ~w21103;
assign w21105 = ~w16905 & w17540;
assign w21106 = pi02530 & ~w21105;
assign w21107 = ~pi02716 & w21105;
assign w21108 = ~w21106 & ~w21107;
assign w21109 = pi02531 & ~w21037;
assign w21110 = ~pi02716 & w21037;
assign w21111 = ~w21109 & ~w21110;
assign w21112 = pi02532 & ~w21041;
assign w21113 = w18813 & w19797;
assign w21114 = ~w21112 & ~w21113;
assign w21115 = ~w16992 & w18526;
assign w21116 = pi02533 & ~w21115;
assign w21117 = w17594 & w18526;
assign w21118 = ~w21116 & ~w21117;
assign w21119 = pi02534 & ~w21041;
assign w21120 = ~pi02718 & w21041;
assign w21121 = ~w21119 & ~w21120;
assign w21122 = ~w16992 & w17556;
assign w21123 = pi02535 & ~w21122;
assign w21124 = ~pi02719 & w21122;
assign w21125 = ~w21123 & ~w21124;
assign w21126 = pi02536 & ~w20867;
assign w21127 = ~pi02718 & w20867;
assign w21128 = ~w21126 & ~w21127;
assign w21129 = pi02537 & ~w21115;
assign w21130 = ~pi02718 & w21115;
assign w21131 = ~w21129 & ~w21130;
assign w21132 = pi02538 & ~w20501;
assign w21133 = ~pi02716 & w20501;
assign w21134 = ~w21132 & ~w21133;
assign w21135 = ~w16892 & w17907;
assign w21136 = pi02539 & ~w21135;
assign w21137 = ~pi02708 & w21135;
assign w21138 = ~w21136 & ~w21137;
assign w21139 = pi02540 & ~w21095;
assign w21140 = ~pi02707 & w21095;
assign w21141 = ~w21139 & ~w21140;
assign w21142 = ~w16928 & w18032;
assign w21143 = pi02541 & ~w21142;
assign w21144 = ~pi02720 & w21142;
assign w21145 = ~w21143 & ~w21144;
assign w21146 = ~w16928 & w17694;
assign w21147 = pi02542 & ~w21146;
assign w21148 = ~pi02720 & w21146;
assign w21149 = ~w21147 & ~w21148;
assign w21150 = ~w16928 & w20566;
assign w21151 = pi02543 & ~w21150;
assign w21152 = ~pi02720 & w21150;
assign w21153 = ~w21151 & ~w21152;
assign w21154 = w16930 & w16938;
assign w21155 = ~w16928 & w21154;
assign w21156 = pi02544 & ~w21155;
assign w21157 = ~pi02720 & w21155;
assign w21158 = ~w21156 & ~w21157;
assign w21159 = pi02545 & ~w20879;
assign w21160 = ~pi02716 & w20879;
assign w21161 = ~w21159 & ~w21160;
assign w21162 = ~w16928 & w19629;
assign w21163 = pi02546 & ~w21162;
assign w21164 = ~pi09961 & w21162;
assign w21165 = ~w21163 & ~w21164;
assign w21166 = ~w16892 & w18027;
assign w21167 = pi02547 & ~w21166;
assign w21168 = ~pi02709 & w21166;
assign w21169 = ~w21167 & ~w21168;
assign w21170 = ~w16905 & w20244;
assign w21171 = pi02548 & ~w21170;
assign w21172 = ~pi02716 & w21170;
assign w21173 = ~w21171 & ~w21172;
assign w21174 = pi02549 & ~w20887;
assign w21175 = ~pi09812 & w20887;
assign w21176 = ~w21174 & ~w21175;
assign w21177 = ~w16928 & w17406;
assign w21178 = pi02550 & ~w21177;
assign w21179 = ~pi09812 & w21177;
assign w21180 = ~w21178 & ~w21179;
assign w21181 = ~w16928 & w20170;
assign w21182 = pi02551 & ~w21181;
assign w21183 = ~pi09812 & w21181;
assign w21184 = ~w21182 & ~w21183;
assign w21185 = ~w16928 & w18422;
assign w21186 = pi02552 & ~w21185;
assign w21187 = ~pi09848 & w21185;
assign w21188 = ~w21186 & ~w21187;
assign w21189 = pi02553 & ~w17227;
assign w21190 = ~pi09961 & w17227;
assign w21191 = ~w21189 & ~w21190;
assign w21192 = ~w16928 & w16961;
assign w21193 = pi02554 & ~w21192;
assign w21194 = w16961 & w17193;
assign w21195 = ~w21193 & ~w21194;
assign w21196 = pi02555 & ~w21155;
assign w21197 = ~pi09812 & w21155;
assign w21198 = ~w21196 & ~w21197;
assign w21199 = pi02556 & ~w21037;
assign w21200 = ~pi02711 & w21037;
assign w21201 = ~w21199 & ~w21200;
assign w21202 = ~w16928 & w17734;
assign w21203 = pi02557 & ~w21202;
assign w21204 = ~pi09954 & w21202;
assign w21205 = ~w21203 & ~w21204;
assign w21206 = pi02558 & ~w21142;
assign w21207 = ~pi09812 & w21142;
assign w21208 = ~w21206 & ~w21207;
assign w21209 = ~w16905 & w19459;
assign w21210 = pi02559 & ~w21209;
assign w21211 = ~pi02713 & w21209;
assign w21212 = ~w21210 & ~w21211;
assign w21213 = pi02560 & ~w17168;
assign w21214 = ~pi02720 & w17168;
assign w21215 = ~w21213 & ~w21214;
assign w21216 = ~w16928 & w17663;
assign w21217 = pi02561 & ~w21216;
assign w21218 = ~pi02720 & w21216;
assign w21219 = ~w21217 & ~w21218;
assign w21220 = ~w16992 & w20170;
assign w21221 = pi02562 & ~w21220;
assign w21222 = ~pi02164 & w21220;
assign w21223 = ~w21221 & ~w21222;
assign w21224 = ~w16928 & w17739;
assign w21225 = pi02563 & ~w21224;
assign w21226 = ~pi09812 & w21224;
assign w21227 = ~w21225 & ~w21226;
assign w21228 = ~w16928 & w17556;
assign w21229 = pi02564 & ~w21228;
assign w21230 = w17513 & w17556;
assign w21231 = ~w21229 & ~w21230;
assign w21232 = ~w16905 & w17279;
assign w21233 = pi02565 & ~w21232;
assign w21234 = ~pi02711 & w21232;
assign w21235 = ~w21233 & ~w21234;
assign w21236 = pi02566 & ~w18210;
assign w21237 = ~pi09848 & w18210;
assign w21238 = ~w21236 & ~w21237;
assign w21239 = ~w16928 & w20470;
assign w21240 = pi02567 & ~w21239;
assign w21241 = ~pi09812 & w21239;
assign w21242 = ~w21240 & ~w21241;
assign w21243 = pi02568 & ~w20621;
assign w21244 = ~pi09848 & w20621;
assign w21245 = ~w21243 & ~w21244;
assign w21246 = w16922 & ~w16928;
assign w21247 = pi02569 & ~w21246;
assign w21248 = ~pi02178 & w21246;
assign w21249 = ~w21247 & ~w21248;
assign w21250 = ~w16928 & w17686;
assign w21251 = pi02570 & ~w21250;
assign w21252 = w17193 & w17686;
assign w21253 = ~w21251 & ~w21252;
assign w21254 = ~w16928 & w18022;
assign w21255 = pi02571 & ~w21254;
assign w21256 = ~pi09812 & w21254;
assign w21257 = ~w21255 & ~w21256;
assign w21258 = ~w16928 & w20561;
assign w21259 = pi02572 & ~w21258;
assign w21260 = ~pi09954 & w21258;
assign w21261 = ~w21259 & ~w21260;
assign w21262 = ~w16928 & w18040;
assign w21263 = pi02573 & ~w21262;
assign w21264 = ~pi09812 & w21262;
assign w21265 = ~w21263 & ~w21264;
assign w21266 = ~w16928 & w17006;
assign w21267 = pi02574 & ~w21266;
assign w21268 = ~pi02178 & w21266;
assign w21269 = ~w21267 & ~w21268;
assign w21270 = ~w16928 & w17053;
assign w21271 = pi02575 & ~w21270;
assign w21272 = w17053 & w17439;
assign w21273 = ~w21271 & ~w21272;
assign w21274 = pi02576 & ~w21270;
assign w21275 = ~pi09812 & w21270;
assign w21276 = ~w21274 & ~w21275;
assign w21277 = ~w16905 & w18781;
assign w21278 = pi02577 & ~w21277;
assign w21279 = ~pi02717 & w21277;
assign w21280 = ~w21278 & ~w21279;
assign w21281 = ~w16892 & w17314;
assign w21282 = pi02578 & ~w21281;
assign w21283 = ~pi02707 & w21281;
assign w21284 = ~w21282 & ~w21283;
assign w21285 = ~w16905 & w18813;
assign w21286 = pi02579 & ~w21285;
assign w21287 = ~pi02713 & w21285;
assign w21288 = ~w21286 & ~w21287;
assign w21289 = ~w16905 & w18422;
assign w21290 = pi02580 & ~w21289;
assign w21291 = ~pi02711 & w21289;
assign w21292 = ~w21290 & ~w21291;
assign w21293 = ~w16992 & w18731;
assign w21294 = pi02581 & ~w21293;
assign w21295 = ~pi02167 & w21293;
assign w21296 = ~w21294 & ~w21295;
assign w21297 = pi02582 & ~w21224;
assign w21298 = ~pi02720 & w21224;
assign w21299 = ~w21297 & ~w21298;
assign w21300 = pi02583 & ~w21258;
assign w21301 = ~pi09812 & w21258;
assign w21302 = ~w21300 & ~w21301;
assign w21303 = ~w16928 & w18300;
assign w21304 = pi02584 & ~w21303;
assign w21305 = ~pi09812 & w21303;
assign w21306 = ~w21304 & ~w21305;
assign w21307 = ~w16928 & w17658;
assign w21308 = pi02585 & ~w21307;
assign w21309 = ~pi09812 & w21307;
assign w21310 = ~w21308 & ~w21309;
assign w21311 = ~w16928 & w17398;
assign w21312 = pi02586 & ~w21311;
assign w21313 = ~pi02720 & w21311;
assign w21314 = ~w21312 & ~w21313;
assign w21315 = pi02587 & ~w21303;
assign w21316 = ~pi02720 & w21303;
assign w21317 = ~w21315 & ~w21316;
assign w21318 = ~w16905 & w17609;
assign w21319 = pi02588 & ~w21318;
assign w21320 = w17317 & w17609;
assign w21321 = ~w21319 & ~w21320;
assign w21322 = ~w16928 & w17907;
assign w21323 = pi02589 & ~w21322;
assign w21324 = w17193 & w17907;
assign w21325 = ~w21323 & ~w21324;
assign w21326 = ~w16928 & w17681;
assign w21327 = pi02590 & ~w21326;
assign w21328 = ~pi09812 & w21326;
assign w21329 = ~w21327 & ~w21328;
assign w21330 = ~w16992 & w17500;
assign w21331 = pi02591 & ~w21330;
assign w21332 = ~pi02719 & w21330;
assign w21333 = ~w21331 & ~w21332;
assign w21334 = pi02592 & ~w20902;
assign w21335 = ~pi09812 & w20902;
assign w21336 = ~w21334 & ~w21335;
assign w21337 = ~w16928 & w17583;
assign w21338 = pi02593 & ~w21337;
assign w21339 = ~pi09812 & w21337;
assign w21340 = ~w21338 & ~w21339;
assign w21341 = ~w16928 & w17917;
assign w21342 = pi02594 & ~w21341;
assign w21343 = ~pi02720 & w21341;
assign w21344 = ~w21342 & ~w21343;
assign w21345 = ~w16992 & w16999;
assign w21346 = pi02595 & ~w21345;
assign w21347 = w16999 & w17594;
assign w21348 = ~w21346 & ~w21347;
assign w21349 = pi02596 & ~w21146;
assign w21350 = ~pi09812 & w21146;
assign w21351 = ~w21349 & ~w21350;
assign w21352 = ~w16928 & w17749;
assign w21353 = pi02597 & ~w21352;
assign w21354 = ~pi02720 & w21352;
assign w21355 = ~w21353 & ~w21354;
assign w21356 = ~w16928 & w17573;
assign w21357 = pi02598 & ~w21356;
assign w21358 = ~pi02704 & w21356;
assign w21359 = ~w21357 & ~w21358;
assign w21360 = ~w16992 & w18370;
assign w21361 = pi02599 & ~w21360;
assign w21362 = ~pi02719 & w21360;
assign w21363 = ~w21361 & ~w21362;
assign w21364 = pi02600 & ~w21352;
assign w21365 = ~pi09812 & w21352;
assign w21366 = ~w21364 & ~w21365;
assign w21367 = ~w16928 & w17775;
assign w21368 = pi02601 & ~w21367;
assign w21369 = ~pi09962 & w21367;
assign w21370 = ~w21368 & ~w21369;
assign w21371 = pi02602 & ~w21345;
assign w21372 = ~pi02718 & w21345;
assign w21373 = ~w21371 & ~w21372;
assign w21374 = ~w16928 & w17641;
assign w21375 = pi02603 & ~w21374;
assign w21376 = ~pi09812 & w21374;
assign w21377 = ~w21375 & ~w21376;
assign w21378 = ~w16928 & w17668;
assign w21379 = pi02604 & ~w21378;
assign w21380 = ~pi09812 & w21378;
assign w21381 = ~w21379 & ~w21380;
assign w21382 = pi02605 & ~w17196;
assign w21383 = w17047 & w17594;
assign w21384 = ~w21382 & ~w21383;
assign w21385 = ~w16928 & w17822;
assign w21386 = pi02606 & ~w21385;
assign w21387 = ~pi02720 & w21385;
assign w21388 = ~w21386 & ~w21387;
assign w21389 = pi02607 & ~w21341;
assign w21390 = ~pi09812 & w21341;
assign w21391 = ~w21389 & ~w21390;
assign w21392 = ~w16928 & w17922;
assign w21393 = pi02608 & ~w21392;
assign w21394 = w17193 & w17922;
assign w21395 = ~w21393 & ~w21394;
assign w21396 = pi02609 & ~w21392;
assign w21397 = ~pi02720 & w21392;
assign w21398 = ~w21396 & ~w21397;
assign w21399 = ~w16928 & w17614;
assign w21400 = pi02610 & ~w21399;
assign w21401 = ~pi02720 & w21399;
assign w21402 = ~w21400 & ~w21401;
assign w21403 = ~w16928 & w17526;
assign w21404 = pi02611 & ~w21403;
assign w21405 = ~pi09812 & w21403;
assign w21406 = ~w21404 & ~w21405;
assign w21407 = ~w16905 & w19379;
assign w21408 = pi02612 & ~w21407;
assign w21409 = ~pi02714 & w21407;
assign w21410 = ~w21408 & ~w21409;
assign w21411 = ~w16892 & w17977;
assign w21412 = pi02613 & ~w21411;
assign w21413 = ~pi02709 & w21411;
assign w21414 = ~w21412 & ~w21413;
assign w21415 = pi02614 & ~w21135;
assign w21416 = ~pi02707 & w21135;
assign w21417 = ~w21415 & ~w21416;
assign w21418 = ~w16905 & w19444;
assign w21419 = pi02615 & ~w21418;
assign w21420 = ~pi02712 & w21418;
assign w21421 = ~w21419 & ~w21420;
assign w21422 = pi02616 & ~w21418;
assign w21423 = w17317 & w19444;
assign w21424 = ~w21422 & ~w21423;
assign w21425 = ~w16992 & w19826;
assign w21426 = pi02617 & ~w21425;
assign w21427 = ~pi02721 & w21425;
assign w21428 = ~w21426 & ~w21427;
assign w21429 = pi02618 & ~w21385;
assign w21430 = ~pi09961 & w21385;
assign w21431 = ~w21429 & ~w21430;
assign w21432 = ~w16928 & w16986;
assign w21433 = pi02619 & ~w21432;
assign w21434 = w16986 & w17193;
assign w21435 = ~w21433 & ~w21434;
assign w21436 = ~w16905 & w19420;
assign w21437 = pi02620 & ~w21436;
assign w21438 = ~pi02712 & w21436;
assign w21439 = ~w21437 & ~w21438;
assign w21440 = pi02621 & ~w21150;
assign w21441 = w17193 & w20566;
assign w21442 = ~w21440 & ~w21441;
assign w21443 = ~w16992 & w18422;
assign w21444 = pi02622 & ~w21443;
assign w21445 = w17594 & w18422;
assign w21446 = ~w21444 & ~w21445;
assign w21447 = pi02623 & ~w21399;
assign w21448 = ~pi09812 & w21399;
assign w21449 = ~w21447 & ~w21448;
assign w21450 = pi02624 & ~w21209;
assign w21451 = ~pi02716 & w21209;
assign w21452 = ~w21450 & ~w21451;
assign w21453 = pi02625 & ~w16987;
assign w21454 = ~pi02717 & w16987;
assign w21455 = ~w21453 & ~w21454;
assign w21456 = ~w16905 & w17325;
assign w21457 = pi02626 & ~w21456;
assign w21458 = ~pi02717 & w21456;
assign w21459 = ~w21457 & ~w21458;
assign w21460 = ~w16992 & w18683;
assign w21461 = pi02627 & ~w21460;
assign w21462 = ~pi02719 & w21460;
assign w21463 = ~w21461 & ~w21462;
assign w21464 = pi02628 & ~w21460;
assign w21465 = ~pi02167 & w21460;
assign w21466 = ~w21464 & ~w21465;
assign w21467 = ~w16905 & w17917;
assign w21468 = pi02629 & ~w21467;
assign w21469 = ~pi02716 & w21467;
assign w21470 = ~w21468 & ~w21469;
assign w21471 = pi02630 & ~w21293;
assign w21472 = ~pi02719 & w21293;
assign w21473 = ~w21471 & ~w21472;
assign w21474 = pi02631 & ~w17269;
assign w21475 = ~pi02713 & w17269;
assign w21476 = ~w21474 & ~w21475;
assign w21477 = ~w16892 & w17300;
assign w21478 = pi02632 & ~w21477;
assign w21479 = ~pi02706 & w21477;
assign w21480 = ~w21478 & ~w21479;
assign w21481 = pi02633 & ~w21443;
assign w21482 = ~pi02169 & w21443;
assign w21483 = ~w21481 & ~w21482;
assign w21484 = ~w16992 & w17039;
assign w21485 = pi02634 & ~w21484;
assign w21486 = ~pi02703 & w21484;
assign w21487 = ~w21485 & ~w21486;
assign w21488 = ~w16928 & w17814;
assign w21489 = pi02635 & ~w21488;
assign w21490 = ~pi09954 & w21488;
assign w21491 = ~w21489 & ~w21490;
assign w21492 = ~w16892 & w17510;
assign w21493 = pi02636 & ~w21492;
assign w21494 = ~pi02710 & w21492;
assign w21495 = ~w21493 & ~w21494;
assign w21496 = ~w16992 & w18772;
assign w21497 = pi02637 & ~w21496;
assign w21498 = w17586 & w18772;
assign w21499 = ~w21497 & ~w21498;
assign w21500 = ~w16892 & w17361;
assign w21501 = pi02638 & ~w21500;
assign w21502 = ~pi02710 & w21500;
assign w21503 = ~w21501 & ~w21502;
assign w21504 = pi02639 & ~w21293;
assign w21505 = ~pi02169 & w21293;
assign w21506 = ~w21504 & ~w21505;
assign w21507 = pi02640 & ~w21052;
assign w21508 = ~pi02712 & w21052;
assign w21509 = ~w21507 & ~w21508;
assign w21510 = ~w16905 & w18370;
assign w21511 = pi02641 & ~w21510;
assign w21512 = ~pi02713 & w21510;
assign w21513 = ~w21511 & ~w21512;
assign w21514 = pi02642 & ~w21496;
assign w21515 = ~pi02167 & w21496;
assign w21516 = ~w21514 & ~w21515;
assign w21517 = ~w16992 & w18554;
assign w21518 = pi02643 & ~w21517;
assign w21519 = ~pi02167 & w21517;
assign w21520 = ~w21518 & ~w21519;
assign w21521 = pi02644 & ~w21407;
assign w21522 = ~pi02170 & w21407;
assign w21523 = ~w21521 & ~w21522;
assign w21524 = pi02645 & ~w21517;
assign w21525 = ~pi02703 & w21517;
assign w21526 = ~w21524 & ~w21525;
assign w21527 = ~w16992 & w20566;
assign w21528 = pi02646 & ~w21527;
assign w21529 = ~pi02169 & w21527;
assign w21530 = ~w21528 & ~w21529;
assign w21531 = pi02647 & ~w17340;
assign w21532 = ~pi02706 & w17340;
assign w21533 = ~w21531 & ~w21532;
assign w21534 = pi02648 & ~w11335;
assign w21535 = ~w11336 & ~w21534;
assign w21536 = pi09805 & ~w14192;
assign w21537 = ~w14193 & ~w21536;
assign w21538 = w11341 & w21537;
assign w21539 = ~w21535 & ~w21538;
assign w21540 = ~w16905 & w17938;
assign w21541 = pi02649 & ~w21540;
assign w21542 = ~pi02170 & w21540;
assign w21543 = ~w21541 & ~w21542;
assign w21544 = ~w16992 & w18563;
assign w21545 = pi02650 & ~w21544;
assign w21546 = ~pi02719 & w21544;
assign w21547 = ~w21545 & ~w21546;
assign w21548 = ~w16905 & w17505;
assign w21549 = pi02651 & ~w21548;
assign w21550 = ~pi02717 & w21548;
assign w21551 = ~w21549 & ~w21550;
assign w21552 = pi02652 & ~w21548;
assign w21553 = ~pi02714 & w21548;
assign w21554 = ~w21552 & ~w21553;
assign w21555 = ~w16992 & w17148;
assign w21556 = pi02653 & ~w21555;
assign w21557 = ~pi02719 & w21555;
assign w21558 = ~w21556 & ~w21557;
assign w21559 = ~w16992 & w17922;
assign w21560 = pi02654 & ~w21559;
assign w21561 = ~pi02169 & w21559;
assign w21562 = ~w21560 & ~w21561;
assign w21563 = ~w16905 & w21154;
assign w21564 = pi02655 & ~w21563;
assign w21565 = ~pi02711 & w21563;
assign w21566 = ~w21564 & ~w21565;
assign w21567 = pi09964 & ~w668;
assign w21568 = ~w502 & ~w21567;
assign w21569 = pi09969 & ~w21568;
assign w21570 = pi09822 & w21569;
assign w21571 = pi02656 & w21570;
assign w21572 = ~pi02656 & ~w21570;
assign w21573 = pi02666 & pi09964;
assign w21574 = w668 & w21573;
assign w21575 = ~pi00037 & ~w21574;
assign w21576 = w507 & w21575;
assign w21577 = ~w21571 & ~w21572;
assign w21578 = w21576 & w21577;
assign w21579 = pi02657 & ~w14136;
assign w21580 = pi01310 & w14136;
assign w21581 = ~w21579 & ~w21580;
assign w21582 = pi02658 & ~w14136;
assign w21583 = pi02657 & w14136;
assign w21584 = ~w21582 & ~w21583;
assign w21585 = pi02659 & ~w14136;
assign w21586 = pi02663 & w14136;
assign w21587 = ~w21585 & ~w21586;
assign w21588 = pi02660 & ~w14136;
assign w21589 = pi10453 & w14136;
assign w21590 = ~w21588 & ~w21589;
assign w21591 = pi02661 & ~w14136;
assign w21592 = ~pi01211 & w14136;
assign w21593 = ~w21591 & ~w21592;
assign w21594 = pi02662 & ~w14136;
assign w21595 = pi02341 & w14136;
assign w21596 = ~w21594 & ~w21595;
assign w21597 = pi02663 & ~w14136;
assign w21598 = pi10001 & w14136;
assign w21599 = ~w21597 & ~w21598;
assign w21600 = ~w16992 & w17658;
assign w21601 = pi02664 & ~w21600;
assign w21602 = ~pi02703 & w21600;
assign w21603 = ~w21601 & ~w21602;
assign w21604 = w321 & ~w386;
assign w21605 = ~w14215 & ~w21604;
assign w21606 = ~pi02666 & ~w21571;
assign w21607 = pi02666 & w21571;
assign w21608 = w21576 & ~w21606;
assign w21609 = ~w21607 & w21608;
assign w21610 = ~w16905 & w19601;
assign w21611 = pi02667 & ~w21610;
assign w21612 = ~pi02715 & w21610;
assign w21613 = ~w21611 & ~w21612;
assign w21614 = pi10632 & ~w16408;
assign w21615 = ~pi02668 & w16408;
assign w21616 = ~w21614 & ~w21615;
assign w21617 = pi10634 & ~w16408;
assign w21618 = ~pi02669 & w16408;
assign w21619 = ~w21617 & ~w21618;
assign w21620 = pi10622 & ~w16408;
assign w21621 = ~pi02670 & w16408;
assign w21622 = ~w21620 & ~w21621;
assign w21623 = pi10637 & ~w16408;
assign w21624 = ~pi02671 & w16408;
assign w21625 = ~w21623 & ~w21624;
assign w21626 = pi10623 & ~w16408;
assign w21627 = ~pi02672 & w16408;
assign w21628 = ~w21626 & ~w21627;
assign w21629 = pi10641 & ~w16408;
assign w21630 = ~pi02673 & w16408;
assign w21631 = ~w21629 & ~w21630;
assign w21632 = pi10645 & ~w16408;
assign w21633 = ~pi02674 & w16408;
assign w21634 = ~w21632 & ~w21633;
assign w21635 = pi10647 & ~w16408;
assign w21636 = ~pi02675 & w16408;
assign w21637 = ~w21635 & ~w21636;
assign w21638 = pi10650 & ~w16408;
assign w21639 = ~pi02676 & w16408;
assign w21640 = ~w21638 & ~w21639;
assign w21641 = pi10624 & ~w16408;
assign w21642 = ~pi02677 & w16408;
assign w21643 = ~w21641 & ~w21642;
assign w21644 = pi10652 & ~w16408;
assign w21645 = ~pi02678 & w16408;
assign w21646 = ~w21644 & ~w21645;
assign w21647 = pi10627 & ~w16408;
assign w21648 = ~pi02679 & w16408;
assign w21649 = ~w21647 & ~w21648;
assign w21650 = pi10626 & ~w16408;
assign w21651 = ~pi02680 & w16408;
assign w21652 = ~w21650 & ~w21651;
assign w21653 = pi10631 & ~w16408;
assign w21654 = ~pi02681 & w16408;
assign w21655 = ~w21653 & ~w21654;
assign w21656 = pi10630 & ~w16408;
assign w21657 = ~pi02682 & w16408;
assign w21658 = ~w21656 & ~w21657;
assign w21659 = pi02683 & ~w16214;
assign w21660 = ~pi10642 & w16214;
assign w21661 = ~w21659 & ~w21660;
assign w21662 = pi02684 & ~w16214;
assign w21663 = ~pi10649 & w16214;
assign w21664 = ~w21662 & ~w21663;
assign w21665 = pi02685 & ~w16251;
assign w21666 = ~pi10636 & w16251;
assign w21667 = ~w21665 & ~w21666;
assign w21668 = pi02686 & ~w16251;
assign w21669 = ~pi10649 & w16251;
assign w21670 = ~w21668 & ~w21669;
assign w21671 = pi02687 & ~w16251;
assign w21672 = ~pi10628 & w16251;
assign w21673 = ~w21671 & ~w21672;
assign w21674 = pi02688 & ~w16251;
assign w21675 = ~pi10626 & w16251;
assign w21676 = ~w21674 & ~w21675;
assign w21677 = pi02689 & ~w16244;
assign w21678 = ~pi10632 & w16244;
assign w21679 = ~w21677 & ~w21678;
assign w21680 = pi02690 & ~w16244;
assign w21681 = ~pi10649 & w16244;
assign w21682 = ~w21680 & ~w21681;
assign w21683 = pi02691 & ~w16229;
assign w21684 = ~pi10649 & w16229;
assign w21685 = ~w21683 & ~w21684;
assign w21686 = pi02692 & ~w16225;
assign w21687 = ~pi10626 & w16225;
assign w21688 = ~w21686 & ~w21687;
assign w21689 = ~w16992 & w17641;
assign w21690 = pi02693 & ~w21689;
assign w21691 = ~pi02721 & w21689;
assign w21692 = ~w21690 & ~w21691;
assign w21693 = pi02694 & ~w16219;
assign w21694 = ~pi10632 & w16219;
assign w21695 = ~w21693 & ~w21694;
assign w21696 = pi02695 & ~w16219;
assign w21697 = ~pi10628 & w16219;
assign w21698 = ~w21696 & ~w21697;
assign w21699 = pi10654 & w19704;
assign w21700 = pi02696 & w19713;
assign w21701 = pi10471 & w19712;
assign w21702 = pi10432 & w19710;
assign w21703 = ~w21699 & ~w21701;
assign w21704 = ~w21702 & w21703;
assign w21705 = ~w21700 & w21704;
assign w21706 = pi10655 & w19704;
assign w21707 = pi02697 & w19713;
assign w21708 = pi10364 & w19712;
assign w21709 = pi02796 & w19710;
assign w21710 = ~w21706 & ~w21708;
assign w21711 = ~w21709 & w21710;
assign w21712 = ~w21707 & w21711;
assign w21713 = pi10656 & w19704;
assign w21714 = pi02698 & w19713;
assign w21715 = pi10374 & w19712;
assign w21716 = pi09867 & w19710;
assign w21717 = ~w21713 & ~w21715;
assign w21718 = ~w21716 & w21717;
assign w21719 = ~w21714 & w21718;
assign w21720 = pi10657 & w19704;
assign w21721 = pi02699 & w19713;
assign w21722 = pi01304 & w19712;
assign w21723 = pi09802 & w19710;
assign w21724 = ~w21720 & ~w21722;
assign w21725 = ~w21723 & w21724;
assign w21726 = ~w21721 & w21725;
assign w21727 = pi10658 & w19704;
assign w21728 = pi02700 & w19713;
assign w21729 = pi01207 & w19712;
assign w21730 = pi01455 & w19710;
assign w21731 = ~w21727 & ~w21729;
assign w21732 = ~w21730 & w21731;
assign w21733 = ~w21728 & w21732;
assign w21734 = pi10659 & w19704;
assign w21735 = pi02701 & w19713;
assign w21736 = pi01311 & w19712;
assign w21737 = pi09866 & w19710;
assign w21738 = ~w21734 & ~w21736;
assign w21739 = ~w21737 & w21738;
assign w21740 = ~w21735 & w21739;
assign w21741 = pi10661 & w19704;
assign w21742 = pi02702 & w19713;
assign w21743 = pi00850 & w19712;
assign w21744 = ~pi01453 & w19710;
assign w21745 = ~w21741 & ~w21743;
assign w21746 = ~w21744 & w21745;
assign w21747 = ~w21742 & w21746;
assign w21748 = pi10590 & w19704;
assign w21749 = ~pi02703 & w19713;
assign w21750 = pi10482 & w19712;
assign w21751 = pi10050 & w19710;
assign w21752 = ~w21748 & ~w21750;
assign w21753 = ~w21751 & w21752;
assign w21754 = ~w21749 & w21753;
assign w21755 = pi10603 & w19704;
assign w21756 = ~pi02704 & w19713;
assign w21757 = ~pi00132 & w19712;
assign w21758 = ~pi00139 & w19710;
assign w21759 = ~w21755 & ~w21757;
assign w21760 = ~w21758 & w21759;
assign w21761 = ~w21756 & w21760;
assign w21762 = pi10606 & w19704;
assign w21763 = ~pi02705 & w19713;
assign w21764 = pi10422 & w19712;
assign w21765 = ~pi00280 & w19710;
assign w21766 = ~w21762 & ~w21764;
assign w21767 = ~w21765 & w21766;
assign w21768 = ~w21763 & w21767;
assign w21769 = pi10607 & w19704;
assign w21770 = ~pi02706 & w19713;
assign w21771 = pi10419 & w19712;
assign w21772 = ~pi00281 & w19710;
assign w21773 = ~w21769 & ~w21771;
assign w21774 = ~w21772 & w21773;
assign w21775 = ~w21770 & w21774;
assign w21776 = pi10608 & w19704;
assign w21777 = ~pi02707 & w19713;
assign w21778 = pi10409 & w19712;
assign w21779 = ~pi00257 & w19710;
assign w21780 = ~w21776 & ~w21778;
assign w21781 = ~w21779 & w21780;
assign w21782 = ~w21777 & w21781;
assign w21783 = pi10611 & w19704;
assign w21784 = ~pi02708 & w19713;
assign w21785 = ~pi02729 & w19712;
assign w21786 = ~pi00260 & w19710;
assign w21787 = ~w21783 & ~w21785;
assign w21788 = ~w21786 & w21787;
assign w21789 = ~w21784 & w21788;
assign w21790 = pi10612 & w19704;
assign w21791 = ~pi02709 & w19713;
assign w21792 = ~pi01212 & w19712;
assign w21793 = ~pi00259 & w19710;
assign w21794 = ~w21790 & ~w21792;
assign w21795 = ~w21793 & w21794;
assign w21796 = ~w21791 & w21795;
assign w21797 = pi10613 & w19704;
assign w21798 = ~pi02710 & w19713;
assign w21799 = ~pi02795 & w19712;
assign w21800 = ~pi00218 & w19710;
assign w21801 = ~w21797 & ~w21799;
assign w21802 = ~w21800 & w21801;
assign w21803 = ~w21798 & w21802;
assign w21804 = pi10614 & w19704;
assign w21805 = ~pi02711 & w19713;
assign w21806 = ~pi01479 & w19712;
assign w21807 = ~pi00196 & w19710;
assign w21808 = ~w21804 & ~w21806;
assign w21809 = ~w21807 & w21808;
assign w21810 = ~w21805 & w21809;
assign w21811 = pi10615 & w19704;
assign w21812 = ~pi02712 & w19713;
assign w21813 = ~pi01250 & w19712;
assign w21814 = ~pi00197 & w19710;
assign w21815 = ~w21811 & ~w21813;
assign w21816 = ~w21814 & w21815;
assign w21817 = ~w21812 & w21816;
assign w21818 = pi10617 & w19704;
assign w21819 = ~pi02713 & w19713;
assign w21820 = ~pi00873 & w19712;
assign w21821 = ~pi00194 & w19710;
assign w21822 = ~w21818 & ~w21820;
assign w21823 = ~w21821 & w21822;
assign w21824 = ~w21819 & w21823;
assign w21825 = pi10618 & w19704;
assign w21826 = ~pi02714 & w19713;
assign w21827 = ~pi02785 & w19712;
assign w21828 = ~pi00174 & w19710;
assign w21829 = ~w21825 & ~w21827;
assign w21830 = ~w21828 & w21829;
assign w21831 = ~w21826 & w21830;
assign w21832 = pi10619 & w19704;
assign w21833 = ~pi02715 & w19713;
assign w21834 = ~pi00866 & w19712;
assign w21835 = ~pi00215 & w19710;
assign w21836 = ~w21832 & ~w21834;
assign w21837 = ~w21835 & w21836;
assign w21838 = ~w21833 & w21837;
assign w21839 = pi10620 & w19704;
assign w21840 = ~pi02716 & w19713;
assign w21841 = ~pi01208 & w19712;
assign w21842 = ~pi00216 & w19710;
assign w21843 = ~w21839 & ~w21841;
assign w21844 = ~w21842 & w21843;
assign w21845 = ~w21840 & w21844;
assign w21846 = pi10621 & w19704;
assign w21847 = ~pi02717 & w19713;
assign w21848 = ~pi00871 & w19712;
assign w21849 = ~pi00195 & w19710;
assign w21850 = ~w21846 & ~w21848;
assign w21851 = ~w21849 & w21850;
assign w21852 = ~w21847 & w21851;
assign w21853 = pi10593 & w19704;
assign w21854 = ~pi02718 & w19713;
assign w21855 = pi10521 & w19712;
assign w21856 = pi00045 & w19710;
assign w21857 = ~w21853 & ~w21855;
assign w21858 = ~w21856 & w21857;
assign w21859 = ~w21854 & w21858;
assign w21860 = pi10597 & w19704;
assign w21861 = ~pi02719 & w19713;
assign w21862 = pi10541 & w19712;
assign w21863 = pi00050 & w19710;
assign w21864 = ~w21860 & ~w21862;
assign w21865 = ~w21863 & w21864;
assign w21866 = ~w21861 & w21865;
assign w21867 = pi10598 & w19704;
assign w21868 = ~pi02720 & w19713;
assign w21869 = pi10538 & w19712;
assign w21870 = pi10476 & w19710;
assign w21871 = ~w21867 & ~w21869;
assign w21872 = ~w21870 & w21871;
assign w21873 = ~w21868 & w21872;
assign w21874 = pi10591 & w19704;
assign w21875 = ~pi02721 & w19713;
assign w21876 = pi10522 & w19712;
assign w21877 = pi10265 & w19710;
assign w21878 = ~w21874 & ~w21876;
assign w21879 = ~w21877 & w21878;
assign w21880 = ~w21875 & w21879;
assign w21881 = pi10596 & w19704;
assign w21882 = ~pi02722 & w19713;
assign w21883 = pi10536 & w19712;
assign w21884 = pi00049 & w19710;
assign w21885 = ~w21881 & ~w21883;
assign w21886 = ~w21884 & w21885;
assign w21887 = ~w21882 & w21886;
assign w21888 = pi10610 & w19704;
assign w21889 = ~pi02723 & w19713;
assign w21890 = pi09999 & w19712;
assign w21891 = ~pi00217 & w19710;
assign w21892 = ~w21888 & ~w21890;
assign w21893 = ~w21891 & w21892;
assign w21894 = ~w21889 & w21893;
assign w21895 = ~pi09810 & ~pi09811;
assign w21896 = pi09854 & ~pi09857;
assign w21897 = ~pi09858 & w21896;
assign w21898 = w21895 & w21897;
assign w21899 = w14250 & w21898;
assign w21900 = pi02724 & ~w21899;
assign w21901 = ~pi00455 & w21899;
assign w21902 = ~w21900 & ~w21901;
assign w21903 = pi00485 & w14250;
assign w21904 = pi02725 & ~w14250;
assign w21905 = ~w21903 & ~w21904;
assign w21906 = ~pi10589 & w14250;
assign w21907 = pi02726 & ~w14250;
assign w21908 = ~w21906 & ~w21907;
assign w21909 = pi00456 & w14250;
assign w21910 = pi02727 & ~w14250;
assign w21911 = ~w21909 & ~w21910;
assign w21912 = pi00466 & w14250;
assign w21913 = pi02728 & ~w14250;
assign w21914 = ~w21912 & ~w21913;
assign w21915 = pi00869 & ~w1429;
assign w21916 = ~pi00869 & pi02729;
assign w21917 = ~w21915 & ~w21916;
assign w21918 = pi00467 & w14250;
assign w21919 = pi02730 & ~w14250;
assign w21920 = ~w21918 & ~w21919;
assign w21921 = ~w16892 & w17153;
assign w21922 = pi02731 & ~w21921;
assign w21923 = ~pi02708 & w21921;
assign w21924 = ~w21922 & ~w21923;
assign w21925 = ~w16892 & w18813;
assign w21926 = pi02732 & ~w21925;
assign w21927 = ~pi02706 & w21925;
assign w21928 = ~w21926 & ~w21927;
assign w21929 = ~w16992 & w17375;
assign w21930 = pi02733 & ~w21929;
assign w21931 = ~pi02719 & w21929;
assign w21932 = ~w21930 & ~w21931;
assign w21933 = ~w16892 & w18745;
assign w21934 = pi02734 & ~w21933;
assign w21935 = ~pi02709 & w21933;
assign w21936 = ~w21934 & ~w21935;
assign w21937 = ~w16892 & w17466;
assign w21938 = pi02735 & ~w21937;
assign w21939 = ~pi02706 & w21937;
assign w21940 = ~w21938 & ~w21939;
assign w21941 = pi02736 & ~w21411;
assign w21942 = ~pi02707 & w21411;
assign w21943 = ~w21941 & ~w21942;
assign w21944 = ~w16892 & w19379;
assign w21945 = pi02737 & ~w21944;
assign w21946 = ~pi02709 & w21944;
assign w21947 = ~w21945 & ~w21946;
assign w21948 = ~w16892 & w18449;
assign w21949 = pi02738 & ~w21948;
assign w21950 = ~pi02706 & w21948;
assign w21951 = ~w21949 & ~w21950;
assign w21952 = pi02739 & ~w21921;
assign w21953 = ~pi02706 & w21921;
assign w21954 = ~w21952 & ~w21953;
assign w21955 = pi02740 & ~w21944;
assign w21956 = ~pi02707 & w21944;
assign w21957 = ~w21955 & ~w21956;
assign w21958 = ~w16928 & w17361;
assign w21959 = pi02741 & ~w21958;
assign w21960 = ~pi02720 & w21958;
assign w21961 = ~w21959 & ~w21960;
assign w21962 = ~w16928 & w19343;
assign w21963 = pi02742 & ~w21962;
assign w21964 = w18861 & w19343;
assign w21965 = ~w21963 & ~w21964;
assign w21966 = pi02743 & ~w21925;
assign w21967 = ~pi02708 & w21925;
assign w21968 = ~w21966 & ~w21967;
assign w21969 = pi02744 & ~w21962;
assign w21970 = ~pi09961 & w21962;
assign w21971 = ~w21969 & ~w21970;
assign w21972 = ~w16892 & w17505;
assign w21973 = pi02745 & ~w21972;
assign w21974 = w17505 & w18689;
assign w21975 = ~w21973 & ~w21974;
assign w21976 = ~w16928 & w19348;
assign w21977 = pi02746 & ~w21976;
assign w21978 = w18861 & w19348;
assign w21979 = ~w21977 & ~w21978;
assign w21980 = pi02747 & ~w21972;
assign w21981 = ~pi02706 & w21972;
assign w21982 = ~w21980 & ~w21981;
assign w21983 = ~w16928 & w19374;
assign w21984 = pi02748 & ~w21983;
assign w21985 = ~pi02178 & w21983;
assign w21986 = ~w21984 & ~w21985;
assign w21987 = pi02749 & ~w21983;
assign w21988 = ~pi09961 & w21983;
assign w21989 = ~w21987 & ~w21988;
assign w21990 = ~w16892 & w18781;
assign w21991 = pi02750 & ~w21990;
assign w21992 = w17925 & w18781;
assign w21993 = ~w21991 & ~w21992;
assign w21994 = ~w16928 & w19012;
assign w21995 = pi02751 & ~w21994;
assign w21996 = ~pi02178 & w21994;
assign w21997 = ~w21995 & ~w21996;
assign w21998 = ~w16992 & w19838;
assign w21999 = pi02752 & ~w21998;
assign w22000 = ~pi02721 & w21998;
assign w22001 = ~w21999 & ~w22000;
assign w22002 = ~w16928 & w19591;
assign w22003 = pi02753 & ~w22002;
assign w22004 = ~pi09961 & w22002;
assign w22005 = ~w22003 & ~w22004;
assign w22006 = pi02754 & ~w22002;
assign w22007 = ~pi02178 & w22002;
assign w22008 = ~w22006 & ~w22007;
assign w22009 = ~w16905 & w19492;
assign w22010 = pi02755 & ~w22009;
assign w22011 = ~pi02713 & w22009;
assign w22012 = ~w22010 & ~w22011;
assign w22013 = ~w16905 & w19480;
assign w22014 = pi02756 & ~w22013;
assign w22015 = w18059 & w19480;
assign w22016 = ~w22014 & ~w22015;
assign w22017 = pi02757 & ~w22013;
assign w22018 = ~pi02712 & w22013;
assign w22019 = ~w22017 & ~w22018;
assign w22020 = ~w16905 & w19518;
assign w22021 = pi02758 & ~w22020;
assign w22022 = w17020 & w19518;
assign w22023 = ~w22021 & ~w22022;
assign w22024 = ~w16992 & w19852;
assign w22025 = pi02759 & ~w22024;
assign w22026 = ~pi02167 & w22024;
assign w22027 = ~w22025 & ~w22026;
assign w22028 = pi02760 & ~w22024;
assign w22029 = ~pi02721 & w22024;
assign w22030 = ~w22028 & ~w22029;
assign w22031 = ~w16905 & w19561;
assign w22032 = pi02761 & ~w22031;
assign w22033 = ~pi02712 & w22031;
assign w22034 = ~w22032 & ~w22033;
assign w22035 = ~w16905 & w19530;
assign w22036 = pi02762 & ~w22035;
assign w22037 = w18059 & w19530;
assign w22038 = ~w22036 & ~w22037;
assign w22039 = pi02763 & ~w22035;
assign w22040 = ~pi02712 & w22035;
assign w22041 = ~w22039 & ~w22040;
assign w22042 = ~w16905 & w19435;
assign w22043 = pi02764 & ~w22042;
assign w22044 = w17020 & w19435;
assign w22045 = ~w22043 & ~w22044;
assign w22046 = ~w16905 & w19552;
assign w22047 = pi02765 & ~w22046;
assign w22048 = ~pi02715 & w22046;
assign w22049 = ~w22047 & ~w22048;
assign w22050 = pi02766 & ~w22046;
assign w22051 = w17020 & w19552;
assign w22052 = ~w22050 & ~w22051;
assign w22053 = ~w16928 & w20465;
assign w22054 = pi02767 & ~w22053;
assign w22055 = ~pi09812 & w22053;
assign w22056 = ~w22054 & ~w22055;
assign w22057 = pi02768 & ~w21610;
assign w22058 = ~pi02712 & w21610;
assign w22059 = ~w22057 & ~w22058;
assign w22060 = ~w16905 & w19606;
assign w22061 = pi02769 & ~w22060;
assign w22062 = w17020 & w19606;
assign w22063 = ~w22061 & ~w22062;
assign w22064 = ~w16905 & w19624;
assign w22065 = pi02770 & ~w22064;
assign w22066 = ~pi02715 & w22064;
assign w22067 = ~w22065 & ~w22066;
assign w22068 = pi02771 & ~w22064;
assign w22069 = ~pi02712 & w22064;
assign w22070 = ~w22068 & ~w22069;
assign w22071 = ~w16905 & w19576;
assign w22072 = pi02772 & ~w22071;
assign w22073 = w18059 & w19576;
assign w22074 = ~w22072 & ~w22073;
assign w22075 = pi02773 & ~w22071;
assign w22076 = ~pi02712 & w22071;
assign w22077 = ~w22075 & ~w22076;
assign w22078 = ~w16905 & w19645;
assign w22079 = pi02774 & ~w22078;
assign w22080 = ~pi02715 & w22078;
assign w22081 = ~w22079 & ~w22080;
assign w22082 = pi02775 & ~w22078;
assign w22083 = ~pi02712 & w22078;
assign w22084 = ~w22082 & ~w22083;
assign w22085 = ~w16992 & w19909;
assign w22086 = pi02776 & ~w22085;
assign w22087 = ~pi02164 & w22085;
assign w22088 = ~w22086 & ~w22087;
assign w22089 = ~w16905 & w19650;
assign w22090 = pi02777 & ~w22089;
assign w22091 = ~pi02712 & w22089;
assign w22092 = ~w22090 & ~w22091;
assign w22093 = pi02778 & ~w22085;
assign w22094 = ~pi02721 & w22085;
assign w22095 = ~w22093 & ~w22094;
assign w22096 = ~w16992 & w19930;
assign w22097 = pi02779 & ~w22096;
assign w22098 = ~pi02721 & w22096;
assign w22099 = ~w22097 & ~w22098;
assign w22100 = ~w16905 & w19679;
assign w22101 = pi02780 & ~w22100;
assign w22102 = w18059 & w19679;
assign w22103 = ~w22101 & ~w22102;
assign w22104 = pi02781 & ~w22100;
assign w22105 = ~pi02712 & w22100;
assign w22106 = ~w22104 & ~w22105;
assign w22107 = ~w16905 & w19660;
assign w22108 = pi02782 & ~w22107;
assign w22109 = ~pi02712 & w22107;
assign w22110 = ~w22108 & ~w22109;
assign w22111 = ~w16905 & w19723;
assign w22112 = pi02783 & ~w22111;
assign w22113 = ~pi02715 & w22111;
assign w22114 = ~w22112 & ~w22113;
assign w22115 = pi02784 & ~w22111;
assign w22116 = ~pi02712 & w22111;
assign w22117 = ~w22115 & ~w22116;
assign w22118 = pi00869 & ~w1475;
assign w22119 = ~pi00869 & pi02785;
assign w22120 = ~w22118 & ~w22119;
assign w22121 = ~w16905 & w19728;
assign w22122 = pi02786 & ~w22121;
assign w22123 = w17020 & w19728;
assign w22124 = ~w22122 & ~w22123;
assign w22125 = pi02787 & ~w19267;
assign w22126 = pi10598 & w19267;
assign w22127 = ~w22125 & ~w22126;
assign w22128 = pi02788 & ~w19267;
assign w22129 = pi10599 & w19267;
assign w22130 = ~w22128 & ~w22129;
assign w22131 = pi02789 & ~w19267;
assign w22132 = pi10602 & w19267;
assign w22133 = ~w22131 & ~w22132;
assign w22134 = pi02790 & ~w19267;
assign w22135 = pi10603 & w19267;
assign w22136 = ~w22134 & ~w22135;
assign w22137 = pi02791 & ~w19267;
assign w22138 = pi10601 & w19267;
assign w22139 = ~w22137 & ~w22138;
assign w22140 = pi02792 & ~w19267;
assign w22141 = pi10605 & w19267;
assign w22142 = ~w22140 & ~w22141;
assign w22143 = pi02793 & ~w21318;
assign w22144 = w17609 & w20209;
assign w22145 = ~w22143 & ~w22144;
assign w22146 = w16931 & ~w16992;
assign w22147 = pi02794 & ~w22146;
assign w22148 = ~pi02722 & w22146;
assign w22149 = ~w22147 & ~w22148;
assign w22150 = pi00869 & ~w1421;
assign w22151 = ~pi00869 & pi02795;
assign w22152 = ~w22150 & ~w22151;
assign w22153 = ~pi02796 & w16786;
assign w22154 = ~w16785 & ~w22153;
assign w22155 = ~pi02796 & ~w16775;
assign w22156 = ~w22154 & ~w22155;
assign w22157 = w1217 & w11485;
assign w22158 = pi02797 & ~w22157;
assign w22159 = pi10590 & w22157;
assign w22160 = ~w22158 & ~w22159;
assign w22161 = pi02798 & ~w22157;
assign w22162 = pi10591 & w22157;
assign w22163 = ~w22161 & ~w22162;
assign w22164 = pi02799 & ~w22157;
assign w22165 = pi10592 & w22157;
assign w22166 = ~w22164 & ~w22165;
assign w22167 = pi02800 & ~w22157;
assign w22168 = pi10593 & w22157;
assign w22169 = ~w22167 & ~w22168;
assign w22170 = pi02801 & ~w22157;
assign w22171 = pi10594 & w22157;
assign w22172 = ~w22170 & ~w22171;
assign w22173 = pi02802 & ~w22157;
assign w22174 = pi10595 & w22157;
assign w22175 = ~w22173 & ~w22174;
assign w22176 = pi02803 & ~w22157;
assign w22177 = pi10596 & w22157;
assign w22178 = ~w22176 & ~w22177;
assign w22179 = pi02804 & ~w22157;
assign w22180 = pi10597 & w22157;
assign w22181 = ~w22179 & ~w22180;
assign w22182 = pi02805 & ~w21080;
assign w22183 = ~pi02713 & w21080;
assign w22184 = ~w22182 & ~w22183;
assign w22185 = ~w16928 & w17108;
assign w22186 = pi02806 & ~w22185;
assign w22187 = ~pi09812 & w22185;
assign w22188 = ~w22186 & ~w22187;
assign w22189 = ~w16892 & w18263;
assign w22190 = pi02807 & ~w22189;
assign w22191 = w18263 & w18364;
assign w22192 = ~w22190 & ~w22191;
assign w22193 = ~w16892 & w18155;
assign w22194 = pi02808 & ~w22193;
assign w22195 = ~pi02707 & w22193;
assign w22196 = ~w22194 & ~w22195;
assign w22197 = pi02809 & ~w22146;
assign w22198 = ~pi02721 & w22146;
assign w22199 = ~w22197 & ~w22198;
assign w22200 = ~pi02810 & ~w16879;
assign w22201 = ~w16881 & ~w22200;
assign w22202 = ~pi00300 & ~pi09871;
assign w22203 = w14260 & w22202;
assign w22204 = ~pi02812 & ~w14845;
assign w22205 = w16880 & ~w22204;
assign w22206 = pi02813 & ~w21962;
assign w22207 = ~pi09954 & w21962;
assign w22208 = ~w22206 & ~w22207;
assign w22209 = pi02814 & ~w21962;
assign w22210 = ~pi02720 & w21962;
assign w22211 = ~w22209 & ~w22210;
assign w22212 = pi02815 & ~w21962;
assign w22213 = ~pi09962 & w21962;
assign w22214 = ~w22212 & ~w22213;
assign w22215 = pi02816 & ~w17381;
assign w22216 = ~pi02705 & w17381;
assign w22217 = ~w22215 & ~w22216;
assign w22218 = pi02817 & ~w17381;
assign w22219 = ~pi02706 & w17381;
assign w22220 = ~w22218 & ~w22219;
assign w22221 = pi02818 & ~w17381;
assign w22222 = ~pi02707 & w17381;
assign w22223 = ~w22221 & ~w22222;
assign w22224 = pi02819 & ~w17381;
assign w22225 = ~pi02160 & w17381;
assign w22226 = ~w22224 & ~w22225;
assign w22227 = pi02820 & ~w17381;
assign w22228 = ~pi02708 & w17381;
assign w22229 = ~w22227 & ~w22228;
assign w22230 = pi02821 & ~w17381;
assign w22231 = ~pi02709 & w17381;
assign w22232 = ~w22230 & ~w22231;
assign w22233 = pi02822 & ~w17381;
assign w22234 = ~pi02710 & w17381;
assign w22235 = ~w22233 & ~w22234;
assign w22236 = pi02823 & ~w16900;
assign w22237 = ~pi02706 & w16900;
assign w22238 = ~w22236 & ~w22237;
assign w22239 = pi02824 & ~w16900;
assign w22240 = w16899 & w18067;
assign w22241 = ~w22239 & ~w22240;
assign w22242 = pi02825 & ~w16900;
assign w22243 = ~pi02160 & w16900;
assign w22244 = ~w22242 & ~w22243;
assign w22245 = pi02826 & ~w16900;
assign w22246 = ~pi02708 & w16900;
assign w22247 = ~w22245 & ~w22246;
assign w22248 = pi02827 & ~w16900;
assign w22249 = ~pi02709 & w16900;
assign w22250 = ~w22248 & ~w22249;
assign w22251 = pi02828 & ~w16900;
assign w22252 = ~pi02710 & w16900;
assign w22253 = ~w22251 & ~w22252;
assign w22254 = pi02829 & ~w17219;
assign w22255 = ~pi02705 & w17219;
assign w22256 = ~w22254 & ~w22255;
assign w22257 = pi02830 & ~w17219;
assign w22258 = ~pi02706 & w17219;
assign w22259 = ~w22257 & ~w22258;
assign w22260 = pi02831 & ~w17219;
assign w22261 = ~pi02707 & w17219;
assign w22262 = ~w22260 & ~w22261;
assign w22263 = pi02832 & ~w17219;
assign w22264 = ~pi02160 & w17219;
assign w22265 = ~w22263 & ~w22264;
assign w22266 = pi02833 & ~w17219;
assign w22267 = ~pi02708 & w17219;
assign w22268 = ~w22266 & ~w22267;
assign w22269 = pi02834 & ~w17219;
assign w22270 = ~pi02709 & w17219;
assign w22271 = ~w22269 & ~w22270;
assign w22272 = pi02835 & ~w17219;
assign w22273 = ~pi02710 & w17219;
assign w22274 = ~w22272 & ~w22273;
assign w22275 = pi02836 & ~w16949;
assign w22276 = ~pi02706 & w16949;
assign w22277 = ~w22275 & ~w22276;
assign w22278 = pi02837 & ~w16949;
assign w22279 = ~pi02707 & w16949;
assign w22280 = ~w22278 & ~w22279;
assign w22281 = pi02838 & ~w16949;
assign w22282 = w16948 & w18234;
assign w22283 = ~w22281 & ~w22282;
assign w22284 = pi02839 & ~w16949;
assign w22285 = ~pi02708 & w16949;
assign w22286 = ~w22284 & ~w22285;
assign w22287 = pi02840 & ~w16949;
assign w22288 = ~pi02709 & w16949;
assign w22289 = ~w22287 & ~w22288;
assign w22290 = pi02841 & ~w16949;
assign w22291 = w16948 & w18364;
assign w22292 = ~w22290 & ~w22291;
assign w22293 = pi02842 & ~w17132;
assign w22294 = ~pi02705 & w17132;
assign w22295 = ~w22293 & ~w22294;
assign w22296 = pi02843 & ~w17132;
assign w22297 = ~pi02706 & w17132;
assign w22298 = ~w22296 & ~w22297;
assign w22299 = pi02844 & ~w17132;
assign w22300 = ~pi02707 & w17132;
assign w22301 = ~w22299 & ~w22300;
assign w22302 = pi02845 & ~w17132;
assign w22303 = ~pi02160 & w17132;
assign w22304 = ~w22302 & ~w22303;
assign w22305 = pi02846 & ~w17132;
assign w22306 = w17131 & w18689;
assign w22307 = ~w22305 & ~w22306;
assign w22308 = pi02847 & ~w17132;
assign w22309 = ~pi02709 & w17132;
assign w22310 = ~w22308 & ~w22309;
assign w22311 = pi02848 & ~w17132;
assign w22312 = ~pi02710 & w17132;
assign w22313 = ~w22311 & ~w22312;
assign w22314 = pi02849 & ~w17061;
assign w22315 = ~pi02706 & w17061;
assign w22316 = ~w22314 & ~w22315;
assign w22317 = pi02850 & ~w17061;
assign w22318 = ~pi02707 & w17061;
assign w22319 = ~w22317 & ~w22318;
assign w22320 = pi02851 & ~w17061;
assign w22321 = ~pi02160 & w17061;
assign w22322 = ~w22320 & ~w22321;
assign w22323 = pi02852 & ~w17061;
assign w22324 = ~pi02708 & w17061;
assign w22325 = ~w22323 & ~w22324;
assign w22326 = pi02853 & ~w17061;
assign w22327 = ~pi02709 & w17061;
assign w22328 = ~w22326 & ~w22327;
assign w22329 = pi02854 & ~w17061;
assign w22330 = ~pi02710 & w17061;
assign w22331 = ~w22329 & ~w22330;
assign w22332 = ~w16892 & w19106;
assign w22333 = pi02855 & ~w22332;
assign w22334 = w18578 & w19106;
assign w22335 = ~w22333 & ~w22334;
assign w22336 = pi02856 & ~w22332;
assign w22337 = w17925 & w19106;
assign w22338 = ~w22336 & ~w22337;
assign w22339 = pi02857 & ~w22332;
assign w22340 = ~pi02707 & w22332;
assign w22341 = ~w22339 & ~w22340;
assign w22342 = pi02858 & ~w22332;
assign w22343 = w18234 & w19106;
assign w22344 = ~w22342 & ~w22343;
assign w22345 = pi02859 & ~w22332;
assign w22346 = ~pi02708 & w22332;
assign w22347 = ~w22345 & ~w22346;
assign w22348 = pi02860 & ~w22332;
assign w22349 = ~pi02709 & w22332;
assign w22350 = ~w22348 & ~w22349;
assign w22351 = pi02861 & ~w22332;
assign w22352 = w18364 & w19106;
assign w22353 = ~w22351 & ~w22352;
assign w22354 = ~w16892 & w19149;
assign w22355 = pi02862 & ~w22354;
assign w22356 = ~pi02706 & w22354;
assign w22357 = ~w22355 & ~w22356;
assign w22358 = pi02863 & ~w22354;
assign w22359 = w18067 & w19149;
assign w22360 = ~w22358 & ~w22359;
assign w22361 = pi02864 & ~w22354;
assign w22362 = w18234 & w19149;
assign w22363 = ~w22361 & ~w22362;
assign w22364 = pi02865 & ~w22354;
assign w22365 = ~pi02708 & w22354;
assign w22366 = ~w22364 & ~w22365;
assign w22367 = pi02866 & ~w22354;
assign w22368 = w18092 & w19149;
assign w22369 = ~w22367 & ~w22368;
assign w22370 = pi02867 & ~w22354;
assign w22371 = ~pi02710 & w22354;
assign w22372 = ~w22370 & ~w22371;
assign w22373 = ~w16892 & w19166;
assign w22374 = pi02868 & ~w22373;
assign w22375 = ~pi02705 & w22373;
assign w22376 = ~w22374 & ~w22375;
assign w22377 = pi02869 & ~w22373;
assign w22378 = ~pi02706 & w22373;
assign w22379 = ~w22377 & ~w22378;
assign w22380 = pi02870 & ~w22373;
assign w22381 = ~pi02707 & w22373;
assign w22382 = ~w22380 & ~w22381;
assign w22383 = pi02871 & ~w22373;
assign w22384 = ~pi02160 & w22373;
assign w22385 = ~w22383 & ~w22384;
assign w22386 = pi02872 & ~w22373;
assign w22387 = ~pi02708 & w22373;
assign w22388 = ~w22386 & ~w22387;
assign w22389 = pi02873 & ~w22373;
assign w22390 = ~pi02709 & w22373;
assign w22391 = ~w22389 & ~w22390;
assign w22392 = pi02874 & ~w22373;
assign w22393 = ~pi02710 & w22373;
assign w22394 = ~w22392 & ~w22393;
assign w22395 = ~w16892 & w19130;
assign w22396 = pi02875 & ~w22395;
assign w22397 = ~pi02706 & w22395;
assign w22398 = ~w22396 & ~w22397;
assign w22399 = pi02876 & ~w22395;
assign w22400 = ~pi02707 & w22395;
assign w22401 = ~w22399 & ~w22400;
assign w22402 = pi02877 & ~w22395;
assign w22403 = ~pi02160 & w22395;
assign w22404 = ~w22402 & ~w22403;
assign w22405 = pi02878 & ~w22395;
assign w22406 = ~pi02708 & w22395;
assign w22407 = ~w22405 & ~w22406;
assign w22408 = pi02879 & ~w22395;
assign w22409 = ~pi02709 & w22395;
assign w22410 = ~w22408 & ~w22409;
assign w22411 = pi02880 & ~w22395;
assign w22412 = ~pi02710 & w22395;
assign w22413 = ~w22411 & ~w22412;
assign w22414 = ~w16892 & w19115;
assign w22415 = pi02881 & ~w22414;
assign w22416 = ~pi02705 & w22414;
assign w22417 = ~w22415 & ~w22416;
assign w22418 = pi02882 & ~w22414;
assign w22419 = ~pi02706 & w22414;
assign w22420 = ~w22418 & ~w22419;
assign w22421 = pi02883 & ~w22414;
assign w22422 = ~pi02707 & w22414;
assign w22423 = ~w22421 & ~w22422;
assign w22424 = pi02884 & ~w22414;
assign w22425 = ~pi02160 & w22414;
assign w22426 = ~w22424 & ~w22425;
assign w22427 = pi02885 & ~w22414;
assign w22428 = ~pi02708 & w22414;
assign w22429 = ~w22427 & ~w22428;
assign w22430 = pi02886 & ~w22414;
assign w22431 = ~pi02709 & w22414;
assign w22432 = ~w22430 & ~w22431;
assign w22433 = pi02887 & ~w22414;
assign w22434 = ~pi02710 & w22414;
assign w22435 = ~w22433 & ~w22434;
assign w22436 = ~w16892 & w19087;
assign w22437 = pi02888 & ~w22436;
assign w22438 = ~pi02706 & w22436;
assign w22439 = ~w22437 & ~w22438;
assign w22440 = pi02889 & ~w22436;
assign w22441 = ~pi02707 & w22436;
assign w22442 = ~w22440 & ~w22441;
assign w22443 = pi02890 & ~w22436;
assign w22444 = ~pi02160 & w22436;
assign w22445 = ~w22443 & ~w22444;
assign w22446 = pi02891 & ~w22436;
assign w22447 = ~pi02708 & w22436;
assign w22448 = ~w22446 & ~w22447;
assign w22449 = pi02892 & ~w22436;
assign w22450 = ~pi02709 & w22436;
assign w22451 = ~w22449 & ~w22450;
assign w22452 = pi02893 & ~w22436;
assign w22453 = ~pi02710 & w22436;
assign w22454 = ~w22452 & ~w22453;
assign w22455 = ~w16892 & w19075;
assign w22456 = pi02894 & ~w22455;
assign w22457 = ~pi02705 & w22455;
assign w22458 = ~w22456 & ~w22457;
assign w22459 = pi02895 & ~w22455;
assign w22460 = ~pi02706 & w22455;
assign w22461 = ~w22459 & ~w22460;
assign w22462 = pi02896 & ~w22455;
assign w22463 = ~pi02707 & w22455;
assign w22464 = ~w22462 & ~w22463;
assign w22465 = pi02897 & ~w22455;
assign w22466 = w18234 & w19075;
assign w22467 = ~w22465 & ~w22466;
assign w22468 = pi02898 & ~w22455;
assign w22469 = w18689 & w19075;
assign w22470 = ~w22468 & ~w22469;
assign w22471 = pi02899 & ~w22455;
assign w22472 = ~pi02709 & w22455;
assign w22473 = ~w22471 & ~w22472;
assign w22474 = pi02900 & ~w22455;
assign w22475 = ~pi02710 & w22455;
assign w22476 = ~w22474 & ~w22475;
assign w22477 = ~w16892 & w18995;
assign w22478 = pi02901 & ~w22477;
assign w22479 = ~pi02706 & w22477;
assign w22480 = ~w22478 & ~w22479;
assign w22481 = pi02902 & ~w22477;
assign w22482 = ~pi02707 & w22477;
assign w22483 = ~w22481 & ~w22482;
assign w22484 = pi02903 & ~w22477;
assign w22485 = ~pi02160 & w22477;
assign w22486 = ~w22484 & ~w22485;
assign w22487 = pi02904 & ~w22477;
assign w22488 = ~pi02708 & w22477;
assign w22489 = ~w22487 & ~w22488;
assign w22490 = pi02905 & ~w22477;
assign w22491 = ~pi02709 & w22477;
assign w22492 = ~w22490 & ~w22491;
assign w22493 = pi02906 & ~w22477;
assign w22494 = w18364 & w18995;
assign w22495 = ~w22493 & ~w22494;
assign w22496 = ~w16892 & w19053;
assign w22497 = pi02907 & ~w22496;
assign w22498 = ~pi02705 & w22496;
assign w22499 = ~w22497 & ~w22498;
assign w22500 = pi02908 & ~w22496;
assign w22501 = w17925 & w19053;
assign w22502 = ~w22500 & ~w22501;
assign w22503 = pi02909 & ~w22496;
assign w22504 = ~pi02707 & w22496;
assign w22505 = ~w22503 & ~w22504;
assign w22506 = pi02910 & ~w22496;
assign w22507 = ~pi02160 & w22496;
assign w22508 = ~w22506 & ~w22507;
assign w22509 = pi02911 & ~w22496;
assign w22510 = ~pi02723 & w22496;
assign w22511 = ~w22509 & ~w22510;
assign w22512 = pi02912 & ~w22496;
assign w22513 = ~pi02708 & w22496;
assign w22514 = ~w22512 & ~w22513;
assign w22515 = pi02913 & ~w22496;
assign w22516 = ~pi02709 & w22496;
assign w22517 = ~w22515 & ~w22516;
assign w22518 = pi02914 & ~w22496;
assign w22519 = ~pi02710 & w22496;
assign w22520 = ~w22518 & ~w22519;
assign w22521 = ~w16892 & w19034;
assign w22522 = pi02915 & ~w22521;
assign w22523 = ~pi02706 & w22521;
assign w22524 = ~w22522 & ~w22523;
assign w22525 = pi02916 & ~w22521;
assign w22526 = ~pi02707 & w22521;
assign w22527 = ~w22525 & ~w22526;
assign w22528 = pi02917 & ~w22521;
assign w22529 = ~pi02160 & w22521;
assign w22530 = ~w22528 & ~w22529;
assign w22531 = pi02918 & ~w22521;
assign w22532 = ~pi02708 & w22521;
assign w22533 = ~w22531 & ~w22532;
assign w22534 = pi02919 & ~w22521;
assign w22535 = ~pi02709 & w22521;
assign w22536 = ~w22534 & ~w22535;
assign w22537 = pi02920 & ~w22521;
assign w22538 = ~pi02710 & w22521;
assign w22539 = ~w22537 & ~w22538;
assign w22540 = ~w16892 & w18986;
assign w22541 = pi02921 & ~w22540;
assign w22542 = ~pi02705 & w22540;
assign w22543 = ~w22541 & ~w22542;
assign w22544 = pi02922 & ~w22540;
assign w22545 = ~pi02706 & w22540;
assign w22546 = ~w22544 & ~w22545;
assign w22547 = pi02923 & ~w22540;
assign w22548 = ~pi02707 & w22540;
assign w22549 = ~w22547 & ~w22548;
assign w22550 = pi02924 & ~w22540;
assign w22551 = ~pi02160 & w22540;
assign w22552 = ~w22550 & ~w22551;
assign w22553 = pi02925 & ~w22540;
assign w22554 = ~pi02708 & w22540;
assign w22555 = ~w22553 & ~w22554;
assign w22556 = pi02926 & ~w22540;
assign w22557 = ~pi02709 & w22540;
assign w22558 = ~w22556 & ~w22557;
assign w22559 = pi02927 & ~w22540;
assign w22560 = ~pi02710 & w22540;
assign w22561 = ~w22559 & ~w22560;
assign w22562 = ~w16892 & w18925;
assign w22563 = pi02928 & ~w22562;
assign w22564 = w17925 & w18925;
assign w22565 = ~w22563 & ~w22564;
assign w22566 = pi02929 & ~w22562;
assign w22567 = ~pi02707 & w22562;
assign w22568 = ~w22566 & ~w22567;
assign w22569 = pi02930 & ~w22562;
assign w22570 = ~pi02160 & w22562;
assign w22571 = ~w22569 & ~w22570;
assign w22572 = pi02931 & ~w22562;
assign w22573 = ~pi02708 & w22562;
assign w22574 = ~w22572 & ~w22573;
assign w22575 = pi02932 & ~w22562;
assign w22576 = ~pi02709 & w22562;
assign w22577 = ~w22575 & ~w22576;
assign w22578 = pi02933 & ~w22562;
assign w22579 = ~pi02710 & w22562;
assign w22580 = ~w22578 & ~w22579;
assign w22581 = ~w16892 & w18944;
assign w22582 = pi02934 & ~w22581;
assign w22583 = ~pi02705 & w22581;
assign w22584 = ~w22582 & ~w22583;
assign w22585 = pi02935 & ~w22581;
assign w22586 = ~pi02706 & w22581;
assign w22587 = ~w22585 & ~w22586;
assign w22588 = pi02936 & ~w22581;
assign w22589 = ~pi02707 & w22581;
assign w22590 = ~w22588 & ~w22589;
assign w22591 = pi02937 & ~w22581;
assign w22592 = ~pi02160 & w22581;
assign w22593 = ~w22591 & ~w22592;
assign w22594 = pi02938 & ~w22581;
assign w22595 = ~pi02708 & w22581;
assign w22596 = ~w22594 & ~w22595;
assign w22597 = pi02939 & ~w22581;
assign w22598 = ~pi02709 & w22581;
assign w22599 = ~w22597 & ~w22598;
assign w22600 = pi02940 & ~w22581;
assign w22601 = ~pi02710 & w22581;
assign w22602 = ~w22600 & ~w22601;
assign w22603 = ~w16892 & w18913;
assign w22604 = pi02941 & ~w22603;
assign w22605 = w17925 & w18913;
assign w22606 = ~w22604 & ~w22605;
assign w22607 = pi02942 & ~w22603;
assign w22608 = ~pi02707 & w22603;
assign w22609 = ~w22607 & ~w22608;
assign w22610 = pi02943 & ~w22603;
assign w22611 = ~pi02160 & w22603;
assign w22612 = ~w22610 & ~w22611;
assign w22613 = pi02944 & ~w22603;
assign w22614 = ~pi02708 & w22603;
assign w22615 = ~w22613 & ~w22614;
assign w22616 = pi02945 & ~w22603;
assign w22617 = ~pi02709 & w22603;
assign w22618 = ~w22616 & ~w22617;
assign w22619 = pi02946 & ~w22603;
assign w22620 = ~pi02710 & w22603;
assign w22621 = ~w22619 & ~w22620;
assign w22622 = ~w16892 & w18897;
assign w22623 = pi02947 & ~w22622;
assign w22624 = w18578 & w18897;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = pi02948 & ~w22622;
assign w22627 = ~pi02706 & w22622;
assign w22628 = ~w22626 & ~w22627;
assign w22629 = pi02949 & ~w22622;
assign w22630 = ~pi02707 & w22622;
assign w22631 = ~w22629 & ~w22630;
assign w22632 = pi02950 & ~w22622;
assign w22633 = ~pi02160 & w22622;
assign w22634 = ~w22632 & ~w22633;
assign w22635 = pi02951 & ~w22622;
assign w22636 = ~pi02708 & w22622;
assign w22637 = ~w22635 & ~w22636;
assign w22638 = pi02952 & ~w22622;
assign w22639 = ~pi02709 & w22622;
assign w22640 = ~w22638 & ~w22639;
assign w22641 = pi02953 & ~w22622;
assign w22642 = ~pi02710 & w22622;
assign w22643 = ~w22641 & ~w22642;
assign w22644 = ~w16892 & w18871;
assign w22645 = pi02954 & ~w22644;
assign w22646 = ~pi02706 & w22644;
assign w22647 = ~w22645 & ~w22646;
assign w22648 = pi02955 & ~w22644;
assign w22649 = ~pi02707 & w22644;
assign w22650 = ~w22648 & ~w22649;
assign w22651 = pi02956 & ~w22644;
assign w22652 = ~pi02160 & w22644;
assign w22653 = ~w22651 & ~w22652;
assign w22654 = pi02957 & ~w22644;
assign w22655 = w18689 & w18871;
assign w22656 = ~w22654 & ~w22655;
assign w22657 = pi02958 & ~w22644;
assign w22658 = ~pi02709 & w22644;
assign w22659 = ~w22657 & ~w22658;
assign w22660 = pi02959 & ~w22644;
assign w22661 = ~pi02710 & w22644;
assign w22662 = ~w22660 & ~w22661;
assign w22663 = ~w16892 & w18831;
assign w22664 = pi02960 & ~w22663;
assign w22665 = ~pi02705 & w22663;
assign w22666 = ~w22664 & ~w22665;
assign w22667 = pi02961 & ~w22663;
assign w22668 = ~pi02706 & w22663;
assign w22669 = ~w22667 & ~w22668;
assign w22670 = pi02962 & ~w22663;
assign w22671 = ~pi02707 & w22663;
assign w22672 = ~w22670 & ~w22671;
assign w22673 = pi02963 & ~w19088;
assign w22674 = ~pi02704 & w19088;
assign w22675 = ~w22673 & ~w22674;
assign w22676 = pi02964 & ~w22663;
assign w22677 = ~pi02723 & w22663;
assign w22678 = ~w22676 & ~w22677;
assign w22679 = pi02965 & ~w22663;
assign w22680 = ~pi02708 & w22663;
assign w22681 = ~w22679 & ~w22680;
assign w22682 = pi02966 & ~w22663;
assign w22683 = ~pi02709 & w22663;
assign w22684 = ~w22682 & ~w22683;
assign w22685 = ~w16892 & w18822;
assign w22686 = pi02967 & ~w22685;
assign w22687 = ~pi02705 & w22685;
assign w22688 = ~w22686 & ~w22687;
assign w22689 = pi02968 & ~w22685;
assign w22690 = ~pi02706 & w22685;
assign w22691 = ~w22689 & ~w22690;
assign w22692 = pi02969 & ~w22685;
assign w22693 = ~pi02707 & w22685;
assign w22694 = ~w22692 & ~w22693;
assign w22695 = pi02970 & ~w22685;
assign w22696 = ~pi02723 & w22685;
assign w22697 = ~w22695 & ~w22696;
assign w22698 = pi02971 & ~w22685;
assign w22699 = ~pi02708 & w22685;
assign w22700 = ~w22698 & ~w22699;
assign w22701 = pi02972 & ~w22685;
assign w22702 = ~pi02709 & w22685;
assign w22703 = ~w22701 & ~w22702;
assign w22704 = pi02973 & ~w22685;
assign w22705 = ~pi02710 & w22685;
assign w22706 = ~w22704 & ~w22705;
assign w22707 = ~w16892 & w18612;
assign w22708 = pi02974 & ~w22707;
assign w22709 = ~pi02705 & w22707;
assign w22710 = ~w22708 & ~w22709;
assign w22711 = pi02975 & ~w22707;
assign w22712 = ~pi02706 & w22707;
assign w22713 = ~w22711 & ~w22712;
assign w22714 = pi02976 & ~w22707;
assign w22715 = w18067 & w18612;
assign w22716 = ~w22714 & ~w22715;
assign w22717 = pi02977 & ~w22707;
assign w22718 = ~pi02723 & w22707;
assign w22719 = ~w22717 & ~w22718;
assign w22720 = pi02978 & ~w22707;
assign w22721 = ~pi02708 & w22707;
assign w22722 = ~w22720 & ~w22721;
assign w22723 = pi02979 & ~w22707;
assign w22724 = ~pi02709 & w22707;
assign w22725 = ~w22723 & ~w22724;
assign w22726 = ~w16892 & w17516;
assign w22727 = pi02980 & ~w22726;
assign w22728 = ~pi02705 & w22726;
assign w22729 = ~w22727 & ~w22728;
assign w22730 = pi02981 & ~w22726;
assign w22731 = ~pi02706 & w22726;
assign w22732 = ~w22730 & ~w22731;
assign w22733 = pi02982 & ~w22726;
assign w22734 = ~pi02707 & w22726;
assign w22735 = ~w22733 & ~w22734;
assign w22736 = pi02983 & ~w22726;
assign w22737 = ~pi02723 & w22726;
assign w22738 = ~w22736 & ~w22737;
assign w22739 = pi02984 & ~w22726;
assign w22740 = ~pi02708 & w22726;
assign w22741 = ~w22739 & ~w22740;
assign w22742 = pi02985 & ~w22726;
assign w22743 = ~pi02709 & w22726;
assign w22744 = ~w22742 & ~w22743;
assign w22745 = pi02986 & ~w22726;
assign w22746 = w17516 & w18364;
assign w22747 = ~w22745 & ~w22746;
assign w22748 = ~w16892 & w18431;
assign w22749 = pi02987 & ~w22748;
assign w22750 = ~pi02705 & w22748;
assign w22751 = ~w22749 & ~w22750;
assign w22752 = pi02988 & ~w22748;
assign w22753 = ~pi02706 & w22748;
assign w22754 = ~w22752 & ~w22753;
assign w22755 = pi02989 & ~w22748;
assign w22756 = ~pi02707 & w22748;
assign w22757 = ~w22755 & ~w22756;
assign w22758 = pi02990 & ~w22748;
assign w22759 = ~pi02723 & w22748;
assign w22760 = ~w22758 & ~w22759;
assign w22761 = pi02991 & ~w22748;
assign w22762 = ~pi02708 & w22748;
assign w22763 = ~w22761 & ~w22762;
assign w22764 = pi02992 & ~w22748;
assign w22765 = ~pi02709 & w22748;
assign w22766 = ~w22764 & ~w22765;
assign w22767 = ~w16892 & w18247;
assign w22768 = pi02993 & ~w22767;
assign w22769 = ~pi02705 & w22767;
assign w22770 = ~w22768 & ~w22769;
assign w22771 = pi02994 & ~w22767;
assign w22772 = ~pi02706 & w22767;
assign w22773 = ~w22771 & ~w22772;
assign w22774 = pi02995 & ~w22767;
assign w22775 = ~pi02707 & w22767;
assign w22776 = ~w22774 & ~w22775;
assign w22777 = pi02996 & ~w22767;
assign w22778 = w17671 & w18247;
assign w22779 = ~w22777 & ~w22778;
assign w22780 = pi02997 & ~w22767;
assign w22781 = ~pi02708 & w22767;
assign w22782 = ~w22780 & ~w22781;
assign w22783 = pi02998 & ~w22767;
assign w22784 = ~pi02709 & w22767;
assign w22785 = ~w22783 & ~w22784;
assign w22786 = pi02999 & ~w22767;
assign w22787 = ~pi02710 & w22767;
assign w22788 = ~w22786 & ~w22787;
assign w22789 = pi03000 & ~w21492;
assign w22790 = ~pi02705 & w21492;
assign w22791 = ~w22789 & ~w22790;
assign w22792 = pi03001 & ~w21492;
assign w22793 = w17510 & w17925;
assign w22794 = ~w22792 & ~w22793;
assign w22795 = pi03002 & ~w21492;
assign w22796 = ~pi02707 & w21492;
assign w22797 = ~w22795 & ~w22796;
assign w22798 = pi03003 & ~w21492;
assign w22799 = ~pi02723 & w21492;
assign w22800 = ~w22798 & ~w22799;
assign w22801 = pi03004 & ~w21492;
assign w22802 = ~pi02708 & w21492;
assign w22803 = ~w22801 & ~w22802;
assign w22804 = pi03005 & ~w21492;
assign w22805 = ~pi02709 & w21492;
assign w22806 = ~w22804 & ~w22805;
assign w22807 = ~w16892 & w18308;
assign w22808 = pi03006 & ~w22807;
assign w22809 = ~pi02705 & w22807;
assign w22810 = ~w22808 & ~w22809;
assign w22811 = pi03007 & ~w22807;
assign w22812 = ~pi02706 & w22807;
assign w22813 = ~w22811 & ~w22812;
assign w22814 = pi03008 & ~w22807;
assign w22815 = ~pi02707 & w22807;
assign w22816 = ~w22814 & ~w22815;
assign w22817 = pi03009 & ~w22807;
assign w22818 = ~pi02723 & w22807;
assign w22819 = ~w22817 & ~w22818;
assign w22820 = pi03010 & ~w22807;
assign w22821 = w18308 & w18689;
assign w22822 = ~w22820 & ~w22821;
assign w22823 = pi03011 & ~w22807;
assign w22824 = ~pi02709 & w22807;
assign w22825 = ~w22823 & ~w22824;
assign w22826 = pi03012 & ~w22807;
assign w22827 = ~pi02710 & w22807;
assign w22828 = ~w22826 & ~w22827;
assign w22829 = pi03013 & ~w22189;
assign w22830 = ~pi02705 & w22189;
assign w22831 = ~w22829 & ~w22830;
assign w22832 = pi03014 & ~w22189;
assign w22833 = ~pi02706 & w22189;
assign w22834 = ~w22832 & ~w22833;
assign w22835 = pi03015 & ~w22189;
assign w22836 = w18067 & w18263;
assign w22837 = ~w22835 & ~w22836;
assign w22838 = pi03016 & ~w22189;
assign w22839 = ~pi02723 & w22189;
assign w22840 = ~w22838 & ~w22839;
assign w22841 = pi03017 & ~w22189;
assign w22842 = ~pi02708 & w22189;
assign w22843 = ~w22841 & ~w22842;
assign w22844 = pi03018 & ~w22189;
assign w22845 = w18092 & w18263;
assign w22846 = ~w22844 & ~w22845;
assign w22847 = pi03019 & ~w19080;
assign w22848 = ~pi09848 & w19080;
assign w22849 = ~w22847 & ~w22848;
assign w22850 = pi03020 & ~w22193;
assign w22851 = ~pi02705 & w22193;
assign w22852 = ~w22850 & ~w22851;
assign w22853 = pi03021 & ~w22193;
assign w22854 = w17925 & w18155;
assign w22855 = ~w22853 & ~w22854;
assign w22856 = pi03022 & ~w22193;
assign w22857 = w18155 & w18234;
assign w22858 = ~w22856 & ~w22857;
assign w22859 = pi03023 & ~w22193;
assign w22860 = w17671 & w18155;
assign w22861 = ~w22859 & ~w22860;
assign w22862 = pi03024 & ~w22193;
assign w22863 = ~pi02708 & w22193;
assign w22864 = ~w22862 & ~w22863;
assign w22865 = pi03025 & ~w22193;
assign w22866 = ~pi02709 & w22193;
assign w22867 = ~w22865 & ~w22866;
assign w22868 = pi03026 & ~w22193;
assign w22869 = w18155 & w18364;
assign w22870 = ~w22868 & ~w22869;
assign w22871 = pi03027 & ~w21095;
assign w22872 = ~pi02705 & w21095;
assign w22873 = ~w22871 & ~w22872;
assign w22874 = pi03028 & ~w21095;
assign w22875 = ~pi02706 & w21095;
assign w22876 = ~w22874 & ~w22875;
assign w22877 = pi03029 & ~w21095;
assign w22878 = ~pi02160 & w21095;
assign w22879 = ~w22877 & ~w22878;
assign w22880 = pi03030 & ~w21095;
assign w22881 = ~pi02723 & w21095;
assign w22882 = ~w22880 & ~w22881;
assign w22883 = pi03031 & ~w21095;
assign w22884 = w18146 & w18689;
assign w22885 = ~w22883 & ~w22884;
assign w22886 = pi03032 & ~w21095;
assign w22887 = ~pi02710 & w21095;
assign w22888 = ~w22886 & ~w22887;
assign w22889 = pi03033 & ~w21018;
assign w22890 = ~pi02705 & w21018;
assign w22891 = ~w22889 & ~w22890;
assign w22892 = pi03034 & ~w21018;
assign w22893 = ~pi02706 & w21018;
assign w22894 = ~w22892 & ~w22893;
assign w22895 = pi03035 & ~w21018;
assign w22896 = ~pi02160 & w21018;
assign w22897 = ~w22895 & ~w22896;
assign w22898 = pi03036 & ~w21018;
assign w22899 = w17671 & w18116;
assign w22900 = ~w22898 & ~w22899;
assign w22901 = pi03037 & ~w21018;
assign w22902 = ~pi02708 & w21018;
assign w22903 = ~w22901 & ~w22902;
assign w22904 = pi03038 & ~w21018;
assign w22905 = ~pi02709 & w21018;
assign w22906 = ~w22904 & ~w22905;
assign w22907 = pi03039 & ~w21018;
assign w22908 = ~pi02710 & w21018;
assign w22909 = ~w22907 & ~w22908;
assign w22910 = pi03040 & ~w20407;
assign w22911 = w18070 & w18578;
assign w22912 = ~w22910 & ~w22911;
assign w22913 = pi03041 & ~w20407;
assign w22914 = ~pi02706 & w20407;
assign w22915 = ~w22913 & ~w22914;
assign w22916 = pi03042 & ~w20407;
assign w22917 = ~pi02160 & w20407;
assign w22918 = ~w22916 & ~w22917;
assign w22919 = pi03043 & ~w20407;
assign w22920 = ~pi02723 & w20407;
assign w22921 = ~w22919 & ~w22920;
assign w22922 = pi03044 & ~w20407;
assign w22923 = ~pi02708 & w20407;
assign w22924 = ~w22922 & ~w22923;
assign w22925 = pi03045 & ~w20407;
assign w22926 = ~pi02710 & w20407;
assign w22927 = ~w22925 & ~w22926;
assign w22928 = pi03046 & ~w20581;
assign w22929 = ~pi02705 & w20581;
assign w22930 = ~w22928 & ~w22929;
assign w22931 = pi03047 & ~w20581;
assign w22932 = ~pi02706 & w20581;
assign w22933 = ~w22931 & ~w22932;
assign w22934 = pi03048 & ~w20581;
assign w22935 = ~pi02160 & w20581;
assign w22936 = ~w22934 & ~w22935;
assign w22937 = pi03049 & ~w20581;
assign w22938 = ~pi02723 & w20581;
assign w22939 = ~w22937 & ~w22938;
assign w22940 = pi03050 & ~w20581;
assign w22941 = ~pi02708 & w20581;
assign w22942 = ~w22940 & ~w22941;
assign w22943 = pi03051 & ~w20581;
assign w22944 = ~pi02709 & w20581;
assign w22945 = ~w22943 & ~w22944;
assign w22946 = pi03052 & ~w20581;
assign w22947 = ~pi02710 & w20581;
assign w22948 = ~w22946 & ~w22947;
assign w22949 = pi03053 & ~w20637;
assign w22950 = ~pi02705 & w20637;
assign w22951 = ~w22949 & ~w22950;
assign w22952 = pi03054 & ~w20637;
assign w22953 = ~pi02706 & w20637;
assign w22954 = ~w22952 & ~w22953;
assign w22955 = pi03055 & ~w20637;
assign w22956 = ~pi02160 & w20637;
assign w22957 = ~w22955 & ~w22956;
assign w22958 = pi03056 & ~w20637;
assign w22959 = ~pi02723 & w20637;
assign w22960 = ~w22958 & ~w22959;
assign w22961 = pi03057 & ~w20637;
assign w22962 = ~pi02708 & w20637;
assign w22963 = ~w22961 & ~w22962;
assign w22964 = pi03058 & ~w20637;
assign w22965 = ~pi02710 & w20637;
assign w22966 = ~w22964 & ~w22965;
assign w22967 = pi03059 & ~w20617;
assign w22968 = ~pi02705 & w20617;
assign w22969 = ~w22967 & ~w22968;
assign w22970 = pi03060 & ~w20617;
assign w22971 = w17445 & w17925;
assign w22972 = ~w22970 & ~w22971;
assign w22973 = pi03061 & ~w20617;
assign w22974 = w17445 & w18234;
assign w22975 = ~w22973 & ~w22974;
assign w22976 = pi03062 & ~w20617;
assign w22977 = ~pi02723 & w20617;
assign w22978 = ~w22976 & ~w22977;
assign w22979 = pi03063 & ~w20617;
assign w22980 = ~pi02708 & w20617;
assign w22981 = ~w22979 & ~w22980;
assign w22982 = pi03064 & ~w20617;
assign w22983 = ~pi02709 & w20617;
assign w22984 = ~w22982 & ~w22983;
assign w22985 = pi03065 & ~w20617;
assign w22986 = w17445 & w18364;
assign w22987 = ~w22985 & ~w22986;
assign w22988 = pi03066 & ~w20411;
assign w22989 = ~pi02705 & w20411;
assign w22990 = ~w22988 & ~w22989;
assign w22991 = pi03067 & ~w20411;
assign w22992 = ~pi02706 & w20411;
assign w22993 = ~w22991 & ~w22992;
assign w22994 = pi03068 & ~w20411;
assign w22995 = ~pi02160 & w20411;
assign w22996 = ~w22994 & ~w22995;
assign w22997 = pi03069 & ~w20411;
assign w22998 = ~pi02723 & w20411;
assign w22999 = ~w22997 & ~w22998;
assign w23000 = pi03070 & ~w20411;
assign w23001 = ~pi02708 & w20411;
assign w23002 = ~w23000 & ~w23001;
assign w23003 = pi03071 & ~w20411;
assign w23004 = ~pi02710 & w20411;
assign w23005 = ~w23003 & ~w23004;
assign w23006 = pi03072 & ~w20549;
assign w23007 = ~pi02705 & w20549;
assign w23008 = ~w23006 & ~w23007;
assign w23009 = pi03073 & ~w20549;
assign w23010 = ~pi02706 & w20549;
assign w23011 = ~w23009 & ~w23010;
assign w23012 = pi03074 & ~w20549;
assign w23013 = ~pi02160 & w20549;
assign w23014 = ~w23012 & ~w23013;
assign w23015 = pi03075 & ~w20549;
assign w23016 = ~pi02723 & w20549;
assign w23017 = ~w23015 & ~w23016;
assign w23018 = pi03076 & ~w20549;
assign w23019 = ~pi02708 & w20549;
assign w23020 = ~w23018 & ~w23019;
assign w23021 = pi03077 & ~w20549;
assign w23022 = ~pi02709 & w20549;
assign w23023 = ~w23021 & ~w23022;
assign w23024 = pi03078 & ~w20549;
assign w23025 = ~pi02710 & w20549;
assign w23026 = ~w23024 & ~w23025;
assign w23027 = pi03079 & ~w20277;
assign w23028 = ~pi02705 & w20277;
assign w23029 = ~w23027 & ~w23028;
assign w23030 = pi03080 & ~w20277;
assign w23031 = ~pi02706 & w20277;
assign w23032 = ~w23030 & ~w23031;
assign w23033 = pi03081 & ~w20277;
assign w23034 = ~pi02160 & w20277;
assign w23035 = ~w23033 & ~w23034;
assign w23036 = pi03082 & ~w20277;
assign w23037 = ~pi02723 & w20277;
assign w23038 = ~w23036 & ~w23037;
assign w23039 = pi03083 & ~w20277;
assign w23040 = ~pi02708 & w20277;
assign w23041 = ~w23039 & ~w23040;
assign w23042 = pi03084 & ~w20277;
assign w23043 = ~pi02710 & w20277;
assign w23044 = ~w23042 & ~w23043;
assign w23045 = pi03085 & ~w20353;
assign w23046 = ~pi02705 & w20353;
assign w23047 = ~w23045 & ~w23046;
assign w23048 = pi03086 & ~w20353;
assign w23049 = ~pi02706 & w20353;
assign w23050 = ~w23048 & ~w23049;
assign w23051 = pi03087 & ~w20353;
assign w23052 = ~pi02160 & w20353;
assign w23053 = ~w23051 & ~w23052;
assign w23054 = pi03088 & ~w20353;
assign w23055 = w17671 & w17965;
assign w23056 = ~w23054 & ~w23055;
assign w23057 = pi03089 & ~w20353;
assign w23058 = w17965 & w18689;
assign w23059 = ~w23057 & ~w23058;
assign w23060 = pi03090 & ~w20353;
assign w23061 = ~pi02709 & w20353;
assign w23062 = ~w23060 & ~w23061;
assign w23063 = pi03091 & ~w20353;
assign w23064 = w17965 & w18364;
assign w23065 = ~w23063 & ~w23064;
assign w23066 = pi03092 & ~w20034;
assign w23067 = w17912 & w18578;
assign w23068 = ~w23066 & ~w23067;
assign w23069 = pi03093 & ~w20034;
assign w23070 = ~pi02706 & w20034;
assign w23071 = ~w23069 & ~w23070;
assign w23072 = pi03094 & ~w20034;
assign w23073 = ~pi02160 & w20034;
assign w23074 = ~w23072 & ~w23073;
assign w23075 = pi03095 & ~w20034;
assign w23076 = ~pi02723 & w20034;
assign w23077 = ~w23075 & ~w23076;
assign w23078 = pi03096 & ~w20034;
assign w23079 = ~pi02708 & w20034;
assign w23080 = ~w23078 & ~w23079;
assign w23081 = pi03097 & ~w20034;
assign w23082 = ~pi02710 & w20034;
assign w23083 = ~w23081 & ~w23082;
assign w23084 = pi03098 & ~w20136;
assign w23085 = ~pi02705 & w20136;
assign w23086 = ~w23084 & ~w23085;
assign w23087 = pi03099 & ~w20136;
assign w23088 = ~pi02706 & w20136;
assign w23089 = ~w23087 & ~w23088;
assign w23090 = pi03100 & ~w20136;
assign w23091 = ~pi02160 & w20136;
assign w23092 = ~w23090 & ~w23091;
assign w23093 = pi03101 & ~w20136;
assign w23094 = ~pi02723 & w20136;
assign w23095 = ~w23093 & ~w23094;
assign w23096 = pi03102 & ~w20136;
assign w23097 = ~pi02708 & w20136;
assign w23098 = ~w23096 & ~w23097;
assign w23099 = pi03103 & ~w20136;
assign w23100 = ~pi02709 & w20136;
assign w23101 = ~w23099 & ~w23100;
assign w23102 = pi03104 & ~w20136;
assign w23103 = ~pi02710 & w20136;
assign w23104 = ~w23102 & ~w23103;
assign w23105 = pi03105 & ~w20120;
assign w23106 = w18578 & w20119;
assign w23107 = ~w23105 & ~w23106;
assign w23108 = pi03106 & ~w20120;
assign w23109 = ~pi02706 & w20120;
assign w23110 = ~w23108 & ~w23109;
assign w23111 = pi03107 & ~w20120;
assign w23112 = ~pi02160 & w20120;
assign w23113 = ~w23111 & ~w23112;
assign w23114 = pi03108 & ~w20120;
assign w23115 = ~pi02723 & w20120;
assign w23116 = ~w23114 & ~w23115;
assign w23117 = pi03109 & ~w20120;
assign w23118 = w18689 & w20119;
assign w23119 = ~w23117 & ~w23118;
assign w23120 = pi03110 & ~w20120;
assign w23121 = ~pi02710 & w20120;
assign w23122 = ~w23120 & ~w23121;
assign w23123 = pi03111 & ~w20115;
assign w23124 = ~pi02705 & w20115;
assign w23125 = ~w23123 & ~w23124;
assign w23126 = pi03112 & ~w20115;
assign w23127 = ~pi02706 & w20115;
assign w23128 = ~w23126 & ~w23127;
assign w23129 = pi03113 & ~w21277;
assign w23130 = ~pi02714 & w21277;
assign w23131 = ~w23129 & ~w23130;
assign w23132 = pi03114 & ~w18848;
assign w23133 = ~pi09848 & w18848;
assign w23134 = ~w23132 & ~w23133;
assign w23135 = pi03115 & ~w20115;
assign w23136 = ~pi02160 & w20115;
assign w23137 = ~w23135 & ~w23136;
assign w23138 = pi03116 & ~w20115;
assign w23139 = ~pi02723 & w20115;
assign w23140 = ~w23138 & ~w23139;
assign w23141 = pi03117 & ~w20115;
assign w23142 = ~pi02708 & w20115;
assign w23143 = ~w23141 & ~w23142;
assign w23144 = pi03118 & ~w20115;
assign w23145 = ~pi02709 & w20115;
assign w23146 = ~w23144 & ~w23145;
assign w23147 = pi03119 & ~w20115;
assign w23148 = ~pi02710 & w20115;
assign w23149 = ~w23147 & ~w23148;
assign w23150 = pi03120 & ~w20097;
assign w23151 = ~pi02705 & w20097;
assign w23152 = ~w23150 & ~w23151;
assign w23153 = pi03121 & ~w20097;
assign w23154 = ~pi02706 & w20097;
assign w23155 = ~w23153 & ~w23154;
assign w23156 = pi03122 & ~w20097;
assign w23157 = ~pi02160 & w20097;
assign w23158 = ~w23156 & ~w23157;
assign w23159 = pi03123 & ~w20097;
assign w23160 = ~pi02723 & w20097;
assign w23161 = ~w23159 & ~w23160;
assign w23162 = pi03124 & ~w20097;
assign w23163 = ~pi02708 & w20097;
assign w23164 = ~w23162 & ~w23163;
assign w23165 = pi03125 & ~w20097;
assign w23166 = ~pi02710 & w20097;
assign w23167 = ~w23165 & ~w23166;
assign w23168 = pi03126 & ~w20080;
assign w23169 = w17078 & w18578;
assign w23170 = ~w23168 & ~w23169;
assign w23171 = pi03127 & ~w20080;
assign w23172 = w17078 & w17925;
assign w23173 = ~w23171 & ~w23172;
assign w23174 = pi03128 & ~w20080;
assign w23175 = w17078 & w18234;
assign w23176 = ~w23174 & ~w23175;
assign w23177 = pi03129 & ~w20080;
assign w23178 = w17078 & w17671;
assign w23179 = ~w23177 & ~w23178;
assign w23180 = pi03130 & ~w20080;
assign w23181 = w17078 & w18689;
assign w23182 = ~w23180 & ~w23181;
assign w23183 = pi03131 & ~w20080;
assign w23184 = w17078 & w18092;
assign w23185 = ~w23183 & ~w23184;
assign w23186 = pi03132 & ~w20080;
assign w23187 = w17078 & w18364;
assign w23188 = ~w23186 & ~w23187;
assign w23189 = pi03133 & ~w20076;
assign w23190 = ~pi02705 & w20076;
assign w23191 = ~w23189 & ~w23190;
assign w23192 = pi03134 & ~w20076;
assign w23193 = ~pi02706 & w20076;
assign w23194 = ~w23192 & ~w23193;
assign w23195 = pi03135 & ~w20076;
assign w23196 = ~pi02160 & w20076;
assign w23197 = ~w23195 & ~w23196;
assign w23198 = pi03136 & ~w20076;
assign w23199 = ~pi02723 & w20076;
assign w23200 = ~w23198 & ~w23199;
assign w23201 = pi03137 & ~w20076;
assign w23202 = ~pi02708 & w20076;
assign w23203 = ~w23201 & ~w23202;
assign w23204 = pi03138 & ~w20076;
assign w23205 = ~pi02710 & w20076;
assign w23206 = ~w23204 & ~w23205;
assign w23207 = pi03139 & ~w20060;
assign w23208 = w18578 & w20059;
assign w23209 = ~w23207 & ~w23208;
assign w23210 = pi03140 & ~w20060;
assign w23211 = ~pi02706 & w20060;
assign w23212 = ~w23210 & ~w23211;
assign w23213 = pi03141 & ~w20060;
assign w23214 = ~pi02160 & w20060;
assign w23215 = ~w23213 & ~w23214;
assign w23216 = pi03142 & ~w20060;
assign w23217 = ~pi02723 & w20060;
assign w23218 = ~w23216 & ~w23217;
assign w23219 = pi03143 & ~w19914;
assign w23220 = ~pi02703 & w19914;
assign w23221 = ~w23219 & ~w23220;
assign w23222 = pi03144 & ~w20060;
assign w23223 = ~pi02708 & w20060;
assign w23224 = ~w23222 & ~w23223;
assign w23225 = pi03145 & ~w20060;
assign w23226 = ~pi02709 & w20060;
assign w23227 = ~w23225 & ~w23226;
assign w23228 = pi03146 & ~w20060;
assign w23229 = ~pi02710 & w20060;
assign w23230 = ~w23228 & ~w23229;
assign w23231 = pi03147 & ~w19914;
assign w23232 = ~pi02721 & w19914;
assign w23233 = ~w23231 & ~w23232;
assign w23234 = pi03148 & ~w19914;
assign w23235 = ~pi02718 & w19914;
assign w23236 = ~w23234 & ~w23235;
assign w23237 = pi03149 & ~w19914;
assign w23238 = ~pi02167 & w19914;
assign w23239 = ~w23237 & ~w23238;
assign w23240 = pi03150 & ~w20015;
assign w23241 = w18578 & w20014;
assign w23242 = ~w23240 & ~w23241;
assign w23243 = pi03151 & ~w20015;
assign w23244 = ~pi02706 & w20015;
assign w23245 = ~w23243 & ~w23244;
assign w23246 = pi03152 & ~w20015;
assign w23247 = w18067 & w20014;
assign w23248 = ~w23246 & ~w23247;
assign w23249 = pi03153 & ~w19914;
assign w23250 = ~pi02722 & w19914;
assign w23251 = ~w23249 & ~w23250;
assign w23252 = pi03154 & ~w20015;
assign w23253 = ~pi02723 & w20015;
assign w23254 = ~w23252 & ~w23253;
assign w23255 = pi03155 & ~w19914;
assign w23256 = ~pi02719 & w19914;
assign w23257 = ~w23255 & ~w23256;
assign w23258 = pi03156 & ~w20015;
assign w23259 = ~pi02708 & w20015;
assign w23260 = ~w23258 & ~w23259;
assign w23261 = pi03157 & ~w20015;
assign w23262 = w18092 & w20014;
assign w23263 = ~w23261 & ~w23262;
assign w23264 = pi03158 & ~w20015;
assign w23265 = ~pi02710 & w20015;
assign w23266 = ~w23264 & ~w23265;
assign w23267 = pi03159 & ~w19996;
assign w23268 = ~pi02703 & w19996;
assign w23269 = ~w23267 & ~w23268;
assign w23270 = pi03160 & ~w19996;
assign w23271 = ~pi02721 & w19996;
assign w23272 = ~w23270 & ~w23271;
assign w23273 = pi03161 & ~w19996;
assign w23274 = ~pi02718 & w19996;
assign w23275 = ~w23273 & ~w23274;
assign w23276 = pi03162 & ~w19996;
assign w23277 = ~pi02167 & w19996;
assign w23278 = ~w23276 & ~w23277;
assign w23279 = pi03163 & ~w19996;
assign w23280 = ~pi02164 & w19996;
assign w23281 = ~w23279 & ~w23280;
assign w23282 = pi03164 & ~w19996;
assign w23283 = ~pi02719 & w19996;
assign w23284 = ~w23282 & ~w23283;
assign w23285 = pi03165 & ~w19989;
assign w23286 = ~pi02705 & w19989;
assign w23287 = ~w23285 & ~w23286;
assign w23288 = pi03166 & ~w19989;
assign w23289 = ~pi02706 & w19989;
assign w23290 = ~w23288 & ~w23289;
assign w23291 = pi03167 & ~w19989;
assign w23292 = ~pi02160 & w19989;
assign w23293 = ~w23291 & ~w23292;
assign w23294 = pi03168 & ~w19989;
assign w23295 = ~pi02723 & w19989;
assign w23296 = ~w23294 & ~w23295;
assign w23297 = pi03169 & ~w19989;
assign w23298 = ~pi02708 & w19989;
assign w23299 = ~w23297 & ~w23298;
assign w23300 = pi03170 & ~w19989;
assign w23301 = w18092 & w19988;
assign w23302 = ~w23300 & ~w23301;
assign w23303 = pi03171 & ~w19989;
assign w23304 = ~pi02710 & w19989;
assign w23305 = ~w23303 & ~w23304;
assign w23306 = pi03172 & ~w19942;
assign w23307 = ~pi02705 & w19942;
assign w23308 = ~w23306 & ~w23307;
assign w23309 = pi03173 & ~w19942;
assign w23310 = ~pi02706 & w19942;
assign w23311 = ~w23309 & ~w23310;
assign w23312 = pi03174 & ~w19942;
assign w23313 = ~pi02160 & w19942;
assign w23314 = ~w23312 & ~w23313;
assign w23315 = pi03175 & ~w19942;
assign w23316 = ~pi02723 & w19942;
assign w23317 = ~w23315 & ~w23316;
assign w23318 = pi03176 & ~w19942;
assign w23319 = ~pi02708 & w19942;
assign w23320 = ~w23318 & ~w23319;
assign w23321 = pi03177 & ~w19942;
assign w23322 = w18364 & w19941;
assign w23323 = ~w23321 & ~w23322;
assign w23324 = pi03178 & ~w19959;
assign w23325 = w17218 & w17532;
assign w23326 = ~w23324 & ~w23325;
assign w23327 = pi03179 & ~w19959;
assign w23328 = w17218 & w17811;
assign w23329 = ~w23327 & ~w23328;
assign w23330 = pi03180 & ~w19959;
assign w23331 = w17218 & w17586;
assign w23332 = ~w23330 & ~w23331;
assign w23333 = pi03181 & ~w19959;
assign w23334 = w17218 & w19273;
assign w23335 = ~w23333 & ~w23334;
assign w23336 = pi03182 & ~w19959;
assign w23337 = w17218 & w17620;
assign w23338 = ~w23336 & ~w23337;
assign w23339 = pi03183 & ~w19959;
assign w23340 = w17218 & w19312;
assign w23341 = ~w23339 & ~w23340;
assign w23342 = pi03184 & ~w19959;
assign w23343 = w17218 & w17594;
assign w23344 = ~w23342 & ~w23343;
assign w23345 = pi03185 & ~w19918;
assign w23346 = w16948 & w17532;
assign w23347 = ~w23345 & ~w23346;
assign w23348 = pi03186 & ~w19918;
assign w23349 = w16948 & w17811;
assign w23350 = ~w23348 & ~w23349;
assign w23351 = pi03187 & ~w19918;
assign w23352 = w16948 & w17586;
assign w23353 = ~w23351 & ~w23352;
assign w23354 = pi03188 & ~w19918;
assign w23355 = ~pi02167 & w19918;
assign w23356 = ~w23354 & ~w23355;
assign w23357 = pi03189 & ~w19918;
assign w23358 = ~pi02164 & w19918;
assign w23359 = ~w23357 & ~w23358;
assign w23360 = pi03190 & ~w19918;
assign w23361 = ~pi02719 & w19918;
assign w23362 = ~w23360 & ~w23361;
assign w23363 = pi03191 & ~w19899;
assign w23364 = ~pi02703 & w19899;
assign w23365 = ~w23363 & ~w23364;
assign w23366 = pi03192 & ~w19931;
assign w23367 = ~pi02705 & w19931;
assign w23368 = ~w23366 & ~w23367;
assign w23369 = pi03193 & ~w19931;
assign w23370 = ~pi02707 & w19931;
assign w23371 = ~w23369 & ~w23370;
assign w23372 = pi03194 & ~w19931;
assign w23373 = ~pi02160 & w19931;
assign w23374 = ~w23372 & ~w23373;
assign w23375 = pi03195 & ~w19899;
assign w23376 = ~pi02721 & w19899;
assign w23377 = ~w23375 & ~w23376;
assign w23378 = pi03196 & ~w19931;
assign w23379 = ~pi02723 & w19931;
assign w23380 = ~w23378 & ~w23379;
assign w23381 = pi03197 & ~w19931;
assign w23382 = w18689 & w19930;
assign w23383 = ~w23381 & ~w23382;
assign w23384 = pi03198 & ~w19931;
assign w23385 = ~pi02709 & w19931;
assign w23386 = ~w23384 & ~w23385;
assign w23387 = pi03199 & ~w19899;
assign w23388 = ~pi02169 & w19899;
assign w23389 = ~w23387 & ~w23388;
assign w23390 = pi03200 & ~w19910;
assign w23391 = ~pi02705 & w19910;
assign w23392 = ~w23390 & ~w23391;
assign w23393 = pi03201 & ~w19899;
assign w23394 = w17131 & w17586;
assign w23395 = ~w23393 & ~w23394;
assign w23396 = pi03202 & ~w19899;
assign w23397 = ~pi02167 & w19899;
assign w23398 = ~w23396 & ~w23397;
assign w23399 = pi03203 & ~w19910;
assign w23400 = ~pi02707 & w19910;
assign w23401 = ~w23399 & ~w23400;
assign w23402 = pi03204 & ~w19910;
assign w23403 = w18234 & w19909;
assign w23404 = ~w23402 & ~w23403;
assign w23405 = pi03205 & ~w19910;
assign w23406 = ~pi02723 & w19910;
assign w23407 = ~w23405 & ~w23406;
assign w23408 = pi03206 & ~w19910;
assign w23409 = ~pi02708 & w19910;
assign w23410 = ~w23408 & ~w23409;
assign w23411 = pi03207 & ~w19910;
assign w23412 = ~pi02709 & w19910;
assign w23413 = ~w23411 & ~w23412;
assign w23414 = pi03208 & ~w19910;
assign w23415 = ~pi02710 & w19910;
assign w23416 = ~w23414 & ~w23415;
assign w23417 = pi03209 & ~w19899;
assign w23418 = ~pi02722 & w19899;
assign w23419 = ~w23417 & ~w23418;
assign w23420 = pi03210 & ~w19899;
assign w23421 = ~pi02719 & w19899;
assign w23422 = ~w23420 & ~w23421;
assign w23423 = pi03211 & ~w19895;
assign w23424 = ~pi02703 & w19895;
assign w23425 = ~w23423 & ~w23424;
assign w23426 = pi03212 & ~w19895;
assign w23427 = ~pi02721 & w19895;
assign w23428 = ~w23426 & ~w23427;
assign w23429 = pi03213 & ~w19895;
assign w23430 = ~pi02718 & w19895;
assign w23431 = ~w23429 & ~w23430;
assign w23432 = pi03214 & ~w19895;
assign w23433 = ~pi02167 & w19895;
assign w23434 = ~w23432 & ~w23433;
assign w23435 = pi03215 & ~w19895;
assign w23436 = ~pi02164 & w19895;
assign w23437 = ~w23435 & ~w23436;
assign w23438 = pi03216 & ~w19895;
assign w23439 = ~pi02719 & w19895;
assign w23440 = ~w23438 & ~w23439;
assign w23441 = pi03217 & ~w19884;
assign w23442 = ~pi02703 & w19884;
assign w23443 = ~w23441 & ~w23442;
assign w23444 = pi03218 & ~w19884;
assign w23445 = w17811 & w19106;
assign w23446 = ~w23444 & ~w23445;
assign w23447 = ~w16992 & w18617;
assign w23448 = pi03219 & ~w23447;
assign w23449 = ~pi02703 & w23447;
assign w23450 = ~w23448 & ~w23449;
assign w23451 = pi03220 & ~w19884;
assign w23452 = w17586 & w19106;
assign w23453 = ~w23451 & ~w23452;
assign w23454 = pi03221 & ~w19884;
assign w23455 = w19106 & w19273;
assign w23456 = ~w23454 & ~w23455;
assign w23457 = pi03222 & ~w19884;
assign w23458 = ~pi02164 & w19884;
assign w23459 = ~w23457 & ~w23458;
assign w23460 = pi03223 & ~w19884;
assign w23461 = ~pi02722 & w19884;
assign w23462 = ~w23460 & ~w23461;
assign w23463 = pi03224 & ~w19884;
assign w23464 = ~pi02719 & w19884;
assign w23465 = ~w23463 & ~w23464;
assign w23466 = pi03225 & ~w19853;
assign w23467 = w18578 & w19852;
assign w23468 = ~w23466 & ~w23467;
assign w23469 = pi03226 & ~w19853;
assign w23470 = w17925 & w19852;
assign w23471 = ~w23469 & ~w23470;
assign w23472 = pi03227 & ~w19853;
assign w23473 = w18234 & w19852;
assign w23474 = ~w23472 & ~w23473;
assign w23475 = pi03228 & ~w19853;
assign w23476 = w17671 & w19852;
assign w23477 = ~w23475 & ~w23476;
assign w23478 = pi03229 & ~w19853;
assign w23479 = w18689 & w19852;
assign w23480 = ~w23478 & ~w23479;
assign w23481 = pi03230 & ~w19853;
assign w23482 = w18364 & w19852;
assign w23483 = ~w23481 & ~w23482;
assign w23484 = pi03231 & ~w19860;
assign w23485 = ~pi02703 & w19860;
assign w23486 = ~w23484 & ~w23485;
assign w23487 = pi03232 & ~w19860;
assign w23488 = ~pi02721 & w19860;
assign w23489 = ~w23487 & ~w23488;
assign w23490 = pi03233 & ~w19860;
assign w23491 = ~pi02718 & w19860;
assign w23492 = ~w23490 & ~w23491;
assign w23493 = pi03234 & ~w19860;
assign w23494 = ~pi02167 & w19860;
assign w23495 = ~w23493 & ~w23494;
assign w23496 = pi03235 & ~w19839;
assign w23497 = ~pi02705 & w19839;
assign w23498 = ~w23496 & ~w23497;
assign w23499 = pi03236 & ~w19839;
assign w23500 = w17925 & w19838;
assign w23501 = ~w23499 & ~w23500;
assign w23502 = pi03237 & ~w19860;
assign w23503 = ~pi02164 & w19860;
assign w23504 = ~w23502 & ~w23503;
assign w23505 = pi03238 & ~w19839;
assign w23506 = ~pi02707 & w19839;
assign w23507 = ~w23505 & ~w23506;
assign w23508 = pi03239 & ~w19860;
assign w23509 = w19149 & w19312;
assign w23510 = ~w23508 & ~w23509;
assign w23511 = pi03240 & ~w19860;
assign w23512 = w17594 & w19149;
assign w23513 = ~w23511 & ~w23512;
assign w23514 = pi03241 & ~w19839;
assign w23515 = ~pi02723 & w19839;
assign w23516 = ~w23514 & ~w23515;
assign w23517 = pi03242 & ~w19839;
assign w23518 = w18689 & w19838;
assign w23519 = ~w23517 & ~w23518;
assign w23520 = pi03243 & ~w19839;
assign w23521 = ~pi02710 & w19839;
assign w23522 = ~w23520 & ~w23521;
assign w23523 = pi03244 & ~w19827;
assign w23524 = ~pi02705 & w19827;
assign w23525 = ~w23523 & ~w23524;
assign w23526 = pi03245 & ~w19827;
assign w23527 = ~pi02706 & w19827;
assign w23528 = ~w23526 & ~w23527;
assign w23529 = ~w16928 & w17565;
assign w23530 = pi03246 & ~w23529;
assign w23531 = ~pi09962 & w23529;
assign w23532 = ~w23530 & ~w23531;
assign w23533 = pi03247 & ~w19827;
assign w23534 = ~pi02160 & w19827;
assign w23535 = ~w23533 & ~w23534;
assign w23536 = pi03248 & ~w19827;
assign w23537 = ~pi02723 & w19827;
assign w23538 = ~w23536 & ~w23537;
assign w23539 = pi03249 & ~w19827;
assign w23540 = ~pi02708 & w19827;
assign w23541 = ~w23539 & ~w23540;
assign w23542 = pi03250 & ~w19827;
assign w23543 = ~pi02709 & w19827;
assign w23544 = ~w23542 & ~w23543;
assign w23545 = pi03251 & ~w19827;
assign w23546 = ~pi02710 & w19827;
assign w23547 = ~w23545 & ~w23546;
assign w23548 = pi03252 & ~w19819;
assign w23549 = ~pi02705 & w19819;
assign w23550 = ~w23548 & ~w23549;
assign w23551 = pi03253 & ~w19819;
assign w23552 = ~pi02706 & w19819;
assign w23553 = ~w23551 & ~w23552;
assign w23554 = pi03254 & ~w19819;
assign w23555 = ~pi02160 & w19819;
assign w23556 = ~w23554 & ~w23555;
assign w23557 = pi03255 & ~w19819;
assign w23558 = ~pi02723 & w19819;
assign w23559 = ~w23557 & ~w23558;
assign w23560 = pi03256 & ~w19819;
assign w23561 = w18689 & w19818;
assign w23562 = ~w23560 & ~w23561;
assign w23563 = pi03257 & ~w19819;
assign w23564 = w18364 & w19818;
assign w23565 = ~w23563 & ~w23564;
assign w23566 = pi03258 & ~w19807;
assign w23567 = ~pi02703 & w19807;
assign w23568 = ~w23566 & ~w23567;
assign w23569 = pi03259 & ~w19807;
assign w23570 = ~pi02721 & w19807;
assign w23571 = ~w23569 & ~w23570;
assign w23572 = pi03260 & ~w19807;
assign w23573 = ~pi02718 & w19807;
assign w23574 = ~w23572 & ~w23573;
assign w23575 = pi03261 & ~w19807;
assign w23576 = ~pi02167 & w19807;
assign w23577 = ~w23575 & ~w23576;
assign w23578 = pi03262 & ~w19807;
assign w23579 = ~pi02164 & w19807;
assign w23580 = ~w23578 & ~w23579;
assign w23581 = pi03263 & ~w19807;
assign w23582 = ~pi02722 & w19807;
assign w23583 = ~w23581 & ~w23582;
assign w23584 = pi03264 & ~w19807;
assign w23585 = ~pi02719 & w19807;
assign w23586 = ~w23584 & ~w23585;
assign w23587 = pi03265 & ~w19773;
assign w23588 = w17532 & w19130;
assign w23589 = ~w23587 & ~w23588;
assign w23590 = pi03266 & ~w19773;
assign w23591 = w17811 & w19130;
assign w23592 = ~w23590 & ~w23591;
assign w23593 = pi03267 & ~w19741;
assign w23594 = w18578 & w19740;
assign w23595 = ~w23593 & ~w23594;
assign w23596 = pi03268 & ~w19773;
assign w23597 = ~pi02718 & w19773;
assign w23598 = ~w23596 & ~w23597;
assign w23599 = pi03269 & ~w19741;
assign w23600 = w17925 & w19740;
assign w23601 = ~w23599 & ~w23600;
assign w23602 = pi03270 & ~w19773;
assign w23603 = ~pi02167 & w19773;
assign w23604 = ~w23602 & ~w23603;
assign w23605 = pi03271 & ~w19741;
assign w23606 = ~pi02160 & w19741;
assign w23607 = ~w23605 & ~w23606;
assign w23608 = pi03272 & ~w19773;
assign w23609 = ~pi02164 & w19773;
assign w23610 = ~w23608 & ~w23609;
assign w23611 = pi03273 & ~w19741;
assign w23612 = ~pi02708 & w19741;
assign w23613 = ~w23611 & ~w23612;
assign w23614 = pi03274 & ~w19741;
assign w23615 = ~pi02709 & w19741;
assign w23616 = ~w23614 & ~w23615;
assign w23617 = pi03275 & ~w19773;
assign w23618 = w19130 & w19312;
assign w23619 = ~w23617 & ~w23618;
assign w23620 = pi03276 & ~w19741;
assign w23621 = ~pi02710 & w19741;
assign w23622 = ~w23620 & ~w23621;
assign w23623 = pi03277 & ~w19729;
assign w23624 = ~pi02705 & w19729;
assign w23625 = ~w23623 & ~w23624;
assign w23626 = pi03278 & ~w19773;
assign w23627 = ~pi02719 & w19773;
assign w23628 = ~w23626 & ~w23627;
assign w23629 = pi03279 & ~w19729;
assign w23630 = ~pi02706 & w19729;
assign w23631 = ~w23629 & ~w23630;
assign w23632 = pi03280 & ~w19729;
assign w23633 = ~pi02160 & w19729;
assign w23634 = ~w23632 & ~w23633;
assign w23635 = pi03281 & ~w19729;
assign w23636 = ~pi02723 & w19729;
assign w23637 = ~w23635 & ~w23636;
assign w23638 = pi03282 & ~w19729;
assign w23639 = ~pi02708 & w19729;
assign w23640 = ~w23638 & ~w23639;
assign w23641 = pi03283 & ~w19729;
assign w23642 = ~pi02710 & w19729;
assign w23643 = ~w23641 & ~w23642;
assign w23644 = pi03284 & ~w19724;
assign w23645 = ~pi02705 & w19724;
assign w23646 = ~w23644 & ~w23645;
assign w23647 = pi03285 & ~w19724;
assign w23648 = ~pi02706 & w19724;
assign w23649 = ~w23647 & ~w23648;
assign w23650 = pi03286 & ~w19724;
assign w23651 = ~pi02160 & w19724;
assign w23652 = ~w23650 & ~w23651;
assign w23653 = pi03287 & ~w19724;
assign w23654 = ~pi02723 & w19724;
assign w23655 = ~w23653 & ~w23654;
assign w23656 = pi03288 & ~w19724;
assign w23657 = ~pi02708 & w19724;
assign w23658 = ~w23656 & ~w23657;
assign w23659 = pi03289 & ~w19724;
assign w23660 = ~pi02709 & w19724;
assign w23661 = ~w23659 & ~w23660;
assign w23662 = pi03290 & ~w19724;
assign w23663 = ~pi02710 & w19724;
assign w23664 = ~w23662 & ~w23663;
assign w23665 = pi03291 & ~w19661;
assign w23666 = w18578 & w19660;
assign w23667 = ~w23665 & ~w23666;
assign w23668 = pi03292 & ~w19661;
assign w23669 = w17925 & w19660;
assign w23670 = ~w23668 & ~w23669;
assign w23671 = pi03293 & ~w19661;
assign w23672 = w18234 & w19660;
assign w23673 = ~w23671 & ~w23672;
assign w23674 = pi03294 & ~w19661;
assign w23675 = w17671 & w19660;
assign w23676 = ~w23674 & ~w23675;
assign w23677 = pi03295 & ~w19661;
assign w23678 = w18689 & w19660;
assign w23679 = ~w23677 & ~w23678;
assign w23680 = pi03296 & ~w19661;
assign w23681 = w18364 & w19660;
assign w23682 = ~w23680 & ~w23681;
assign w23683 = pi03297 & ~w19680;
assign w23684 = w18578 & w19679;
assign w23685 = ~w23683 & ~w23684;
assign w23686 = pi03298 & ~w19680;
assign w23687 = ~pi02706 & w19680;
assign w23688 = ~w23686 & ~w23687;
assign w23689 = pi03299 & ~w19680;
assign w23690 = ~pi02160 & w19680;
assign w23691 = ~w23689 & ~w23690;
assign w23692 = pi03300 & ~w19680;
assign w23693 = ~pi02723 & w19680;
assign w23694 = ~w23692 & ~w23693;
assign w23695 = pi03301 & ~w19680;
assign w23696 = ~pi02708 & w19680;
assign w23697 = ~w23695 & ~w23696;
assign w23698 = pi03302 & ~w19680;
assign w23699 = ~pi02709 & w19680;
assign w23700 = ~w23698 & ~w23699;
assign w23701 = pi03303 & ~w19680;
assign w23702 = ~pi02710 & w19680;
assign w23703 = ~w23701 & ~w23702;
assign w23704 = pi03304 & ~w19651;
assign w23705 = ~pi02705 & w19651;
assign w23706 = ~w23704 & ~w23705;
assign w23707 = pi03305 & ~w19651;
assign w23708 = ~pi02706 & w19651;
assign w23709 = ~w23707 & ~w23708;
assign w23710 = pi03306 & ~w19651;
assign w23711 = w18234 & w19650;
assign w23712 = ~w23710 & ~w23711;
assign w23713 = pi03307 & ~w19651;
assign w23714 = ~pi02723 & w19651;
assign w23715 = ~w23713 & ~w23714;
assign w23716 = pi03308 & ~w19651;
assign w23717 = ~pi02708 & w19651;
assign w23718 = ~w23716 & ~w23717;
assign w23719 = pi03309 & ~w19651;
assign w23720 = ~pi02710 & w19651;
assign w23721 = ~w23719 & ~w23720;
assign w23722 = pi03310 & ~w19646;
assign w23723 = ~pi02705 & w19646;
assign w23724 = ~w23722 & ~w23723;
assign w23725 = pi03311 & ~w19646;
assign w23726 = ~pi02706 & w19646;
assign w23727 = ~w23725 & ~w23726;
assign w23728 = pi03312 & ~w19646;
assign w23729 = w18234 & w19645;
assign w23730 = ~w23728 & ~w23729;
assign w23731 = pi03313 & ~w19646;
assign w23732 = ~pi02723 & w19646;
assign w23733 = ~w23731 & ~w23732;
assign w23734 = pi03314 & ~w19646;
assign w23735 = w18689 & w19645;
assign w23736 = ~w23734 & ~w23735;
assign w23737 = pi03315 & ~w19646;
assign w23738 = ~pi02709 & w19646;
assign w23739 = ~w23737 & ~w23738;
assign w23740 = pi03316 & ~w19646;
assign w23741 = ~pi02710 & w19646;
assign w23742 = ~w23740 & ~w23741;
assign w23743 = pi03317 & ~w19577;
assign w23744 = ~pi02705 & w19577;
assign w23745 = ~w23743 & ~w23744;
assign w23746 = pi03318 & ~w19577;
assign w23747 = ~pi02706 & w19577;
assign w23748 = ~w23746 & ~w23747;
assign w23749 = pi03319 & ~w19577;
assign w23750 = ~pi02160 & w19577;
assign w23751 = ~w23749 & ~w23750;
assign w23752 = pi03320 & ~w19577;
assign w23753 = ~pi02723 & w19577;
assign w23754 = ~w23752 & ~w23753;
assign w23755 = pi03321 & ~w19577;
assign w23756 = ~pi02708 & w19577;
assign w23757 = ~w23755 & ~w23756;
assign w23758 = pi03322 & ~w19577;
assign w23759 = ~pi02710 & w19577;
assign w23760 = ~w23758 & ~w23759;
assign w23761 = pi03323 & ~w19625;
assign w23762 = ~pi02705 & w19625;
assign w23763 = ~w23761 & ~w23762;
assign w23764 = pi03324 & ~w19167;
assign w23765 = ~pi09812 & w19167;
assign w23766 = ~w23764 & ~w23765;
assign w23767 = pi03325 & ~w21170;
assign w23768 = ~pi02712 & w21170;
assign w23769 = ~w23767 & ~w23768;
assign w23770 = pi03326 & ~w19625;
assign w23771 = ~pi02707 & w19625;
assign w23772 = ~w23770 & ~w23771;
assign w23773 = pi03327 & ~w19625;
assign w23774 = ~pi02160 & w19625;
assign w23775 = ~w23773 & ~w23774;
assign w23776 = pi03328 & ~w19625;
assign w23777 = ~pi02723 & w19625;
assign w23778 = ~w23776 & ~w23777;
assign w23779 = pi03329 & ~w19625;
assign w23780 = ~pi02708 & w19625;
assign w23781 = ~w23779 & ~w23780;
assign w23782 = pi03330 & ~w19625;
assign w23783 = ~pi02709 & w19625;
assign w23784 = ~w23782 & ~w23783;
assign w23785 = pi03331 & ~w19625;
assign w23786 = ~pi02710 & w19625;
assign w23787 = ~w23785 & ~w23786;
assign w23788 = pi03332 & ~w19607;
assign w23789 = ~pi02705 & w19607;
assign w23790 = ~w23788 & ~w23789;
assign w23791 = pi03333 & ~w19607;
assign w23792 = ~pi02707 & w19607;
assign w23793 = ~w23791 & ~w23792;
assign w23794 = pi03334 & ~w19607;
assign w23795 = ~pi02160 & w19607;
assign w23796 = ~w23794 & ~w23795;
assign w23797 = pi03335 & ~w19607;
assign w23798 = ~pi02723 & w19607;
assign w23799 = ~w23797 & ~w23798;
assign w23800 = pi03336 & ~w19607;
assign w23801 = ~pi02709 & w19607;
assign w23802 = ~w23800 & ~w23801;
assign w23803 = pi03337 & ~w19607;
assign w23804 = ~pi02710 & w19607;
assign w23805 = ~w23803 & ~w23804;
assign w23806 = pi03338 & ~w19602;
assign w23807 = ~pi02705 & w19602;
assign w23808 = ~w23806 & ~w23807;
assign w23809 = pi03339 & ~w19602;
assign w23810 = ~pi02707 & w19602;
assign w23811 = ~w23809 & ~w23810;
assign w23812 = pi03340 & ~w19602;
assign w23813 = w18234 & w19601;
assign w23814 = ~w23812 & ~w23813;
assign w23815 = pi03341 & ~w19602;
assign w23816 = ~pi02723 & w19602;
assign w23817 = ~w23815 & ~w23816;
assign w23818 = pi03342 & ~w19602;
assign w23819 = ~pi02708 & w19602;
assign w23820 = ~w23818 & ~w23819;
assign w23821 = pi03343 & ~w19602;
assign w23822 = ~pi02709 & w19602;
assign w23823 = ~w23821 & ~w23822;
assign w23824 = pi03344 & ~w19602;
assign w23825 = w18364 & w19601;
assign w23826 = ~w23824 & ~w23825;
assign w23827 = pi03345 & ~w19584;
assign w23828 = ~pi02703 & w19584;
assign w23829 = ~w23827 & ~w23828;
assign w23830 = pi03346 & ~w19584;
assign w23831 = ~pi02169 & w19584;
assign w23832 = ~w23830 & ~w23831;
assign w23833 = pi03347 & ~w19584;
assign w23834 = ~pi02718 & w19584;
assign w23835 = ~w23833 & ~w23834;
assign w23836 = pi03348 & ~w19584;
assign w23837 = ~pi02167 & w19584;
assign w23838 = ~w23836 & ~w23837;
assign w23839 = pi03349 & ~w19584;
assign w23840 = ~pi02722 & w19584;
assign w23841 = ~w23839 & ~w23840;
assign w23842 = pi03350 & ~w19584;
assign w23843 = ~pi02719 & w19584;
assign w23844 = ~w23842 & ~w23843;
assign w23845 = pi03351 & ~w19572;
assign w23846 = ~pi02703 & w19572;
assign w23847 = ~w23845 & ~w23846;
assign w23848 = pi03352 & ~w19572;
assign w23849 = ~pi02169 & w19572;
assign w23850 = ~w23848 & ~w23849;
assign w23851 = pi03353 & ~w19572;
assign w23852 = ~pi02718 & w19572;
assign w23853 = ~w23851 & ~w23852;
assign w23854 = pi03354 & ~w19572;
assign w23855 = ~pi02167 & w19572;
assign w23856 = ~w23854 & ~w23855;
assign w23857 = pi03355 & ~w19572;
assign w23858 = ~pi02164 & w19572;
assign w23859 = ~w23857 & ~w23858;
assign w23860 = pi03356 & ~w19572;
assign w23861 = ~pi02722 & w19572;
assign w23862 = ~w23860 & ~w23861;
assign w23863 = pi03357 & ~w19572;
assign w23864 = ~pi02719 & w19572;
assign w23865 = ~w23863 & ~w23864;
assign w23866 = pi03358 & ~w19562;
assign w23867 = ~pi02705 & w19562;
assign w23868 = ~w23866 & ~w23867;
assign w23869 = pi03359 & ~w19562;
assign w23870 = ~pi02707 & w19562;
assign w23871 = ~w23869 & ~w23870;
assign w23872 = pi03360 & ~w19562;
assign w23873 = w18234 & w19561;
assign w23874 = ~w23872 & ~w23873;
assign w23875 = pi03361 & ~w19562;
assign w23876 = ~pi02723 & w19562;
assign w23877 = ~w23875 & ~w23876;
assign w23878 = pi03362 & ~w19562;
assign w23879 = ~pi02708 & w19562;
assign w23880 = ~w23878 & ~w23879;
assign w23881 = pi03363 & ~w19562;
assign w23882 = ~pi02709 & w19562;
assign w23883 = ~w23881 & ~w23882;
assign w23884 = pi03364 & ~w19562;
assign w23885 = ~pi02710 & w19562;
assign w23886 = ~w23884 & ~w23885;
assign w23887 = pi03365 & ~w19557;
assign w23888 = ~pi02169 & w19557;
assign w23889 = ~w23887 & ~w23888;
assign w23890 = pi03366 & ~w19553;
assign w23891 = ~pi02705 & w19553;
assign w23892 = ~w23890 & ~w23891;
assign w23893 = pi03367 & ~w19557;
assign w23894 = ~pi02718 & w19557;
assign w23895 = ~w23893 & ~w23894;
assign w23896 = pi03368 & ~w19553;
assign w23897 = ~pi02706 & w19553;
assign w23898 = ~w23896 & ~w23897;
assign w23899 = pi03369 & ~w19553;
assign w23900 = ~pi02707 & w19553;
assign w23901 = ~w23899 & ~w23900;
assign w23902 = pi03370 & ~w19557;
assign w23903 = ~pi02167 & w19557;
assign w23904 = ~w23902 & ~w23903;
assign w23905 = pi03371 & ~w19553;
assign w23906 = ~pi02160 & w19553;
assign w23907 = ~w23905 & ~w23906;
assign w23908 = pi03372 & ~w19553;
assign w23909 = ~pi02723 & w19553;
assign w23910 = ~w23908 & ~w23909;
assign w23911 = pi03373 & ~w19557;
assign w23912 = ~pi02722 & w19557;
assign w23913 = ~w23911 & ~w23912;
assign w23914 = pi03374 & ~w19553;
assign w23915 = w18689 & w19552;
assign w23916 = ~w23914 & ~w23915;
assign w23917 = pi03375 & ~w19553;
assign w23918 = w18364 & w19552;
assign w23919 = ~w23917 & ~w23918;
assign w23920 = pi03376 & ~w19557;
assign w23921 = ~pi02719 & w19557;
assign w23922 = ~w23920 & ~w23921;
assign w23923 = pi03377 & ~w19436;
assign w23924 = ~pi02705 & w19436;
assign w23925 = ~w23923 & ~w23924;
assign w23926 = pi03378 & ~w19436;
assign w23927 = ~pi02707 & w19436;
assign w23928 = ~w23926 & ~w23927;
assign w23929 = pi03379 & ~w19436;
assign w23930 = ~pi02160 & w19436;
assign w23931 = ~w23929 & ~w23930;
assign w23932 = pi03380 & ~w19436;
assign w23933 = ~pi02723 & w19436;
assign w23934 = ~w23932 & ~w23933;
assign w23935 = pi03381 & ~w19436;
assign w23936 = ~pi02708 & w19436;
assign w23937 = ~w23935 & ~w23936;
assign w23938 = pi03382 & ~w19436;
assign w23939 = ~pi02709 & w19436;
assign w23940 = ~w23938 & ~w23939;
assign w23941 = pi03383 & ~w19436;
assign w23942 = ~pi02710 & w19436;
assign w23943 = ~w23941 & ~w23942;
assign w23944 = pi03384 & ~w19531;
assign w23945 = ~pi02705 & w19531;
assign w23946 = ~w23944 & ~w23945;
assign w23947 = pi03385 & ~w19531;
assign w23948 = ~pi02707 & w19531;
assign w23949 = ~w23947 & ~w23948;
assign w23950 = pi03386 & ~w19531;
assign w23951 = ~pi02160 & w19531;
assign w23952 = ~w23950 & ~w23951;
assign w23953 = pi03387 & ~w19531;
assign w23954 = ~pi02723 & w19531;
assign w23955 = ~w23953 & ~w23954;
assign w23956 = pi03388 & ~w19531;
assign w23957 = ~pi02709 & w19531;
assign w23958 = ~w23956 & ~w23957;
assign w23959 = pi03389 & ~w19531;
assign w23960 = ~pi02710 & w19531;
assign w23961 = ~w23959 & ~w23960;
assign w23962 = pi03390 & ~w19501;
assign w23963 = w17532 & w18995;
assign w23964 = ~w23962 & ~w23963;
assign w23965 = pi03391 & ~w19519;
assign w23966 = w17925 & w19518;
assign w23967 = ~w23965 & ~w23966;
assign w23968 = pi03392 & ~w19519;
assign w23969 = w18067 & w19518;
assign w23970 = ~w23968 & ~w23969;
assign w23971 = pi03393 & ~w19519;
assign w23972 = w18234 & w19518;
assign w23973 = ~w23971 & ~w23972;
assign w23974 = pi03394 & ~w19501;
assign w23975 = ~pi02721 & w19501;
assign w23976 = ~w23974 & ~w23975;
assign w23977 = pi03395 & ~w19519;
assign w23978 = w17671 & w19518;
assign w23979 = ~w23977 & ~w23978;
assign w23980 = pi03396 & ~w19519;
assign w23981 = w18689 & w19518;
assign w23982 = ~w23980 & ~w23981;
assign w23983 = pi03397 & ~w19519;
assign w23984 = w18092 & w19518;
assign w23985 = ~w23983 & ~w23984;
assign w23986 = pi03398 & ~w19519;
assign w23987 = w18364 & w19518;
assign w23988 = ~w23986 & ~w23987;
assign w23989 = pi03399 & ~w19501;
assign w23990 = ~pi02718 & w19501;
assign w23991 = ~w23989 & ~w23990;
assign w23992 = pi03400 & ~w19501;
assign w23993 = w18995 & w19273;
assign w23994 = ~w23992 & ~w23993;
assign w23995 = pi03401 & ~w19501;
assign w23996 = ~pi02722 & w19501;
assign w23997 = ~w23995 & ~w23996;
assign w23998 = pi03402 & ~w19501;
assign w23999 = w17594 & w18995;
assign w24000 = ~w23998 & ~w23999;
assign w24001 = pi03403 & ~w19416;
assign w24002 = ~pi02703 & w19416;
assign w24003 = ~w24001 & ~w24002;
assign w24004 = ~w16928 & w17837;
assign w24005 = pi03404 & ~w24004;
assign w24006 = ~pi09954 & w24004;
assign w24007 = ~w24005 & ~w24006;
assign w24008 = pi03405 & ~w19416;
assign w24009 = ~pi02169 & w19416;
assign w24010 = ~w24008 & ~w24009;
assign w24011 = pi03406 & ~w19416;
assign w24012 = ~pi02718 & w19416;
assign w24013 = ~w24011 & ~w24012;
assign w24014 = pi03407 & ~w19416;
assign w24015 = ~pi02167 & w19416;
assign w24016 = ~w24014 & ~w24015;
assign w24017 = pi03408 & ~w19416;
assign w24018 = ~pi02164 & w19416;
assign w24019 = ~w24017 & ~w24018;
assign w24020 = pi03409 & ~w19416;
assign w24021 = ~pi02722 & w19416;
assign w24022 = ~w24020 & ~w24021;
assign w24023 = pi03410 & ~w19493;
assign w24024 = ~pi02705 & w19493;
assign w24025 = ~w24023 & ~w24024;
assign w24026 = pi03411 & ~w19493;
assign w24027 = w17925 & w19492;
assign w24028 = ~w24026 & ~w24027;
assign w24029 = pi03412 & ~w19493;
assign w24030 = ~pi02707 & w19493;
assign w24031 = ~w24029 & ~w24030;
assign w24032 = pi03413 & ~w19493;
assign w24033 = ~pi02160 & w19493;
assign w24034 = ~w24032 & ~w24033;
assign w24035 = pi03414 & ~w19493;
assign w24036 = ~pi02723 & w19493;
assign w24037 = ~w24035 & ~w24036;
assign w24038 = pi03415 & ~w19493;
assign w24039 = ~pi02709 & w19493;
assign w24040 = ~w24038 & ~w24039;
assign w24041 = pi03416 & ~w19493;
assign w24042 = w18364 & w19492;
assign w24043 = ~w24041 & ~w24042;
assign w24044 = pi03417 & ~w19481;
assign w24045 = ~pi02705 & w19481;
assign w24046 = ~w24044 & ~w24045;
assign w24047 = pi03418 & ~w19481;
assign w24048 = ~pi02707 & w19481;
assign w24049 = ~w24047 & ~w24048;
assign w24050 = pi03419 & ~w19481;
assign w24051 = ~pi02160 & w19481;
assign w24052 = ~w24050 & ~w24051;
assign w24053 = pi03420 & ~w19481;
assign w24054 = ~pi02723 & w19481;
assign w24055 = ~w24053 & ~w24054;
assign w24056 = pi03421 & ~w19481;
assign w24057 = ~pi02708 & w19481;
assign w24058 = ~w24056 & ~w24057;
assign w24059 = pi03422 & ~w19481;
assign w24060 = ~pi02709 & w19481;
assign w24061 = ~w24059 & ~w24060;
assign w24062 = pi03423 & ~w19481;
assign w24063 = w18364 & w19480;
assign w24064 = ~w24062 & ~w24063;
assign w24065 = pi03424 & ~w19460;
assign w24066 = ~pi02705 & w19460;
assign w24067 = ~w24065 & ~w24066;
assign w24068 = pi03425 & ~w19460;
assign w24069 = ~pi02707 & w19460;
assign w24070 = ~w24068 & ~w24069;
assign w24071 = pi03426 & ~w19460;
assign w24072 = ~pi02160 & w19460;
assign w24073 = ~w24071 & ~w24072;
assign w24074 = pi03427 & ~w19460;
assign w24075 = ~pi02723 & w19460;
assign w24076 = ~w24074 & ~w24075;
assign w24077 = pi03428 & ~w19460;
assign w24078 = ~pi02709 & w19460;
assign w24079 = ~w24077 & ~w24078;
assign w24080 = pi03429 & ~w19460;
assign w24081 = ~pi02710 & w19460;
assign w24082 = ~w24080 & ~w24081;
assign w24083 = pi03430 & ~w19421;
assign w24084 = w18578 & w19420;
assign w24085 = ~w24083 & ~w24084;
assign w24086 = pi03431 & ~w19421;
assign w24087 = ~pi02707 & w19421;
assign w24088 = ~w24086 & ~w24087;
assign w24089 = pi03432 & ~w19421;
assign w24090 = ~pi02160 & w19421;
assign w24091 = ~w24089 & ~w24090;
assign w24092 = pi03433 & ~w19421;
assign w24093 = ~pi02723 & w19421;
assign w24094 = ~w24092 & ~w24093;
assign w24095 = pi03434 & ~w19421;
assign w24096 = ~pi02708 & w19421;
assign w24097 = ~w24095 & ~w24096;
assign w24098 = pi03435 & ~w19421;
assign w24099 = ~pi02709 & w19421;
assign w24100 = ~w24098 & ~w24099;
assign w24101 = pi03436 & ~w19421;
assign w24102 = ~pi02710 & w19421;
assign w24103 = ~w24101 & ~w24102;
assign w24104 = pi03437 & ~w19445;
assign w24105 = ~pi02705 & w19445;
assign w24106 = ~w24104 & ~w24105;
assign w24107 = pi03438 & ~w19445;
assign w24108 = ~pi02707 & w19445;
assign w24109 = ~w24107 & ~w24108;
assign w24110 = pi03439 & ~w19445;
assign w24111 = ~pi02160 & w19445;
assign w24112 = ~w24110 & ~w24111;
assign w24113 = pi03440 & ~w19445;
assign w24114 = ~pi02723 & w19445;
assign w24115 = ~w24113 & ~w24114;
assign w24116 = pi03441 & ~w19445;
assign w24117 = ~pi02709 & w19445;
assign w24118 = ~w24116 & ~w24117;
assign w24119 = pi03442 & ~w19445;
assign w24120 = ~pi02710 & w19445;
assign w24121 = ~w24119 & ~w24120;
assign w24122 = pi03443 & ~w19328;
assign w24123 = ~pi02705 & w19328;
assign w24124 = ~w24122 & ~w24123;
assign w24125 = pi03444 & ~w19328;
assign w24126 = ~pi02707 & w19328;
assign w24127 = ~w24125 & ~w24126;
assign w24128 = pi03445 & ~w19328;
assign w24129 = ~pi02160 & w19328;
assign w24130 = ~w24128 & ~w24129;
assign w24131 = pi03446 & ~w19388;
assign w24132 = ~pi02703 & w19388;
assign w24133 = ~w24131 & ~w24132;
assign w24134 = pi03447 & ~w19328;
assign w24135 = ~pi02723 & w19328;
assign w24136 = ~w24134 & ~w24135;
assign w24137 = pi03448 & ~w19328;
assign w24138 = ~pi02708 & w19328;
assign w24139 = ~w24137 & ~w24138;
assign w24140 = pi03449 & ~w19328;
assign w24141 = ~pi02709 & w19328;
assign w24142 = ~w24140 & ~w24141;
assign w24143 = pi03450 & ~w19388;
assign w24144 = ~pi02721 & w19388;
assign w24145 = ~w24143 & ~w24144;
assign w24146 = pi03451 & ~w19388;
assign w24147 = ~pi02169 & w19388;
assign w24148 = ~w24146 & ~w24147;
assign w24149 = pi03452 & ~w19388;
assign w24150 = ~pi02718 & w19388;
assign w24151 = ~w24149 & ~w24150;
assign w24152 = pi03453 & ~w19388;
assign w24153 = ~pi02167 & w19388;
assign w24154 = ~w24152 & ~w24153;
assign w24155 = ~w16892 & w19591;
assign w24156 = pi03454 & ~w24155;
assign w24157 = ~pi02705 & w24155;
assign w24158 = ~w24156 & ~w24157;
assign w24159 = pi03455 & ~w24155;
assign w24160 = ~pi02706 & w24155;
assign w24161 = ~w24159 & ~w24160;
assign w24162 = pi03456 & ~w19388;
assign w24163 = ~pi02722 & w19388;
assign w24164 = ~w24162 & ~w24163;
assign w24165 = pi03457 & ~w24155;
assign w24166 = ~pi02707 & w24155;
assign w24167 = ~w24165 & ~w24166;
assign w24168 = pi03458 & ~w24155;
assign w24169 = ~pi02160 & w24155;
assign w24170 = ~w24168 & ~w24169;
assign w24171 = pi03459 & ~w24155;
assign w24172 = ~pi02723 & w24155;
assign w24173 = ~w24171 & ~w24172;
assign w24174 = pi03460 & ~w24155;
assign w24175 = ~pi02708 & w24155;
assign w24176 = ~w24174 & ~w24175;
assign w24177 = pi03461 & ~w24155;
assign w24178 = ~pi02709 & w24155;
assign w24179 = ~w24177 & ~w24178;
assign w24180 = pi03462 & ~w24155;
assign w24181 = ~pi02710 & w24155;
assign w24182 = ~w24180 & ~w24181;
assign w24183 = pi03463 & ~w19384;
assign w24184 = ~pi02705 & w19384;
assign w24185 = ~w24183 & ~w24184;
assign w24186 = pi03464 & ~w19384;
assign w24187 = ~pi02707 & w19384;
assign w24188 = ~w24186 & ~w24187;
assign w24189 = pi03465 & ~w19384;
assign w24190 = ~pi02160 & w19384;
assign w24191 = ~w24189 & ~w24190;
assign w24192 = pi03466 & ~w19384;
assign w24193 = ~pi02723 & w19384;
assign w24194 = ~w24192 & ~w24193;
assign w24195 = pi03467 & ~w19384;
assign w24196 = ~pi02709 & w19384;
assign w24197 = ~w24195 & ~w24196;
assign w24198 = pi03468 & ~w19384;
assign w24199 = ~pi02710 & w19384;
assign w24200 = ~w24198 & ~w24199;
assign w24201 = pi03469 & ~w19375;
assign w24202 = ~pi02705 & w19375;
assign w24203 = ~w24201 & ~w24202;
assign w24204 = pi03470 & ~w19375;
assign w24205 = ~pi02707 & w19375;
assign w24206 = ~w24204 & ~w24205;
assign w24207 = pi03471 & ~w19375;
assign w24208 = w18234 & w19374;
assign w24209 = ~w24207 & ~w24208;
assign w24210 = pi03472 & ~w19359;
assign w24211 = ~pi02703 & w19359;
assign w24212 = ~w24210 & ~w24211;
assign w24213 = pi03473 & ~w19375;
assign w24214 = ~pi02723 & w19375;
assign w24215 = ~w24213 & ~w24214;
assign w24216 = pi03474 & ~w19375;
assign w24217 = ~pi02708 & w19375;
assign w24218 = ~w24216 & ~w24217;
assign w24219 = pi03475 & ~w19375;
assign w24220 = ~pi02709 & w19375;
assign w24221 = ~w24219 & ~w24220;
assign w24222 = pi03476 & ~w19375;
assign w24223 = ~pi02710 & w19375;
assign w24224 = ~w24222 & ~w24223;
assign w24225 = pi03477 & ~w19359;
assign w24226 = ~pi02721 & w19359;
assign w24227 = ~w24225 & ~w24226;
assign w24228 = pi03478 & ~w19349;
assign w24229 = ~pi02706 & w19349;
assign w24230 = ~w24228 & ~w24229;
assign w24231 = pi03479 & ~w19359;
assign w24232 = ~pi02169 & w19359;
assign w24233 = ~w24231 & ~w24232;
assign w24234 = pi03480 & ~w19359;
assign w24235 = ~pi02718 & w19359;
assign w24236 = ~w24234 & ~w24235;
assign w24237 = pi03481 & ~w19349;
assign w24238 = ~pi02160 & w19349;
assign w24239 = ~w24237 & ~w24238;
assign w24240 = pi03482 & ~w19349;
assign w24241 = ~pi02723 & w19349;
assign w24242 = ~w24240 & ~w24241;
assign w24243 = ~w16928 & w17114;
assign w24244 = pi03483 & ~w24243;
assign w24245 = ~pi09812 & w24243;
assign w24246 = ~w24244 & ~w24245;
assign w24247 = pi03484 & ~w19349;
assign w24248 = ~pi02708 & w19349;
assign w24249 = ~w24247 & ~w24248;
assign w24250 = pi03485 & ~w19349;
assign w24251 = ~pi02709 & w19349;
assign w24252 = ~w24250 & ~w24251;
assign w24253 = pi03486 & ~w19349;
assign w24254 = ~pi02710 & w19349;
assign w24255 = ~w24253 & ~w24254;
assign w24256 = pi03487 & ~w19359;
assign w24257 = w17620 & w18986;
assign w24258 = ~w24256 & ~w24257;
assign w24259 = pi03488 & ~w19359;
assign w24260 = ~pi02722 & w19359;
assign w24261 = ~w24259 & ~w24260;
assign w24262 = pi03489 & ~w19359;
assign w24263 = ~pi02719 & w19359;
assign w24264 = ~w24262 & ~w24263;
assign w24265 = pi03490 & ~w19339;
assign w24266 = ~pi02703 & w19339;
assign w24267 = ~w24265 & ~w24266;
assign w24268 = pi03491 & ~w19339;
assign w24269 = ~pi02169 & w19339;
assign w24270 = ~w24268 & ~w24269;
assign w24271 = pi03492 & ~w19339;
assign w24272 = w17586 & w18925;
assign w24273 = ~w24271 & ~w24272;
assign w24274 = pi03493 & ~w19339;
assign w24275 = ~pi02167 & w19339;
assign w24276 = ~w24274 & ~w24275;
assign w24277 = pi03494 & ~w19339;
assign w24278 = w18925 & w19312;
assign w24279 = ~w24277 & ~w24278;
assign w24280 = pi03495 & ~w19339;
assign w24281 = ~pi02719 & w19339;
assign w24282 = ~w24280 & ~w24281;
assign w24283 = pi03496 & ~w19344;
assign w24284 = ~pi02705 & w19344;
assign w24285 = ~w24283 & ~w24284;
assign w24286 = pi03497 & ~w19344;
assign w24287 = ~pi02707 & w19344;
assign w24288 = ~w24286 & ~w24287;
assign w24289 = pi03498 & ~w19344;
assign w24290 = ~pi02160 & w19344;
assign w24291 = ~w24289 & ~w24290;
assign w24292 = pi03499 & ~w19344;
assign w24293 = ~pi02723 & w19344;
assign w24294 = ~w24292 & ~w24293;
assign w24295 = pi03500 & ~w19344;
assign w24296 = w18689 & w19343;
assign w24297 = ~w24295 & ~w24296;
assign w24298 = pi03501 & ~w19344;
assign w24299 = ~pi02709 & w19344;
assign w24300 = ~w24298 & ~w24299;
assign w24301 = pi03502 & ~w19344;
assign w24302 = ~pi02710 & w19344;
assign w24303 = ~w24301 & ~w24302;
assign w24304 = pi03503 & ~w19298;
assign w24305 = w17532 & w18944;
assign w24306 = ~w24304 & ~w24305;
assign w24307 = pi03504 & ~w19319;
assign w24308 = ~pi02712 & w19319;
assign w24309 = ~w24307 & ~w24308;
assign w24310 = pi03505 & ~w19298;
assign w24311 = w17811 & w18944;
assign w24312 = ~w24310 & ~w24311;
assign w24313 = pi03506 & ~w19319;
assign w24314 = ~pi02170 & w19319;
assign w24315 = ~w24313 & ~w24314;
assign w24316 = pi03507 & ~w19319;
assign w24317 = ~pi02713 & w19319;
assign w24318 = ~w24316 & ~w24317;
assign w24319 = pi03508 & ~w19298;
assign w24320 = ~pi02718 & w19298;
assign w24321 = ~w24319 & ~w24320;
assign w24322 = pi03509 & ~w19319;
assign w24323 = ~pi02714 & w19319;
assign w24324 = ~w24322 & ~w24323;
assign w24325 = pi03510 & ~w19298;
assign w24326 = ~pi02167 & w19298;
assign w24327 = ~w24325 & ~w24326;
assign w24328 = pi03511 & ~w19319;
assign w24329 = ~pi02716 & w19319;
assign w24330 = ~w24328 & ~w24329;
assign w24331 = pi03512 & ~w19319;
assign w24332 = ~pi02717 & w19319;
assign w24333 = ~w24331 & ~w24332;
assign w24334 = pi03513 & ~w19315;
assign w24335 = ~pi02711 & w19315;
assign w24336 = ~w24334 & ~w24335;
assign w24337 = pi03514 & ~w19298;
assign w24338 = ~pi02164 & w19298;
assign w24339 = ~w24337 & ~w24338;
assign w24340 = pi03515 & ~w19315;
assign w24341 = ~pi02712 & w19315;
assign w24342 = ~w24340 & ~w24341;
assign w24343 = pi03516 & ~w19315;
assign w24344 = ~pi02170 & w19315;
assign w24345 = ~w24343 & ~w24344;
assign w24346 = pi03517 & ~w19315;
assign w24347 = ~pi02713 & w19315;
assign w24348 = ~w24346 & ~w24347;
assign w24349 = pi03518 & ~w19315;
assign w24350 = ~pi02714 & w19315;
assign w24351 = ~w24349 & ~w24350;
assign w24352 = pi03519 & ~w19298;
assign w24353 = ~pi02719 & w19298;
assign w24354 = ~w24352 & ~w24353;
assign w24355 = pi03520 & ~w19315;
assign w24356 = ~pi02716 & w19315;
assign w24357 = ~w24355 & ~w24356;
assign w24358 = pi03521 & ~w19302;
assign w24359 = ~pi02703 & w19302;
assign w24360 = ~w24358 & ~w24359;
assign w24361 = pi03522 & ~w19315;
assign w24362 = ~pi02717 & w19315;
assign w24363 = ~w24361 & ~w24362;
assign w24364 = pi03523 & ~w19302;
assign w24365 = ~pi02169 & w19302;
assign w24366 = ~w24364 & ~w24365;
assign w24367 = pi03524 & ~w19302;
assign w24368 = ~pi02718 & w19302;
assign w24369 = ~w24367 & ~w24368;
assign w24370 = pi03525 & ~w19302;
assign w24371 = ~pi02167 & w19302;
assign w24372 = ~w24370 & ~w24371;
assign w24373 = pi03526 & ~w19302;
assign w24374 = w17620 & w18913;
assign w24375 = ~w24373 & ~w24374;
assign w24376 = pi03527 & ~w19302;
assign w24377 = ~pi02722 & w19302;
assign w24378 = ~w24376 & ~w24377;
assign w24379 = pi03528 & ~w19302;
assign w24380 = w17594 & w18913;
assign w24381 = ~w24379 & ~w24380;
assign w24382 = pi03529 & ~w19287;
assign w24383 = ~pi02711 & w19287;
assign w24384 = ~w24382 & ~w24383;
assign w24385 = pi03530 & ~w19287;
assign w24386 = ~pi02170 & w19287;
assign w24387 = ~w24385 & ~w24386;
assign w24388 = pi03531 & ~w19287;
assign w24389 = ~pi02713 & w19287;
assign w24390 = ~w24388 & ~w24389;
assign w24391 = pi03532 & ~w19287;
assign w24392 = ~pi02714 & w19287;
assign w24393 = ~w24391 & ~w24392;
assign w24394 = pi03533 & ~w19287;
assign w24395 = ~pi02716 & w19287;
assign w24396 = ~w24394 & ~w24395;
assign w24397 = pi03534 & ~w19287;
assign w24398 = ~pi02717 & w19287;
assign w24399 = ~w24397 & ~w24398;
assign w24400 = pi03535 & ~w19291;
assign w24401 = ~pi02711 & w19291;
assign w24402 = ~w24400 & ~w24401;
assign w24403 = ~w16928 & w18001;
assign w24404 = pi03536 & ~w24403;
assign w24405 = w18001 & w19365;
assign w24406 = ~w24404 & ~w24405;
assign w24407 = pi03537 & ~w19291;
assign w24408 = ~pi02170 & w19291;
assign w24409 = ~w24407 & ~w24408;
assign w24410 = pi03538 & ~w19291;
assign w24411 = ~pi02713 & w19291;
assign w24412 = ~w24410 & ~w24411;
assign w24413 = pi03539 & ~w19291;
assign w24414 = ~pi02714 & w19291;
assign w24415 = ~w24413 & ~w24414;
assign w24416 = pi03540 & ~w19291;
assign w24417 = ~pi02715 & w19291;
assign w24418 = ~w24416 & ~w24417;
assign w24419 = pi03541 & ~w19291;
assign w24420 = ~pi02716 & w19291;
assign w24421 = ~w24419 & ~w24420;
assign w24422 = pi03542 & ~w19271;
assign w24423 = ~pi02703 & w19271;
assign w24424 = ~w24422 & ~w24423;
assign w24425 = pi03543 & ~w19291;
assign w24426 = ~pi02717 & w19291;
assign w24427 = ~w24425 & ~w24426;
assign w24428 = pi03544 & ~w19271;
assign w24429 = ~pi02169 & w19271;
assign w24430 = ~w24428 & ~w24429;
assign w24431 = pi03545 & ~w19271;
assign w24432 = ~pi02718 & w19271;
assign w24433 = ~w24431 & ~w24432;
assign w24434 = pi03546 & ~w19253;
assign w24435 = ~pi02711 & w19253;
assign w24436 = ~w24434 & ~w24435;
assign w24437 = pi03547 & ~w19253;
assign w24438 = w17020 & w17131;
assign w24439 = ~w24437 & ~w24438;
assign w24440 = pi03548 & ~w19271;
assign w24441 = ~pi02164 & w19271;
assign w24442 = ~w24440 & ~w24441;
assign w24443 = pi03549 & ~w19253;
assign w24444 = ~pi02170 & w19253;
assign w24445 = ~w24443 & ~w24444;
assign w24446 = pi03550 & ~w19271;
assign w24447 = ~pi02722 & w19271;
assign w24448 = ~w24446 & ~w24447;
assign w24449 = pi03551 & ~w19253;
assign w24450 = ~pi02714 & w19253;
assign w24451 = ~w24449 & ~w24450;
assign w24452 = pi03552 & ~w19271;
assign w24453 = ~pi02719 & w19271;
assign w24454 = ~w24452 & ~w24453;
assign w24455 = pi03553 & ~w19253;
assign w24456 = ~pi02715 & w19253;
assign w24457 = ~w24455 & ~w24456;
assign w24458 = pi03554 & ~w19253;
assign w24459 = ~pi02716 & w19253;
assign w24460 = ~w24458 & ~w24459;
assign w24461 = pi03555 & ~w19253;
assign w24462 = ~pi02717 & w19253;
assign w24463 = ~w24461 & ~w24462;
assign w24464 = pi03556 & ~w19242;
assign w24465 = w17060 & w17603;
assign w24466 = ~w24464 & ~w24465;
assign w24467 = pi03557 & ~w19242;
assign w24468 = w17060 & w20209;
assign w24469 = ~w24467 & ~w24468;
assign w24470 = pi03558 & ~w19242;
assign w24471 = w17060 & w17929;
assign w24472 = ~w24470 & ~w24471;
assign w24473 = pi03559 & ~w19242;
assign w24474 = w17060 & w17742;
assign w24475 = ~w24473 & ~w24474;
assign w24476 = pi03560 & ~w19242;
assign w24477 = ~pi02716 & w19242;
assign w24478 = ~w24476 & ~w24477;
assign w24479 = pi03561 & ~w19242;
assign w24480 = w16973 & w17060;
assign w24481 = ~w24479 & ~w24480;
assign w24482 = pi03562 & ~w19238;
assign w24483 = ~pi02711 & w19238;
assign w24484 = ~w24482 & ~w24483;
assign w24485 = pi03563 & ~w19228;
assign w24486 = ~pi02703 & w19228;
assign w24487 = ~w24485 & ~w24486;
assign w24488 = pi03564 & ~w19238;
assign w24489 = w19106 & w20209;
assign w24490 = ~w24488 & ~w24489;
assign w24491 = pi03565 & ~w19228;
assign w24492 = ~pi02721 & w19228;
assign w24493 = ~w24491 & ~w24492;
assign w24494 = pi03566 & ~w19238;
assign w24495 = ~pi02713 & w19238;
assign w24496 = ~w24494 & ~w24495;
assign w24497 = pi03567 & ~w19228;
assign w24498 = ~pi02169 & w19228;
assign w24499 = ~w24497 & ~w24498;
assign w24500 = pi03568 & ~w19238;
assign w24501 = w17742 & w19106;
assign w24502 = ~w24500 & ~w24501;
assign w24503 = pi03569 & ~w19238;
assign w24504 = w18059 & w19106;
assign w24505 = ~w24503 & ~w24504;
assign w24506 = pi03570 & ~w19238;
assign w24507 = w17317 & w19106;
assign w24508 = ~w24506 & ~w24507;
assign w24509 = pi03571 & ~w19238;
assign w24510 = ~pi02717 & w19238;
assign w24511 = ~w24509 & ~w24510;
assign w24512 = pi03572 & ~w19228;
assign w24513 = ~pi02167 & w19228;
assign w24514 = ~w24512 & ~w24513;
assign w24515 = pi03573 & ~w19228;
assign w24516 = ~pi02722 & w19228;
assign w24517 = ~w24515 & ~w24516;
assign w24518 = pi03574 & ~w19228;
assign w24519 = ~pi02719 & w19228;
assign w24520 = ~w24518 & ~w24519;
assign w24521 = pi03575 & ~w19224;
assign w24522 = ~pi02711 & w19224;
assign w24523 = ~w24521 & ~w24522;
assign w24524 = pi03576 & ~w19224;
assign w24525 = ~pi02170 & w19224;
assign w24526 = ~w24524 & ~w24525;
assign w24527 = pi03577 & ~w19224;
assign w24528 = ~pi02713 & w19224;
assign w24529 = ~w24527 & ~w24528;
assign w24530 = pi03578 & ~w19224;
assign w24531 = ~pi02714 & w19224;
assign w24532 = ~w24530 & ~w24531;
assign w24533 = pi03579 & ~w19224;
assign w24534 = ~pi02715 & w19224;
assign w24535 = ~w24533 & ~w24534;
assign w24536 = pi03580 & ~w19224;
assign w24537 = ~pi02716 & w19224;
assign w24538 = ~w24536 & ~w24537;
assign w24539 = pi03581 & ~w19224;
assign w24540 = ~pi02717 & w19224;
assign w24541 = ~w24539 & ~w24540;
assign w24542 = pi03582 & ~w19217;
assign w24543 = ~pi02703 & w19217;
assign w24544 = ~w24542 & ~w24543;
assign w24545 = pi03583 & ~w19217;
assign w24546 = ~pi02169 & w19217;
assign w24547 = ~w24545 & ~w24546;
assign w24548 = pi03584 & ~w19192;
assign w24549 = ~pi02711 & w19192;
assign w24550 = ~w24548 & ~w24549;
assign w24551 = pi03585 & ~w19217;
assign w24552 = ~pi02718 & w19217;
assign w24553 = ~w24551 & ~w24552;
assign w24554 = pi03586 & ~w19192;
assign w24555 = ~pi02170 & w19192;
assign w24556 = ~w24554 & ~w24555;
assign w24557 = pi03587 & ~w19217;
assign w24558 = ~pi02167 & w19217;
assign w24559 = ~w24557 & ~w24558;
assign w24560 = pi03588 & ~w19192;
assign w24561 = ~pi02713 & w19192;
assign w24562 = ~w24560 & ~w24561;
assign w24563 = pi03589 & ~w19217;
assign w24564 = w17620 & w18831;
assign w24565 = ~w24563 & ~w24564;
assign w24566 = pi03590 & ~w19192;
assign w24567 = ~pi02715 & w19192;
assign w24568 = ~w24566 & ~w24567;
assign w24569 = pi03591 & ~w19217;
assign w24570 = ~pi02722 & w19217;
assign w24571 = ~w24569 & ~w24570;
assign w24572 = pi03592 & ~w19192;
assign w24573 = ~pi02716 & w19192;
assign w24574 = ~w24572 & ~w24573;
assign w24575 = pi03593 & ~w19217;
assign w24576 = ~pi02719 & w19217;
assign w24577 = ~w24575 & ~w24576;
assign w24578 = pi03594 & ~w19192;
assign w24579 = ~pi02717 & w19192;
assign w24580 = ~w24578 & ~w24579;
assign w24581 = pi03595 & ~w19206;
assign w24582 = ~pi02711 & w19206;
assign w24583 = ~w24581 & ~w24582;
assign w24584 = pi03596 & ~w19188;
assign w24585 = ~pi02703 & w19188;
assign w24586 = ~w24584 & ~w24585;
assign w24587 = pi03597 & ~w19206;
assign w24588 = ~pi02170 & w19206;
assign w24589 = ~w24587 & ~w24588;
assign w24590 = pi03598 & ~w19206;
assign w24591 = ~pi02713 & w19206;
assign w24592 = ~w24590 & ~w24591;
assign w24593 = pi03599 & ~w19206;
assign w24594 = ~pi02714 & w19206;
assign w24595 = ~w24593 & ~w24594;
assign w24596 = pi03600 & ~w19206;
assign w24597 = ~pi02715 & w19206;
assign w24598 = ~w24596 & ~w24597;
assign w24599 = pi03601 & ~w19206;
assign w24600 = ~pi02716 & w19206;
assign w24601 = ~w24599 & ~w24600;
assign w24602 = pi03602 & ~w19206;
assign w24603 = ~pi02717 & w19206;
assign w24604 = ~w24602 & ~w24603;
assign w24605 = pi03603 & ~w19188;
assign w24606 = ~pi02718 & w19188;
assign w24607 = ~w24605 & ~w24606;
assign w24608 = pi03604 & ~w19188;
assign w24609 = ~pi02167 & w19188;
assign w24610 = ~w24608 & ~w24609;
assign w24611 = pi03605 & ~w19188;
assign w24612 = ~pi02164 & w19188;
assign w24613 = ~w24611 & ~w24612;
assign w24614 = pi03606 & ~w19188;
assign w24615 = ~pi02722 & w19188;
assign w24616 = ~w24614 & ~w24615;
assign w24617 = pi03607 & ~w19188;
assign w24618 = ~pi02719 & w19188;
assign w24619 = ~w24617 & ~w24618;
assign w24620 = pi03608 & ~w19162;
assign w24621 = ~pi02703 & w19162;
assign w24622 = ~w24620 & ~w24621;
assign w24623 = pi03609 & ~w19162;
assign w24624 = ~pi02169 & w19162;
assign w24625 = ~w24623 & ~w24624;
assign w24626 = pi03610 & ~w19162;
assign w24627 = w17586 & w18612;
assign w24628 = ~w24626 & ~w24627;
assign w24629 = pi03611 & ~w19162;
assign w24630 = ~pi02167 & w19162;
assign w24631 = ~w24629 & ~w24630;
assign w24632 = pi03612 & ~w19162;
assign w24633 = w18612 & w19312;
assign w24634 = ~w24632 & ~w24633;
assign w24635 = pi03613 & ~w19162;
assign w24636 = ~pi02719 & w19162;
assign w24637 = ~w24635 & ~w24636;
assign w24638 = pi03614 & ~w19181;
assign w24639 = ~pi02703 & w19181;
assign w24640 = ~w24638 & ~w24639;
assign w24641 = pi03615 & ~w19181;
assign w24642 = w17516 & w19797;
assign w24643 = ~w24641 & ~w24642;
assign w24644 = pi03616 & ~w19181;
assign w24645 = ~pi02718 & w19181;
assign w24646 = ~w24644 & ~w24645;
assign w24647 = pi03617 & ~w19181;
assign w24648 = ~pi02167 & w19181;
assign w24649 = ~w24647 & ~w24648;
assign w24650 = pi03618 & ~w19181;
assign w24651 = ~pi02164 & w19181;
assign w24652 = ~w24650 & ~w24651;
assign w24653 = pi03619 & ~w19181;
assign w24654 = ~pi02722 & w19181;
assign w24655 = ~w24653 & ~w24654;
assign w24656 = pi03620 & ~w19181;
assign w24657 = ~pi02719 & w19181;
assign w24658 = ~w24656 & ~w24657;
assign w24659 = pi03621 & ~w19158;
assign w24660 = ~pi02703 & w19158;
assign w24661 = ~w24659 & ~w24660;
assign w24662 = pi03622 & ~w19158;
assign w24663 = ~pi02169 & w19158;
assign w24664 = ~w24662 & ~w24663;
assign w24665 = pi03623 & ~w19158;
assign w24666 = ~pi02718 & w19158;
assign w24667 = ~w24665 & ~w24666;
assign w24668 = pi03624 & ~w19158;
assign w24669 = ~pi02167 & w19158;
assign w24670 = ~w24668 & ~w24669;
assign w24671 = pi03625 & ~w19158;
assign w24672 = w18431 & w19312;
assign w24673 = ~w24671 & ~w24672;
assign w24674 = pi03626 & ~w19158;
assign w24675 = ~pi02719 & w19158;
assign w24676 = ~w24674 & ~w24675;
assign w24677 = pi03627 & ~w19017;
assign w24678 = ~pi02703 & w19017;
assign w24679 = ~w24677 & ~w24678;
assign w24680 = pi03628 & ~w19017;
assign w24681 = w18247 & w19797;
assign w24682 = ~w24680 & ~w24681;
assign w24683 = pi03629 & ~w19017;
assign w24684 = ~pi02718 & w19017;
assign w24685 = ~w24683 & ~w24684;
assign w24686 = pi03630 & ~w19017;
assign w24687 = ~pi02167 & w19017;
assign w24688 = ~w24686 & ~w24687;
assign w24689 = pi03631 & ~w19017;
assign w24690 = ~pi02164 & w19017;
assign w24691 = ~w24689 & ~w24690;
assign w24692 = pi03632 & ~w19017;
assign w24693 = ~pi02722 & w19017;
assign w24694 = ~w24692 & ~w24693;
assign w24695 = pi03633 & ~w19017;
assign w24696 = ~pi02719 & w19017;
assign w24697 = ~w24695 & ~w24696;
assign w24698 = pi03634 & ~w19120;
assign w24699 = ~pi02703 & w19120;
assign w24700 = ~w24698 & ~w24699;
assign w24701 = pi03635 & ~w19120;
assign w24702 = ~pi02169 & w19120;
assign w24703 = ~w24701 & ~w24702;
assign w24704 = pi03636 & ~w19120;
assign w24705 = ~pi02718 & w19120;
assign w24706 = ~w24704 & ~w24705;
assign w24707 = pi03637 & ~w19120;
assign w24708 = w17510 & w19273;
assign w24709 = ~w24707 & ~w24708;
assign w24710 = ~w16905 & w19115;
assign w24711 = pi03638 & ~w24710;
assign w24712 = w17603 & w19115;
assign w24713 = ~w24711 & ~w24712;
assign w24714 = pi03639 & ~w24710;
assign w24715 = ~pi02712 & w24710;
assign w24716 = ~w24714 & ~w24715;
assign w24717 = pi03640 & ~w19120;
assign w24718 = ~pi02722 & w19120;
assign w24719 = ~w24717 & ~w24718;
assign w24720 = pi03641 & ~w24710;
assign w24721 = ~pi02170 & w24710;
assign w24722 = ~w24720 & ~w24721;
assign w24723 = pi03642 & ~w24710;
assign w24724 = ~pi02713 & w24710;
assign w24725 = ~w24723 & ~w24724;
assign w24726 = pi03643 & ~w24710;
assign w24727 = ~pi02714 & w24710;
assign w24728 = ~w24726 & ~w24727;
assign w24729 = pi03644 & ~w24710;
assign w24730 = ~pi02715 & w24710;
assign w24731 = ~w24729 & ~w24730;
assign w24732 = pi03645 & ~w24710;
assign w24733 = ~pi02716 & w24710;
assign w24734 = ~w24732 & ~w24733;
assign w24735 = pi03646 & ~w24710;
assign w24736 = ~pi02717 & w24710;
assign w24737 = ~w24735 & ~w24736;
assign w24738 = pi03647 & ~w19092;
assign w24739 = ~pi02711 & w19092;
assign w24740 = ~w24738 & ~w24739;
assign w24741 = pi03648 & ~w19092;
assign w24742 = ~pi02170 & w19092;
assign w24743 = ~w24741 & ~w24742;
assign w24744 = pi03649 & ~w19092;
assign w24745 = ~pi02713 & w19092;
assign w24746 = ~w24744 & ~w24745;
assign w24747 = pi03650 & ~w19092;
assign w24748 = ~pi02714 & w19092;
assign w24749 = ~w24747 & ~w24748;
assign w24750 = pi03651 & ~w19092;
assign w24751 = ~pi02716 & w19092;
assign w24752 = ~w24750 & ~w24751;
assign w24753 = pi03652 & ~w19092;
assign w24754 = ~pi02717 & w19092;
assign w24755 = ~w24753 & ~w24754;
assign w24756 = pi03653 & ~w19096;
assign w24757 = ~pi02703 & w19096;
assign w24758 = ~w24756 & ~w24757;
assign w24759 = pi03654 & ~w19096;
assign w24760 = ~pi02169 & w19096;
assign w24761 = ~w24759 & ~w24760;
assign w24762 = pi03655 & ~w19096;
assign w24763 = ~pi02718 & w19096;
assign w24764 = ~w24762 & ~w24763;
assign w24765 = pi03656 & ~w19096;
assign w24766 = ~pi02167 & w19096;
assign w24767 = ~w24765 & ~w24766;
assign w24768 = pi03657 & ~w19096;
assign w24769 = ~pi02164 & w19096;
assign w24770 = ~w24768 & ~w24769;
assign w24771 = pi03658 & ~w19096;
assign w24772 = ~pi02722 & w19096;
assign w24773 = ~w24771 & ~w24772;
assign w24774 = pi03659 & ~w19096;
assign w24775 = ~pi02719 & w19096;
assign w24776 = ~w24774 & ~w24775;
assign w24777 = pi03660 & ~w19076;
assign w24778 = ~pi02711 & w19076;
assign w24779 = ~w24777 & ~w24778;
assign w24780 = pi03661 & ~w19076;
assign w24781 = ~pi02170 & w19076;
assign w24782 = ~w24780 & ~w24781;
assign w24783 = pi03662 & ~w19076;
assign w24784 = ~pi02713 & w19076;
assign w24785 = ~w24783 & ~w24784;
assign w24786 = pi03663 & ~w19076;
assign w24787 = ~pi02714 & w19076;
assign w24788 = ~w24786 & ~w24787;
assign w24789 = pi03664 & ~w19076;
assign w24790 = ~pi02716 & w19076;
assign w24791 = ~w24789 & ~w24790;
assign w24792 = pi03665 & ~w19004;
assign w24793 = ~pi02703 & w19004;
assign w24794 = ~w24792 & ~w24793;
assign w24795 = pi03666 & ~w19076;
assign w24796 = ~pi02717 & w19076;
assign w24797 = ~w24795 & ~w24796;
assign w24798 = pi03667 & ~w19004;
assign w24799 = ~pi02169 & w19004;
assign w24800 = ~w24798 & ~w24799;
assign w24801 = pi03668 & ~w19004;
assign w24802 = ~pi02718 & w19004;
assign w24803 = ~w24801 & ~w24802;
assign w24804 = pi03669 & ~w19004;
assign w24805 = ~pi02167 & w19004;
assign w24806 = ~w24804 & ~w24805;
assign w24807 = pi03670 & ~w19004;
assign w24808 = ~pi02164 & w19004;
assign w24809 = ~w24807 & ~w24808;
assign w24810 = pi03671 & ~w19065;
assign w24811 = ~pi02711 & w19065;
assign w24812 = ~w24810 & ~w24811;
assign w24813 = pi03672 & ~w19065;
assign w24814 = ~pi02712 & w19065;
assign w24815 = ~w24813 & ~w24814;
assign w24816 = pi03673 & ~w19004;
assign w24817 = ~pi02722 & w19004;
assign w24818 = ~w24816 & ~w24817;
assign w24819 = pi03674 & ~w19065;
assign w24820 = ~pi02170 & w19065;
assign w24821 = ~w24819 & ~w24820;
assign w24822 = pi03675 & ~w19065;
assign w24823 = ~pi02713 & w19065;
assign w24824 = ~w24822 & ~w24823;
assign w24825 = pi03676 & ~w19065;
assign w24826 = ~pi02714 & w19065;
assign w24827 = ~w24825 & ~w24826;
assign w24828 = pi03677 & ~w19065;
assign w24829 = ~pi02716 & w19065;
assign w24830 = ~w24828 & ~w24829;
assign w24831 = pi03678 & ~w19065;
assign w24832 = w16973 & w18995;
assign w24833 = ~w24831 & ~w24832;
assign w24834 = pi03679 & ~w19061;
assign w24835 = ~pi02711 & w19061;
assign w24836 = ~w24834 & ~w24835;
assign w24837 = pi03680 & ~w19061;
assign w24838 = ~pi02170 & w19061;
assign w24839 = ~w24837 & ~w24838;
assign w24840 = pi03681 & ~w19061;
assign w24841 = ~pi02713 & w19061;
assign w24842 = ~w24840 & ~w24841;
assign w24843 = pi03682 & ~w19061;
assign w24844 = ~pi02714 & w19061;
assign w24845 = ~w24843 & ~w24844;
assign w24846 = pi03683 & ~w19061;
assign w24847 = ~pi02715 & w19061;
assign w24848 = ~w24846 & ~w24847;
assign w24849 = pi03684 & ~w19061;
assign w24850 = ~pi02716 & w19061;
assign w24851 = ~w24849 & ~w24850;
assign w24852 = pi03685 & ~w19061;
assign w24853 = ~pi02717 & w19061;
assign w24854 = ~w24852 & ~w24853;
assign w24855 = pi03686 & ~w18991;
assign w24856 = ~pi02703 & w18991;
assign w24857 = ~w24855 & ~w24856;
assign w24858 = pi03687 & ~w18991;
assign w24859 = ~pi02169 & w18991;
assign w24860 = ~w24858 & ~w24859;
assign w24861 = pi03688 & ~w18991;
assign w24862 = ~pi02718 & w18991;
assign w24863 = ~w24861 & ~w24862;
assign w24864 = pi03689 & ~w18991;
assign w24865 = ~pi02167 & w18991;
assign w24866 = ~w24864 & ~w24865;
assign w24867 = pi03690 & ~w18991;
assign w24868 = ~pi02722 & w18991;
assign w24869 = ~w24867 & ~w24868;
assign w24870 = pi03691 & ~w18991;
assign w24871 = ~pi02719 & w18991;
assign w24872 = ~w24870 & ~w24871;
assign w24873 = pi03692 & ~w19035;
assign w24874 = ~pi02711 & w19035;
assign w24875 = ~w24873 & ~w24874;
assign w24876 = pi03693 & ~w19035;
assign w24877 = w19034 & w20209;
assign w24878 = ~w24876 & ~w24877;
assign w24879 = pi03694 & ~w19035;
assign w24880 = ~pi02713 & w19035;
assign w24881 = ~w24879 & ~w24880;
assign w24882 = pi03695 & ~w19035;
assign w24883 = w17742 & w19034;
assign w24884 = ~w24882 & ~w24883;
assign w24885 = pi03696 & ~w19035;
assign w24886 = ~pi02715 & w19035;
assign w24887 = ~w24885 & ~w24886;
assign w24888 = pi03697 & ~w19035;
assign w24889 = ~pi02716 & w19035;
assign w24890 = ~w24888 & ~w24889;
assign w24891 = pi03698 & ~w19035;
assign w24892 = ~pi02717 & w19035;
assign w24893 = ~w24891 & ~w24892;
assign w24894 = pi03699 & ~w18987;
assign w24895 = ~pi02711 & w18987;
assign w24896 = ~w24894 & ~w24895;
assign w24897 = pi03700 & ~w18987;
assign w24898 = ~pi02170 & w18987;
assign w24899 = ~w24897 & ~w24898;
assign w24900 = pi03701 & ~w18987;
assign w24901 = ~pi02713 & w18987;
assign w24902 = ~w24900 & ~w24901;
assign w24903 = pi03702 & ~w18987;
assign w24904 = ~pi02714 & w18987;
assign w24905 = ~w24903 & ~w24904;
assign w24906 = pi03703 & ~w18987;
assign w24907 = ~pi02716 & w18987;
assign w24908 = ~w24906 & ~w24907;
assign w24909 = pi03704 & ~w18864;
assign w24910 = ~pi02703 & w18864;
assign w24911 = ~w24909 & ~w24910;
assign w24912 = pi03705 & ~w18987;
assign w24913 = w16973 & w18986;
assign w24914 = ~w24912 & ~w24913;
assign w24915 = pi03706 & ~w18864;
assign w24916 = ~pi02169 & w18864;
assign w24917 = ~w24915 & ~w24916;
assign w24918 = pi03707 & ~w18864;
assign w24919 = w17586 & w18146;
assign w24920 = ~w24918 & ~w24919;
assign w24921 = pi03708 & ~w18864;
assign w24922 = ~pi02167 & w18864;
assign w24923 = ~w24921 & ~w24922;
assign w24924 = pi03709 & ~w18978;
assign w24925 = ~pi02711 & w18978;
assign w24926 = ~w24924 & ~w24925;
assign w24927 = pi03710 & ~w18978;
assign w24928 = ~pi02712 & w18978;
assign w24929 = ~w24927 & ~w24928;
assign w24930 = pi03711 & ~w18864;
assign w24931 = ~pi02164 & w18864;
assign w24932 = ~w24930 & ~w24931;
assign w24933 = pi03712 & ~w18978;
assign w24934 = ~pi02170 & w18978;
assign w24935 = ~w24933 & ~w24934;
assign w24936 = pi03713 & ~w18864;
assign w24937 = ~pi02722 & w18864;
assign w24938 = ~w24936 & ~w24937;
assign w24939 = pi03714 & ~w18978;
assign w24940 = ~pi02714 & w18978;
assign w24941 = ~w24939 & ~w24940;
assign w24942 = pi03715 & ~w18978;
assign w24943 = ~pi02715 & w18978;
assign w24944 = ~w24942 & ~w24943;
assign w24945 = pi03716 & ~w18978;
assign w24946 = ~pi02716 & w18978;
assign w24947 = ~w24945 & ~w24946;
assign w24948 = pi03717 & ~w18978;
assign w24949 = ~pi02717 & w18978;
assign w24950 = ~w24948 & ~w24949;
assign w24951 = pi03718 & ~w18967;
assign w24952 = ~pi02703 & w18967;
assign w24953 = ~w24951 & ~w24952;
assign w24954 = pi03719 & ~w18967;
assign w24955 = ~pi02169 & w18967;
assign w24956 = ~w24954 & ~w24955;
assign w24957 = pi03720 & ~w18967;
assign w24958 = ~pi02718 & w18967;
assign w24959 = ~w24957 & ~w24958;
assign w24960 = pi03721 & ~w18967;
assign w24961 = ~pi02167 & w18967;
assign w24962 = ~w24960 & ~w24961;
assign w24963 = pi03722 & ~w18967;
assign w24964 = w17620 & w18116;
assign w24965 = ~w24963 & ~w24964;
assign w24966 = pi03723 & ~w18967;
assign w24967 = ~pi02722 & w18967;
assign w24968 = ~w24966 & ~w24967;
assign w24969 = pi03724 & ~w18967;
assign w24970 = ~pi02719 & w18967;
assign w24971 = ~w24969 & ~w24970;
assign w24972 = pi03725 & ~w18945;
assign w24973 = ~pi02711 & w18945;
assign w24974 = ~w24972 & ~w24973;
assign w24975 = pi03726 & ~w18945;
assign w24976 = ~pi02170 & w18945;
assign w24977 = ~w24975 & ~w24976;
assign w24978 = pi03727 & ~w18945;
assign w24979 = ~pi02713 & w18945;
assign w24980 = ~w24978 & ~w24979;
assign w24981 = pi03728 & ~w18945;
assign w24982 = ~pi02714 & w18945;
assign w24983 = ~w24981 & ~w24982;
assign w24984 = pi03729 & ~w18945;
assign w24985 = ~pi02716 & w18945;
assign w24986 = ~w24984 & ~w24985;
assign w24987 = pi03730 & ~w18945;
assign w24988 = ~pi02717 & w18945;
assign w24989 = ~w24987 & ~w24988;
assign w24990 = pi03731 & ~w18940;
assign w24991 = w17603 & w18913;
assign w24992 = ~w24990 & ~w24991;
assign w24993 = pi03732 & ~w18940;
assign w24994 = ~pi02170 & w18940;
assign w24995 = ~w24993 & ~w24994;
assign w24996 = pi03733 & ~w18940;
assign w24997 = ~pi02713 & w18940;
assign w24998 = ~w24996 & ~w24997;
assign w24999 = pi03734 & ~w18940;
assign w25000 = ~pi02714 & w18940;
assign w25001 = ~w24999 & ~w25000;
assign w25002 = pi03735 & ~w18940;
assign w25003 = ~pi02715 & w18940;
assign w25004 = ~w25002 & ~w25003;
assign w25005 = pi03736 & ~w18940;
assign w25006 = ~pi02716 & w18940;
assign w25007 = ~w25005 & ~w25006;
assign w25008 = pi03737 & ~w18940;
assign w25009 = ~pi02717 & w18940;
assign w25010 = ~w25008 & ~w25009;
assign w25011 = pi03738 & ~w18898;
assign w25012 = ~pi02711 & w18898;
assign w25013 = ~w25011 & ~w25012;
assign w25014 = pi03739 & ~w18898;
assign w25015 = ~pi02170 & w18898;
assign w25016 = ~w25014 & ~w25015;
assign w25017 = pi03740 & ~w18898;
assign w25018 = ~pi02713 & w18898;
assign w25019 = ~w25017 & ~w25018;
assign w25020 = pi03741 & ~w18898;
assign w25021 = w17742 & w18897;
assign w25022 = ~w25020 & ~w25021;
assign w25023 = pi03742 & ~w18898;
assign w25024 = ~pi02716 & w18898;
assign w25025 = ~w25023 & ~w25024;
assign w25026 = pi03743 & ~w18898;
assign w25027 = ~pi02717 & w18898;
assign w25028 = ~w25026 & ~w25027;
assign w25029 = pi03744 & ~w18909;
assign w25030 = ~pi02703 & w18909;
assign w25031 = ~w25029 & ~w25030;
assign w25032 = pi03745 & ~w18909;
assign w25033 = ~pi02169 & w18909;
assign w25034 = ~w25032 & ~w25033;
assign w25035 = pi03746 & ~w18909;
assign w25036 = ~pi02718 & w18909;
assign w25037 = ~w25035 & ~w25036;
assign w25038 = pi03747 & ~w18909;
assign w25039 = w18070 & w19273;
assign w25040 = ~w25038 & ~w25039;
assign w25041 = pi03748 & ~w18909;
assign w25042 = ~pi02164 & w18909;
assign w25043 = ~w25041 & ~w25042;
assign w25044 = pi03749 & ~w18909;
assign w25045 = w18070 & w19312;
assign w25046 = ~w25044 & ~w25045;
assign w25047 = pi03750 & ~w18909;
assign w25048 = ~pi02719 & w18909;
assign w25049 = ~w25047 & ~w25048;
assign w25050 = pi03751 & ~w18872;
assign w25051 = ~pi02711 & w18872;
assign w25052 = ~w25050 & ~w25051;
assign w25053 = pi03752 & ~w18872;
assign w25054 = w18871 & w20209;
assign w25055 = ~w25053 & ~w25054;
assign w25056 = pi03753 & ~w18872;
assign w25057 = ~pi02713 & w18872;
assign w25058 = ~w25056 & ~w25057;
assign w25059 = pi03754 & ~w18872;
assign w25060 = w17742 & w18871;
assign w25061 = ~w25059 & ~w25060;
assign w25062 = pi03755 & ~w18872;
assign w25063 = ~pi02716 & w18872;
assign w25064 = ~w25062 & ~w25063;
assign w25065 = pi03756 & ~w18872;
assign w25066 = ~pi02717 & w18872;
assign w25067 = ~w25065 & ~w25066;
assign w25068 = pi03757 & ~w18786;
assign w25069 = ~pi02703 & w18786;
assign w25070 = ~w25068 & ~w25069;
assign w25071 = pi03758 & ~w18786;
assign w25072 = ~pi02169 & w18786;
assign w25073 = ~w25071 & ~w25072;
assign w25074 = pi03759 & ~w18786;
assign w25075 = ~pi02718 & w18786;
assign w25076 = ~w25074 & ~w25075;
assign w25077 = pi03760 & ~w18786;
assign w25078 = ~pi02167 & w18786;
assign w25079 = ~w25077 & ~w25078;
assign w25080 = pi03761 & ~w18786;
assign w25081 = ~pi02164 & w18786;
assign w25082 = ~w25080 & ~w25081;
assign w25083 = pi03762 & ~w18786;
assign w25084 = ~pi02722 & w18786;
assign w25085 = ~w25083 & ~w25084;
assign w25086 = pi03763 & ~w18786;
assign w25087 = ~pi02719 & w18786;
assign w25088 = ~w25086 & ~w25087;
assign w25089 = pi03764 & ~w18832;
assign w25090 = ~pi02711 & w18832;
assign w25091 = ~w25089 & ~w25090;
assign w25092 = pi03765 & ~w18832;
assign w25093 = ~pi02170 & w18832;
assign w25094 = ~w25092 & ~w25093;
assign w25095 = pi03766 & ~w18832;
assign w25096 = ~pi02713 & w18832;
assign w25097 = ~w25095 & ~w25096;
assign w25098 = pi03767 & ~w18832;
assign w25099 = ~pi02714 & w18832;
assign w25100 = ~w25098 & ~w25099;
assign w25101 = pi03768 & ~w18832;
assign w25102 = ~pi02716 & w18832;
assign w25103 = ~w25101 & ~w25102;
assign w25104 = pi03769 & ~w18832;
assign w25105 = ~pi02717 & w18832;
assign w25106 = ~w25104 & ~w25105;
assign w25107 = pi03770 & ~w18823;
assign w25108 = ~pi02711 & w18823;
assign w25109 = ~w25107 & ~w25108;
assign w25110 = pi03771 & ~w18823;
assign w25111 = ~pi02170 & w18823;
assign w25112 = ~w25110 & ~w25111;
assign w25113 = pi03772 & ~w18823;
assign w25114 = ~pi02713 & w18823;
assign w25115 = ~w25113 & ~w25114;
assign w25116 = pi03773 & ~w18823;
assign w25117 = ~pi02714 & w18823;
assign w25118 = ~w25116 & ~w25117;
assign w25119 = pi03774 & ~w18823;
assign w25120 = ~pi02715 & w18823;
assign w25121 = ~w25119 & ~w25120;
assign w25122 = pi03775 & ~w18823;
assign w25123 = ~pi02716 & w18823;
assign w25124 = ~w25122 & ~w25123;
assign w25125 = pi03776 & ~w18823;
assign w25126 = ~pi02717 & w18823;
assign w25127 = ~w25125 & ~w25126;
assign w25128 = pi03777 & ~w18613;
assign w25129 = ~pi02711 & w18613;
assign w25130 = ~w25128 & ~w25129;
assign w25131 = pi03778 & ~w18613;
assign w25132 = ~pi02712 & w18613;
assign w25133 = ~w25131 & ~w25132;
assign w25134 = pi03779 & ~w18613;
assign w25135 = w18612 & w20209;
assign w25136 = ~w25134 & ~w25135;
assign w25137 = pi03780 & ~w18503;
assign w25138 = ~pi02721 & w18503;
assign w25139 = ~w25137 & ~w25138;
assign w25140 = pi03781 & ~w18613;
assign w25141 = ~pi02714 & w18613;
assign w25142 = ~w25140 & ~w25141;
assign w25143 = pi03782 & ~w18503;
assign w25144 = ~pi02169 & w18503;
assign w25145 = ~w25143 & ~w25144;
assign w25146 = pi03783 & ~w18613;
assign w25147 = ~pi02715 & w18613;
assign w25148 = ~w25146 & ~w25147;
assign w25149 = pi03784 & ~w18503;
assign w25150 = ~pi02718 & w18503;
assign w25151 = ~w25149 & ~w25150;
assign w25152 = pi03785 & ~w18613;
assign w25153 = ~pi02717 & w18613;
assign w25154 = ~w25152 & ~w25153;
assign w25155 = pi03786 & ~w17517;
assign w25156 = ~pi02711 & w17517;
assign w25157 = ~w25155 & ~w25156;
assign w25158 = pi03787 & ~w17517;
assign w25159 = ~pi02712 & w17517;
assign w25160 = ~w25158 & ~w25159;
assign w25161 = pi03788 & ~w18503;
assign w25162 = ~pi02167 & w18503;
assign w25163 = ~w25161 & ~w25162;
assign w25164 = pi03789 & ~w17517;
assign w25165 = ~pi02170 & w17517;
assign w25166 = ~w25164 & ~w25165;
assign w25167 = pi03790 & ~w17517;
assign w25168 = ~pi02713 & w17517;
assign w25169 = ~w25167 & ~w25168;
assign w25170 = pi03791 & ~w17517;
assign w25171 = ~pi02714 & w17517;
assign w25172 = ~w25170 & ~w25171;
assign w25173 = pi03792 & ~w17517;
assign w25174 = w17516 & w18059;
assign w25175 = ~w25173 & ~w25174;
assign w25176 = pi03793 & ~w18503;
assign w25177 = ~pi02722 & w18503;
assign w25178 = ~w25176 & ~w25177;
assign w25179 = pi03794 & ~w17517;
assign w25180 = ~pi02717 & w17517;
assign w25181 = ~w25179 & ~w25180;
assign w25182 = pi03795 & ~w18432;
assign w25183 = ~pi02711 & w18432;
assign w25184 = ~w25182 & ~w25183;
assign w25185 = pi03796 & ~w18503;
assign w25186 = w17594 & w18051;
assign w25187 = ~w25185 & ~w25186;
assign w25188 = pi03797 & ~w18432;
assign w25189 = ~pi02170 & w18432;
assign w25190 = ~w25188 & ~w25189;
assign w25191 = pi03798 & ~w18432;
assign w25192 = ~pi02713 & w18432;
assign w25193 = ~w25191 & ~w25192;
assign w25194 = pi03799 & ~w18432;
assign w25195 = ~pi02714 & w18432;
assign w25196 = ~w25194 & ~w25195;
assign w25197 = pi03800 & ~w18432;
assign w25198 = w18059 & w18431;
assign w25199 = ~w25197 & ~w25198;
assign w25200 = pi03801 & ~w18432;
assign w25201 = ~pi02716 & w18432;
assign w25202 = ~w25200 & ~w25201;
assign w25203 = pi03802 & ~w18432;
assign w25204 = ~pi02717 & w18432;
assign w25205 = ~w25203 & ~w25204;
assign w25206 = pi03803 & ~w18248;
assign w25207 = ~pi02711 & w18248;
assign w25208 = ~w25206 & ~w25207;
assign w25209 = pi03804 & ~w18248;
assign w25210 = ~pi02170 & w18248;
assign w25211 = ~w25209 & ~w25210;
assign w25212 = pi03805 & ~w18248;
assign w25213 = ~pi02713 & w18248;
assign w25214 = ~w25212 & ~w25213;
assign w25215 = pi03806 & ~w18248;
assign w25216 = ~pi02714 & w18248;
assign w25217 = ~w25215 & ~w25216;
assign w25218 = pi03807 & ~w18248;
assign w25219 = ~pi02716 & w18248;
assign w25220 = ~w25218 & ~w25219;
assign w25221 = pi03808 & ~w18248;
assign w25222 = ~pi02717 & w18248;
assign w25223 = ~w25221 & ~w25222;
assign w25224 = pi03809 & ~w18319;
assign w25225 = w17510 & w17603;
assign w25226 = ~w25224 & ~w25225;
assign w25227 = pi03810 & ~w18319;
assign w25228 = ~pi02170 & w18319;
assign w25229 = ~w25227 & ~w25228;
assign w25230 = pi03811 & ~w18319;
assign w25231 = ~pi02713 & w18319;
assign w25232 = ~w25230 & ~w25231;
assign w25233 = pi03812 & ~w18319;
assign w25234 = w17510 & w17742;
assign w25235 = ~w25233 & ~w25234;
assign w25236 = pi03813 & ~w18319;
assign w25237 = ~pi02715 & w18319;
assign w25238 = ~w25236 & ~w25237;
assign w25239 = pi03814 & ~w18319;
assign w25240 = ~pi02716 & w18319;
assign w25241 = ~w25239 & ~w25240;
assign w25242 = pi03815 & ~w18319;
assign w25243 = ~pi02717 & w18319;
assign w25244 = ~w25242 & ~w25243;
assign w25245 = pi03816 & ~w18309;
assign w25246 = ~pi02711 & w18309;
assign w25247 = ~w25245 & ~w25246;
assign w25248 = pi03817 & ~w18309;
assign w25249 = ~pi02170 & w18309;
assign w25250 = ~w25248 & ~w25249;
assign w25251 = pi03818 & ~w18309;
assign w25252 = ~pi02713 & w18309;
assign w25253 = ~w25251 & ~w25252;
assign w25254 = pi03819 & ~w18309;
assign w25255 = ~pi02714 & w18309;
assign w25256 = ~w25254 & ~w25255;
assign w25257 = pi03820 & ~w18309;
assign w25258 = ~pi02716 & w18309;
assign w25259 = ~w25257 & ~w25258;
assign w25260 = pi03821 & ~w18309;
assign w25261 = ~pi02717 & w18309;
assign w25262 = ~w25260 & ~w25261;
assign w25263 = pi03822 & ~w18264;
assign w25264 = ~pi02711 & w18264;
assign w25265 = ~w25263 & ~w25264;
assign w25266 = pi03823 & ~w18264;
assign w25267 = ~pi02170 & w18264;
assign w25268 = ~w25266 & ~w25267;
assign w25269 = pi03824 & ~w18264;
assign w25270 = ~pi02713 & w18264;
assign w25271 = ~w25269 & ~w25270;
assign w25272 = pi03825 & ~w18264;
assign w25273 = ~pi02714 & w18264;
assign w25274 = ~w25272 & ~w25273;
assign w25275 = pi03826 & ~w18264;
assign w25276 = w18059 & w18263;
assign w25277 = ~w25275 & ~w25276;
assign w25278 = pi03827 & ~w18264;
assign w25279 = ~pi02716 & w18264;
assign w25280 = ~w25278 & ~w25279;
assign w25281 = pi03828 & ~w18264;
assign w25282 = ~pi02717 & w18264;
assign w25283 = ~w25281 & ~w25282;
assign w25284 = pi03829 & ~w18156;
assign w25285 = w17603 & w18155;
assign w25286 = ~w25284 & ~w25285;
assign w25287 = pi03830 & ~w18156;
assign w25288 = w18155 & w20209;
assign w25289 = ~w25287 & ~w25288;
assign w25290 = pi03831 & ~w18156;
assign w25291 = w17929 & w18155;
assign w25292 = ~w25290 & ~w25291;
assign w25293 = pi03832 & ~w18156;
assign w25294 = w17742 & w18155;
assign w25295 = ~w25293 & ~w25294;
assign w25296 = pi03833 & ~w18156;
assign w25297 = w17317 & w18155;
assign w25298 = ~w25296 & ~w25297;
assign w25299 = pi03834 & ~w18156;
assign w25300 = w16973 & w18155;
assign w25301 = ~w25299 & ~w25300;
assign w25302 = pi03835 & ~w18147;
assign w25303 = ~pi02711 & w18147;
assign w25304 = ~w25302 & ~w25303;
assign w25305 = pi03836 & ~w18147;
assign w25306 = ~pi02170 & w18147;
assign w25307 = ~w25305 & ~w25306;
assign w25308 = pi03837 & ~w18147;
assign w25309 = w17929 & w18146;
assign w25310 = ~w25308 & ~w25309;
assign w25311 = pi03838 & ~w18147;
assign w25312 = w17742 & w18146;
assign w25313 = ~w25311 & ~w25312;
assign w25314 = pi03839 & ~w18147;
assign w25315 = ~pi02715 & w18147;
assign w25316 = ~w25314 & ~w25315;
assign w25317 = pi03840 & ~w18147;
assign w25318 = w17317 & w18146;
assign w25319 = ~w25317 & ~w25318;
assign w25320 = pi03841 & ~w18147;
assign w25321 = ~pi02717 & w18147;
assign w25322 = ~w25320 & ~w25321;
assign w25323 = pi03842 & ~w18117;
assign w25324 = ~pi02711 & w18117;
assign w25325 = ~w25323 & ~w25324;
assign w25326 = pi03843 & ~w18117;
assign w25327 = ~pi02170 & w18117;
assign w25328 = ~w25326 & ~w25327;
assign w25329 = pi03844 & ~w18117;
assign w25330 = ~pi02713 & w18117;
assign w25331 = ~w25329 & ~w25330;
assign w25332 = pi03845 & ~w18117;
assign w25333 = ~pi02714 & w18117;
assign w25334 = ~w25332 & ~w25333;
assign w25335 = pi03846 & ~w18117;
assign w25336 = ~pi02716 & w18117;
assign w25337 = ~w25335 & ~w25336;
assign w25338 = pi03847 & ~w18117;
assign w25339 = ~pi02717 & w18117;
assign w25340 = ~w25338 & ~w25339;
assign w25341 = pi03848 & ~w18071;
assign w25342 = w17603 & w18070;
assign w25343 = ~w25341 & ~w25342;
assign w25344 = pi03849 & ~w18071;
assign w25345 = ~pi02170 & w18071;
assign w25346 = ~w25344 & ~w25345;
assign w25347 = pi03850 & ~w18071;
assign w25348 = w17929 & w18070;
assign w25349 = ~w25347 & ~w25348;
assign w25350 = pi03851 & ~w18071;
assign w25351 = w17742 & w18070;
assign w25352 = ~w25350 & ~w25351;
assign w25353 = pi03852 & ~w18071;
assign w25354 = ~pi02715 & w18071;
assign w25355 = ~w25353 & ~w25354;
assign w25356 = pi03853 & ~w18071;
assign w25357 = ~pi02716 & w18071;
assign w25358 = ~w25356 & ~w25357;
assign w25359 = pi03854 & ~w18071;
assign w25360 = w16973 & w18070;
assign w25361 = ~w25359 & ~w25360;
assign w25362 = pi03855 & ~w18057;
assign w25363 = ~pi02711 & w18057;
assign w25364 = ~w25362 & ~w25363;
assign w25365 = pi03856 & ~w18057;
assign w25366 = ~pi02170 & w18057;
assign w25367 = ~w25365 & ~w25366;
assign w25368 = pi03857 & ~w18057;
assign w25369 = ~pi02713 & w18057;
assign w25370 = ~w25368 & ~w25369;
assign w25371 = pi03858 & ~w18057;
assign w25372 = ~pi02714 & w18057;
assign w25373 = ~w25371 & ~w25372;
assign w25374 = pi03859 & ~w18057;
assign w25375 = ~pi02716 & w18057;
assign w25376 = ~w25374 & ~w25375;
assign w25377 = pi03860 & ~w18057;
assign w25378 = ~pi02717 & w18057;
assign w25379 = ~w25377 & ~w25378;
assign w25380 = pi03861 & ~w18052;
assign w25381 = ~pi02711 & w18052;
assign w25382 = ~w25380 & ~w25381;
assign w25383 = pi03862 & ~w18052;
assign w25384 = ~pi02170 & w18052;
assign w25385 = ~w25383 & ~w25384;
assign w25386 = pi03863 & ~w18052;
assign w25387 = ~pi02713 & w18052;
assign w25388 = ~w25386 & ~w25387;
assign w25389 = pi03864 & ~w18052;
assign w25390 = ~pi02714 & w18052;
assign w25391 = ~w25389 & ~w25390;
assign w25392 = pi03865 & ~w18052;
assign w25393 = ~pi02715 & w18052;
assign w25394 = ~w25392 & ~w25393;
assign w25395 = pi03866 & ~w18052;
assign w25396 = ~pi02716 & w18052;
assign w25397 = ~w25395 & ~w25396;
assign w25398 = pi03867 & ~w18052;
assign w25399 = ~pi02717 & w18052;
assign w25400 = ~w25398 & ~w25399;
assign w25401 = pi03868 & ~w17889;
assign w25402 = ~pi02703 & w17889;
assign w25403 = ~w25401 & ~w25402;
assign w25404 = pi03869 & ~w17889;
assign w25405 = ~pi02169 & w17889;
assign w25406 = ~w25404 & ~w25405;
assign w25407 = pi03870 & ~w17889;
assign w25408 = ~pi02718 & w17889;
assign w25409 = ~w25407 & ~w25408;
assign w25410 = pi03871 & ~w17889;
assign w25411 = ~pi02167 & w17889;
assign w25412 = ~w25410 & ~w25411;
assign w25413 = pi03872 & ~w17889;
assign w25414 = ~pi02722 & w17889;
assign w25415 = ~w25413 & ~w25414;
assign w25416 = pi03873 & ~w17889;
assign w25417 = ~pi02719 & w17889;
assign w25418 = ~w25416 & ~w25417;
assign w25419 = pi03874 & ~w17730;
assign w25420 = w17017 & w17532;
assign w25421 = ~w25419 & ~w25420;
assign w25422 = pi03875 & ~w17730;
assign w25423 = ~pi02169 & w17730;
assign w25424 = ~w25422 & ~w25423;
assign w25425 = pi03876 & ~w17730;
assign w25426 = ~pi02718 & w17730;
assign w25427 = ~w25425 & ~w25426;
assign w25428 = pi03877 & ~w17730;
assign w25429 = w17017 & w19273;
assign w25430 = ~w25428 & ~w25429;
assign w25431 = pi03878 & ~w17730;
assign w25432 = ~pi02164 & w17730;
assign w25433 = ~w25431 & ~w25432;
assign w25434 = pi03879 & ~w17730;
assign w25435 = ~pi02722 & w17730;
assign w25436 = ~w25434 & ~w25435;
assign w25437 = pi03880 & ~w17730;
assign w25438 = ~pi02719 & w17730;
assign w25439 = ~w25437 & ~w25438;
assign w25440 = pi03881 & ~w17578;
assign w25441 = ~pi02703 & w17578;
assign w25442 = ~w25440 & ~w25441;
assign w25443 = pi03882 & ~w17578;
assign w25444 = ~pi02169 & w17578;
assign w25445 = ~w25443 & ~w25444;
assign w25446 = pi03883 & ~w17578;
assign w25447 = ~pi02718 & w17578;
assign w25448 = ~w25446 & ~w25447;
assign w25449 = pi03884 & ~w17578;
assign w25450 = ~pi02167 & w17578;
assign w25451 = ~w25449 & ~w25450;
assign w25452 = pi03885 & ~w17578;
assign w25453 = ~pi02722 & w17578;
assign w25454 = ~w25452 & ~w25453;
assign w25455 = pi03886 & ~w17578;
assign w25456 = ~pi02719 & w17578;
assign w25457 = ~w25455 & ~w25456;
assign w25458 = pi03887 & ~w17446;
assign w25459 = ~pi02711 & w17446;
assign w25460 = ~w25458 & ~w25459;
assign w25461 = pi03888 & ~w17446;
assign w25462 = ~pi02170 & w17446;
assign w25463 = ~w25461 & ~w25462;
assign w25464 = pi03889 & ~w17446;
assign w25465 = ~pi02713 & w17446;
assign w25466 = ~w25464 & ~w25465;
assign w25467 = pi03890 & ~w17446;
assign w25468 = ~pi02714 & w17446;
assign w25469 = ~w25467 & ~w25468;
assign w25470 = pi03891 & ~w17446;
assign w25471 = w17445 & w18059;
assign w25472 = ~w25470 & ~w25471;
assign w25473 = pi03892 & ~w17446;
assign w25474 = ~pi02716 & w17446;
assign w25475 = ~w25473 & ~w25474;
assign w25476 = pi03893 & ~w17446;
assign w25477 = ~pi02717 & w17446;
assign w25478 = ~w25476 & ~w25477;
assign w25479 = pi03894 & ~w17018;
assign w25480 = ~pi02711 & w17018;
assign w25481 = ~w25479 & ~w25480;
assign w25482 = pi03895 & ~w17018;
assign w25483 = ~pi02170 & w17018;
assign w25484 = ~w25482 & ~w25483;
assign w25485 = pi03896 & ~w17018;
assign w25486 = ~pi02713 & w17018;
assign w25487 = ~w25485 & ~w25486;
assign w25488 = pi03897 & ~w17018;
assign w25489 = ~pi02714 & w17018;
assign w25490 = ~w25488 & ~w25489;
assign w25491 = pi03898 & ~w17018;
assign w25492 = ~pi02716 & w17018;
assign w25493 = ~w25491 & ~w25492;
assign w25494 = pi03899 & ~w17018;
assign w25495 = ~pi02717 & w17018;
assign w25496 = ~w25494 & ~w25495;
assign w25497 = pi03900 & ~w17138;
assign w25498 = ~pi02711 & w17138;
assign w25499 = ~w25497 & ~w25498;
assign w25500 = ~w16928 & w19327;
assign w25501 = pi03901 & ~w25500;
assign w25502 = ~pi02178 & w25500;
assign w25503 = ~w25501 & ~w25502;
assign w25504 = pi03902 & ~w17138;
assign w25505 = ~pi02170 & w17138;
assign w25506 = ~w25504 & ~w25505;
assign w25507 = pi03903 & ~w17138;
assign w25508 = ~pi02713 & w17138;
assign w25509 = ~w25507 & ~w25508;
assign w25510 = pi03904 & ~w17138;
assign w25511 = ~pi02714 & w17138;
assign w25512 = ~w25510 & ~w25511;
assign w25513 = pi03905 & ~w17138;
assign w25514 = ~pi02715 & w17138;
assign w25515 = ~w25513 & ~w25514;
assign w25516 = pi03906 & ~w17138;
assign w25517 = ~pi02716 & w17138;
assign w25518 = ~w25516 & ~w25517;
assign w25519 = pi03907 & ~w17138;
assign w25520 = ~pi02717 & w17138;
assign w25521 = ~w25519 & ~w25520;
assign w25522 = pi03908 & ~w16995;
assign w25523 = ~pi02703 & w16995;
assign w25524 = ~w25522 & ~w25523;
assign w25525 = pi03909 & ~w16995;
assign w25526 = w16994 & w19797;
assign w25527 = ~w25525 & ~w25526;
assign w25528 = pi03910 & ~w16995;
assign w25529 = ~pi02718 & w16995;
assign w25530 = ~w25528 & ~w25529;
assign w25531 = pi03911 & ~w16995;
assign w25532 = ~pi02167 & w16995;
assign w25533 = ~w25531 & ~w25532;
assign w25534 = pi03912 & ~w16995;
assign w25535 = ~pi02164 & w16995;
assign w25536 = ~w25534 & ~w25535;
assign w25537 = pi03913 & ~w17071;
assign w25538 = ~pi02712 & w17071;
assign w25539 = ~w25537 & ~w25538;
assign w25540 = pi03914 & ~w17071;
assign w25541 = ~pi02170 & w17071;
assign w25542 = ~w25540 & ~w25541;
assign w25543 = pi03915 & ~w17071;
assign w25544 = ~pi02713 & w17071;
assign w25545 = ~w25543 & ~w25544;
assign w25546 = pi03916 & ~w17071;
assign w25547 = ~pi02714 & w17071;
assign w25548 = ~w25546 & ~w25547;
assign w25549 = pi03917 & ~w16995;
assign w25550 = ~pi02719 & w16995;
assign w25551 = ~w25549 & ~w25550;
assign w25552 = pi03918 & ~w17071;
assign w25553 = ~pi02715 & w17071;
assign w25554 = ~w25552 & ~w25553;
assign w25555 = pi03919 & ~w17071;
assign w25556 = ~pi02716 & w17071;
assign w25557 = ~w25555 & ~w25556;
assign w25558 = ~w16992 & w17965;
assign w25559 = pi03920 & ~w25558;
assign w25560 = w17532 & w17965;
assign w25561 = ~w25559 & ~w25560;
assign w25562 = pi03921 & ~w17071;
assign w25563 = ~pi02717 & w17071;
assign w25564 = ~w25562 & ~w25563;
assign w25565 = ~w16905 & w17965;
assign w25566 = pi03922 & ~w25565;
assign w25567 = w17020 & w17965;
assign w25568 = ~w25566 & ~w25567;
assign w25569 = pi03923 & ~w25558;
assign w25570 = w17811 & w17965;
assign w25571 = ~w25569 & ~w25570;
assign w25572 = pi03924 & ~w25565;
assign w25573 = w17965 & w20209;
assign w25574 = ~w25572 & ~w25573;
assign w25575 = pi03925 & ~w25558;
assign w25576 = ~pi02169 & w25558;
assign w25577 = ~w25575 & ~w25576;
assign w25578 = pi03926 & ~w25565;
assign w25579 = ~pi02714 & w25565;
assign w25580 = ~w25578 & ~w25579;
assign w25581 = pi03927 & ~w25565;
assign w25582 = ~pi02715 & w25565;
assign w25583 = ~w25581 & ~w25582;
assign w25584 = pi03928 & ~w25565;
assign w25585 = ~pi02716 & w25565;
assign w25586 = ~w25584 & ~w25585;
assign w25587 = pi03929 & ~w25565;
assign w25588 = ~pi02717 & w25565;
assign w25589 = ~w25587 & ~w25588;
assign w25590 = pi03930 & ~w25558;
assign w25591 = ~pi02167 & w25558;
assign w25592 = ~w25590 & ~w25591;
assign w25593 = pi03931 & ~w25558;
assign w25594 = ~pi02164 & w25558;
assign w25595 = ~w25593 & ~w25594;
assign w25596 = pi03932 & ~w25558;
assign w25597 = ~pi02722 & w25558;
assign w25598 = ~w25596 & ~w25597;
assign w25599 = pi03933 & ~w25558;
assign w25600 = ~pi02719 & w25558;
assign w25601 = ~w25599 & ~w25600;
assign w25602 = ~w16905 & w17912;
assign w25603 = pi03934 & ~w25602;
assign w25604 = ~pi02711 & w25602;
assign w25605 = ~w25603 & ~w25604;
assign w25606 = pi03935 & ~w25602;
assign w25607 = ~pi02170 & w25602;
assign w25608 = ~w25606 & ~w25607;
assign w25609 = pi03936 & ~w25602;
assign w25610 = ~pi02713 & w25602;
assign w25611 = ~w25609 & ~w25610;
assign w25612 = pi03937 & ~w25602;
assign w25613 = ~pi02714 & w25602;
assign w25614 = ~w25612 & ~w25613;
assign w25615 = pi03938 & ~w25602;
assign w25616 = ~pi02716 & w25602;
assign w25617 = ~w25615 & ~w25616;
assign w25618 = pi03939 & ~w25602;
assign w25619 = ~pi02717 & w25602;
assign w25620 = ~w25618 & ~w25619;
assign w25621 = ~w16992 & w17912;
assign w25622 = pi03940 & ~w25621;
assign w25623 = ~pi02703 & w25621;
assign w25624 = ~w25622 & ~w25623;
assign w25625 = pi03941 & ~w25621;
assign w25626 = ~pi02169 & w25621;
assign w25627 = ~w25625 & ~w25626;
assign w25628 = pi03942 & ~w25621;
assign w25629 = ~pi02718 & w25621;
assign w25630 = ~w25628 & ~w25629;
assign w25631 = pi03943 & ~w25621;
assign w25632 = ~pi02167 & w25621;
assign w25633 = ~w25631 & ~w25632;
assign w25634 = pi03944 & ~w25621;
assign w25635 = ~pi02164 & w25621;
assign w25636 = ~w25634 & ~w25635;
assign w25637 = pi03945 & ~w25621;
assign w25638 = ~pi02722 & w25621;
assign w25639 = ~w25637 & ~w25638;
assign w25640 = pi03946 & ~w25621;
assign w25641 = w17594 & w17912;
assign w25642 = ~w25640 & ~w25641;
assign w25643 = ~w16905 & w17626;
assign w25644 = pi03947 & ~w25643;
assign w25645 = ~pi02711 & w25643;
assign w25646 = ~w25644 & ~w25645;
assign w25647 = pi03948 & ~w25643;
assign w25648 = ~pi02170 & w25643;
assign w25649 = ~w25647 & ~w25648;
assign w25650 = pi03949 & ~w25643;
assign w25651 = ~pi02713 & w25643;
assign w25652 = ~w25650 & ~w25651;
assign w25653 = pi03950 & ~w25643;
assign w25654 = ~pi02714 & w25643;
assign w25655 = ~w25653 & ~w25654;
assign w25656 = pi03951 & ~w25643;
assign w25657 = ~pi02716 & w25643;
assign w25658 = ~w25656 & ~w25657;
assign w25659 = pi03952 & ~w25643;
assign w25660 = ~pi02717 & w25643;
assign w25661 = ~w25659 & ~w25660;
assign w25662 = ~w16905 & w20119;
assign w25663 = pi03953 & ~w25662;
assign w25664 = ~pi02711 & w25662;
assign w25665 = ~w25663 & ~w25664;
assign w25666 = pi03954 & ~w25662;
assign w25667 = w20119 & w20209;
assign w25668 = ~w25666 & ~w25667;
assign w25669 = pi03955 & ~w25662;
assign w25670 = ~pi02713 & w25662;
assign w25671 = ~w25669 & ~w25670;
assign w25672 = pi03956 & ~w25662;
assign w25673 = ~pi02714 & w25662;
assign w25674 = ~w25672 & ~w25673;
assign w25675 = pi03957 & ~w25662;
assign w25676 = ~pi02715 & w25662;
assign w25677 = ~w25675 & ~w25676;
assign w25678 = pi03958 & ~w25662;
assign w25679 = ~pi02716 & w25662;
assign w25680 = ~w25678 & ~w25679;
assign w25681 = pi03959 & ~w25662;
assign w25682 = ~pi02717 & w25662;
assign w25683 = ~w25681 & ~w25682;
assign w25684 = ~w16905 & w16954;
assign w25685 = pi03960 & ~w25684;
assign w25686 = ~pi02711 & w25684;
assign w25687 = ~w25685 & ~w25686;
assign w25688 = pi03961 & ~w25684;
assign w25689 = ~pi02170 & w25684;
assign w25690 = ~w25688 & ~w25689;
assign w25691 = pi03962 & ~w25684;
assign w25692 = ~pi02713 & w25684;
assign w25693 = ~w25691 & ~w25692;
assign w25694 = pi03963 & ~w25684;
assign w25695 = ~pi02714 & w25684;
assign w25696 = ~w25694 & ~w25695;
assign w25697 = pi03964 & ~w25684;
assign w25698 = ~pi02716 & w25684;
assign w25699 = ~w25697 & ~w25698;
assign w25700 = pi03965 & ~w25684;
assign w25701 = ~pi02717 & w25684;
assign w25702 = ~w25700 & ~w25701;
assign w25703 = ~w16992 & w17626;
assign w25704 = pi03966 & ~w25703;
assign w25705 = w17532 & w17626;
assign w25706 = ~w25704 & ~w25705;
assign w25707 = pi03967 & ~w25703;
assign w25708 = ~pi02169 & w25703;
assign w25709 = ~w25707 & ~w25708;
assign w25710 = ~w16905 & w17103;
assign w25711 = pi03968 & ~w25710;
assign w25712 = w17103 & w17603;
assign w25713 = ~w25711 & ~w25712;
assign w25714 = pi03969 & ~w25703;
assign w25715 = ~pi02718 & w25703;
assign w25716 = ~w25714 & ~w25715;
assign w25717 = pi03970 & ~w25703;
assign w25718 = ~pi02167 & w25703;
assign w25719 = ~w25717 & ~w25718;
assign w25720 = pi03971 & ~w25710;
assign w25721 = w17020 & w17103;
assign w25722 = ~w25720 & ~w25721;
assign w25723 = pi03972 & ~w25710;
assign w25724 = ~pi02170 & w25710;
assign w25725 = ~w25723 & ~w25724;
assign w25726 = pi03973 & ~w25703;
assign w25727 = ~pi02164 & w25703;
assign w25728 = ~w25726 & ~w25727;
assign w25729 = pi03974 & ~w25710;
assign w25730 = w17103 & w17742;
assign w25731 = ~w25729 & ~w25730;
assign w25732 = pi03975 & ~w25703;
assign w25733 = w17626 & w19312;
assign w25734 = ~w25732 & ~w25733;
assign w25735 = pi03976 & ~w25710;
assign w25736 = w17103 & w18059;
assign w25737 = ~w25735 & ~w25736;
assign w25738 = pi03977 & ~w25703;
assign w25739 = ~pi02719 & w25703;
assign w25740 = ~w25738 & ~w25739;
assign w25741 = pi03978 & ~w25710;
assign w25742 = w16973 & w17103;
assign w25743 = ~w25741 & ~w25742;
assign w25744 = ~w16905 & w17078;
assign w25745 = pi03979 & ~w25744;
assign w25746 = w17078 & w17603;
assign w25747 = ~w25745 & ~w25746;
assign w25748 = pi03980 & ~w25744;
assign w25749 = ~pi02170 & w25744;
assign w25750 = ~w25748 & ~w25749;
assign w25751 = pi03981 & ~w25744;
assign w25752 = w17078 & w17929;
assign w25753 = ~w25751 & ~w25752;
assign w25754 = pi03982 & ~w25744;
assign w25755 = w17078 & w17742;
assign w25756 = ~w25754 & ~w25755;
assign w25757 = pi03983 & ~w25744;
assign w25758 = w17078 & w18059;
assign w25759 = ~w25757 & ~w25758;
assign w25760 = pi03984 & ~w25744;
assign w25761 = ~pi02716 & w25744;
assign w25762 = ~w25760 & ~w25761;
assign w25763 = pi03985 & ~w25744;
assign w25764 = w16973 & w17078;
assign w25765 = ~w25763 & ~w25764;
assign w25766 = ~w16992 & w20119;
assign w25767 = pi03986 & ~w25766;
assign w25768 = ~pi02703 & w25766;
assign w25769 = ~w25767 & ~w25768;
assign w25770 = pi03987 & ~w25766;
assign w25771 = ~pi02169 & w25766;
assign w25772 = ~w25770 & ~w25771;
assign w25773 = pi03988 & ~w25766;
assign w25774 = ~pi02718 & w25766;
assign w25775 = ~w25773 & ~w25774;
assign w25776 = pi03989 & ~w25766;
assign w25777 = ~pi02167 & w25766;
assign w25778 = ~w25776 & ~w25777;
assign w25779 = pi03990 & ~w25766;
assign w25780 = ~pi02722 & w25766;
assign w25781 = ~w25779 & ~w25780;
assign w25782 = pi03991 & ~w25766;
assign w25783 = ~pi02719 & w25766;
assign w25784 = ~w25782 & ~w25783;
assign w25785 = w16954 & ~w16992;
assign w25786 = pi03992 & ~w25785;
assign w25787 = ~pi02703 & w25785;
assign w25788 = ~w25786 & ~w25787;
assign w25789 = pi03993 & ~w25785;
assign w25790 = w16954 & w19797;
assign w25791 = ~w25789 & ~w25790;
assign w25792 = pi03994 & ~w25785;
assign w25793 = ~pi02718 & w25785;
assign w25794 = ~w25792 & ~w25793;
assign w25795 = pi03995 & ~w25785;
assign w25796 = ~pi02167 & w25785;
assign w25797 = ~w25795 & ~w25796;
assign w25798 = pi03996 & ~w25785;
assign w25799 = ~pi02164 & w25785;
assign w25800 = ~w25798 & ~w25799;
assign w25801 = pi03997 & ~w25785;
assign w25802 = ~pi02722 & w25785;
assign w25803 = ~w25801 & ~w25802;
assign w25804 = pi03998 & ~w25785;
assign w25805 = ~pi02719 & w25785;
assign w25806 = ~w25804 & ~w25805;
assign w25807 = ~w16905 & w20075;
assign w25808 = pi03999 & ~w25807;
assign w25809 = ~pi02711 & w25807;
assign w25810 = ~w25808 & ~w25809;
assign w25811 = pi04000 & ~w25807;
assign w25812 = ~pi02170 & w25807;
assign w25813 = ~w25811 & ~w25812;
assign w25814 = pi04001 & ~w25807;
assign w25815 = ~pi02713 & w25807;
assign w25816 = ~w25814 & ~w25815;
assign w25817 = pi04002 & ~w25807;
assign w25818 = ~pi02714 & w25807;
assign w25819 = ~w25817 & ~w25818;
assign w25820 = pi04003 & ~w25807;
assign w25821 = ~pi02716 & w25807;
assign w25822 = ~w25820 & ~w25821;
assign w25823 = pi04004 & ~w25807;
assign w25824 = ~pi02717 & w25807;
assign w25825 = ~w25823 & ~w25824;
assign w25826 = ~w16905 & w20059;
assign w25827 = pi04005 & ~w25826;
assign w25828 = ~pi02711 & w25826;
assign w25829 = ~w25827 & ~w25828;
assign w25830 = pi04006 & ~w25826;
assign w25831 = ~pi02170 & w25826;
assign w25832 = ~w25830 & ~w25831;
assign w25833 = pi04007 & ~w25826;
assign w25834 = ~pi02713 & w25826;
assign w25835 = ~w25833 & ~w25834;
assign w25836 = pi04008 & ~w25826;
assign w25837 = ~pi02714 & w25826;
assign w25838 = ~w25836 & ~w25837;
assign w25839 = pi04009 & ~w25826;
assign w25840 = ~pi02715 & w25826;
assign w25841 = ~w25839 & ~w25840;
assign w25842 = pi04010 & ~w25826;
assign w25843 = ~pi02716 & w25826;
assign w25844 = ~w25842 & ~w25843;
assign w25845 = pi04011 & ~w25826;
assign w25846 = w16973 & w20059;
assign w25847 = ~w25845 & ~w25846;
assign w25848 = ~w16905 & w20014;
assign w25849 = pi04012 & ~w25848;
assign w25850 = ~pi02711 & w25848;
assign w25851 = ~w25849 & ~w25850;
assign w25852 = pi04013 & ~w25848;
assign w25853 = ~pi02170 & w25848;
assign w25854 = ~w25852 & ~w25853;
assign w25855 = pi04014 & ~w25848;
assign w25856 = w17929 & w20014;
assign w25857 = ~w25855 & ~w25856;
assign w25858 = pi04015 & ~w25848;
assign w25859 = ~pi02714 & w25848;
assign w25860 = ~w25858 & ~w25859;
assign w25861 = pi04016 & ~w25848;
assign w25862 = w17317 & w20014;
assign w25863 = ~w25861 & ~w25862;
assign w25864 = pi04017 & ~w25848;
assign w25865 = w16973 & w20014;
assign w25866 = ~w25864 & ~w25865;
assign w25867 = ~w16992 & w17103;
assign w25868 = pi04018 & ~w25867;
assign w25869 = ~pi02703 & w25867;
assign w25870 = ~w25868 & ~w25869;
assign w25871 = ~w16905 & w19988;
assign w25872 = pi04019 & ~w25871;
assign w25873 = ~pi02711 & w25871;
assign w25874 = ~w25872 & ~w25873;
assign w25875 = pi04020 & ~w25867;
assign w25876 = w17103 & w19797;
assign w25877 = ~w25875 & ~w25876;
assign w25878 = pi04021 & ~w25871;
assign w25879 = ~pi02712 & w25871;
assign w25880 = ~w25878 & ~w25879;
assign w25881 = pi04022 & ~w25871;
assign w25882 = ~pi02170 & w25871;
assign w25883 = ~w25881 & ~w25882;
assign w25884 = pi04023 & ~w25867;
assign w25885 = ~pi02718 & w25867;
assign w25886 = ~w25884 & ~w25885;
assign w25887 = pi04024 & ~w25871;
assign w25888 = w17929 & w19988;
assign w25889 = ~w25887 & ~w25888;
assign w25890 = pi04025 & ~w25867;
assign w25891 = ~pi02167 & w25867;
assign w25892 = ~w25890 & ~w25891;
assign w25893 = pi04026 & ~w25867;
assign w25894 = w17103 & w17620;
assign w25895 = ~w25893 & ~w25894;
assign w25896 = pi04027 & ~w25867;
assign w25897 = ~pi02722 & w25867;
assign w25898 = ~w25896 & ~w25897;
assign w25899 = pi04028 & ~w25871;
assign w25900 = ~pi02715 & w25871;
assign w25901 = ~w25899 & ~w25900;
assign w25902 = pi04029 & ~w25871;
assign w25903 = ~pi02717 & w25871;
assign w25904 = ~w25902 & ~w25903;
assign w25905 = pi04030 & ~w25867;
assign w25906 = ~pi02719 & w25867;
assign w25907 = ~w25905 & ~w25906;
assign w25908 = ~w16992 & w17078;
assign w25909 = pi04031 & ~w25908;
assign w25910 = ~pi02703 & w25908;
assign w25911 = ~w25909 & ~w25910;
assign w25912 = ~w16992 & w18645;
assign w25913 = pi04032 & ~w25912;
assign w25914 = ~pi02719 & w25912;
assign w25915 = ~w25913 & ~w25914;
assign w25916 = pi04033 & ~w25908;
assign w25917 = ~pi02169 & w25908;
assign w25918 = ~w25916 & ~w25917;
assign w25919 = ~w16905 & w19941;
assign w25920 = pi04034 & ~w25919;
assign w25921 = w17603 & w19941;
assign w25922 = ~w25920 & ~w25921;
assign w25923 = pi04035 & ~w25919;
assign w25924 = ~pi02712 & w25919;
assign w25925 = ~w25923 & ~w25924;
assign w25926 = pi04036 & ~w25919;
assign w25927 = ~pi02170 & w25919;
assign w25928 = ~w25926 & ~w25927;
assign w25929 = pi04037 & ~w25908;
assign w25930 = ~pi02718 & w25908;
assign w25931 = ~w25929 & ~w25930;
assign w25932 = pi04038 & ~w25919;
assign w25933 = ~pi02713 & w25919;
assign w25934 = ~w25932 & ~w25933;
assign w25935 = pi04039 & ~w25919;
assign w25936 = ~pi02714 & w25919;
assign w25937 = ~w25935 & ~w25936;
assign w25938 = pi04040 & ~w25919;
assign w25939 = ~pi02715 & w25919;
assign w25940 = ~w25938 & ~w25939;
assign w25941 = pi04041 & ~w25908;
assign w25942 = w17078 & w17620;
assign w25943 = ~w25941 & ~w25942;
assign w25944 = pi04042 & ~w25919;
assign w25945 = ~pi02716 & w25919;
assign w25946 = ~w25944 & ~w25945;
assign w25947 = pi04043 & ~w25908;
assign w25948 = w17078 & w17594;
assign w25949 = ~w25947 & ~w25948;
assign w25950 = pi04044 & ~w25919;
assign w25951 = ~pi02717 & w25919;
assign w25952 = ~w25950 & ~w25951;
assign w25953 = ~w16905 & w19930;
assign w25954 = pi04045 & ~w25953;
assign w25955 = ~pi02711 & w25953;
assign w25956 = ~w25954 & ~w25955;
assign w25957 = pi04046 & ~w25953;
assign w25958 = ~pi02170 & w25953;
assign w25959 = ~w25957 & ~w25958;
assign w25960 = pi04047 & ~w25953;
assign w25961 = w17929 & w19930;
assign w25962 = ~w25960 & ~w25961;
assign w25963 = pi04048 & ~w25953;
assign w25964 = ~pi02714 & w25953;
assign w25965 = ~w25963 & ~w25964;
assign w25966 = pi04049 & ~w25953;
assign w25967 = ~pi02715 & w25953;
assign w25968 = ~w25966 & ~w25967;
assign w25969 = pi04050 & ~w25953;
assign w25970 = ~pi02716 & w25953;
assign w25971 = ~w25969 & ~w25970;
assign w25972 = pi04051 & ~w25953;
assign w25973 = ~pi02717 & w25953;
assign w25974 = ~w25972 & ~w25973;
assign w25975 = ~w16905 & w19909;
assign w25976 = pi04052 & ~w25975;
assign w25977 = ~pi02711 & w25975;
assign w25978 = ~w25976 & ~w25977;
assign w25979 = pi04053 & ~w25975;
assign w25980 = ~pi02170 & w25975;
assign w25981 = ~w25979 & ~w25980;
assign w25982 = pi04054 & ~w25975;
assign w25983 = ~pi02713 & w25975;
assign w25984 = ~w25982 & ~w25983;
assign w25985 = pi04055 & ~w25975;
assign w25986 = ~pi02714 & w25975;
assign w25987 = ~w25985 & ~w25986;
assign w25988 = pi04056 & ~w25975;
assign w25989 = ~pi02716 & w25975;
assign w25990 = ~w25988 & ~w25989;
assign w25991 = pi04057 & ~w25975;
assign w25992 = w16973 & w19909;
assign w25993 = ~w25991 & ~w25992;
assign w25994 = ~w16992 & w20075;
assign w25995 = pi04058 & ~w25994;
assign w25996 = ~pi02703 & w25994;
assign w25997 = ~w25995 & ~w25996;
assign w25998 = pi04059 & ~w25994;
assign w25999 = ~pi02169 & w25994;
assign w26000 = ~w25998 & ~w25999;
assign w26001 = pi04060 & ~w25994;
assign w26002 = ~pi02718 & w25994;
assign w26003 = ~w26001 & ~w26002;
assign w26004 = pi04061 & ~w25994;
assign w26005 = ~pi02167 & w25994;
assign w26006 = ~w26004 & ~w26005;
assign w26007 = pi04062 & ~w25994;
assign w26008 = ~pi02164 & w25994;
assign w26009 = ~w26007 & ~w26008;
assign w26010 = pi04063 & ~w25994;
assign w26011 = ~pi02722 & w25994;
assign w26012 = ~w26010 & ~w26011;
assign w26013 = pi04064 & ~w25994;
assign w26014 = ~pi02719 & w25994;
assign w26015 = ~w26013 & ~w26014;
assign w26016 = ~w16992 & w20059;
assign w26017 = pi04065 & ~w26016;
assign w26018 = ~pi02703 & w26016;
assign w26019 = ~w26017 & ~w26018;
assign w26020 = pi04066 & ~w26016;
assign w26021 = ~pi02169 & w26016;
assign w26022 = ~w26020 & ~w26021;
assign w26023 = pi04067 & ~w26016;
assign w26024 = ~pi02718 & w26016;
assign w26025 = ~w26023 & ~w26024;
assign w26026 = pi04068 & ~w26016;
assign w26027 = ~pi02167 & w26016;
assign w26028 = ~w26026 & ~w26027;
assign w26029 = pi04069 & ~w26016;
assign w26030 = ~pi02722 & w26016;
assign w26031 = ~w26029 & ~w26030;
assign w26032 = pi04070 & ~w26016;
assign w26033 = ~pi02719 & w26016;
assign w26034 = ~w26032 & ~w26033;
assign w26035 = ~w16992 & w20014;
assign w26036 = pi04071 & ~w26035;
assign w26037 = ~pi02703 & w26035;
assign w26038 = ~w26036 & ~w26037;
assign w26039 = pi04072 & ~w26035;
assign w26040 = ~pi02169 & w26035;
assign w26041 = ~w26039 & ~w26040;
assign w26042 = pi04073 & ~w26035;
assign w26043 = ~pi02718 & w26035;
assign w26044 = ~w26042 & ~w26043;
assign w26045 = pi04074 & ~w26035;
assign w26046 = ~pi02167 & w26035;
assign w26047 = ~w26045 & ~w26046;
assign w26048 = pi04075 & ~w26035;
assign w26049 = ~pi02164 & w26035;
assign w26050 = ~w26048 & ~w26049;
assign w26051 = pi04076 & ~w26035;
assign w26052 = ~pi02722 & w26035;
assign w26053 = ~w26051 & ~w26052;
assign w26054 = pi04077 & ~w26035;
assign w26055 = ~pi02719 & w26035;
assign w26056 = ~w26054 & ~w26055;
assign w26057 = ~w16905 & w19852;
assign w26058 = pi04078 & ~w26057;
assign w26059 = ~pi02711 & w26057;
assign w26060 = ~w26058 & ~w26059;
assign w26061 = pi04079 & ~w26057;
assign w26062 = ~pi02170 & w26057;
assign w26063 = ~w26061 & ~w26062;
assign w26064 = pi04080 & ~w26057;
assign w26065 = ~pi02713 & w26057;
assign w26066 = ~w26064 & ~w26065;
assign w26067 = pi04081 & ~w26057;
assign w26068 = ~pi02714 & w26057;
assign w26069 = ~w26067 & ~w26068;
assign w26070 = pi04082 & ~w26057;
assign w26071 = ~pi02716 & w26057;
assign w26072 = ~w26070 & ~w26071;
assign w26073 = pi04083 & ~w26057;
assign w26074 = ~pi02717 & w26057;
assign w26075 = ~w26073 & ~w26074;
assign w26076 = ~w16905 & w19838;
assign w26077 = pi04084 & ~w26076;
assign w26078 = ~pi02711 & w26076;
assign w26079 = ~w26077 & ~w26078;
assign w26080 = pi04085 & ~w26076;
assign w26081 = ~pi02170 & w26076;
assign w26082 = ~w26080 & ~w26081;
assign w26083 = pi04086 & ~w26076;
assign w26084 = ~pi02713 & w26076;
assign w26085 = ~w26083 & ~w26084;
assign w26086 = pi04087 & ~w26076;
assign w26087 = ~pi02714 & w26076;
assign w26088 = ~w26086 & ~w26087;
assign w26089 = pi04088 & ~w26076;
assign w26090 = w18059 & w19838;
assign w26091 = ~w26089 & ~w26090;
assign w26092 = pi04089 & ~w26076;
assign w26093 = ~pi02716 & w26076;
assign w26094 = ~w26092 & ~w26093;
assign w26095 = pi04090 & ~w26076;
assign w26096 = ~pi02717 & w26076;
assign w26097 = ~w26095 & ~w26096;
assign w26098 = ~w16992 & w19988;
assign w26099 = pi04091 & ~w26098;
assign w26100 = ~pi02703 & w26098;
assign w26101 = ~w26099 & ~w26100;
assign w26102 = ~w16905 & w19826;
assign w26103 = pi04092 & ~w26102;
assign w26104 = ~pi02711 & w26102;
assign w26105 = ~w26103 & ~w26104;
assign w26106 = pi04093 & ~w26102;
assign w26107 = ~pi02712 & w26102;
assign w26108 = ~w26106 & ~w26107;
assign w26109 = pi04094 & ~w26102;
assign w26110 = w19826 & w20209;
assign w26111 = ~w26109 & ~w26110;
assign w26112 = pi04095 & ~w26102;
assign w26113 = w17742 & w19826;
assign w26114 = ~w26112 & ~w26113;
assign w26115 = pi04096 & ~w26098;
assign w26116 = ~pi02169 & w26098;
assign w26117 = ~w26115 & ~w26116;
assign w26118 = pi04097 & ~w26098;
assign w26119 = ~pi02718 & w26098;
assign w26120 = ~w26118 & ~w26119;
assign w26121 = pi04098 & ~w26102;
assign w26122 = ~pi02716 & w26102;
assign w26123 = ~w26121 & ~w26122;
assign w26124 = pi04099 & ~w26098;
assign w26125 = ~pi02167 & w26098;
assign w26126 = ~w26124 & ~w26125;
assign w26127 = pi04100 & ~w26102;
assign w26128 = ~pi02717 & w26102;
assign w26129 = ~w26127 & ~w26128;
assign w26130 = pi04101 & ~w26098;
assign w26131 = ~pi02164 & w26098;
assign w26132 = ~w26130 & ~w26131;
assign w26133 = pi04102 & ~w26098;
assign w26134 = ~pi02722 & w26098;
assign w26135 = ~w26133 & ~w26134;
assign w26136 = pi04103 & ~w26098;
assign w26137 = ~pi02719 & w26098;
assign w26138 = ~w26136 & ~w26137;
assign w26139 = ~w16905 & w19818;
assign w26140 = pi04104 & ~w26139;
assign w26141 = ~pi02711 & w26139;
assign w26142 = ~w26140 & ~w26141;
assign w26143 = pi04105 & ~w26139;
assign w26144 = ~pi02170 & w26139;
assign w26145 = ~w26143 & ~w26144;
assign w26146 = pi04106 & ~w26139;
assign w26147 = w17929 & w19818;
assign w26148 = ~w26146 & ~w26147;
assign w26149 = pi04107 & ~w26139;
assign w26150 = ~pi02714 & w26139;
assign w26151 = ~w26149 & ~w26150;
assign w26152 = pi04108 & ~w26139;
assign w26153 = ~pi02716 & w26139;
assign w26154 = ~w26152 & ~w26153;
assign w26155 = pi04109 & ~w26139;
assign w26156 = ~pi02717 & w26139;
assign w26157 = ~w26155 & ~w26156;
assign w26158 = ~w16992 & w19941;
assign w26159 = pi04110 & ~w26158;
assign w26160 = w17532 & w19941;
assign w26161 = ~w26159 & ~w26160;
assign w26162 = ~w16905 & w17167;
assign w26163 = pi04111 & ~w26162;
assign w26164 = ~pi02714 & w26162;
assign w26165 = ~w26163 & ~w26164;
assign w26166 = pi04112 & ~w26158;
assign w26167 = ~pi02169 & w26158;
assign w26168 = ~w26166 & ~w26167;
assign w26169 = pi04113 & ~w26158;
assign w26170 = ~pi02718 & w26158;
assign w26171 = ~w26169 & ~w26170;
assign w26172 = pi04114 & ~w26158;
assign w26173 = w19273 & w19941;
assign w26174 = ~w26172 & ~w26173;
assign w26175 = pi04115 & ~w26158;
assign w26176 = w17620 & w19941;
assign w26177 = ~w26175 & ~w26176;
assign w26178 = pi04116 & ~w26158;
assign w26179 = w19312 & w19941;
assign w26180 = ~w26178 & ~w26179;
assign w26181 = pi04117 & ~w26158;
assign w26182 = w17594 & w19941;
assign w26183 = ~w26181 & ~w26182;
assign w26184 = ~w16905 & w19740;
assign w26185 = pi04118 & ~w26184;
assign w26186 = w17603 & w19740;
assign w26187 = ~w26185 & ~w26186;
assign w26188 = pi04119 & ~w26184;
assign w26189 = ~pi02170 & w26184;
assign w26190 = ~w26188 & ~w26189;
assign w26191 = pi04120 & ~w26184;
assign w26192 = ~pi02713 & w26184;
assign w26193 = ~w26191 & ~w26192;
assign w26194 = pi04121 & ~w26184;
assign w26195 = w17742 & w19740;
assign w26196 = ~w26194 & ~w26195;
assign w26197 = pi04122 & ~w26184;
assign w26198 = ~pi02716 & w26184;
assign w26199 = ~w26197 & ~w26198;
assign w26200 = pi04123 & ~w26184;
assign w26201 = ~pi02717 & w26184;
assign w26202 = ~w26200 & ~w26201;
assign w26203 = pi04124 & ~w22121;
assign w26204 = w17603 & w19728;
assign w26205 = ~w26203 & ~w26204;
assign w26206 = pi04125 & ~w22121;
assign w26207 = ~pi02170 & w22121;
assign w26208 = ~w26206 & ~w26207;
assign w26209 = pi04126 & ~w22121;
assign w26210 = ~pi02713 & w22121;
assign w26211 = ~w26209 & ~w26210;
assign w26212 = pi04127 & ~w22121;
assign w26213 = ~pi02714 & w22121;
assign w26214 = ~w26212 & ~w26213;
assign w26215 = pi04128 & ~w22121;
assign w26216 = ~pi02715 & w22121;
assign w26217 = ~w26215 & ~w26216;
assign w26218 = pi04129 & ~w22121;
assign w26219 = w17317 & w19728;
assign w26220 = ~w26218 & ~w26219;
assign w26221 = pi04130 & ~w22121;
assign w26222 = ~pi02717 & w22121;
assign w26223 = ~w26221 & ~w26222;
assign w26224 = pi04131 & ~w22111;
assign w26225 = w17603 & w19723;
assign w26226 = ~w26224 & ~w26225;
assign w26227 = pi04132 & ~w22111;
assign w26228 = ~pi02170 & w22111;
assign w26229 = ~w26227 & ~w26228;
assign w26230 = pi04133 & ~w22111;
assign w26231 = ~pi02713 & w22111;
assign w26232 = ~w26230 & ~w26231;
assign w26233 = pi04134 & ~w22111;
assign w26234 = ~pi02714 & w22111;
assign w26235 = ~w26233 & ~w26234;
assign w26236 = pi04135 & ~w22111;
assign w26237 = ~pi02716 & w22111;
assign w26238 = ~w26236 & ~w26237;
assign w26239 = pi04136 & ~w22111;
assign w26240 = ~pi02717 & w22111;
assign w26241 = ~w26239 & ~w26240;
assign w26242 = pi04137 & ~w22107;
assign w26243 = ~pi02711 & w22107;
assign w26244 = ~w26242 & ~w26243;
assign w26245 = pi04138 & ~w22107;
assign w26246 = ~pi02170 & w22107;
assign w26247 = ~w26245 & ~w26246;
assign w26248 = pi04139 & ~w22107;
assign w26249 = w17929 & w19660;
assign w26250 = ~w26248 & ~w26249;
assign w26251 = pi04140 & ~w22107;
assign w26252 = ~pi02714 & w22107;
assign w26253 = ~w26251 & ~w26252;
assign w26254 = pi04141 & ~w22107;
assign w26255 = w18059 & w19660;
assign w26256 = ~w26254 & ~w26255;
assign w26257 = pi04142 & ~w22107;
assign w26258 = ~pi02716 & w22107;
assign w26259 = ~w26257 & ~w26258;
assign w26260 = pi04143 & ~w22107;
assign w26261 = ~pi02717 & w22107;
assign w26262 = ~w26260 & ~w26261;
assign w26263 = pi04144 & ~w22100;
assign w26264 = w17603 & w19679;
assign w26265 = ~w26263 & ~w26264;
assign w26266 = pi04145 & ~w22100;
assign w26267 = ~pi02170 & w22100;
assign w26268 = ~w26266 & ~w26267;
assign w26269 = pi04146 & ~w22100;
assign w26270 = ~pi02713 & w22100;
assign w26271 = ~w26269 & ~w26270;
assign w26272 = pi04147 & ~w22100;
assign w26273 = ~pi02714 & w22100;
assign w26274 = ~w26272 & ~w26273;
assign w26275 = pi04148 & ~w22100;
assign w26276 = ~pi02716 & w22100;
assign w26277 = ~w26275 & ~w26276;
assign w26278 = pi04149 & ~w22100;
assign w26279 = ~pi02717 & w22100;
assign w26280 = ~w26278 & ~w26279;
assign w26281 = pi04150 & ~w22096;
assign w26282 = w17532 & w19930;
assign w26283 = ~w26281 & ~w26282;
assign w26284 = pi04151 & ~w22096;
assign w26285 = ~pi02169 & w22096;
assign w26286 = ~w26284 & ~w26285;
assign w26287 = pi04152 & ~w22096;
assign w26288 = ~pi02718 & w22096;
assign w26289 = ~w26287 & ~w26288;
assign w26290 = pi04153 & ~w22096;
assign w26291 = ~pi02167 & w22096;
assign w26292 = ~w26290 & ~w26291;
assign w26293 = pi04154 & ~w22096;
assign w26294 = ~pi02164 & w22096;
assign w26295 = ~w26293 & ~w26294;
assign w26296 = pi04155 & ~w22096;
assign w26297 = w19312 & w19930;
assign w26298 = ~w26296 & ~w26297;
assign w26299 = pi04156 & ~w22096;
assign w26300 = ~pi02719 & w22096;
assign w26301 = ~w26299 & ~w26300;
assign w26302 = pi04157 & ~w22085;
assign w26303 = ~pi02703 & w22085;
assign w26304 = ~w26302 & ~w26303;
assign w26305 = pi04158 & ~w22085;
assign w26306 = ~pi02169 & w22085;
assign w26307 = ~w26305 & ~w26306;
assign w26308 = pi04159 & ~w22085;
assign w26309 = ~pi02718 & w22085;
assign w26310 = ~w26308 & ~w26309;
assign w26311 = pi04160 & ~w22085;
assign w26312 = ~pi02167 & w22085;
assign w26313 = ~w26311 & ~w26312;
assign w26314 = pi04161 & ~w22085;
assign w26315 = ~pi02722 & w22085;
assign w26316 = ~w26314 & ~w26315;
assign w26317 = pi04162 & ~w22085;
assign w26318 = ~pi02719 & w22085;
assign w26319 = ~w26317 & ~w26318;
assign w26320 = pi04163 & ~w22089;
assign w26321 = ~pi02711 & w22089;
assign w26322 = ~w26320 & ~w26321;
assign w26323 = pi04164 & ~w22089;
assign w26324 = ~pi02170 & w22089;
assign w26325 = ~w26323 & ~w26324;
assign w26326 = pi04165 & ~w22089;
assign w26327 = ~pi02713 & w22089;
assign w26328 = ~w26326 & ~w26327;
assign w26329 = pi04166 & ~w22089;
assign w26330 = w17742 & w19650;
assign w26331 = ~w26329 & ~w26330;
assign w26332 = pi04167 & ~w22089;
assign w26333 = ~pi02715 & w22089;
assign w26334 = ~w26332 & ~w26333;
assign w26335 = pi04168 & ~w22089;
assign w26336 = w17317 & w19650;
assign w26337 = ~w26335 & ~w26336;
assign w26338 = pi04169 & ~w22089;
assign w26339 = ~pi02717 & w22089;
assign w26340 = ~w26338 & ~w26339;
assign w26341 = pi04170 & ~w22078;
assign w26342 = ~pi02711 & w22078;
assign w26343 = ~w26341 & ~w26342;
assign w26344 = pi04171 & ~w22078;
assign w26345 = ~pi02170 & w22078;
assign w26346 = ~w26344 & ~w26345;
assign w26347 = pi04172 & ~w22078;
assign w26348 = ~pi02713 & w22078;
assign w26349 = ~w26347 & ~w26348;
assign w26350 = pi04173 & ~w22078;
assign w26351 = ~pi02714 & w22078;
assign w26352 = ~w26350 & ~w26351;
assign w26353 = pi04174 & ~w22078;
assign w26354 = ~pi02716 & w22078;
assign w26355 = ~w26353 & ~w26354;
assign w26356 = pi04175 & ~w22078;
assign w26357 = ~pi02717 & w22078;
assign w26358 = ~w26356 & ~w26357;
assign w26359 = pi04176 & ~w22071;
assign w26360 = ~pi02711 & w22071;
assign w26361 = ~w26359 & ~w26360;
assign w26362 = pi04177 & ~w24004;
assign w26363 = ~pi09848 & w24004;
assign w26364 = ~w26362 & ~w26363;
assign w26365 = pi04178 & ~w22071;
assign w26366 = ~pi02170 & w22071;
assign w26367 = ~w26365 & ~w26366;
assign w26368 = pi04179 & ~w22071;
assign w26369 = ~pi02713 & w22071;
assign w26370 = ~w26368 & ~w26369;
assign w26371 = pi04180 & ~w22071;
assign w26372 = ~pi02714 & w22071;
assign w26373 = ~w26371 & ~w26372;
assign w26374 = pi04181 & ~w22071;
assign w26375 = ~pi02716 & w22071;
assign w26376 = ~w26374 & ~w26375;
assign w26377 = pi04182 & ~w22071;
assign w26378 = ~pi02717 & w22071;
assign w26379 = ~w26377 & ~w26378;
assign w26380 = pi04183 & ~w22064;
assign w26381 = ~pi02711 & w22064;
assign w26382 = ~w26380 & ~w26381;
assign w26383 = pi04184 & ~w22064;
assign w26384 = w19624 & w20209;
assign w26385 = ~w26383 & ~w26384;
assign w26386 = pi04185 & ~w22064;
assign w26387 = w17929 & w19624;
assign w26388 = ~w26386 & ~w26387;
assign w26389 = pi04186 & ~w22064;
assign w26390 = ~pi02714 & w22064;
assign w26391 = ~w26389 & ~w26390;
assign w26392 = pi04187 & ~w22064;
assign w26393 = ~pi02716 & w22064;
assign w26394 = ~w26392 & ~w26393;
assign w26395 = pi04188 & ~w22064;
assign w26396 = ~pi02717 & w22064;
assign w26397 = ~w26395 & ~w26396;
assign w26398 = pi04189 & ~w22060;
assign w26399 = ~pi02711 & w22060;
assign w26400 = ~w26398 & ~w26399;
assign w26401 = pi04190 & ~w22060;
assign w26402 = ~pi02170 & w22060;
assign w26403 = ~w26401 & ~w26402;
assign w26404 = pi04191 & ~w22060;
assign w26405 = ~pi02713 & w22060;
assign w26406 = ~w26404 & ~w26405;
assign w26407 = pi04192 & ~w22060;
assign w26408 = ~pi02714 & w22060;
assign w26409 = ~w26407 & ~w26408;
assign w26410 = pi04193 & ~w22060;
assign w26411 = w18059 & w19606;
assign w26412 = ~w26410 & ~w26411;
assign w26413 = pi04194 & ~w22060;
assign w26414 = ~pi02716 & w22060;
assign w26415 = ~w26413 & ~w26414;
assign w26416 = pi04195 & ~w22060;
assign w26417 = ~pi02717 & w22060;
assign w26418 = ~w26416 & ~w26417;
assign w26419 = pi04196 & ~w21610;
assign w26420 = ~pi02711 & w21610;
assign w26421 = ~w26419 & ~w26420;
assign w26422 = pi04197 & ~w21610;
assign w26423 = ~pi02170 & w21610;
assign w26424 = ~w26422 & ~w26423;
assign w26425 = pi04198 & ~w21610;
assign w26426 = ~pi02713 & w21610;
assign w26427 = ~w26425 & ~w26426;
assign w26428 = pi04199 & ~w21610;
assign w26429 = w17742 & w19601;
assign w26430 = ~w26428 & ~w26429;
assign w26431 = pi04200 & ~w21610;
assign w26432 = ~pi02716 & w21610;
assign w26433 = ~w26431 & ~w26432;
assign w26434 = pi04201 & ~w21610;
assign w26435 = ~pi02717 & w21610;
assign w26436 = ~w26434 & ~w26435;
assign w26437 = pi04202 & ~w22031;
assign w26438 = ~pi02711 & w22031;
assign w26439 = ~w26437 & ~w26438;
assign w26440 = pi04203 & ~w22031;
assign w26441 = w19561 & w20209;
assign w26442 = ~w26440 & ~w26441;
assign w26443 = pi04204 & ~w22031;
assign w26444 = ~pi02713 & w22031;
assign w26445 = ~w26443 & ~w26444;
assign w26446 = pi04205 & ~w22031;
assign w26447 = ~pi02714 & w22031;
assign w26448 = ~w26446 & ~w26447;
assign w26449 = pi04206 & ~w22031;
assign w26450 = ~pi02715 & w22031;
assign w26451 = ~w26449 & ~w26450;
assign w26452 = pi04207 & ~w22031;
assign w26453 = ~pi02716 & w22031;
assign w26454 = ~w26452 & ~w26453;
assign w26455 = pi04208 & ~w22031;
assign w26456 = ~pi02717 & w22031;
assign w26457 = ~w26455 & ~w26456;
assign w26458 = pi04209 & ~w22046;
assign w26459 = w17603 & w19552;
assign w26460 = ~w26458 & ~w26459;
assign w26461 = pi04210 & ~w22046;
assign w26462 = ~pi02170 & w22046;
assign w26463 = ~w26461 & ~w26462;
assign w26464 = pi04211 & ~w22046;
assign w26465 = ~pi02713 & w22046;
assign w26466 = ~w26464 & ~w26465;
assign w26467 = pi04212 & ~w22046;
assign w26468 = w17742 & w19552;
assign w26469 = ~w26467 & ~w26468;
assign w26470 = pi04213 & ~w22046;
assign w26471 = ~pi02716 & w22046;
assign w26472 = ~w26470 & ~w26471;
assign w26473 = pi04214 & ~w22046;
assign w26474 = ~pi02717 & w22046;
assign w26475 = ~w26473 & ~w26474;
assign w26476 = pi04215 & ~w22042;
assign w26477 = ~pi02711 & w22042;
assign w26478 = ~w26476 & ~w26477;
assign w26479 = pi04216 & ~w22042;
assign w26480 = ~pi02170 & w22042;
assign w26481 = ~w26479 & ~w26480;
assign w26482 = pi04217 & ~w22042;
assign w26483 = ~pi02713 & w22042;
assign w26484 = ~w26482 & ~w26483;
assign w26485 = pi04218 & ~w22042;
assign w26486 = ~pi02714 & w22042;
assign w26487 = ~w26485 & ~w26486;
assign w26488 = pi04219 & ~w22042;
assign w26489 = ~pi02715 & w22042;
assign w26490 = ~w26488 & ~w26489;
assign w26491 = pi04220 & ~w22042;
assign w26492 = w17317 & w19435;
assign w26493 = ~w26491 & ~w26492;
assign w26494 = pi04221 & ~w22042;
assign w26495 = ~pi02717 & w22042;
assign w26496 = ~w26494 & ~w26495;
assign w26497 = pi04222 & ~w22035;
assign w26498 = ~pi02711 & w22035;
assign w26499 = ~w26497 & ~w26498;
assign w26500 = pi04223 & ~w22035;
assign w26501 = ~pi02170 & w22035;
assign w26502 = ~w26500 & ~w26501;
assign w26503 = pi04224 & ~w22035;
assign w26504 = ~pi02713 & w22035;
assign w26505 = ~w26503 & ~w26504;
assign w26506 = pi04225 & ~w22035;
assign w26507 = ~pi02714 & w22035;
assign w26508 = ~w26506 & ~w26507;
assign w26509 = pi04226 & ~w22035;
assign w26510 = ~pi02716 & w22035;
assign w26511 = ~w26509 & ~w26510;
assign w26512 = pi04227 & ~w22035;
assign w26513 = ~pi02717 & w22035;
assign w26514 = ~w26512 & ~w26513;
assign w26515 = pi04228 & ~w22020;
assign w26516 = ~pi02711 & w22020;
assign w26517 = ~w26515 & ~w26516;
assign w26518 = pi04229 & ~w22020;
assign w26519 = ~pi02170 & w22020;
assign w26520 = ~w26518 & ~w26519;
assign w26521 = pi04230 & ~w22020;
assign w26522 = ~pi02713 & w22020;
assign w26523 = ~w26521 & ~w26522;
assign w26524 = pi04231 & ~w22020;
assign w26525 = ~pi02714 & w22020;
assign w26526 = ~w26524 & ~w26525;
assign w26527 = pi04232 & ~w22020;
assign w26528 = ~pi02715 & w22020;
assign w26529 = ~w26527 & ~w26528;
assign w26530 = pi04233 & ~w22020;
assign w26531 = ~pi02716 & w22020;
assign w26532 = ~w26530 & ~w26531;
assign w26533 = pi04234 & ~w22020;
assign w26534 = ~pi02717 & w22020;
assign w26535 = ~w26533 & ~w26534;
assign w26536 = pi04235 & ~w22024;
assign w26537 = w17532 & w19852;
assign w26538 = ~w26536 & ~w26537;
assign w26539 = pi04236 & ~w22024;
assign w26540 = w19797 & w19852;
assign w26541 = ~w26539 & ~w26540;
assign w26542 = pi04237 & ~w22024;
assign w26543 = ~pi02718 & w22024;
assign w26544 = ~w26542 & ~w26543;
assign w26545 = pi04238 & ~w22009;
assign w26546 = ~pi02711 & w22009;
assign w26547 = ~w26545 & ~w26546;
assign w26548 = pi04239 & ~w22009;
assign w26549 = ~pi02712 & w22009;
assign w26550 = ~w26548 & ~w26549;
assign w26551 = pi04240 & ~w22009;
assign w26552 = ~pi02170 & w22009;
assign w26553 = ~w26551 & ~w26552;
assign w26554 = pi04241 & ~w22024;
assign w26555 = ~pi02164 & w22024;
assign w26556 = ~w26554 & ~w26555;
assign w26557 = pi04242 & ~w22009;
assign w26558 = w17742 & w19492;
assign w26559 = ~w26557 & ~w26558;
assign w26560 = pi04243 & ~w22024;
assign w26561 = ~pi02722 & w22024;
assign w26562 = ~w26560 & ~w26561;
assign w26563 = pi04244 & ~w22009;
assign w26564 = ~pi02715 & w22009;
assign w26565 = ~w26563 & ~w26564;
assign w26566 = pi04245 & ~w22009;
assign w26567 = w17317 & w19492;
assign w26568 = ~w26566 & ~w26567;
assign w26569 = pi04246 & ~w22024;
assign w26570 = ~pi02719 & w22024;
assign w26571 = ~w26569 & ~w26570;
assign w26572 = pi04247 & ~w22009;
assign w26573 = ~pi02717 & w22009;
assign w26574 = ~w26572 & ~w26573;
assign w26575 = pi04248 & ~w22013;
assign w26576 = w17603 & w19480;
assign w26577 = ~w26575 & ~w26576;
assign w26578 = pi04249 & ~w22013;
assign w26579 = w19480 & w20209;
assign w26580 = ~w26578 & ~w26579;
assign w26581 = pi04250 & ~w22013;
assign w26582 = ~pi02713 & w22013;
assign w26583 = ~w26581 & ~w26582;
assign w26584 = pi04251 & ~w22013;
assign w26585 = w17742 & w19480;
assign w26586 = ~w26584 & ~w26585;
assign w26587 = pi04252 & ~w22013;
assign w26588 = ~pi02716 & w22013;
assign w26589 = ~w26587 & ~w26588;
assign w26590 = pi04253 & ~w22013;
assign w26591 = w16973 & w19480;
assign w26592 = ~w26590 & ~w26591;
assign w26593 = pi04254 & ~w21998;
assign w26594 = w17532 & w19838;
assign w26595 = ~w26593 & ~w26594;
assign w26596 = pi04255 & ~w21998;
assign w26597 = ~pi02169 & w21998;
assign w26598 = ~w26596 & ~w26597;
assign w26599 = pi04256 & ~w21998;
assign w26600 = ~pi02718 & w21998;
assign w26601 = ~w26599 & ~w26600;
assign w26602 = pi04257 & ~w21209;
assign w26603 = ~pi02711 & w21209;
assign w26604 = ~w26602 & ~w26603;
assign w26605 = pi04258 & ~w21998;
assign w26606 = ~pi02167 & w21998;
assign w26607 = ~w26605 & ~w26606;
assign w26608 = pi04259 & ~w21209;
assign w26609 = ~pi02712 & w21209;
assign w26610 = ~w26608 & ~w26609;
assign w26611 = pi04260 & ~w21209;
assign w26612 = ~pi02170 & w21209;
assign w26613 = ~w26611 & ~w26612;
assign w26614 = pi04261 & ~w21998;
assign w26615 = ~pi02164 & w21998;
assign w26616 = ~w26614 & ~w26615;
assign w26617 = pi04262 & ~w21209;
assign w26618 = w17742 & w19459;
assign w26619 = ~w26617 & ~w26618;
assign w26620 = pi04263 & ~w21998;
assign w26621 = ~pi02722 & w21998;
assign w26622 = ~w26620 & ~w26621;
assign w26623 = pi04264 & ~w21209;
assign w26624 = ~pi02715 & w21209;
assign w26625 = ~w26623 & ~w26624;
assign w26626 = pi04265 & ~w21998;
assign w26627 = ~pi02719 & w21998;
assign w26628 = ~w26626 & ~w26627;
assign w26629 = pi04266 & ~w21209;
assign w26630 = ~pi02717 & w21209;
assign w26631 = ~w26629 & ~w26630;
assign w26632 = pi04267 & ~w21436;
assign w26633 = ~pi02711 & w21436;
assign w26634 = ~w26632 & ~w26633;
assign w26635 = ~w16992 & w18662;
assign w26636 = pi04268 & ~w26635;
assign w26637 = w18662 & w19273;
assign w26638 = ~w26636 & ~w26637;
assign w26639 = pi04269 & ~w21436;
assign w26640 = ~pi02170 & w21436;
assign w26641 = ~w26639 & ~w26640;
assign w26642 = pi04270 & ~w21436;
assign w26643 = ~pi02713 & w21436;
assign w26644 = ~w26642 & ~w26643;
assign w26645 = pi04271 & ~w21436;
assign w26646 = ~pi02714 & w21436;
assign w26647 = ~w26645 & ~w26646;
assign w26648 = pi04272 & ~w21436;
assign w26649 = ~pi02715 & w21436;
assign w26650 = ~w26648 & ~w26649;
assign w26651 = pi04273 & ~w21436;
assign w26652 = ~pi02716 & w21436;
assign w26653 = ~w26651 & ~w26652;
assign w26654 = pi04274 & ~w21436;
assign w26655 = ~pi02717 & w21436;
assign w26656 = ~w26654 & ~w26655;
assign w26657 = pi04275 & ~w21418;
assign w26658 = ~pi02711 & w21418;
assign w26659 = ~w26657 & ~w26658;
assign w26660 = pi04276 & ~w21425;
assign w26661 = ~pi02703 & w21425;
assign w26662 = ~w26660 & ~w26661;
assign w26663 = pi04277 & ~w21418;
assign w26664 = ~pi02170 & w21418;
assign w26665 = ~w26663 & ~w26664;
assign w26666 = pi04278 & ~w21418;
assign w26667 = w17929 & w19444;
assign w26668 = ~w26666 & ~w26667;
assign w26669 = pi04279 & ~w21418;
assign w26670 = ~pi02714 & w21418;
assign w26671 = ~w26669 & ~w26670;
assign w26672 = pi04280 & ~w21418;
assign w26673 = w18059 & w19444;
assign w26674 = ~w26672 & ~w26673;
assign w26675 = pi04281 & ~w21425;
assign w26676 = w19797 & w19826;
assign w26677 = ~w26675 & ~w26676;
assign w26678 = pi04282 & ~w21418;
assign w26679 = ~pi02717 & w21418;
assign w26680 = ~w26678 & ~w26679;
assign w26681 = pi04283 & ~w20879;
assign w26682 = ~pi02711 & w20879;
assign w26683 = ~w26681 & ~w26682;
assign w26684 = pi04284 & ~w21425;
assign w26685 = ~pi02718 & w21425;
assign w26686 = ~w26684 & ~w26685;
assign w26687 = pi04285 & ~w20879;
assign w26688 = w17020 & w19327;
assign w26689 = ~w26687 & ~w26688;
assign w26690 = pi04286 & ~w21425;
assign w26691 = ~pi02167 & w21425;
assign w26692 = ~w26690 & ~w26691;
assign w26693 = pi04287 & ~w20879;
assign w26694 = ~pi02170 & w20879;
assign w26695 = ~w26693 & ~w26694;
assign w26696 = pi04288 & ~w20879;
assign w26697 = ~pi02713 & w20879;
assign w26698 = ~w26696 & ~w26697;
assign w26699 = pi04289 & ~w21425;
assign w26700 = ~pi02164 & w21425;
assign w26701 = ~w26699 & ~w26700;
assign w26702 = pi04290 & ~w21425;
assign w26703 = ~pi02722 & w21425;
assign w26704 = ~w26702 & ~w26703;
assign w26705 = pi04291 & ~w20879;
assign w26706 = ~pi02715 & w20879;
assign w26707 = ~w26705 & ~w26706;
assign w26708 = pi04292 & ~w21425;
assign w26709 = ~pi02719 & w21425;
assign w26710 = ~w26708 & ~w26709;
assign w26711 = pi04293 & ~w20879;
assign w26712 = ~pi02717 & w20879;
assign w26713 = ~w26711 & ~w26712;
assign w26714 = pi04294 & ~w21084;
assign w26715 = ~pi02711 & w21084;
assign w26716 = ~w26714 & ~w26715;
assign w26717 = pi04295 & ~w21084;
assign w26718 = w19591 & w20209;
assign w26719 = ~w26717 & ~w26718;
assign w26720 = pi04296 & ~w21084;
assign w26721 = ~pi02713 & w21084;
assign w26722 = ~w26720 & ~w26721;
assign w26723 = pi04297 & ~w21084;
assign w26724 = ~pi02714 & w21084;
assign w26725 = ~w26723 & ~w26724;
assign w26726 = pi04298 & ~w21084;
assign w26727 = ~pi02715 & w21084;
assign w26728 = ~w26726 & ~w26727;
assign w26729 = pi04299 & ~w21084;
assign w26730 = w17317 & w19591;
assign w26731 = ~w26729 & ~w26730;
assign w26732 = pi04300 & ~w21084;
assign w26733 = ~pi02717 & w21084;
assign w26734 = ~w26732 & ~w26733;
assign w26735 = pi04301 & ~w20891;
assign w26736 = ~pi02711 & w20891;
assign w26737 = ~w26735 & ~w26736;
assign w26738 = pi04302 & ~w21026;
assign w26739 = w17532 & w19818;
assign w26740 = ~w26738 & ~w26739;
assign w26741 = pi04303 & ~w20891;
assign w26742 = ~pi02170 & w20891;
assign w26743 = ~w26741 & ~w26742;
assign w26744 = pi04304 & ~w20891;
assign w26745 = ~pi02713 & w20891;
assign w26746 = ~w26744 & ~w26745;
assign w26747 = pi04305 & ~w20891;
assign w26748 = ~pi02714 & w20891;
assign w26749 = ~w26747 & ~w26748;
assign w26750 = pi04306 & ~w20891;
assign w26751 = ~pi02715 & w20891;
assign w26752 = ~w26750 & ~w26751;
assign w26753 = pi04307 & ~w21026;
assign w26754 = w19797 & w19818;
assign w26755 = ~w26753 & ~w26754;
assign w26756 = pi04308 & ~w20891;
assign w26757 = ~pi02717 & w20891;
assign w26758 = ~w26756 & ~w26757;
assign w26759 = pi04309 & ~w20604;
assign w26760 = ~pi02711 & w20604;
assign w26761 = ~w26759 & ~w26760;
assign w26762 = pi04310 & ~w21026;
assign w26763 = ~pi02718 & w21026;
assign w26764 = ~w26762 & ~w26763;
assign w26765 = pi04311 & ~w20604;
assign w26766 = ~pi02712 & w20604;
assign w26767 = ~w26765 & ~w26766;
assign w26768 = pi04312 & ~w20604;
assign w26769 = ~pi02170 & w20604;
assign w26770 = ~w26768 & ~w26769;
assign w26771 = pi04313 & ~w21026;
assign w26772 = ~pi02167 & w21026;
assign w26773 = ~w26771 & ~w26772;
assign w26774 = pi04314 & ~w20604;
assign w26775 = ~pi02713 & w20604;
assign w26776 = ~w26774 & ~w26775;
assign w26777 = pi04315 & ~w21026;
assign w26778 = ~pi02164 & w21026;
assign w26779 = ~w26777 & ~w26778;
assign w26780 = pi04316 & ~w20604;
assign w26781 = ~pi02715 & w20604;
assign w26782 = ~w26780 & ~w26781;
assign w26783 = pi04317 & ~w21026;
assign w26784 = ~pi02722 & w21026;
assign w26785 = ~w26783 & ~w26784;
assign w26786 = pi04318 & ~w21026;
assign w26787 = ~pi02719 & w21026;
assign w26788 = ~w26786 & ~w26787;
assign w26789 = pi04319 & ~w20604;
assign w26790 = ~pi02717 & w20604;
assign w26791 = ~w26789 & ~w26790;
assign w26792 = pi04320 & ~w20633;
assign w26793 = w17603 & w19348;
assign w26794 = ~w26792 & ~w26793;
assign w26795 = pi04321 & ~w25912;
assign w26796 = w18645 & w19797;
assign w26797 = ~w26795 & ~w26796;
assign w26798 = pi04322 & ~w20633;
assign w26799 = w19348 & w20209;
assign w26800 = ~w26798 & ~w26799;
assign w26801 = pi04323 & ~w20633;
assign w26802 = ~pi02713 & w20633;
assign w26803 = ~w26801 & ~w26802;
assign w26804 = pi04324 & ~w20633;
assign w26805 = w17742 & w19348;
assign w26806 = ~w26804 & ~w26805;
assign w26807 = pi04325 & ~w20633;
assign w26808 = w18059 & w19348;
assign w26809 = ~w26807 & ~w26808;
assign w26810 = pi04326 & ~w20633;
assign w26811 = ~pi02716 & w20633;
assign w26812 = ~w26810 & ~w26811;
assign w26813 = pi04327 & ~w20633;
assign w26814 = w16973 & w19348;
assign w26815 = ~w26813 & ~w26814;
assign w26816 = pi04328 & ~w20592;
assign w26817 = ~pi02711 & w20592;
assign w26818 = ~w26816 & ~w26817;
assign w26819 = pi04329 & ~w20592;
assign w26820 = ~pi02713 & w20592;
assign w26821 = ~w26819 & ~w26820;
assign w26822 = pi04330 & ~w20592;
assign w26823 = ~pi02714 & w20592;
assign w26824 = ~w26822 & ~w26823;
assign w26825 = pi04331 & ~w20592;
assign w26826 = ~pi02715 & w20592;
assign w26827 = ~w26825 & ~w26826;
assign w26828 = pi04332 & ~w20592;
assign w26829 = ~pi02717 & w20592;
assign w26830 = ~w26828 & ~w26829;
assign w26831 = pi04333 & ~w20592;
assign w26832 = ~pi02170 & w20592;
assign w26833 = ~w26831 & ~w26832;
assign w26834 = pi04334 & ~w20557;
assign w26835 = w17532 & w19740;
assign w26836 = ~w26834 & ~w26835;
assign w26837 = pi04335 & ~w20557;
assign w26838 = ~pi02169 & w20557;
assign w26839 = ~w26837 & ~w26838;
assign w26840 = pi04336 & ~w20557;
assign w26841 = ~pi02718 & w20557;
assign w26842 = ~w26840 & ~w26841;
assign w26843 = pi04337 & ~w20557;
assign w26844 = ~pi02167 & w20557;
assign w26845 = ~w26843 & ~w26844;
assign w26846 = pi04338 & ~w20557;
assign w26847 = ~pi02164 & w20557;
assign w26848 = ~w26846 & ~w26847;
assign w26849 = pi04339 & ~w20557;
assign w26850 = ~pi02722 & w20557;
assign w26851 = ~w26849 & ~w26850;
assign w26852 = pi04340 & ~w20557;
assign w26853 = ~pi02719 & w20557;
assign w26854 = ~w26852 & ~w26853;
assign w26855 = pi04341 & ~w20497;
assign w26856 = ~pi02703 & w20497;
assign w26857 = ~w26855 & ~w26856;
assign w26858 = pi04342 & ~w20497;
assign w26859 = ~pi02169 & w20497;
assign w26860 = ~w26858 & ~w26859;
assign w26861 = pi04343 & ~w20497;
assign w26862 = ~pi02718 & w20497;
assign w26863 = ~w26861 & ~w26862;
assign w26864 = pi04344 & ~w20497;
assign w26865 = ~pi02167 & w20497;
assign w26866 = ~w26864 & ~w26865;
assign w26867 = pi04345 & ~w20497;
assign w26868 = ~pi02722 & w20497;
assign w26869 = ~w26867 & ~w26868;
assign w26870 = pi04346 & ~w20497;
assign w26871 = ~pi02719 & w20497;
assign w26872 = ~w26870 & ~w26871;
assign w26873 = pi04347 & ~w20253;
assign w26874 = w17532 & w19723;
assign w26875 = ~w26873 & ~w26874;
assign w26876 = pi04348 & ~w20253;
assign w26877 = ~pi02169 & w20253;
assign w26878 = ~w26876 & ~w26877;
assign w26879 = pi04349 & ~w20253;
assign w26880 = ~pi02718 & w20253;
assign w26881 = ~w26879 & ~w26880;
assign w26882 = pi04350 & ~w20253;
assign w26883 = ~pi02167 & w20253;
assign w26884 = ~w26882 & ~w26883;
assign w26885 = pi04351 & ~w20253;
assign w26886 = ~pi02164 & w20253;
assign w26887 = ~w26885 & ~w26886;
assign w26888 = pi04352 & ~w20253;
assign w26889 = ~pi02722 & w20253;
assign w26890 = ~w26888 & ~w26889;
assign w26891 = pi04353 & ~w20253;
assign w26892 = ~pi02719 & w20253;
assign w26893 = ~w26891 & ~w26892;
assign w26894 = pi04354 & ~w20038;
assign w26895 = ~pi02703 & w20038;
assign w26896 = ~w26894 & ~w26895;
assign w26897 = pi04355 & ~w20038;
assign w26898 = ~pi02169 & w20038;
assign w26899 = ~w26897 & ~w26898;
assign w26900 = pi04356 & ~w20038;
assign w26901 = ~pi02718 & w20038;
assign w26902 = ~w26900 & ~w26901;
assign w26903 = pi04357 & ~w20038;
assign w26904 = ~pi02167 & w20038;
assign w26905 = ~w26903 & ~w26904;
assign w26906 = pi04358 & ~w20038;
assign w26907 = ~pi02722 & w20038;
assign w26908 = ~w26906 & ~w26907;
assign w26909 = pi04359 & ~w20038;
assign w26910 = ~pi02719 & w20038;
assign w26911 = ~w26909 & ~w26910;
assign w26912 = pi04360 & ~w20140;
assign w26913 = w17532 & w19679;
assign w26914 = ~w26912 & ~w26913;
assign w26915 = pi04361 & ~w20140;
assign w26916 = ~pi02169 & w20140;
assign w26917 = ~w26915 & ~w26916;
assign w26918 = pi04362 & ~w20140;
assign w26919 = ~pi02718 & w20140;
assign w26920 = ~w26918 & ~w26919;
assign w26921 = pi04363 & ~w20140;
assign w26922 = ~pi02167 & w20140;
assign w26923 = ~w26921 & ~w26922;
assign w26924 = pi04364 & ~w20140;
assign w26925 = ~pi02164 & w20140;
assign w26926 = ~w26924 & ~w26925;
assign w26927 = pi04365 & ~w20140;
assign w26928 = w19312 & w19679;
assign w26929 = ~w26927 & ~w26928;
assign w26930 = pi04366 & ~w20140;
assign w26931 = ~pi02719 & w20140;
assign w26932 = ~w26930 & ~w26931;
assign w26933 = pi04367 & ~w20104;
assign w26934 = w17532 & w19650;
assign w26935 = ~w26933 & ~w26934;
assign w26936 = pi04368 & ~w20104;
assign w26937 = ~pi02169 & w20104;
assign w26938 = ~w26936 & ~w26937;
assign w26939 = pi04369 & ~w20104;
assign w26940 = ~pi02718 & w20104;
assign w26941 = ~w26939 & ~w26940;
assign w26942 = pi04370 & ~w20104;
assign w26943 = w19273 & w19650;
assign w26944 = ~w26942 & ~w26943;
assign w26945 = pi04371 & ~w20104;
assign w26946 = ~pi02722 & w20104;
assign w26947 = ~w26945 & ~w26946;
assign w26948 = pi04372 & ~w20104;
assign w26949 = ~pi02719 & w20104;
assign w26950 = ~w26948 & ~w26949;
assign w26951 = pi04373 & ~w20045;
assign w26952 = ~pi02703 & w20045;
assign w26953 = ~w26951 & ~w26952;
assign w26954 = pi04374 & ~w26635;
assign w26955 = w17532 & w18662;
assign w26956 = ~w26954 & ~w26955;
assign w26957 = pi04375 & ~w20045;
assign w26958 = w17586 & w19645;
assign w26959 = ~w26957 & ~w26958;
assign w26960 = pi04376 & ~w20045;
assign w26961 = ~pi02169 & w20045;
assign w26962 = ~w26960 & ~w26961;
assign w26963 = pi04377 & ~w20045;
assign w26964 = ~pi02167 & w20045;
assign w26965 = ~w26963 & ~w26964;
assign w26966 = pi04378 & ~w20045;
assign w26967 = ~pi02164 & w20045;
assign w26968 = ~w26966 & ~w26967;
assign w26969 = pi04379 & ~w20045;
assign w26970 = ~pi02719 & w20045;
assign w26971 = ~w26969 & ~w26970;
assign w26972 = pi04380 & ~w20045;
assign w26973 = ~pi02722 & w20045;
assign w26974 = ~w26972 & ~w26973;
assign w26975 = pi04381 & ~w20052;
assign w26976 = ~pi02703 & w20052;
assign w26977 = ~w26975 & ~w26976;
assign w26978 = pi04382 & ~w20052;
assign w26979 = ~pi02721 & w20052;
assign w26980 = ~w26978 & ~w26979;
assign w26981 = pi04383 & ~w20052;
assign w26982 = ~pi02169 & w20052;
assign w26983 = ~w26981 & ~w26982;
assign w26984 = pi04384 & ~w20052;
assign w26985 = ~pi02718 & w20052;
assign w26986 = ~w26984 & ~w26985;
assign w26987 = pi04385 & ~w20052;
assign w26988 = ~pi02167 & w20052;
assign w26989 = ~w26987 & ~w26988;
assign w26990 = pi04386 & ~w20052;
assign w26991 = ~pi02722 & w20052;
assign w26992 = ~w26990 & ~w26991;
assign w26993 = pi04387 & ~w20052;
assign w26994 = ~pi02719 & w20052;
assign w26995 = ~w26993 & ~w26994;
assign w26996 = pi04388 & ~w20064;
assign w26997 = w17532 & w19624;
assign w26998 = ~w26996 & ~w26997;
assign w26999 = pi04389 & ~w20064;
assign w27000 = ~pi02718 & w20064;
assign w27001 = ~w26999 & ~w27000;
assign w27002 = pi04390 & ~w20064;
assign w27003 = ~pi02169 & w20064;
assign w27004 = ~w27002 & ~w27003;
assign w27005 = pi04391 & ~w20064;
assign w27006 = ~pi02167 & w20064;
assign w27007 = ~w27005 & ~w27006;
assign w27008 = pi04392 & ~w20064;
assign w27009 = ~pi02164 & w20064;
assign w27010 = ~w27008 & ~w27009;
assign w27011 = pi04393 & ~w20064;
assign w27012 = ~pi02719 & w20064;
assign w27013 = ~w27011 & ~w27012;
assign w27014 = pi04394 & ~w20064;
assign w27015 = ~pi02722 & w20064;
assign w27016 = ~w27014 & ~w27015;
assign w27017 = pi04395 & ~w20007;
assign w27018 = ~pi02703 & w20007;
assign w27019 = ~w27017 & ~w27018;
assign w27020 = pi04396 & ~w20007;
assign w27021 = ~pi02169 & w20007;
assign w27022 = ~w27020 & ~w27021;
assign w27023 = pi04397 & ~w20007;
assign w27024 = w17586 & w19606;
assign w27025 = ~w27023 & ~w27024;
assign w27026 = pi04398 & ~w20007;
assign w27027 = ~pi02167 & w20007;
assign w27028 = ~w27026 & ~w27027;
assign w27029 = pi04399 & ~w20007;
assign w27030 = ~pi02722 & w20007;
assign w27031 = ~w27029 & ~w27030;
assign w27032 = pi04400 & ~w20007;
assign w27033 = ~pi02719 & w20007;
assign w27034 = ~w27032 & ~w27033;
assign w27035 = pi04401 & ~w19978;
assign w27036 = ~pi02703 & w19978;
assign w27037 = ~w27035 & ~w27036;
assign w27038 = ~w16928 & w18217;
assign w27039 = pi04402 & ~w27038;
assign w27040 = ~pi09812 & w27038;
assign w27041 = ~w27039 & ~w27040;
assign w27042 = pi04403 & ~w19978;
assign w27043 = ~pi02169 & w19978;
assign w27044 = ~w27042 & ~w27043;
assign w27045 = pi04404 & ~w19978;
assign w27046 = ~pi02718 & w19978;
assign w27047 = ~w27045 & ~w27046;
assign w27048 = pi04405 & ~w19978;
assign w27049 = ~pi02167 & w19978;
assign w27050 = ~w27048 & ~w27049;
assign w27051 = pi04406 & ~w19978;
assign w27052 = ~pi02164 & w19978;
assign w27053 = ~w27051 & ~w27052;
assign w27054 = pi04407 & ~w19978;
assign w27055 = ~pi02722 & w19978;
assign w27056 = ~w27054 & ~w27055;
assign w27057 = pi04408 & ~w19978;
assign w27058 = ~pi02719 & w19978;
assign w27059 = ~w27057 & ~w27058;
assign w27060 = pi04409 & ~w19922;
assign w27061 = w17532 & w19561;
assign w27062 = ~w27060 & ~w27061;
assign w27063 = pi04410 & ~w19922;
assign w27064 = w19561 & w19797;
assign w27065 = ~w27063 & ~w27064;
assign w27066 = pi04411 & ~w19922;
assign w27067 = w17586 & w19561;
assign w27068 = ~w27066 & ~w27067;
assign w27069 = pi04412 & ~w19922;
assign w27070 = w19273 & w19561;
assign w27071 = ~w27069 & ~w27070;
assign w27072 = pi04413 & ~w19922;
assign w27073 = w19312 & w19561;
assign w27074 = ~w27072 & ~w27073;
assign w27075 = pi04414 & ~w19922;
assign w27076 = w17594 & w19561;
assign w27077 = ~w27075 & ~w27076;
assign w27078 = pi04415 & ~w19946;
assign w27079 = ~pi02703 & w19946;
assign w27080 = ~w27078 & ~w27079;
assign w27081 = pi04416 & ~w19946;
assign w27082 = ~pi02169 & w19946;
assign w27083 = ~w27081 & ~w27082;
assign w27084 = pi04417 & ~w19946;
assign w27085 = ~pi02718 & w19946;
assign w27086 = ~w27084 & ~w27085;
assign w27087 = pi04418 & ~w19946;
assign w27088 = ~pi02167 & w19946;
assign w27089 = ~w27087 & ~w27088;
assign w27090 = pi04419 & ~w19946;
assign w27091 = ~pi02164 & w19946;
assign w27092 = ~w27090 & ~w27091;
assign w27093 = pi04420 & ~w19946;
assign w27094 = ~pi02722 & w19946;
assign w27095 = ~w27093 & ~w27094;
assign w27096 = pi04421 & ~w19946;
assign w27097 = ~pi02719 & w19946;
assign w27098 = ~w27096 & ~w27097;
assign w27099 = pi04422 & ~w19783;
assign w27100 = ~pi02703 & w19783;
assign w27101 = ~w27099 & ~w27100;
assign w27102 = pi04423 & ~w19783;
assign w27103 = ~pi02169 & w19783;
assign w27104 = ~w27102 & ~w27103;
assign w27105 = pi04424 & ~w19783;
assign w27106 = ~pi02718 & w19783;
assign w27107 = ~w27105 & ~w27106;
assign w27108 = pi04425 & ~w19783;
assign w27109 = ~pi02167 & w19783;
assign w27110 = ~w27108 & ~w27109;
assign w27111 = pi04426 & ~w19783;
assign w27112 = w19312 & w19435;
assign w27113 = ~w27111 & ~w27112;
assign w27114 = pi04427 & ~w19783;
assign w27115 = ~pi02719 & w19783;
assign w27116 = ~w27114 & ~w27115;
assign w27117 = pi04428 & ~w19888;
assign w27118 = ~pi02703 & w19888;
assign w27119 = ~w27117 & ~w27118;
assign w27120 = pi04429 & ~w19888;
assign w27121 = ~pi02169 & w19888;
assign w27122 = ~w27120 & ~w27121;
assign w27123 = pi04430 & ~w19888;
assign w27124 = ~pi02718 & w19888;
assign w27125 = ~w27123 & ~w27124;
assign w27126 = pi04431 & ~w19888;
assign w27127 = ~pi02167 & w19888;
assign w27128 = ~w27126 & ~w27127;
assign w27129 = pi04432 & ~w19888;
assign w27130 = ~pi02164 & w19888;
assign w27131 = ~w27129 & ~w27130;
assign w27132 = pi04433 & ~w19888;
assign w27133 = w19312 & w19530;
assign w27134 = ~w27132 & ~w27133;
assign w27135 = pi04434 & ~w19888;
assign w27136 = ~pi02719 & w19888;
assign w27137 = ~w27135 & ~w27136;
assign w27138 = pi04435 & ~w19831;
assign w27139 = ~pi02703 & w19831;
assign w27140 = ~w27138 & ~w27139;
assign w27141 = pi04436 & ~w19831;
assign w27142 = ~pi02169 & w19831;
assign w27143 = ~w27141 & ~w27142;
assign w27144 = pi04437 & ~w19831;
assign w27145 = ~pi02718 & w19831;
assign w27146 = ~w27144 & ~w27145;
assign w27147 = pi04438 & ~w19831;
assign w27148 = ~pi02167 & w19831;
assign w27149 = ~w27147 & ~w27148;
assign w27150 = pi04439 & ~w19831;
assign w27151 = w17594 & w19518;
assign w27152 = ~w27150 & ~w27151;
assign w27153 = pi04440 & ~w19831;
assign w27154 = w19312 & w19518;
assign w27155 = ~w27153 & ~w27154;
assign w27156 = pi04441 & ~w19795;
assign w27157 = w17532 & w19492;
assign w27158 = ~w27156 & ~w27157;
assign w27159 = pi04442 & ~w19795;
assign w27160 = w17811 & w19492;
assign w27161 = ~w27159 & ~w27160;
assign w27162 = pi04443 & ~w19795;
assign w27163 = w17586 & w19492;
assign w27164 = ~w27162 & ~w27163;
assign w27165 = pi04444 & ~w19795;
assign w27166 = w19273 & w19492;
assign w27167 = ~w27165 & ~w27166;
assign w27168 = pi04445 & ~w19795;
assign w27169 = w17620 & w19492;
assign w27170 = ~w27168 & ~w27169;
assign w27171 = pi04446 & ~w19795;
assign w27172 = w19312 & w19492;
assign w27173 = ~w27171 & ~w27172;
assign w27174 = pi04447 & ~w19795;
assign w27175 = w17594 & w19492;
assign w27176 = ~w27174 & ~w27175;
assign w27177 = pi04448 & ~w19690;
assign w27178 = w17532 & w19480;
assign w27179 = ~w27177 & ~w27178;
assign w27180 = pi04449 & ~w19690;
assign w27181 = w19480 & w19797;
assign w27182 = ~w27180 & ~w27181;
assign w27183 = pi04450 & ~w19690;
assign w27184 = ~pi02167 & w19690;
assign w27185 = ~w27183 & ~w27184;
assign w27186 = pi04451 & ~w19690;
assign w27187 = ~pi02718 & w19690;
assign w27188 = ~w27186 & ~w27187;
assign w27189 = pi04452 & ~w19690;
assign w27190 = w19312 & w19480;
assign w27191 = ~w27189 & ~w27190;
assign w27192 = pi04453 & ~w19690;
assign w27193 = ~pi02719 & w19690;
assign w27194 = ~w27192 & ~w27193;
assign w27195 = pi04454 & ~w19755;
assign w27196 = ~pi02721 & w19755;
assign w27197 = ~w27195 & ~w27196;
assign w27198 = pi04455 & ~w19755;
assign w27199 = ~pi02169 & w19755;
assign w27200 = ~w27198 & ~w27199;
assign w27201 = pi04456 & ~w19755;
assign w27202 = ~pi02718 & w19755;
assign w27203 = ~w27201 & ~w27202;
assign w27204 = pi04457 & ~w19755;
assign w27205 = ~pi02167 & w19755;
assign w27206 = ~w27204 & ~w27205;
assign w27207 = pi04458 & ~w19755;
assign w27208 = ~pi02164 & w19755;
assign w27209 = ~w27207 & ~w27208;
assign w27210 = pi04459 & ~w19755;
assign w27211 = w19312 & w19459;
assign w27212 = ~w27210 & ~w27211;
assign w27213 = pi04460 & ~w19755;
assign w27214 = w17594 & w19459;
assign w27215 = ~w27213 & ~w27214;
assign w27216 = pi04461 & ~w19638;
assign w27217 = ~pi02703 & w19638;
assign w27218 = ~w27216 & ~w27217;
assign w27219 = pi04462 & ~w19638;
assign w27220 = ~pi02169 & w19638;
assign w27221 = ~w27219 & ~w27220;
assign w27222 = pi04463 & ~w19638;
assign w27223 = ~pi02718 & w19638;
assign w27224 = ~w27222 & ~w27223;
assign w27225 = pi04464 & ~w19638;
assign w27226 = ~pi02167 & w19638;
assign w27227 = ~w27225 & ~w27226;
assign w27228 = pi04465 & ~w19638;
assign w27229 = ~pi02722 & w19638;
assign w27230 = ~w27228 & ~w27229;
assign w27231 = pi04466 & ~w19638;
assign w27232 = ~pi02719 & w19638;
assign w27233 = ~w27231 & ~w27232;
assign w27234 = pi04467 & ~w19675;
assign w27235 = w17532 & w19444;
assign w27236 = ~w27234 & ~w27235;
assign w27237 = pi04468 & ~w19675;
assign w27238 = w19444 & w19797;
assign w27239 = ~w27237 & ~w27238;
assign w27240 = pi04469 & ~w19675;
assign w27241 = w17586 & w19444;
assign w27242 = ~w27240 & ~w27241;
assign w27243 = pi04470 & ~w19675;
assign w27244 = w19273 & w19444;
assign w27245 = ~w27243 & ~w27244;
assign w27246 = pi04471 & ~w19675;
assign w27247 = w17620 & w19444;
assign w27248 = ~w27246 & ~w27247;
assign w27249 = pi04472 & ~w19675;
assign w27250 = w19312 & w19444;
assign w27251 = ~w27249 & ~w27250;
assign w27252 = pi04473 & ~w19675;
assign w27253 = w17594 & w19444;
assign w27254 = ~w27252 & ~w27253;
assign w27255 = pi04474 & ~w19611;
assign w27256 = ~pi02703 & w19611;
assign w27257 = ~w27255 & ~w27256;
assign w27258 = pi04475 & ~w19611;
assign w27259 = ~pi02169 & w19611;
assign w27260 = ~w27258 & ~w27259;
assign w27261 = pi04476 & ~w19611;
assign w27262 = ~pi02718 & w19611;
assign w27263 = ~w27261 & ~w27262;
assign w27264 = pi04477 & ~w19611;
assign w27265 = ~pi02167 & w19611;
assign w27266 = ~w27264 & ~w27265;
assign w27267 = pi04478 & ~w19611;
assign w27268 = ~pi02722 & w19611;
assign w27269 = ~w27267 & ~w27268;
assign w27270 = pi04479 & ~w19611;
assign w27271 = ~pi02719 & w19611;
assign w27272 = ~w27270 & ~w27271;
assign w27273 = pi04480 & ~w19592;
assign w27274 = w17532 & w19591;
assign w27275 = ~w27273 & ~w27274;
assign w27276 = pi04481 & ~w19592;
assign w27277 = w19591 & w19797;
assign w27278 = ~w27276 & ~w27277;
assign w27279 = pi04482 & ~w19592;
assign w27280 = w17586 & w19591;
assign w27281 = ~w27279 & ~w27280;
assign w27282 = pi04483 & ~w19592;
assign w27283 = w19273 & w19591;
assign w27284 = ~w27282 & ~w27283;
assign w27285 = pi04484 & ~w19592;
assign w27286 = w17620 & w19591;
assign w27287 = ~w27285 & ~w27286;
assign w27288 = pi04485 & ~w19592;
assign w27289 = w17594 & w19591;
assign w27290 = ~w27288 & ~w27289;
assign w27291 = pi04486 & ~w19592;
assign w27292 = w19312 & w19591;
assign w27293 = ~w27291 & ~w27292;
assign w27294 = pi04487 & ~w19013;
assign w27295 = ~pi02703 & w19013;
assign w27296 = ~w27294 & ~w27295;
assign w27297 = pi04488 & ~w19013;
assign w27298 = ~pi02169 & w19013;
assign w27299 = ~w27297 & ~w27298;
assign w27300 = pi04489 & ~w19013;
assign w27301 = ~pi02718 & w19013;
assign w27302 = ~w27300 & ~w27301;
assign w27303 = pi04490 & ~w19013;
assign w27304 = ~pi02167 & w19013;
assign w27305 = ~w27303 & ~w27304;
assign w27306 = pi04491 & ~w19013;
assign w27307 = ~pi02722 & w19013;
assign w27308 = ~w27306 & ~w27307;
assign w27309 = pi04492 & ~w19013;
assign w27310 = ~pi02719 & w19013;
assign w27311 = ~w27309 & ~w27310;
assign w27312 = pi04493 & ~w19508;
assign w27313 = ~pi02703 & w19508;
assign w27314 = ~w27312 & ~w27313;
assign w27315 = pi04494 & ~w19508;
assign w27316 = ~pi02169 & w19508;
assign w27317 = ~w27315 & ~w27316;
assign w27318 = pi04495 & ~w19508;
assign w27319 = ~pi02718 & w19508;
assign w27320 = ~w27318 & ~w27319;
assign w27321 = pi04496 & ~w19508;
assign w27322 = w19273 & w19374;
assign w27323 = ~w27321 & ~w27322;
assign w27324 = pi04497 & ~w19508;
assign w27325 = ~pi02164 & w19508;
assign w27326 = ~w27324 & ~w27325;
assign w27327 = pi04498 & ~w19508;
assign w27328 = ~pi02722 & w19508;
assign w27329 = ~w27327 & ~w27328;
assign w27330 = pi04499 & ~w19508;
assign w27331 = ~pi02719 & w19508;
assign w27332 = ~w27330 & ~w27331;
assign w27333 = pi04500 & ~w19440;
assign w27334 = ~pi02703 & w19440;
assign w27335 = ~w27333 & ~w27334;
assign w27336 = pi04501 & ~w19440;
assign w27337 = ~pi02169 & w19440;
assign w27338 = ~w27336 & ~w27337;
assign w27339 = pi04502 & ~w19440;
assign w27340 = ~pi02718 & w19440;
assign w27341 = ~w27339 & ~w27340;
assign w27342 = pi04503 & ~w19440;
assign w27343 = ~pi02167 & w19440;
assign w27344 = ~w27342 & ~w27343;
assign w27345 = pi04504 & ~w19440;
assign w27346 = ~pi02722 & w19440;
assign w27347 = ~w27345 & ~w27346;
assign w27348 = pi04505 & ~w19440;
assign w27349 = ~pi02719 & w19440;
assign w27350 = ~w27348 & ~w27349;
assign w27351 = pi04506 & ~w19428;
assign w27352 = ~pi02703 & w19428;
assign w27353 = ~w27351 & ~w27352;
assign w27354 = pi04507 & ~w19428;
assign w27355 = ~pi02169 & w19428;
assign w27356 = ~w27354 & ~w27355;
assign w27357 = pi04508 & ~w19428;
assign w27358 = ~pi02718 & w19428;
assign w27359 = ~w27357 & ~w27358;
assign w27360 = pi04509 & ~w19428;
assign w27361 = ~pi02167 & w19428;
assign w27362 = ~w27360 & ~w27361;
assign w27363 = pi04510 & ~w19428;
assign w27364 = ~pi02164 & w19428;
assign w27365 = ~w27363 & ~w27364;
assign w27366 = pi04511 & ~w19428;
assign w27367 = ~pi02722 & w19428;
assign w27368 = ~w27366 & ~w27367;
assign w27369 = pi04512 & ~w19428;
assign w27370 = ~pi02719 & w19428;
assign w27371 = ~w27369 & ~w27370;
assign w27372 = pi04513 & ~w19363;
assign w27373 = w17186 & w17380;
assign w27374 = ~w27372 & ~w27373;
assign w27375 = pi04514 & ~w19363;
assign w27376 = w17193 & w17380;
assign w27377 = ~w27375 & ~w27376;
assign w27378 = pi04515 & ~w19363;
assign w27379 = w17311 & w17380;
assign w27380 = ~w27378 & ~w27379;
assign w27381 = pi04516 & ~w19363;
assign w27382 = w17380 & w18861;
assign w27383 = ~w27381 & ~w27382;
assign w27384 = pi04517 & ~w19363;
assign w27385 = w17128 & w17380;
assign w27386 = ~w27384 & ~w27385;
assign w27387 = pi04518 & ~w19363;
assign w27388 = w17380 & w17439;
assign w27389 = ~w27387 & ~w27388;
assign w27390 = pi04519 & ~w19395;
assign w27391 = ~pi09961 & w19395;
assign w27392 = ~w27390 & ~w27391;
assign w27393 = pi04520 & ~w19395;
assign w27394 = ~pi09812 & w19395;
assign w27395 = ~w27393 & ~w27394;
assign w27396 = pi04521 & ~w19395;
assign w27397 = ~pi02704 & w19395;
assign w27398 = ~w27396 & ~w27397;
assign w27399 = pi04522 & ~w19395;
assign w27400 = ~pi02178 & w19395;
assign w27401 = ~w27399 & ~w27400;
assign w27402 = pi04523 & ~w19395;
assign w27403 = ~pi09954 & w19395;
assign w27404 = ~w27402 & ~w27403;
assign w27405 = pi04524 & ~w19395;
assign w27406 = ~pi02720 & w19395;
assign w27407 = ~w27405 & ~w27406;
assign w27408 = pi04525 & ~w19395;
assign w27409 = ~pi09962 & w19395;
assign w27410 = ~w27408 & ~w27409;
assign w27411 = pi04526 & ~w19335;
assign w27412 = ~pi09848 & w19335;
assign w27413 = ~w27411 & ~w27412;
assign w27414 = pi04527 & ~w19335;
assign w27415 = ~pi09812 & w19335;
assign w27416 = ~w27414 & ~w27415;
assign w27417 = pi04528 & ~w19335;
assign w27418 = w17218 & w17311;
assign w27419 = ~w27417 & ~w27418;
assign w27420 = pi04529 & ~w19335;
assign w27421 = ~pi02178 & w19335;
assign w27422 = ~w27420 & ~w27421;
assign w27423 = pi04530 & ~w19335;
assign w27424 = w17128 & w17218;
assign w27425 = ~w27423 & ~w27424;
assign w27426 = pi04531 & ~w19335;
assign w27427 = ~pi09962 & w19335;
assign w27428 = ~w27426 & ~w27427;
assign w27429 = pi04532 & ~w19323;
assign w27430 = ~pi09961 & w19323;
assign w27431 = ~w27429 & ~w27430;
assign w27432 = ~w16905 & w17500;
assign w27433 = pi04533 & ~w27432;
assign w27434 = ~pi02713 & w27432;
assign w27435 = ~w27433 & ~w27434;
assign w27436 = pi04534 & ~w21311;
assign w27437 = ~pi09812 & w21311;
assign w27438 = ~w27436 & ~w27437;
assign w27439 = pi04535 & ~w19323;
assign w27440 = ~pi09812 & w19323;
assign w27441 = ~w27439 & ~w27440;
assign w27442 = pi04536 & ~w19323;
assign w27443 = ~pi02704 & w19323;
assign w27444 = ~w27442 & ~w27443;
assign w27445 = pi04537 & ~w19323;
assign w27446 = ~pi02178 & w19323;
assign w27447 = ~w27445 & ~w27446;
assign w27448 = pi04538 & ~w19323;
assign w27449 = ~pi09954 & w19323;
assign w27450 = ~w27448 & ~w27449;
assign w27451 = pi04539 & ~w19323;
assign w27452 = ~pi02720 & w19323;
assign w27453 = ~w27451 & ~w27452;
assign w27454 = pi04540 & ~w19323;
assign w27455 = ~pi09962 & w19323;
assign w27456 = ~w27454 & ~w27455;
assign w27457 = pi04541 & ~w19008;
assign w27458 = w17131 & w19365;
assign w27459 = ~w27457 & ~w27458;
assign w27460 = pi04542 & ~w19008;
assign w27461 = ~pi09812 & w19008;
assign w27462 = ~w27460 & ~w27461;
assign w27463 = pi04543 & ~w19008;
assign w27464 = ~pi02178 & w19008;
assign w27465 = ~w27463 & ~w27464;
assign w27466 = pi04544 & ~w19008;
assign w27467 = ~pi02704 & w19008;
assign w27468 = ~w27466 & ~w27467;
assign w27469 = pi04545 & ~w19008;
assign w27470 = ~pi02720 & w19008;
assign w27471 = ~w27469 & ~w27470;
assign w27472 = pi04546 & ~w19008;
assign w27473 = w17131 & w17439;
assign w27474 = ~w27472 & ~w27473;
assign w27475 = pi04547 & ~w19249;
assign w27476 = w17060 & w19365;
assign w27477 = ~w27475 & ~w27476;
assign w27478 = pi04548 & ~w19249;
assign w27479 = ~pi09812 & w19249;
assign w27480 = ~w27478 & ~w27479;
assign w27481 = pi04549 & ~w19249;
assign w27482 = ~pi02178 & w19249;
assign w27483 = ~w27481 & ~w27482;
assign w27484 = pi04550 & ~w19249;
assign w27485 = ~pi02720 & w19249;
assign w27486 = ~w27484 & ~w27485;
assign w27487 = pi04551 & ~w19249;
assign w27488 = ~pi09962 & w19249;
assign w27489 = ~w27487 & ~w27488;
assign w27490 = pi04552 & ~w19107;
assign w27491 = ~pi09961 & w19107;
assign w27492 = ~w27490 & ~w27491;
assign w27493 = pi04553 & ~w19107;
assign w27494 = ~pi09848 & w19107;
assign w27495 = ~w27493 & ~w27494;
assign w27496 = pi04554 & ~w19107;
assign w27497 = ~pi09812 & w19107;
assign w27498 = ~w27496 & ~w27497;
assign w27499 = pi04555 & ~w19107;
assign w27500 = ~pi02178 & w19107;
assign w27501 = ~w27499 & ~w27500;
assign w27502 = pi04556 & ~w19107;
assign w27503 = ~pi02720 & w19107;
assign w27504 = ~w27502 & ~w27503;
assign w27505 = pi04557 & ~w19107;
assign w27506 = ~pi09962 & w19107;
assign w27507 = ~w27505 & ~w27506;
assign w27508 = pi04558 & ~w19150;
assign w27509 = ~pi09848 & w19150;
assign w27510 = ~w27508 & ~w27509;
assign w27511 = pi04559 & ~w19150;
assign w27512 = w17193 & w19149;
assign w27513 = ~w27511 & ~w27512;
assign w27514 = pi04560 & ~w19150;
assign w27515 = ~pi02704 & w19150;
assign w27516 = ~w27514 & ~w27515;
assign w27517 = pi04561 & ~w19150;
assign w27518 = ~pi09954 & w19150;
assign w27519 = ~w27517 & ~w27518;
assign w27520 = pi04562 & ~w19150;
assign w27521 = ~pi02720 & w19150;
assign w27522 = ~w27520 & ~w27521;
assign w27523 = pi04563 & ~w19150;
assign w27524 = ~pi09962 & w19150;
assign w27525 = ~w27523 & ~w27524;
assign w27526 = pi04564 & ~w19167;
assign w27527 = w19166 & w19365;
assign w27528 = ~w27526 & ~w27527;
assign w27529 = pi04565 & ~w19167;
assign w27530 = ~pi09848 & w19167;
assign w27531 = ~w27529 & ~w27530;
assign w27532 = pi04566 & ~w19167;
assign w27533 = ~pi02704 & w19167;
assign w27534 = ~w27532 & ~w27533;
assign w27535 = pi04567 & ~w19167;
assign w27536 = ~pi02178 & w19167;
assign w27537 = ~w27535 & ~w27536;
assign w27538 = pi04568 & ~w19167;
assign w27539 = ~pi02720 & w19167;
assign w27540 = ~w27538 & ~w27539;
assign w27541 = pi04569 & ~w19249;
assign w27542 = ~pi09954 & w19249;
assign w27543 = ~w27541 & ~w27542;
assign w27544 = pi04570 & ~w19167;
assign w27545 = ~pi09962 & w19167;
assign w27546 = ~w27544 & ~w27545;
assign w27547 = pi04571 & ~w19131;
assign w27548 = ~pi09848 & w19131;
assign w27549 = ~w27547 & ~w27548;
assign w27550 = pi04572 & ~w19131;
assign w27551 = ~pi09812 & w19131;
assign w27552 = ~w27550 & ~w27551;
assign w27553 = pi04573 & ~w19131;
assign w27554 = ~pi02704 & w19131;
assign w27555 = ~w27553 & ~w27554;
assign w27556 = pi04574 & ~w19131;
assign w27557 = ~pi02720 & w19131;
assign w27558 = ~w27556 & ~w27557;
assign w27559 = pi04575 & ~w19131;
assign w27560 = ~pi09962 & w19131;
assign w27561 = ~w27559 & ~w27560;
assign w27562 = pi04576 & ~w19249;
assign w27563 = ~pi02704 & w19249;
assign w27564 = ~w27562 & ~w27563;
assign w27565 = pi04577 & ~w19116;
assign w27566 = w17186 & w19115;
assign w27567 = ~w27565 & ~w27566;
assign w27568 = pi04578 & ~w19116;
assign w27569 = ~pi09961 & w19116;
assign w27570 = ~w27568 & ~w27569;
assign w27571 = pi04579 & ~w19116;
assign w27572 = ~pi09812 & w19116;
assign w27573 = ~w27571 & ~w27572;
assign w27574 = pi04580 & ~w19116;
assign w27575 = w17311 & w19115;
assign w27576 = ~w27574 & ~w27575;
assign w27577 = pi04581 & ~w19116;
assign w27578 = ~pi09954 & w19116;
assign w27579 = ~w27577 & ~w27578;
assign w27580 = pi04582 & ~w19116;
assign w27581 = ~pi02720 & w19116;
assign w27582 = ~w27580 & ~w27581;
assign w27583 = pi04583 & ~w19116;
assign w27584 = ~pi09962 & w19116;
assign w27585 = ~w27583 & ~w27584;
assign w27586 = pi04584 & ~w19088;
assign w27587 = ~pi09961 & w19088;
assign w27588 = ~w27586 & ~w27587;
assign w27589 = pi04585 & ~w19088;
assign w27590 = ~pi09848 & w19088;
assign w27591 = ~w27589 & ~w27590;
assign w27592 = pi04586 & ~w19088;
assign w27593 = ~pi09812 & w19088;
assign w27594 = ~w27592 & ~w27593;
assign w27595 = ~w16905 & w18032;
assign w27596 = pi04587 & ~w27595;
assign w27597 = ~pi02717 & w27595;
assign w27598 = ~w27596 & ~w27597;
assign w27599 = pi04588 & ~w19088;
assign w27600 = w17513 & w19087;
assign w27601 = ~w27599 & ~w27600;
assign w27602 = pi04589 & ~w19088;
assign w27603 = w17128 & w19087;
assign w27604 = ~w27602 & ~w27603;
assign w27605 = pi04590 & ~w19088;
assign w27606 = ~pi09962 & w19088;
assign w27607 = ~w27605 & ~w27606;
assign w27608 = pi04591 & ~w19080;
assign w27609 = ~pi09961 & w19080;
assign w27610 = ~w27608 & ~w27609;
assign w27611 = pi04592 & ~w19080;
assign w27612 = w17193 & w19075;
assign w27613 = ~w27611 & ~w27612;
assign w27614 = pi04593 & ~w19080;
assign w27615 = ~pi02704 & w19080;
assign w27616 = ~w27614 & ~w27615;
assign w27617 = pi04594 & ~w19080;
assign w27618 = ~pi02178 & w19080;
assign w27619 = ~w27617 & ~w27618;
assign w27620 = pi04595 & ~w19080;
assign w27621 = ~pi02720 & w19080;
assign w27622 = ~w27620 & ~w27621;
assign w27623 = pi04596 & ~w19080;
assign w27624 = w17439 & w19075;
assign w27625 = ~w27623 & ~w27624;
assign w27626 = pi04597 & ~w18996;
assign w27627 = ~pi09961 & w18996;
assign w27628 = ~w27626 & ~w27627;
assign w27629 = pi04598 & ~w18996;
assign w27630 = ~pi09812 & w18996;
assign w27631 = ~w27629 & ~w27630;
assign w27632 = pi04599 & ~w18996;
assign w27633 = ~pi02704 & w18996;
assign w27634 = ~w27632 & ~w27633;
assign w27635 = pi04600 & ~w18996;
assign w27636 = ~pi02178 & w18996;
assign w27637 = ~w27635 & ~w27636;
assign w27638 = pi04601 & ~w18996;
assign w27639 = ~pi02720 & w18996;
assign w27640 = ~w27638 & ~w27639;
assign w27641 = pi04602 & ~w18996;
assign w27642 = ~pi09962 & w18996;
assign w27643 = ~w27641 & ~w27642;
assign w27644 = pi04603 & ~w19054;
assign w27645 = ~pi09961 & w19054;
assign w27646 = ~w27644 & ~w27645;
assign w27647 = pi04604 & ~w19054;
assign w27648 = w17186 & w19053;
assign w27649 = ~w27647 & ~w27648;
assign w27650 = pi04605 & ~w19054;
assign w27651 = ~pi09812 & w19054;
assign w27652 = ~w27650 & ~w27651;
assign w27653 = pi04606 & ~w19054;
assign w27654 = ~pi02704 & w19054;
assign w27655 = ~w27653 & ~w27654;
assign w27656 = pi04607 & ~w19054;
assign w27657 = ~pi02178 & w19054;
assign w27658 = ~w27656 & ~w27657;
assign w27659 = pi04608 & ~w19054;
assign w27660 = ~pi02720 & w19054;
assign w27661 = ~w27659 & ~w27660;
assign w27662 = pi04609 & ~w19054;
assign w27663 = ~pi09962 & w19054;
assign w27664 = ~w27662 & ~w27663;
assign w27665 = pi04610 & ~w19043;
assign w27666 = ~pi09961 & w19043;
assign w27667 = ~w27665 & ~w27666;
assign w27668 = pi04611 & ~w19043;
assign w27669 = ~pi09812 & w19043;
assign w27670 = ~w27668 & ~w27669;
assign w27671 = pi04612 & ~w19043;
assign w27672 = ~pi02704 & w19043;
assign w27673 = ~w27671 & ~w27672;
assign w27674 = pi04613 & ~w19043;
assign w27675 = ~pi02178 & w19043;
assign w27676 = ~w27674 & ~w27675;
assign w27677 = pi04614 & ~w19043;
assign w27678 = ~pi02720 & w19043;
assign w27679 = ~w27677 & ~w27678;
assign w27680 = pi04615 & ~w19043;
assign w27681 = ~pi09962 & w19043;
assign w27682 = ~w27680 & ~w27681;
assign w27683 = pi04616 & ~w19027;
assign w27684 = ~pi09961 & w19027;
assign w27685 = ~w27683 & ~w27684;
assign w27686 = pi04617 & ~w19027;
assign w27687 = ~pi09848 & w19027;
assign w27688 = ~w27686 & ~w27687;
assign w27689 = pi04618 & ~w19027;
assign w27690 = ~pi09812 & w19027;
assign w27691 = ~w27689 & ~w27690;
assign w27692 = pi04619 & ~w19027;
assign w27693 = ~pi02704 & w19027;
assign w27694 = ~w27692 & ~w27693;
assign w27695 = pi04620 & ~w19027;
assign w27696 = ~pi02178 & w19027;
assign w27697 = ~w27695 & ~w27696;
assign w27698 = pi04621 & ~w19027;
assign w27699 = ~pi02720 & w19027;
assign w27700 = ~w27698 & ~w27699;
assign w27701 = pi04622 & ~w19027;
assign w27702 = ~pi09962 & w19027;
assign w27703 = ~w27701 & ~w27702;
assign w27704 = pi04623 & ~w18926;
assign w27705 = ~pi09961 & w18926;
assign w27706 = ~w27704 & ~w27705;
assign w27707 = pi04624 & ~w18926;
assign w27708 = ~pi09812 & w18926;
assign w27709 = ~w27707 & ~w27708;
assign w27710 = pi04625 & ~w18926;
assign w27711 = ~pi02704 & w18926;
assign w27712 = ~w27710 & ~w27711;
assign w27713 = pi04626 & ~w18926;
assign w27714 = ~pi02178 & w18926;
assign w27715 = ~w27713 & ~w27714;
assign w27716 = pi04627 & ~w18926;
assign w27717 = ~pi02720 & w18926;
assign w27718 = ~w27716 & ~w27717;
assign w27719 = pi04628 & ~w18926;
assign w27720 = ~pi09962 & w18926;
assign w27721 = ~w27719 & ~w27720;
assign w27722 = pi04629 & ~w18954;
assign w27723 = ~pi09961 & w18954;
assign w27724 = ~w27722 & ~w27723;
assign w27725 = pi04630 & ~w18954;
assign w27726 = ~pi09848 & w18954;
assign w27727 = ~w27725 & ~w27726;
assign w27728 = pi04631 & ~w18954;
assign w27729 = ~pi09812 & w18954;
assign w27730 = ~w27728 & ~w27729;
assign w27731 = pi04632 & ~w18954;
assign w27732 = ~pi02704 & w18954;
assign w27733 = ~w27731 & ~w27732;
assign w27734 = pi04633 & ~w18954;
assign w27735 = ~pi02178 & w18954;
assign w27736 = ~w27734 & ~w27735;
assign w27737 = pi04634 & ~w18954;
assign w27738 = ~pi02720 & w18954;
assign w27739 = ~w27737 & ~w27738;
assign w27740 = pi04635 & ~w18954;
assign w27741 = ~pi09962 & w18954;
assign w27742 = ~w27740 & ~w27741;
assign w27743 = pi04636 & ~w18914;
assign w27744 = w18913 & w19365;
assign w27745 = ~w27743 & ~w27744;
assign w27746 = pi04637 & ~w18914;
assign w27747 = ~pi09812 & w18914;
assign w27748 = ~w27746 & ~w27747;
assign w27749 = pi04638 & ~w18914;
assign w27750 = ~pi02704 & w18914;
assign w27751 = ~w27749 & ~w27750;
assign w27752 = pi04639 & ~w18914;
assign w27753 = ~pi02178 & w18914;
assign w27754 = ~w27752 & ~w27753;
assign w27755 = pi04640 & ~w18914;
assign w27756 = ~pi02720 & w18914;
assign w27757 = ~w27755 & ~w27756;
assign w27758 = pi04641 & ~w18914;
assign w27759 = ~pi09962 & w18914;
assign w27760 = ~w27758 & ~w27759;
assign w27761 = pi04642 & ~w18936;
assign w27762 = ~pi09961 & w18936;
assign w27763 = ~w27761 & ~w27762;
assign w27764 = pi04643 & ~w18936;
assign w27765 = ~pi09848 & w18936;
assign w27766 = ~w27764 & ~w27765;
assign w27767 = pi04644 & ~w18936;
assign w27768 = ~pi09812 & w18936;
assign w27769 = ~w27767 & ~w27768;
assign w27770 = pi04645 & ~w18936;
assign w27771 = ~pi02704 & w18936;
assign w27772 = ~w27770 & ~w27771;
assign w27773 = pi04646 & ~w18936;
assign w27774 = w18861 & w18897;
assign w27775 = ~w27773 & ~w27774;
assign w27776 = pi04647 & ~w18936;
assign w27777 = ~pi02720 & w18936;
assign w27778 = ~w27776 & ~w27777;
assign w27779 = pi04648 & ~w18936;
assign w27780 = ~pi09962 & w18936;
assign w27781 = ~w27779 & ~w27780;
assign w27782 = pi04649 & ~w18905;
assign w27783 = ~pi09961 & w18905;
assign w27784 = ~w27782 & ~w27783;
assign w27785 = pi04650 & ~w18905;
assign w27786 = ~pi09812 & w18905;
assign w27787 = ~w27785 & ~w27786;
assign w27788 = pi04651 & ~w18905;
assign w27789 = w17311 & w18871;
assign w27790 = ~w27788 & ~w27789;
assign w27791 = pi04652 & ~w18905;
assign w27792 = ~pi02178 & w18905;
assign w27793 = ~w27791 & ~w27792;
assign w27794 = pi04653 & ~w18905;
assign w27795 = ~pi02720 & w18905;
assign w27796 = ~w27794 & ~w27795;
assign w27797 = pi04654 & ~w18905;
assign w27798 = ~pi09962 & w18905;
assign w27799 = ~w27797 & ~w27798;
assign w27800 = pi04655 & ~w18889;
assign w27801 = ~pi09961 & w18889;
assign w27802 = ~w27800 & ~w27801;
assign w27803 = pi04656 & ~w18889;
assign w27804 = ~pi09848 & w18889;
assign w27805 = ~w27803 & ~w27804;
assign w27806 = pi04657 & ~w18889;
assign w27807 = ~pi09812 & w18889;
assign w27808 = ~w27806 & ~w27807;
assign w27809 = pi04658 & ~w18889;
assign w27810 = ~pi02704 & w18889;
assign w27811 = ~w27809 & ~w27810;
assign w27812 = pi04659 & ~w18889;
assign w27813 = ~pi02178 & w18889;
assign w27814 = ~w27812 & ~w27813;
assign w27815 = pi04660 & ~w18889;
assign w27816 = ~pi02720 & w18889;
assign w27817 = ~w27815 & ~w27816;
assign w27818 = pi04661 & ~w18889;
assign w27819 = ~pi09962 & w18889;
assign w27820 = ~w27818 & ~w27819;
assign w27821 = pi04662 & ~w18856;
assign w27822 = ~pi09961 & w18856;
assign w27823 = ~w27821 & ~w27822;
assign w27824 = pi04663 & ~w18856;
assign w27825 = ~pi09812 & w18856;
assign w27826 = ~w27824 & ~w27825;
assign w27827 = pi04664 & ~w18856;
assign w27828 = ~pi02704 & w18856;
assign w27829 = ~w27827 & ~w27828;
assign w27830 = pi04665 & ~w18856;
assign w27831 = ~pi02178 & w18856;
assign w27832 = ~w27830 & ~w27831;
assign w27833 = pi04666 & ~w18856;
assign w27834 = ~pi02720 & w18856;
assign w27835 = ~w27833 & ~w27834;
assign w27836 = pi04667 & ~w18856;
assign w27837 = ~pi09962 & w18856;
assign w27838 = ~w27836 & ~w27837;
assign w27839 = pi04668 & ~w18852;
assign w27840 = ~pi09961 & w18852;
assign w27841 = ~w27839 & ~w27840;
assign w27842 = pi04669 & ~w18852;
assign w27843 = w17186 & w18612;
assign w27844 = ~w27842 & ~w27843;
assign w27845 = pi04670 & ~w18852;
assign w27846 = ~pi09812 & w18852;
assign w27847 = ~w27845 & ~w27846;
assign w27848 = pi04671 & ~w18852;
assign w27849 = ~pi02704 & w18852;
assign w27850 = ~w27848 & ~w27849;
assign w27851 = pi04672 & ~w18852;
assign w27852 = ~pi02178 & w18852;
assign w27853 = ~w27851 & ~w27852;
assign w27854 = pi04673 & ~w18852;
assign w27855 = ~pi02720 & w18852;
assign w27856 = ~w27854 & ~w27855;
assign w27857 = pi04674 & ~w18852;
assign w27858 = w17439 & w18612;
assign w27859 = ~w27857 & ~w27858;
assign w27860 = pi04675 & ~w18818;
assign w27861 = ~pi09961 & w18818;
assign w27862 = ~w27860 & ~w27861;
assign w27863 = pi04676 & ~w18818;
assign w27864 = w17193 & w17516;
assign w27865 = ~w27863 & ~w27864;
assign w27866 = pi04677 & ~w18818;
assign w27867 = ~pi02704 & w18818;
assign w27868 = ~w27866 & ~w27867;
assign w27869 = pi04678 & ~w18818;
assign w27870 = ~pi02178 & w18818;
assign w27871 = ~w27869 & ~w27870;
assign w27872 = pi04679 & ~w18818;
assign w27873 = ~pi02720 & w18818;
assign w27874 = ~w27872 & ~w27873;
assign w27875 = pi04680 & ~w18818;
assign w27876 = ~pi09962 & w18818;
assign w27877 = ~w27875 & ~w27876;
assign w27878 = pi04681 & ~w18790;
assign w27879 = ~pi09961 & w18790;
assign w27880 = ~w27878 & ~w27879;
assign w27881 = pi04682 & ~w18790;
assign w27882 = ~pi09848 & w18790;
assign w27883 = ~w27881 & ~w27882;
assign w27884 = pi04683 & ~w18790;
assign w27885 = ~pi09812 & w18790;
assign w27886 = ~w27884 & ~w27885;
assign w27887 = pi04684 & ~w18790;
assign w27888 = ~pi02704 & w18790;
assign w27889 = ~w27887 & ~w27888;
assign w27890 = pi04685 & ~w18790;
assign w27891 = ~pi02178 & w18790;
assign w27892 = ~w27890 & ~w27891;
assign w27893 = pi04686 & ~w18790;
assign w27894 = ~pi02720 & w18790;
assign w27895 = ~w27893 & ~w27894;
assign w27896 = pi04687 & ~w18790;
assign w27897 = ~pi09962 & w18790;
assign w27898 = ~w27896 & ~w27897;
assign w27899 = pi04688 & ~w18710;
assign w27900 = ~pi09961 & w18710;
assign w27901 = ~w27899 & ~w27900;
assign w27902 = pi04689 & ~w18710;
assign w27903 = ~pi09812 & w18710;
assign w27904 = ~w27902 & ~w27903;
assign w27905 = pi04690 & ~w18710;
assign w27906 = ~pi02704 & w18710;
assign w27907 = ~w27905 & ~w27906;
assign w27908 = pi04691 & ~w18710;
assign w27909 = ~pi02178 & w18710;
assign w27910 = ~w27908 & ~w27909;
assign w27911 = pi04692 & ~w18710;
assign w27912 = ~pi02720 & w18710;
assign w27913 = ~w27911 & ~w27912;
assign w27914 = pi04693 & ~w18710;
assign w27915 = ~pi09962 & w18710;
assign w27916 = ~w27914 & ~w27915;
assign w27917 = pi04694 & ~w17511;
assign w27918 = ~pi09961 & w17511;
assign w27919 = ~w27917 & ~w27918;
assign w27920 = pi04695 & ~w17511;
assign w27921 = w17186 & w17510;
assign w27922 = ~w27920 & ~w27921;
assign w27923 = pi04696 & ~w17511;
assign w27924 = w17193 & w17510;
assign w27925 = ~w27923 & ~w27924;
assign w27926 = pi04697 & ~w17511;
assign w27927 = ~pi02704 & w17511;
assign w27928 = ~w27926 & ~w27927;
assign w27929 = pi04698 & ~w17511;
assign w27930 = w17510 & w18861;
assign w27931 = ~w27929 & ~w27930;
assign w27932 = pi04699 & ~w17511;
assign w27933 = w17128 & w17510;
assign w27934 = ~w27932 & ~w27933;
assign w27935 = pi04700 & ~w17511;
assign w27936 = w17439 & w17510;
assign w27937 = ~w27935 & ~w27936;
assign w27938 = pi04701 & ~w18404;
assign w27939 = ~pi09961 & w18404;
assign w27940 = ~w27938 & ~w27939;
assign w27941 = pi04702 & ~w18404;
assign w27942 = ~pi09812 & w18404;
assign w27943 = ~w27941 & ~w27942;
assign w27944 = pi04703 & ~w18404;
assign w27945 = ~pi02704 & w18404;
assign w27946 = ~w27944 & ~w27945;
assign w27947 = pi04704 & ~w18404;
assign w27948 = ~pi02178 & w18404;
assign w27949 = ~w27947 & ~w27948;
assign w27950 = pi04705 & ~w18404;
assign w27951 = ~pi02720 & w18404;
assign w27952 = ~w27950 & ~w27951;
assign w27953 = pi04706 & ~w18404;
assign w27954 = w17439 & w18308;
assign w27955 = ~w27953 & ~w27954;
assign w27956 = pi04707 & ~w18482;
assign w27957 = ~pi09961 & w18482;
assign w27958 = ~w27956 & ~w27957;
assign w27959 = pi04708 & ~w18482;
assign w27960 = ~pi09848 & w18482;
assign w27961 = ~w27959 & ~w27960;
assign w27962 = pi04709 & ~w18482;
assign w27963 = ~pi09812 & w18482;
assign w27964 = ~w27962 & ~w27963;
assign w27965 = pi04710 & ~w18482;
assign w27966 = ~pi02704 & w18482;
assign w27967 = ~w27965 & ~w27966;
assign w27968 = pi04711 & ~w18482;
assign w27969 = ~pi02178 & w18482;
assign w27970 = ~w27968 & ~w27969;
assign w27971 = pi04712 & ~w18482;
assign w27972 = w17128 & w18263;
assign w27973 = ~w27971 & ~w27972;
assign w27974 = pi04713 & ~w18482;
assign w27975 = ~pi09962 & w18482;
assign w27976 = ~w27974 & ~w27975;
assign w27977 = pi04714 & ~w18439;
assign w27978 = ~pi09961 & w18439;
assign w27979 = ~w27977 & ~w27978;
assign w27980 = pi04715 & ~w18439;
assign w27981 = ~pi09812 & w18439;
assign w27982 = ~w27980 & ~w27981;
assign w27983 = pi04716 & ~w18439;
assign w27984 = ~pi02704 & w18439;
assign w27985 = ~w27983 & ~w27984;
assign w27986 = pi04717 & ~w18439;
assign w27987 = ~pi02178 & w18439;
assign w27988 = ~w27986 & ~w27987;
assign w27989 = pi04718 & ~w18439;
assign w27990 = ~pi02720 & w18439;
assign w27991 = ~w27989 & ~w27990;
assign w27992 = pi04719 & ~w18439;
assign w27993 = ~pi09962 & w18439;
assign w27994 = ~w27992 & ~w27993;
assign w27995 = pi04720 & ~w18326;
assign w27996 = w18146 & w19365;
assign w27997 = ~w27995 & ~w27996;
assign w27998 = pi04721 & ~w18326;
assign w27999 = ~pi09848 & w18326;
assign w28000 = ~w27998 & ~w27999;
assign w28001 = pi04722 & ~w18326;
assign w28002 = ~pi09812 & w18326;
assign w28003 = ~w28001 & ~w28002;
assign w28004 = pi04723 & ~w18326;
assign w28005 = w17311 & w18146;
assign w28006 = ~w28004 & ~w28005;
assign w28007 = pi04724 & ~w18326;
assign w28008 = ~pi02178 & w18326;
assign w28009 = ~w28007 & ~w28008;
assign w28010 = pi04725 & ~w18326;
assign w28011 = ~pi02720 & w18326;
assign w28012 = ~w28010 & ~w28011;
assign w28013 = pi04726 & ~w18326;
assign w28014 = ~pi09962 & w18326;
assign w28015 = ~w28013 & ~w28014;
assign w28016 = pi04727 & ~w18337;
assign w28017 = ~pi09961 & w18337;
assign w28018 = ~w28016 & ~w28017;
assign w28019 = pi04728 & ~w18337;
assign w28020 = ~pi09812 & w18337;
assign w28021 = ~w28019 & ~w28020;
assign w28022 = pi04729 & ~w18337;
assign w28023 = ~pi02704 & w18337;
assign w28024 = ~w28022 & ~w28023;
assign w28025 = pi04730 & ~w18337;
assign w28026 = ~pi02178 & w18337;
assign w28027 = ~w28025 & ~w28026;
assign w28028 = pi04731 & ~w18337;
assign w28029 = ~pi02720 & w18337;
assign w28030 = ~w28028 & ~w28029;
assign w28031 = pi04732 & ~w18337;
assign w28032 = ~pi09962 & w18337;
assign w28033 = ~w28031 & ~w28032;
assign w28034 = pi04733 & ~w18344;
assign w28035 = ~pi09961 & w18344;
assign w28036 = ~w28034 & ~w28035;
assign w28037 = pi04734 & ~w18344;
assign w28038 = ~pi09848 & w18344;
assign w28039 = ~w28037 & ~w28038;
assign w28040 = pi04735 & ~w18344;
assign w28041 = ~pi09812 & w18344;
assign w28042 = ~w28040 & ~w28041;
assign w28043 = pi04736 & ~w18344;
assign w28044 = ~pi02704 & w18344;
assign w28045 = ~w28043 & ~w28044;
assign w28046 = pi04737 & ~w18344;
assign w28047 = ~pi02178 & w18344;
assign w28048 = ~w28046 & ~w28047;
assign w28049 = pi04738 & ~w18344;
assign w28050 = w17128 & w18070;
assign w28051 = ~w28049 & ~w28050;
assign w28052 = pi04739 & ~w18344;
assign w28053 = ~pi09962 & w18344;
assign w28054 = ~w28052 & ~w28053;
assign w28055 = pi04740 & ~w18296;
assign w28056 = ~pi09961 & w18296;
assign w28057 = ~w28055 & ~w28056;
assign w28058 = pi04741 & ~w18296;
assign w28059 = ~pi09812 & w18296;
assign w28060 = ~w28058 & ~w28059;
assign w28061 = pi04742 & ~w18296;
assign w28062 = ~pi02704 & w18296;
assign w28063 = ~w28061 & ~w28062;
assign w28064 = pi04743 & ~w18296;
assign w28065 = w18056 & w18861;
assign w28066 = ~w28064 & ~w28065;
assign w28067 = pi04744 & ~w18296;
assign w28068 = ~pi02720 & w18296;
assign w28069 = ~w28067 & ~w28068;
assign w28070 = pi04745 & ~w18296;
assign w28071 = ~pi09962 & w18296;
assign w28072 = ~w28070 & ~w28071;
assign w28073 = pi04746 & ~w18252;
assign w28074 = ~pi09961 & w18252;
assign w28075 = ~w28073 & ~w28074;
assign w28076 = pi04747 & ~w18252;
assign w28077 = ~pi09848 & w18252;
assign w28078 = ~w28076 & ~w28077;
assign w28079 = pi04748 & ~w18252;
assign w28080 = w17193 & w18051;
assign w28081 = ~w28079 & ~w28080;
assign w28082 = pi04749 & ~w18252;
assign w28083 = ~pi02704 & w18252;
assign w28084 = ~w28082 & ~w28083;
assign w28085 = pi04750 & ~w18252;
assign w28086 = ~pi02178 & w18252;
assign w28087 = ~w28085 & ~w28086;
assign w28088 = pi04751 & ~w18252;
assign w28089 = w17128 & w18051;
assign w28090 = ~w28088 & ~w28089;
assign w28091 = pi04752 & ~w18252;
assign w28092 = ~pi09962 & w18252;
assign w28093 = ~w28091 & ~w28092;
assign w28094 = pi04753 & ~w18138;
assign w28095 = ~pi09961 & w18138;
assign w28096 = ~w28094 & ~w28095;
assign w28097 = pi04754 & ~w18138;
assign w28098 = ~pi09812 & w18138;
assign w28099 = ~w28097 & ~w28098;
assign w28100 = pi04755 & ~w18138;
assign w28101 = w17311 & w17445;
assign w28102 = ~w28100 & ~w28101;
assign w28103 = pi04756 & ~w18138;
assign w28104 = ~pi02178 & w18138;
assign w28105 = ~w28103 & ~w28104;
assign w28106 = pi04757 & ~w18138;
assign w28107 = ~pi02720 & w18138;
assign w28108 = ~w28106 & ~w28107;
assign w28109 = pi04758 & ~w18138;
assign w28110 = ~pi09962 & w18138;
assign w28111 = ~w28109 & ~w28110;
assign w28112 = pi04759 & ~w18194;
assign w28113 = ~pi09961 & w18194;
assign w28114 = ~w28112 & ~w28113;
assign w28115 = pi04760 & ~w18194;
assign w28116 = w17017 & w17186;
assign w28117 = ~w28115 & ~w28116;
assign w28118 = pi04761 & ~w18194;
assign w28119 = ~pi09812 & w18194;
assign w28120 = ~w28118 & ~w28119;
assign w28121 = pi04762 & ~w18194;
assign w28122 = ~pi02704 & w18194;
assign w28123 = ~w28121 & ~w28122;
assign w28124 = pi04763 & ~w18194;
assign w28125 = ~pi02178 & w18194;
assign w28126 = ~w28124 & ~w28125;
assign w28127 = pi04764 & ~w18194;
assign w28128 = ~pi02720 & w18194;
assign w28129 = ~w28127 & ~w28128;
assign w28130 = pi04765 & ~w18194;
assign w28131 = ~pi09962 & w18194;
assign w28132 = ~w28130 & ~w28131;
assign w28133 = pi04766 & ~w18160;
assign w28134 = ~pi09961 & w18160;
assign w28135 = ~w28133 & ~w28134;
assign w28136 = pi04767 & ~w18160;
assign w28137 = ~pi09812 & w18160;
assign w28138 = ~w28136 & ~w28137;
assign w28139 = pi04768 & ~w18160;
assign w28140 = ~pi02704 & w18160;
assign w28141 = ~w28139 & ~w28140;
assign w28142 = pi04769 & ~w18160;
assign w28143 = ~pi02178 & w18160;
assign w28144 = ~w28142 & ~w28143;
assign w28145 = pi04770 & ~w21563;
assign w28146 = ~pi02713 & w21563;
assign w28147 = ~w28145 & ~w28146;
assign w28148 = pi04771 & ~w18160;
assign w28149 = ~pi02720 & w18160;
assign w28150 = ~w28148 & ~w28149;
assign w28151 = pi04772 & ~w18160;
assign w28152 = ~pi09962 & w18160;
assign w28153 = ~w28151 & ~w28152;
assign w28154 = pi04773 & ~w18018;
assign w28155 = w16994 & w19365;
assign w28156 = ~w28154 & ~w28155;
assign w28157 = pi04774 & ~w18018;
assign w28158 = ~pi09848 & w18018;
assign w28159 = ~w28157 & ~w28158;
assign w28160 = pi04775 & ~w18018;
assign w28161 = ~pi09812 & w18018;
assign w28162 = ~w28160 & ~w28161;
assign w28163 = pi04776 & ~w18018;
assign w28164 = ~pi02704 & w18018;
assign w28165 = ~w28163 & ~w28164;
assign w28166 = pi04777 & ~w18018;
assign w28167 = ~pi02178 & w18018;
assign w28168 = ~w28166 & ~w28167;
assign w28169 = pi04778 & ~w18018;
assign w28170 = ~pi02720 & w18018;
assign w28171 = ~w28169 & ~w28170;
assign w28172 = pi04779 & ~w18018;
assign w28173 = w16994 & w17439;
assign w28174 = ~w28172 & ~w28173;
assign w28175 = pi04780 & ~w17966;
assign w28176 = ~pi09961 & w17966;
assign w28177 = ~w28175 & ~w28176;
assign w28178 = pi04781 & ~w17966;
assign w28179 = ~pi09812 & w17966;
assign w28180 = ~w28178 & ~w28179;
assign w28181 = pi04782 & ~w17966;
assign w28182 = ~pi02704 & w17966;
assign w28183 = ~w28181 & ~w28182;
assign w28184 = pi04783 & ~w17966;
assign w28185 = ~pi02178 & w17966;
assign w28186 = ~w28184 & ~w28185;
assign w28187 = pi04784 & ~w17966;
assign w28188 = ~pi02720 & w17966;
assign w28189 = ~w28187 & ~w28188;
assign w28190 = pi04785 & ~w17966;
assign w28191 = w17439 & w17965;
assign w28192 = ~w28190 & ~w28191;
assign w28193 = pi04786 & ~w17913;
assign w28194 = w17912 & w19365;
assign w28195 = ~w28193 & ~w28194;
assign w28196 = pi04787 & ~w17913;
assign w28197 = w17186 & w17912;
assign w28198 = ~w28196 & ~w28197;
assign w28199 = pi04788 & ~w17913;
assign w28200 = ~pi09812 & w17913;
assign w28201 = ~w28199 & ~w28200;
assign w28202 = pi04789 & ~w17913;
assign w28203 = ~pi02704 & w17913;
assign w28204 = ~w28202 & ~w28203;
assign w28205 = pi04790 & ~w17913;
assign w28206 = ~pi02178 & w17913;
assign w28207 = ~w28205 & ~w28206;
assign w28208 = pi04791 & ~w17913;
assign w28209 = ~pi02720 & w17913;
assign w28210 = ~w28208 & ~w28209;
assign w28211 = pi04792 & ~w17913;
assign w28212 = ~pi09962 & w17913;
assign w28213 = ~w28211 & ~w28212;
assign w28214 = pi04793 & ~w17627;
assign w28215 = ~pi09961 & w17627;
assign w28216 = ~w28214 & ~w28215;
assign w28217 = pi04794 & ~w17627;
assign w28218 = ~pi09812 & w17627;
assign w28219 = ~w28217 & ~w28218;
assign w28220 = pi04795 & ~w17627;
assign w28221 = ~pi02704 & w17627;
assign w28222 = ~w28220 & ~w28221;
assign w28223 = pi04796 & ~w17627;
assign w28224 = ~pi02178 & w17627;
assign w28225 = ~w28223 & ~w28224;
assign w28226 = pi04797 & ~w17627;
assign w28227 = w17128 & w17626;
assign w28228 = ~w28226 & ~w28227;
assign w28229 = pi04798 & ~w17627;
assign w28230 = ~pi09962 & w17627;
assign w28231 = ~w28229 & ~w28230;
assign w28232 = ~w16928 & w20119;
assign w28233 = pi04799 & ~w28232;
assign w28234 = ~pi09961 & w28232;
assign w28235 = ~w28233 & ~w28234;
assign w28236 = pi04800 & ~w28232;
assign w28237 = ~pi09848 & w28232;
assign w28238 = ~w28236 & ~w28237;
assign w28239 = pi04801 & ~w28232;
assign w28240 = ~pi09812 & w28232;
assign w28241 = ~w28239 & ~w28240;
assign w28242 = pi04802 & ~w28232;
assign w28243 = ~pi02704 & w28232;
assign w28244 = ~w28242 & ~w28243;
assign w28245 = pi04803 & ~w28232;
assign w28246 = ~pi02178 & w28232;
assign w28247 = ~w28245 & ~w28246;
assign w28248 = pi04804 & ~w28232;
assign w28249 = ~pi09954 & w28232;
assign w28250 = ~w28248 & ~w28249;
assign w28251 = pi04805 & ~w28232;
assign w28252 = ~pi02720 & w28232;
assign w28253 = ~w28251 & ~w28252;
assign w28254 = pi04806 & ~w28232;
assign w28255 = ~pi09962 & w28232;
assign w28256 = ~w28254 & ~w28255;
assign w28257 = pi04807 & ~w16955;
assign w28258 = ~pi09961 & w16955;
assign w28259 = ~w28257 & ~w28258;
assign w28260 = pi04808 & ~w16955;
assign w28261 = ~pi09812 & w16955;
assign w28262 = ~w28260 & ~w28261;
assign w28263 = pi04809 & ~w16955;
assign w28264 = ~pi02704 & w16955;
assign w28265 = ~w28263 & ~w28264;
assign w28266 = pi04810 & ~w16955;
assign w28267 = ~pi02178 & w16955;
assign w28268 = ~w28266 & ~w28267;
assign w28269 = pi04811 & ~w16955;
assign w28270 = ~pi02720 & w16955;
assign w28271 = ~w28269 & ~w28270;
assign w28272 = pi04812 & ~w16955;
assign w28273 = w16954 & w17439;
assign w28274 = ~w28272 & ~w28273;
assign w28275 = pi04813 & ~w17104;
assign w28276 = ~pi09961 & w17104;
assign w28277 = ~w28275 & ~w28276;
assign w28278 = pi04814 & ~w17104;
assign w28279 = ~pi09848 & w17104;
assign w28280 = ~w28278 & ~w28279;
assign w28281 = pi04815 & ~w17104;
assign w28282 = ~pi09812 & w17104;
assign w28283 = ~w28281 & ~w28282;
assign w28284 = pi04816 & ~w17104;
assign w28285 = w17103 & w17311;
assign w28286 = ~w28284 & ~w28285;
assign w28287 = pi04817 & ~w17104;
assign w28288 = ~pi02178 & w17104;
assign w28289 = ~w28287 & ~w28288;
assign w28290 = pi04818 & ~w17104;
assign w28291 = ~pi02720 & w17104;
assign w28292 = ~w28290 & ~w28291;
assign w28293 = pi04819 & ~w17104;
assign w28294 = ~pi09962 & w17104;
assign w28295 = ~w28293 & ~w28294;
assign w28296 = pi04820 & ~w17079;
assign w28297 = ~pi09961 & w17079;
assign w28298 = ~w28296 & ~w28297;
assign w28299 = pi04821 & ~w17079;
assign w28300 = w17078 & w17193;
assign w28301 = ~w28299 & ~w28300;
assign w28302 = pi04822 & ~w17079;
assign w28303 = w17078 & w17311;
assign w28304 = ~w28302 & ~w28303;
assign w28305 = pi04823 & ~w17079;
assign w28306 = ~pi02178 & w17079;
assign w28307 = ~w28305 & ~w28306;
assign w28308 = pi04824 & ~w23529;
assign w28309 = ~pi02704 & w23529;
assign w28310 = ~w28308 & ~w28309;
assign w28311 = pi04825 & ~w17079;
assign w28312 = ~pi02720 & w17079;
assign w28313 = ~w28311 & ~w28312;
assign w28314 = pi04826 & ~w17079;
assign w28315 = ~pi09962 & w17079;
assign w28316 = ~w28314 & ~w28315;
assign w28317 = pi04827 & ~w20505;
assign w28318 = ~pi09961 & w20505;
assign w28319 = ~w28317 & ~w28318;
assign w28320 = pi04828 & ~w20505;
assign w28321 = ~pi09848 & w20505;
assign w28322 = ~w28320 & ~w28321;
assign w28323 = pi04829 & ~w20505;
assign w28324 = ~pi09812 & w20505;
assign w28325 = ~w28323 & ~w28324;
assign w28326 = pi04830 & ~w20505;
assign w28327 = ~pi02704 & w20505;
assign w28328 = ~w28326 & ~w28327;
assign w28329 = pi04831 & ~w20505;
assign w28330 = ~pi02178 & w20505;
assign w28331 = ~w28329 & ~w28330;
assign w28332 = pi04832 & ~w20505;
assign w28333 = ~pi02720 & w20505;
assign w28334 = ~w28332 & ~w28333;
assign w28335 = pi04833 & ~w20505;
assign w28336 = ~pi09962 & w20505;
assign w28337 = ~w28335 & ~w28336;
assign w28338 = ~w16928 & w20059;
assign w28339 = pi04834 & ~w28338;
assign w28340 = ~pi09961 & w28338;
assign w28341 = ~w28339 & ~w28340;
assign w28342 = pi04835 & ~w28338;
assign w28343 = ~pi09812 & w28338;
assign w28344 = ~w28342 & ~w28343;
assign w28345 = pi04836 & ~w28338;
assign w28346 = ~pi02704 & w28338;
assign w28347 = ~w28345 & ~w28346;
assign w28348 = pi04837 & ~w28338;
assign w28349 = w18861 & w20059;
assign w28350 = ~w28348 & ~w28349;
assign w28351 = pi04838 & ~w28338;
assign w28352 = ~pi02720 & w28338;
assign w28353 = ~w28351 & ~w28352;
assign w28354 = pi04839 & ~w28338;
assign w28355 = ~pi09962 & w28338;
assign w28356 = ~w28354 & ~w28355;
assign w28357 = ~w16928 & w20014;
assign w28358 = pi04840 & ~w28357;
assign w28359 = ~pi09961 & w28357;
assign w28360 = ~w28358 & ~w28359;
assign w28361 = pi04841 & ~w28357;
assign w28362 = ~pi09848 & w28357;
assign w28363 = ~w28361 & ~w28362;
assign w28364 = pi04842 & ~w28357;
assign w28365 = ~pi09812 & w28357;
assign w28366 = ~w28364 & ~w28365;
assign w28367 = pi04843 & ~w28357;
assign w28368 = w17311 & w20014;
assign w28369 = ~w28367 & ~w28368;
assign w28370 = pi04844 & ~w28357;
assign w28371 = ~pi02178 & w28357;
assign w28372 = ~w28370 & ~w28371;
assign w28373 = pi04845 & ~w28357;
assign w28374 = ~pi02720 & w28357;
assign w28375 = ~w28373 & ~w28374;
assign w28376 = pi04846 & ~w28357;
assign w28377 = ~pi09962 & w28357;
assign w28378 = ~w28376 & ~w28377;
assign w28379 = ~w16928 & w19988;
assign w28380 = pi04847 & ~w28379;
assign w28381 = ~pi09961 & w28379;
assign w28382 = ~w28380 & ~w28381;
assign w28383 = pi04848 & ~w28379;
assign w28384 = ~pi09812 & w28379;
assign w28385 = ~w28383 & ~w28384;
assign w28386 = pi04849 & ~w28379;
assign w28387 = ~pi02704 & w28379;
assign w28388 = ~w28386 & ~w28387;
assign w28389 = pi04850 & ~w28379;
assign w28390 = ~pi02178 & w28379;
assign w28391 = ~w28389 & ~w28390;
assign w28392 = pi04851 & ~w28379;
assign w28393 = ~pi02720 & w28379;
assign w28394 = ~w28392 & ~w28393;
assign w28395 = pi04852 & ~w28379;
assign w28396 = ~pi09962 & w28379;
assign w28397 = ~w28395 & ~w28396;
assign w28398 = ~w16928 & w19941;
assign w28399 = pi04853 & ~w28398;
assign w28400 = ~pi09961 & w28398;
assign w28401 = ~w28399 & ~w28400;
assign w28402 = pi04854 & ~w28398;
assign w28403 = ~pi09848 & w28398;
assign w28404 = ~w28402 & ~w28403;
assign w28405 = pi04855 & ~w28398;
assign w28406 = ~pi09812 & w28398;
assign w28407 = ~w28405 & ~w28406;
assign w28408 = pi04856 & ~w28398;
assign w28409 = w17311 & w19941;
assign w28410 = ~w28408 & ~w28409;
assign w28411 = pi04857 & ~w28398;
assign w28412 = ~pi02178 & w28398;
assign w28413 = ~w28411 & ~w28412;
assign w28414 = pi04858 & ~w28398;
assign w28415 = ~pi02720 & w28398;
assign w28416 = ~w28414 & ~w28415;
assign w28417 = pi04859 & ~w28398;
assign w28418 = ~pi09962 & w28398;
assign w28419 = ~w28417 & ~w28418;
assign w28420 = ~w16928 & w19930;
assign w28421 = pi04860 & ~w28420;
assign w28422 = ~pi09961 & w28420;
assign w28423 = ~w28421 & ~w28422;
assign w28424 = pi04861 & ~w28420;
assign w28425 = ~pi09812 & w28420;
assign w28426 = ~w28424 & ~w28425;
assign w28427 = pi04862 & ~w28420;
assign w28428 = ~pi02704 & w28420;
assign w28429 = ~w28427 & ~w28428;
assign w28430 = pi04863 & ~w28420;
assign w28431 = ~pi02178 & w28420;
assign w28432 = ~w28430 & ~w28431;
assign w28433 = pi04864 & ~w28420;
assign w28434 = ~pi02720 & w28420;
assign w28435 = ~w28433 & ~w28434;
assign w28436 = pi04865 & ~w28420;
assign w28437 = ~pi09962 & w28420;
assign w28438 = ~w28436 & ~w28437;
assign w28439 = ~w16928 & w19909;
assign w28440 = pi04866 & ~w28439;
assign w28441 = ~pi09961 & w28439;
assign w28442 = ~w28440 & ~w28441;
assign w28443 = pi04867 & ~w28439;
assign w28444 = ~pi09848 & w28439;
assign w28445 = ~w28443 & ~w28444;
assign w28446 = pi04868 & ~w28439;
assign w28447 = ~pi09812 & w28439;
assign w28448 = ~w28446 & ~w28447;
assign w28449 = pi04869 & ~w28439;
assign w28450 = ~pi02704 & w28439;
assign w28451 = ~w28449 & ~w28450;
assign w28452 = pi04870 & ~w28439;
assign w28453 = ~pi02178 & w28439;
assign w28454 = ~w28452 & ~w28453;
assign w28455 = pi04871 & ~w28439;
assign w28456 = ~pi02720 & w28439;
assign w28457 = ~w28455 & ~w28456;
assign w28458 = pi04872 & ~w28439;
assign w28459 = ~pi09962 & w28439;
assign w28460 = ~w28458 & ~w28459;
assign w28461 = pi04873 & ~w19131;
assign w28462 = ~pi09954 & w19131;
assign w28463 = ~w28461 & ~w28462;
assign w28464 = ~w16928 & w19852;
assign w28465 = pi04874 & ~w28464;
assign w28466 = ~pi09848 & w28464;
assign w28467 = ~w28465 & ~w28466;
assign w28468 = pi04875 & ~w28464;
assign w28469 = ~pi09812 & w28464;
assign w28470 = ~w28468 & ~w28469;
assign w28471 = pi04876 & ~w28464;
assign w28472 = ~pi02704 & w28464;
assign w28473 = ~w28471 & ~w28472;
assign w28474 = pi04877 & ~w28464;
assign w28475 = w17513 & w19852;
assign w28476 = ~w28474 & ~w28475;
assign w28477 = pi04878 & ~w28464;
assign w28478 = ~pi02720 & w28464;
assign w28479 = ~w28477 & ~w28478;
assign w28480 = pi04879 & ~w28464;
assign w28481 = ~pi09962 & w28464;
assign w28482 = ~w28480 & ~w28481;
assign w28483 = ~w16928 & w19838;
assign w28484 = pi04880 & ~w28483;
assign w28485 = ~pi09961 & w28483;
assign w28486 = ~w28484 & ~w28485;
assign w28487 = pi04881 & ~w28483;
assign w28488 = ~pi09848 & w28483;
assign w28489 = ~w28487 & ~w28488;
assign w28490 = pi04882 & ~w28483;
assign w28491 = ~pi09812 & w28483;
assign w28492 = ~w28490 & ~w28491;
assign w28493 = pi04883 & ~w28483;
assign w28494 = ~pi02704 & w28483;
assign w28495 = ~w28493 & ~w28494;
assign w28496 = pi04884 & ~w28483;
assign w28497 = ~pi09954 & w28483;
assign w28498 = ~w28496 & ~w28497;
assign w28499 = pi04885 & ~w28483;
assign w28500 = ~pi02720 & w28483;
assign w28501 = ~w28499 & ~w28500;
assign w28502 = pi04886 & ~w28483;
assign w28503 = ~pi09962 & w28483;
assign w28504 = ~w28502 & ~w28503;
assign w28505 = ~w16928 & w19826;
assign w28506 = pi04887 & ~w28505;
assign w28507 = ~pi09848 & w28505;
assign w28508 = ~w28506 & ~w28507;
assign w28509 = pi04888 & ~w28505;
assign w28510 = ~pi09812 & w28505;
assign w28511 = ~w28509 & ~w28510;
assign w28512 = pi04889 & ~w28505;
assign w28513 = ~pi02704 & w28505;
assign w28514 = ~w28512 & ~w28513;
assign w28515 = pi04890 & ~w28505;
assign w28516 = ~pi09954 & w28505;
assign w28517 = ~w28515 & ~w28516;
assign w28518 = pi04891 & ~w28505;
assign w28519 = ~pi02720 & w28505;
assign w28520 = ~w28518 & ~w28519;
assign w28521 = pi04892 & ~w28505;
assign w28522 = ~pi09962 & w28505;
assign w28523 = ~w28521 & ~w28522;
assign w28524 = ~w16928 & w19818;
assign w28525 = pi04893 & ~w28524;
assign w28526 = ~pi09961 & w28524;
assign w28527 = ~w28525 & ~w28526;
assign w28528 = pi04894 & ~w28524;
assign w28529 = ~pi09848 & w28524;
assign w28530 = ~w28528 & ~w28529;
assign w28531 = pi04895 & ~w28524;
assign w28532 = ~pi09812 & w28524;
assign w28533 = ~w28531 & ~w28532;
assign w28534 = pi04896 & ~w28524;
assign w28535 = ~pi02704 & w28524;
assign w28536 = ~w28534 & ~w28535;
assign w28537 = pi04897 & ~w28524;
assign w28538 = ~pi09954 & w28524;
assign w28539 = ~w28537 & ~w28538;
assign w28540 = pi04898 & ~w28524;
assign w28541 = ~pi02720 & w28524;
assign w28542 = ~w28540 & ~w28541;
assign w28543 = pi04899 & ~w28524;
assign w28544 = ~pi09962 & w28524;
assign w28545 = ~w28543 & ~w28544;
assign w28546 = ~w16928 & w19740;
assign w28547 = pi04900 & ~w28546;
assign w28548 = ~pi09848 & w28546;
assign w28549 = ~w28547 & ~w28548;
assign w28550 = pi04901 & ~w28546;
assign w28551 = ~pi09812 & w28546;
assign w28552 = ~w28550 & ~w28551;
assign w28553 = pi04902 & ~w28546;
assign w28554 = ~pi02704 & w28546;
assign w28555 = ~w28553 & ~w28554;
assign w28556 = pi04903 & ~w28546;
assign w28557 = ~pi09954 & w28546;
assign w28558 = ~w28556 & ~w28557;
assign w28559 = pi04904 & ~w28546;
assign w28560 = ~pi02720 & w28546;
assign w28561 = ~w28559 & ~w28560;
assign w28562 = pi04905 & ~w28546;
assign w28563 = ~pi09962 & w28546;
assign w28564 = ~w28562 & ~w28563;
assign w28565 = ~w16928 & w19728;
assign w28566 = pi04906 & ~w28565;
assign w28567 = w19365 & w19728;
assign w28568 = ~w28566 & ~w28567;
assign w28569 = pi04907 & ~w28565;
assign w28570 = ~pi09848 & w28565;
assign w28571 = ~w28569 & ~w28570;
assign w28572 = pi04908 & ~w28565;
assign w28573 = ~pi09812 & w28565;
assign w28574 = ~w28572 & ~w28573;
assign w28575 = pi04909 & ~w28565;
assign w28576 = w17311 & w19728;
assign w28577 = ~w28575 & ~w28576;
assign w28578 = pi04910 & ~w28565;
assign w28579 = w17513 & w19728;
assign w28580 = ~w28578 & ~w28579;
assign w28581 = pi04911 & ~w28565;
assign w28582 = w17128 & w19728;
assign w28583 = ~w28581 & ~w28582;
assign w28584 = pi04912 & ~w28565;
assign w28585 = ~pi09962 & w28565;
assign w28586 = ~w28584 & ~w28585;
assign w28587 = ~w16928 & w19723;
assign w28588 = pi04913 & ~w28587;
assign w28589 = ~pi09848 & w28587;
assign w28590 = ~w28588 & ~w28589;
assign w28591 = pi04914 & ~w28587;
assign w28592 = w17193 & w19723;
assign w28593 = ~w28591 & ~w28592;
assign w28594 = pi04915 & ~w28587;
assign w28595 = ~pi02704 & w28587;
assign w28596 = ~w28594 & ~w28595;
assign w28597 = pi04916 & ~w28587;
assign w28598 = ~pi09954 & w28587;
assign w28599 = ~w28597 & ~w28598;
assign w28600 = pi04917 & ~w28587;
assign w28601 = ~pi02720 & w28587;
assign w28602 = ~w28600 & ~w28601;
assign w28603 = pi04918 & ~w28587;
assign w28604 = ~pi09962 & w28587;
assign w28605 = ~w28603 & ~w28604;
assign w28606 = ~w16928 & w19660;
assign w28607 = pi04919 & ~w28606;
assign w28608 = ~pi09961 & w28606;
assign w28609 = ~w28607 & ~w28608;
assign w28610 = pi04920 & ~w28606;
assign w28611 = ~pi09848 & w28606;
assign w28612 = ~w28610 & ~w28611;
assign w28613 = pi04921 & ~w28606;
assign w28614 = ~pi09812 & w28606;
assign w28615 = ~w28613 & ~w28614;
assign w28616 = pi04922 & ~w28606;
assign w28617 = ~pi02704 & w28606;
assign w28618 = ~w28616 & ~w28617;
assign w28619 = pi04923 & ~w28606;
assign w28620 = ~pi09954 & w28606;
assign w28621 = ~w28619 & ~w28620;
assign w28622 = pi04924 & ~w28606;
assign w28623 = ~pi02720 & w28606;
assign w28624 = ~w28622 & ~w28623;
assign w28625 = pi04925 & ~w28606;
assign w28626 = ~pi09962 & w28606;
assign w28627 = ~w28625 & ~w28626;
assign w28628 = ~w16928 & w19679;
assign w28629 = pi04926 & ~w28628;
assign w28630 = ~pi09848 & w28628;
assign w28631 = ~w28629 & ~w28630;
assign w28632 = pi04927 & ~w28628;
assign w28633 = ~pi09812 & w28628;
assign w28634 = ~w28632 & ~w28633;
assign w28635 = pi04928 & ~w28628;
assign w28636 = ~pi02704 & w28628;
assign w28637 = ~w28635 & ~w28636;
assign w28638 = pi04929 & ~w28628;
assign w28639 = ~pi09954 & w28628;
assign w28640 = ~w28638 & ~w28639;
assign w28641 = pi04930 & ~w28628;
assign w28642 = ~pi02720 & w28628;
assign w28643 = ~w28641 & ~w28642;
assign w28644 = pi04931 & ~w28628;
assign w28645 = ~pi09962 & w28628;
assign w28646 = ~w28644 & ~w28645;
assign w28647 = ~w16928 & w19650;
assign w28648 = pi04932 & ~w28647;
assign w28649 = ~pi09961 & w28647;
assign w28650 = ~w28648 & ~w28649;
assign w28651 = pi04933 & ~w28647;
assign w28652 = ~pi09848 & w28647;
assign w28653 = ~w28651 & ~w28652;
assign w28654 = pi04934 & ~w28647;
assign w28655 = ~pi09812 & w28647;
assign w28656 = ~w28654 & ~w28655;
assign w28657 = pi04935 & ~w28647;
assign w28658 = ~pi02704 & w28647;
assign w28659 = ~w28657 & ~w28658;
assign w28660 = pi04936 & ~w28647;
assign w28661 = ~pi09954 & w28647;
assign w28662 = ~w28660 & ~w28661;
assign w28663 = pi04937 & ~w28647;
assign w28664 = ~pi02720 & w28647;
assign w28665 = ~w28663 & ~w28664;
assign w28666 = pi04938 & ~w28647;
assign w28667 = ~pi09962 & w28647;
assign w28668 = ~w28666 & ~w28667;
assign w28669 = ~w16928 & w19645;
assign w28670 = pi04939 & ~w28669;
assign w28671 = w17186 & w19645;
assign w28672 = ~w28670 & ~w28671;
assign w28673 = pi04940 & ~w28669;
assign w28674 = ~pi09812 & w28669;
assign w28675 = ~w28673 & ~w28674;
assign w28676 = pi04941 & ~w28669;
assign w28677 = ~pi02704 & w28669;
assign w28678 = ~w28676 & ~w28677;
assign w28679 = pi04942 & ~w28669;
assign w28680 = w17513 & w19645;
assign w28681 = ~w28679 & ~w28680;
assign w28682 = pi04943 & ~w28669;
assign w28683 = ~pi02720 & w28669;
assign w28684 = ~w28682 & ~w28683;
assign w28685 = pi04944 & ~w28669;
assign w28686 = ~pi09962 & w28669;
assign w28687 = ~w28685 & ~w28686;
assign w28688 = ~w16928 & w19576;
assign w28689 = pi04945 & ~w28688;
assign w28690 = ~pi09961 & w28688;
assign w28691 = ~w28689 & ~w28690;
assign w28692 = pi04946 & ~w28688;
assign w28693 = ~pi09848 & w28688;
assign w28694 = ~w28692 & ~w28693;
assign w28695 = pi04947 & ~w28688;
assign w28696 = ~pi09812 & w28688;
assign w28697 = ~w28695 & ~w28696;
assign w28698 = pi04948 & ~w28688;
assign w28699 = ~pi02704 & w28688;
assign w28700 = ~w28698 & ~w28699;
assign w28701 = pi04949 & ~w28688;
assign w28702 = ~pi09954 & w28688;
assign w28703 = ~w28701 & ~w28702;
assign w28704 = pi04950 & ~w28688;
assign w28705 = ~pi02720 & w28688;
assign w28706 = ~w28704 & ~w28705;
assign w28707 = pi04951 & ~w28688;
assign w28708 = ~pi09962 & w28688;
assign w28709 = ~w28707 & ~w28708;
assign w28710 = ~w16928 & w19624;
assign w28711 = pi04952 & ~w28710;
assign w28712 = w17186 & w19624;
assign w28713 = ~w28711 & ~w28712;
assign w28714 = pi04953 & ~w28710;
assign w28715 = ~pi09812 & w28710;
assign w28716 = ~w28714 & ~w28715;
assign w28717 = pi04954 & ~w28710;
assign w28718 = ~pi02704 & w28710;
assign w28719 = ~w28717 & ~w28718;
assign w28720 = pi04955 & ~w28710;
assign w28721 = ~pi09954 & w28710;
assign w28722 = ~w28720 & ~w28721;
assign w28723 = pi04956 & ~w28710;
assign w28724 = ~pi02720 & w28710;
assign w28725 = ~w28723 & ~w28724;
assign w28726 = pi04957 & ~w28710;
assign w28727 = ~pi09962 & w28710;
assign w28728 = ~w28726 & ~w28727;
assign w28729 = ~w16928 & w19606;
assign w28730 = pi04958 & ~w28729;
assign w28731 = ~pi09961 & w28729;
assign w28732 = ~w28730 & ~w28731;
assign w28733 = pi04959 & ~w28729;
assign w28734 = ~pi09848 & w28729;
assign w28735 = ~w28733 & ~w28734;
assign w28736 = pi04960 & ~w28729;
assign w28737 = ~pi09812 & w28729;
assign w28738 = ~w28736 & ~w28737;
assign w28739 = pi04961 & ~w28729;
assign w28740 = ~pi02704 & w28729;
assign w28741 = ~w28739 & ~w28740;
assign w28742 = pi04962 & ~w28729;
assign w28743 = ~pi09954 & w28729;
assign w28744 = ~w28742 & ~w28743;
assign w28745 = pi04963 & ~w28729;
assign w28746 = ~pi02720 & w28729;
assign w28747 = ~w28745 & ~w28746;
assign w28748 = pi04964 & ~w28729;
assign w28749 = ~pi09962 & w28729;
assign w28750 = ~w28748 & ~w28749;
assign w28751 = ~w16928 & w19601;
assign w28752 = pi04965 & ~w28751;
assign w28753 = w17186 & w19601;
assign w28754 = ~w28752 & ~w28753;
assign w28755 = pi04966 & ~w28751;
assign w28756 = ~pi09812 & w28751;
assign w28757 = ~w28755 & ~w28756;
assign w28758 = pi04967 & ~w28751;
assign w28759 = ~pi02704 & w28751;
assign w28760 = ~w28758 & ~w28759;
assign w28761 = pi04968 & ~w28751;
assign w28762 = ~pi09954 & w28751;
assign w28763 = ~w28761 & ~w28762;
assign w28764 = pi04969 & ~w28751;
assign w28765 = ~pi02720 & w28751;
assign w28766 = ~w28764 & ~w28765;
assign w28767 = pi04970 & ~w28751;
assign w28768 = ~pi09962 & w28751;
assign w28769 = ~w28767 & ~w28768;
assign w28770 = ~w16928 & w19561;
assign w28771 = pi04971 & ~w28770;
assign w28772 = ~pi09961 & w28770;
assign w28773 = ~w28771 & ~w28772;
assign w28774 = pi04972 & ~w28770;
assign w28775 = ~pi09848 & w28770;
assign w28776 = ~w28774 & ~w28775;
assign w28777 = pi04973 & ~w28770;
assign w28778 = ~pi09812 & w28770;
assign w28779 = ~w28777 & ~w28778;
assign w28780 = pi04974 & ~w28770;
assign w28781 = ~pi02704 & w28770;
assign w28782 = ~w28780 & ~w28781;
assign w28783 = pi04975 & ~w28770;
assign w28784 = ~pi09954 & w28770;
assign w28785 = ~w28783 & ~w28784;
assign w28786 = pi04976 & ~w28770;
assign w28787 = ~pi02720 & w28770;
assign w28788 = ~w28786 & ~w28787;
assign w28789 = pi04977 & ~w28770;
assign w28790 = ~pi09962 & w28770;
assign w28791 = ~w28789 & ~w28790;
assign w28792 = ~w16928 & w19552;
assign w28793 = pi04978 & ~w28792;
assign w28794 = ~pi09848 & w28792;
assign w28795 = ~w28793 & ~w28794;
assign w28796 = pi04979 & ~w28792;
assign w28797 = ~pi09812 & w28792;
assign w28798 = ~w28796 & ~w28797;
assign w28799 = pi04980 & ~w28792;
assign w28800 = ~pi02704 & w28792;
assign w28801 = ~w28799 & ~w28800;
assign w28802 = pi04981 & ~w28792;
assign w28803 = ~pi09954 & w28792;
assign w28804 = ~w28802 & ~w28803;
assign w28805 = pi04982 & ~w28792;
assign w28806 = ~pi02720 & w28792;
assign w28807 = ~w28805 & ~w28806;
assign w28808 = pi04983 & ~w28792;
assign w28809 = ~pi09962 & w28792;
assign w28810 = ~w28808 & ~w28809;
assign w28811 = ~w16928 & w19435;
assign w28812 = pi04984 & ~w28811;
assign w28813 = ~pi09961 & w28811;
assign w28814 = ~w28812 & ~w28813;
assign w28815 = pi04985 & ~w28811;
assign w28816 = ~pi09848 & w28811;
assign w28817 = ~w28815 & ~w28816;
assign w28818 = pi04986 & ~w28811;
assign w28819 = ~pi09812 & w28811;
assign w28820 = ~w28818 & ~w28819;
assign w28821 = pi04987 & ~w28811;
assign w28822 = ~pi02704 & w28811;
assign w28823 = ~w28821 & ~w28822;
assign w28824 = pi04988 & ~w28811;
assign w28825 = w17513 & w19435;
assign w28826 = ~w28824 & ~w28825;
assign w28827 = pi04989 & ~w28811;
assign w28828 = ~pi02720 & w28811;
assign w28829 = ~w28827 & ~w28828;
assign w28830 = pi04990 & ~w28811;
assign w28831 = ~pi09962 & w28811;
assign w28832 = ~w28830 & ~w28831;
assign w28833 = ~w16928 & w19530;
assign w28834 = pi04991 & ~w28833;
assign w28835 = ~pi09848 & w28833;
assign w28836 = ~w28834 & ~w28835;
assign w28837 = pi04992 & ~w28833;
assign w28838 = ~pi09812 & w28833;
assign w28839 = ~w28837 & ~w28838;
assign w28840 = pi04993 & ~w28833;
assign w28841 = ~pi02704 & w28833;
assign w28842 = ~w28840 & ~w28841;
assign w28843 = pi04994 & ~w28833;
assign w28844 = ~pi09954 & w28833;
assign w28845 = ~w28843 & ~w28844;
assign w28846 = pi04995 & ~w28833;
assign w28847 = ~pi02720 & w28833;
assign w28848 = ~w28846 & ~w28847;
assign w28849 = pi04996 & ~w28833;
assign w28850 = ~pi09962 & w28833;
assign w28851 = ~w28849 & ~w28850;
assign w28852 = ~w16928 & w19518;
assign w28853 = pi04997 & ~w28852;
assign w28854 = ~pi09961 & w28852;
assign w28855 = ~w28853 & ~w28854;
assign w28856 = pi04998 & ~w28852;
assign w28857 = ~pi09848 & w28852;
assign w28858 = ~w28856 & ~w28857;
assign w28859 = pi04999 & ~w28852;
assign w28860 = ~pi09812 & w28852;
assign w28861 = ~w28859 & ~w28860;
assign w28862 = pi05000 & ~w28852;
assign w28863 = w17311 & w19518;
assign w28864 = ~w28862 & ~w28863;
assign w28865 = pi05001 & ~w28852;
assign w28866 = ~pi09954 & w28852;
assign w28867 = ~w28865 & ~w28866;
assign w28868 = pi05002 & ~w28852;
assign w28869 = ~pi02720 & w28852;
assign w28870 = ~w28868 & ~w28869;
assign w28871 = pi05003 & ~w28852;
assign w28872 = ~pi09962 & w28852;
assign w28873 = ~w28871 & ~w28872;
assign w28874 = ~w16928 & w19492;
assign w28875 = pi05004 & ~w28874;
assign w28876 = ~pi09848 & w28874;
assign w28877 = ~w28875 & ~w28876;
assign w28878 = pi05005 & ~w28874;
assign w28879 = w17193 & w19492;
assign w28880 = ~w28878 & ~w28879;
assign w28881 = pi05006 & ~w28874;
assign w28882 = w17311 & w19492;
assign w28883 = ~w28881 & ~w28882;
assign w28884 = pi05007 & ~w28874;
assign w28885 = ~pi09954 & w28874;
assign w28886 = ~w28884 & ~w28885;
assign w28887 = pi05008 & ~w28874;
assign w28888 = ~pi02720 & w28874;
assign w28889 = ~w28887 & ~w28888;
assign w28890 = pi05009 & ~w28874;
assign w28891 = ~pi09962 & w28874;
assign w28892 = ~w28890 & ~w28891;
assign w28893 = ~w16928 & w19480;
assign w28894 = pi05010 & ~w28893;
assign w28895 = ~pi09961 & w28893;
assign w28896 = ~w28894 & ~w28895;
assign w28897 = pi05011 & ~w28893;
assign w28898 = ~pi09848 & w28893;
assign w28899 = ~w28897 & ~w28898;
assign w28900 = pi05012 & ~w28893;
assign w28901 = ~pi09812 & w28893;
assign w28902 = ~w28900 & ~w28901;
assign w28903 = pi05013 & ~w28893;
assign w28904 = ~pi02704 & w28893;
assign w28905 = ~w28903 & ~w28904;
assign w28906 = pi05014 & ~w28893;
assign w28907 = w18861 & w19480;
assign w28908 = ~w28906 & ~w28907;
assign w28909 = pi05015 & ~w28893;
assign w28910 = ~pi09954 & w28893;
assign w28911 = ~w28909 & ~w28910;
assign w28912 = pi05016 & ~w28893;
assign w28913 = ~pi02720 & w28893;
assign w28914 = ~w28912 & ~w28913;
assign w28915 = pi05017 & ~w28893;
assign w28916 = ~pi09962 & w28893;
assign w28917 = ~w28915 & ~w28916;
assign w28918 = ~w16928 & w19459;
assign w28919 = pi05018 & ~w28918;
assign w28920 = w17186 & w19459;
assign w28921 = ~w28919 & ~w28920;
assign w28922 = pi05019 & ~w28918;
assign w28923 = w17193 & w19459;
assign w28924 = ~w28922 & ~w28923;
assign w28925 = pi05020 & ~w28918;
assign w28926 = ~pi02704 & w28918;
assign w28927 = ~w28925 & ~w28926;
assign w28928 = pi05021 & ~w28918;
assign w28929 = w17513 & w19459;
assign w28930 = ~w28928 & ~w28929;
assign w28931 = pi05022 & ~w28918;
assign w28932 = w17128 & w19459;
assign w28933 = ~w28931 & ~w28932;
assign w28934 = pi05023 & ~w28918;
assign w28935 = w17439 & w19459;
assign w28936 = ~w28934 & ~w28935;
assign w28937 = ~w16928 & w19420;
assign w28938 = pi05024 & ~w28937;
assign w28939 = ~pi09961 & w28937;
assign w28940 = ~w28938 & ~w28939;
assign w28941 = pi05025 & ~w28937;
assign w28942 = ~pi09848 & w28937;
assign w28943 = ~w28941 & ~w28942;
assign w28944 = pi05026 & ~w28937;
assign w28945 = ~pi09812 & w28937;
assign w28946 = ~w28944 & ~w28945;
assign w28947 = pi05027 & ~w28937;
assign w28948 = ~pi02704 & w28937;
assign w28949 = ~w28947 & ~w28948;
assign w28950 = pi05028 & ~w28937;
assign w28951 = ~pi09954 & w28937;
assign w28952 = ~w28950 & ~w28951;
assign w28953 = pi05029 & ~w28937;
assign w28954 = ~pi02720 & w28937;
assign w28955 = ~w28953 & ~w28954;
assign w28956 = pi05030 & ~w28937;
assign w28957 = ~pi09962 & w28937;
assign w28958 = ~w28956 & ~w28957;
assign w28959 = ~w16928 & w19444;
assign w28960 = pi05031 & ~w28959;
assign w28961 = ~pi09848 & w28959;
assign w28962 = ~w28960 & ~w28961;
assign w28963 = pi05032 & ~w28959;
assign w28964 = ~pi09812 & w28959;
assign w28965 = ~w28963 & ~w28964;
assign w28966 = pi05033 & ~w28959;
assign w28967 = w17311 & w19444;
assign w28968 = ~w28966 & ~w28967;
assign w28969 = pi05034 & ~w28959;
assign w28970 = ~pi09954 & w28959;
assign w28971 = ~w28969 & ~w28970;
assign w28972 = pi05035 & ~w28959;
assign w28973 = ~pi02720 & w28959;
assign w28974 = ~w28972 & ~w28973;
assign w28975 = pi05036 & ~w28959;
assign w28976 = w17439 & w19444;
assign w28977 = ~w28975 & ~w28976;
assign w28978 = pi05037 & ~w25500;
assign w28979 = ~pi09961 & w25500;
assign w28980 = ~w28978 & ~w28979;
assign w28981 = pi05038 & ~w25500;
assign w28982 = ~pi09848 & w25500;
assign w28983 = ~w28981 & ~w28982;
assign w28984 = pi05039 & ~w25500;
assign w28985 = ~pi09812 & w25500;
assign w28986 = ~w28984 & ~w28985;
assign w28987 = pi05040 & ~w25500;
assign w28988 = ~pi02704 & w25500;
assign w28989 = ~w28987 & ~w28988;
assign w28990 = pi05041 & ~w25500;
assign w28991 = ~pi09954 & w25500;
assign w28992 = ~w28990 & ~w28991;
assign w28993 = pi05042 & ~w25500;
assign w28994 = ~pi02720 & w25500;
assign w28995 = ~w28993 & ~w28994;
assign w28996 = pi05043 & ~w25500;
assign w28997 = ~pi09962 & w25500;
assign w28998 = ~w28996 & ~w28997;
assign w28999 = pi05044 & ~w22002;
assign w29000 = ~pi09848 & w22002;
assign w29001 = ~w28999 & ~w29000;
assign w29002 = pi05045 & ~w22002;
assign w29003 = ~pi09812 & w22002;
assign w29004 = ~w29002 & ~w29003;
assign w29005 = pi05046 & ~w22002;
assign w29006 = ~pi02704 & w22002;
assign w29007 = ~w29005 & ~w29006;
assign w29008 = pi05047 & ~w22002;
assign w29009 = ~pi09954 & w22002;
assign w29010 = ~w29008 & ~w29009;
assign w29011 = pi05048 & ~w22002;
assign w29012 = ~pi02720 & w22002;
assign w29013 = ~w29011 & ~w29012;
assign w29014 = pi05049 & ~w22002;
assign w29015 = ~pi09962 & w22002;
assign w29016 = ~w29014 & ~w29015;
assign w29017 = pi05050 & ~w21994;
assign w29018 = ~pi09961 & w21994;
assign w29019 = ~w29017 & ~w29018;
assign w29020 = pi05051 & ~w21994;
assign w29021 = ~pi09848 & w21994;
assign w29022 = ~w29020 & ~w29021;
assign w29023 = pi05052 & ~w21994;
assign w29024 = w17193 & w19012;
assign w29025 = ~w29023 & ~w29024;
assign w29026 = pi05053 & ~w21994;
assign w29027 = ~pi02704 & w21994;
assign w29028 = ~w29026 & ~w29027;
assign w29029 = pi05054 & ~w21994;
assign w29030 = ~pi09954 & w21994;
assign w29031 = ~w29029 & ~w29030;
assign w29032 = pi05055 & ~w21994;
assign w29033 = ~pi02720 & w21994;
assign w29034 = ~w29032 & ~w29033;
assign w29035 = pi05056 & ~w21994;
assign w29036 = ~pi09962 & w21994;
assign w29037 = ~w29035 & ~w29036;
assign w29038 = pi05057 & ~w21983;
assign w29039 = w17186 & w19374;
assign w29040 = ~w29038 & ~w29039;
assign w29041 = pi05058 & ~w21983;
assign w29042 = ~pi09812 & w21983;
assign w29043 = ~w29041 & ~w29042;
assign w29044 = pi05059 & ~w21983;
assign w29045 = ~pi02704 & w21983;
assign w29046 = ~w29044 & ~w29045;
assign w29047 = pi05060 & ~w21983;
assign w29048 = ~pi09954 & w21983;
assign w29049 = ~w29047 & ~w29048;
assign w29050 = pi05061 & ~w21983;
assign w29051 = ~pi02720 & w21983;
assign w29052 = ~w29050 & ~w29051;
assign w29053 = pi05062 & ~w21983;
assign w29054 = ~pi09962 & w21983;
assign w29055 = ~w29053 & ~w29054;
assign w29056 = pi05063 & ~w21976;
assign w29057 = ~pi09961 & w21976;
assign w29058 = ~w29056 & ~w29057;
assign w29059 = pi05064 & ~w21976;
assign w29060 = ~pi09848 & w21976;
assign w29061 = ~w29059 & ~w29060;
assign w29062 = pi05065 & ~w21976;
assign w29063 = w17193 & w19348;
assign w29064 = ~w29062 & ~w29063;
assign w29065 = pi05066 & ~w21976;
assign w29066 = w17311 & w19348;
assign w29067 = ~w29065 & ~w29066;
assign w29068 = pi05067 & ~w21976;
assign w29069 = ~pi09954 & w21976;
assign w29070 = ~w29068 & ~w29069;
assign w29071 = pi05068 & ~w21976;
assign w29072 = ~pi02720 & w21976;
assign w29073 = ~w29071 & ~w29072;
assign w29074 = pi05069 & ~w21976;
assign w29075 = ~pi09962 & w21976;
assign w29076 = ~w29074 & ~w29075;
assign w29077 = pi05070 & ~w21962;
assign w29078 = ~pi09848 & w21962;
assign w29079 = ~w29077 & ~w29078;
assign w29080 = pi05071 & ~w21962;
assign w29081 = ~pi09812 & w21962;
assign w29082 = ~w29080 & ~w29081;
assign w29083 = pi05072 & ~w21962;
assign w29084 = ~pi02704 & w21962;
assign w29085 = ~w29083 & ~w29084;
assign w29086 = pi05073 & ~w21958;
assign w29087 = ~pi09961 & w21958;
assign w29088 = ~w29086 & ~w29087;
assign w29089 = pi05074 & ~w21177;
assign w29090 = ~pi09954 & w21177;
assign w29091 = ~w29089 & ~w29090;
assign w29092 = pi05075 & ~w21958;
assign w29093 = ~pi09848 & w21958;
assign w29094 = ~w29092 & ~w29093;
assign w29095 = pi05076 & ~w21958;
assign w29096 = ~pi09812 & w21958;
assign w29097 = ~w29095 & ~w29096;
assign w29098 = pi05077 & ~w21958;
assign w29099 = w17311 & w17361;
assign w29100 = ~w29098 & ~w29099;
assign w29101 = pi05078 & ~w21958;
assign w29102 = ~pi02178 & w21958;
assign w29103 = ~w29101 & ~w29102;
assign w29104 = pi05079 & ~w21958;
assign w29105 = ~pi09954 & w21958;
assign w29106 = ~w29104 & ~w29105;
assign w29107 = pi05080 & ~w21958;
assign w29108 = w17361 & w17439;
assign w29109 = ~w29107 & ~w29108;
assign w29110 = pi05081 & ~w21944;
assign w29111 = ~pi02705 & w21944;
assign w29112 = ~w29110 & ~w29111;
assign w29113 = pi05082 & ~w21944;
assign w29114 = ~pi02706 & w21944;
assign w29115 = ~w29113 & ~w29114;
assign w29116 = pi05083 & ~w21944;
assign w29117 = ~pi02160 & w21944;
assign w29118 = ~w29116 & ~w29117;
assign w29119 = pi05084 & ~w21944;
assign w29120 = ~pi02723 & w21944;
assign w29121 = ~w29119 & ~w29120;
assign w29122 = pi05085 & ~w21944;
assign w29123 = w18689 & w19379;
assign w29124 = ~w29122 & ~w29123;
assign w29125 = pi05086 & ~w21944;
assign w29126 = ~pi02710 & w21944;
assign w29127 = ~w29125 & ~w29126;
assign w29128 = pi05087 & ~w21933;
assign w29129 = ~pi02705 & w21933;
assign w29130 = ~w29128 & ~w29129;
assign w29131 = pi05088 & ~w21933;
assign w29132 = ~pi02706 & w21933;
assign w29133 = ~w29131 & ~w29132;
assign w29134 = pi05089 & ~w21933;
assign w29135 = ~pi02707 & w21933;
assign w29136 = ~w29134 & ~w29135;
assign w29137 = pi05090 & ~w21933;
assign w29138 = ~pi02160 & w21933;
assign w29139 = ~w29137 & ~w29138;
assign w29140 = pi05091 & ~w21933;
assign w29141 = ~pi02723 & w21933;
assign w29142 = ~w29140 & ~w29141;
assign w29143 = pi05092 & ~w21933;
assign w29144 = ~pi02708 & w21933;
assign w29145 = ~w29143 & ~w29144;
assign w29146 = pi05093 & ~w21933;
assign w29147 = ~pi02710 & w21933;
assign w29148 = ~w29146 & ~w29147;
assign w29149 = pi05094 & ~w21411;
assign w29150 = ~pi02705 & w21411;
assign w29151 = ~w29149 & ~w29150;
assign w29152 = pi05095 & ~w21411;
assign w29153 = ~pi02706 & w21411;
assign w29154 = ~w29152 & ~w29153;
assign w29155 = pi05096 & ~w21411;
assign w29156 = ~pi02160 & w21411;
assign w29157 = ~w29155 & ~w29156;
assign w29158 = pi05097 & ~w21411;
assign w29159 = ~pi02723 & w21411;
assign w29160 = ~w29158 & ~w29159;
assign w29161 = pi05098 & ~w21411;
assign w29162 = ~pi02708 & w21411;
assign w29163 = ~w29161 & ~w29162;
assign w29164 = pi05099 & ~w21411;
assign w29165 = ~pi02710 & w21411;
assign w29166 = ~w29164 & ~w29165;
assign w29167 = pi05100 & ~w21166;
assign w29168 = ~pi02705 & w21166;
assign w29169 = ~w29167 & ~w29168;
assign w29170 = pi05101 & ~w21166;
assign w29171 = ~pi02706 & w21166;
assign w29172 = ~w29170 & ~w29171;
assign w29173 = pi05102 & ~w21166;
assign w29174 = ~pi02707 & w21166;
assign w29175 = ~w29173 & ~w29174;
assign w29176 = pi05103 & ~w21166;
assign w29177 = ~pi02160 & w21166;
assign w29178 = ~w29176 & ~w29177;
assign w29179 = pi05104 & ~w21166;
assign w29180 = ~pi02723 & w21166;
assign w29181 = ~w29179 & ~w29180;
assign w29182 = pi05105 & ~w21166;
assign w29183 = ~pi02708 & w21166;
assign w29184 = ~w29182 & ~w29183;
assign w29185 = pi05106 & ~w21166;
assign w29186 = w18027 & w18364;
assign w29187 = ~w29185 & ~w29186;
assign w29188 = pi05107 & ~w21060;
assign w29189 = w17996 & w18578;
assign w29190 = ~w29188 & ~w29189;
assign w29191 = pi05108 & ~w21060;
assign w29192 = ~pi02706 & w21060;
assign w29193 = ~w29191 & ~w29192;
assign w29194 = pi05109 & ~w21060;
assign w29195 = ~pi02160 & w21060;
assign w29196 = ~w29194 & ~w29195;
assign w29197 = pi05110 & ~w21060;
assign w29198 = ~pi02723 & w21060;
assign w29199 = ~w29197 & ~w29198;
assign w29200 = pi05111 & ~w21060;
assign w29201 = ~pi02708 & w21060;
assign w29202 = ~w29200 & ~w29201;
assign w29203 = ~w16992 & w18278;
assign w29204 = pi05112 & ~w29203;
assign w29205 = ~pi02703 & w29203;
assign w29206 = ~w29204 & ~w29205;
assign w29207 = pi05113 & ~w21060;
assign w29208 = w17996 & w18364;
assign w29209 = ~w29207 & ~w29208;
assign w29210 = pi05114 & ~w20450;
assign w29211 = ~pi02705 & w20450;
assign w29212 = ~w29210 & ~w29211;
assign w29213 = pi05115 & ~w20450;
assign w29214 = ~pi02706 & w20450;
assign w29215 = ~w29213 & ~w29214;
assign w29216 = pi05116 & ~w20450;
assign w29217 = w17231 & w18067;
assign w29218 = ~w29216 & ~w29217;
assign w29219 = pi05117 & ~w20450;
assign w29220 = ~pi02160 & w20450;
assign w29221 = ~w29219 & ~w29220;
assign w29222 = pi05118 & ~w20450;
assign w29223 = ~pi02723 & w20450;
assign w29224 = ~w29222 & ~w29223;
assign w29225 = pi05119 & ~w20450;
assign w29226 = ~pi02708 & w20450;
assign w29227 = ~w29225 & ~w29226;
assign w29228 = pi05120 & ~w20450;
assign w29229 = ~pi02710 & w20450;
assign w29230 = ~w29228 & ~w29229;
assign w29231 = pi05121 & ~w20702;
assign w29232 = ~pi02705 & w20702;
assign w29233 = ~w29231 & ~w29232;
assign w29234 = pi05122 & ~w20702;
assign w29235 = ~pi02706 & w20702;
assign w29236 = ~w29234 & ~w29235;
assign w29237 = pi05123 & ~w20702;
assign w29238 = ~pi02160 & w20702;
assign w29239 = ~w29237 & ~w29238;
assign w29240 = pi05124 & ~w20702;
assign w29241 = ~pi02723 & w20702;
assign w29242 = ~w29240 & ~w29241;
assign w29243 = pi05125 & ~w20702;
assign w29244 = ~pi02708 & w20702;
assign w29245 = ~w29243 & ~w29244;
assign w29246 = pi05126 & ~w20702;
assign w29247 = ~pi02710 & w20702;
assign w29248 = ~w29246 & ~w29247;
assign w29249 = pi05127 & ~w20684;
assign w29250 = ~pi02705 & w20684;
assign w29251 = ~w29249 & ~w29250;
assign w29252 = pi05128 & ~w20684;
assign w29253 = ~pi02706 & w20684;
assign w29254 = ~w29252 & ~w29253;
assign w29255 = pi05129 & ~w20684;
assign w29256 = ~pi02707 & w20684;
assign w29257 = ~w29255 & ~w29256;
assign w29258 = pi05130 & ~w20684;
assign w29259 = ~pi02160 & w20684;
assign w29260 = ~w29258 & ~w29259;
assign w29261 = pi05131 & ~w20684;
assign w29262 = ~pi02723 & w20684;
assign w29263 = ~w29261 & ~w29262;
assign w29264 = pi05132 & ~w20684;
assign w29265 = ~pi02708 & w20684;
assign w29266 = ~w29264 & ~w29265;
assign w29267 = pi05133 & ~w20684;
assign w29268 = ~pi02710 & w20684;
assign w29269 = ~w29267 & ~w29268;
assign w29270 = pi05134 & ~w20660;
assign w29271 = ~pi02705 & w20660;
assign w29272 = ~w29270 & ~w29271;
assign w29273 = pi05135 & ~w20660;
assign w29274 = ~pi02706 & w20660;
assign w29275 = ~w29273 & ~w29274;
assign w29276 = pi05136 & ~w20660;
assign w29277 = ~pi02160 & w20660;
assign w29278 = ~w29276 & ~w29277;
assign w29279 = pi05137 & ~w20660;
assign w29280 = ~pi02723 & w20660;
assign w29281 = ~w29279 & ~w29280;
assign w29282 = pi05138 & ~w20660;
assign w29283 = ~pi02708 & w20660;
assign w29284 = ~w29282 & ~w29283;
assign w29285 = pi05139 & ~w20660;
assign w29286 = ~pi02710 & w20660;
assign w29287 = ~w29285 & ~w29286;
assign w29288 = pi05140 & ~w20629;
assign w29289 = ~pi02705 & w20629;
assign w29290 = ~w29288 & ~w29289;
assign w29291 = pi05141 & ~w20629;
assign w29292 = ~pi02706 & w20629;
assign w29293 = ~w29291 & ~w29292;
assign w29294 = pi05142 & ~w20629;
assign w29295 = ~pi02707 & w20629;
assign w29296 = ~w29294 & ~w29295;
assign w29297 = pi05143 & ~w20629;
assign w29298 = ~pi02160 & w20629;
assign w29299 = ~w29297 & ~w29298;
assign w29300 = pi05144 & ~w20629;
assign w29301 = ~pi02723 & w20629;
assign w29302 = ~w29300 & ~w29301;
assign w29303 = pi05145 & ~w20629;
assign w29304 = ~pi02708 & w20629;
assign w29305 = ~w29303 & ~w29304;
assign w29306 = pi05146 & ~w20629;
assign w29307 = ~pi02710 & w20629;
assign w29308 = ~w29306 & ~w29307;
assign w29309 = pi05147 & ~w18848;
assign w29310 = ~pi09954 & w18848;
assign w29311 = ~w29309 & ~w29310;
assign w29312 = pi05148 & ~w20588;
assign w29313 = ~pi02705 & w20588;
assign w29314 = ~w29312 & ~w29313;
assign w29315 = pi05149 & ~w20588;
assign w29316 = ~pi02707 & w20588;
assign w29317 = ~w29315 & ~w29316;
assign w29318 = pi05150 & ~w20588;
assign w29319 = ~pi02160 & w20588;
assign w29320 = ~w29318 & ~w29319;
assign w29321 = pi05151 & ~w20588;
assign w29322 = ~pi02723 & w20588;
assign w29323 = ~w29321 & ~w29322;
assign w29324 = pi05152 & ~w20588;
assign w29325 = ~pi02709 & w20588;
assign w29326 = ~w29324 & ~w29325;
assign w29327 = pi05153 & ~w20588;
assign w29328 = w16941 & w18364;
assign w29329 = ~w29327 & ~w29328;
assign w29330 = pi05154 & ~w20545;
assign w29331 = ~pi02705 & w20545;
assign w29332 = ~w29330 & ~w29331;
assign w29333 = pi05155 & ~w20545;
assign w29334 = ~pi02706 & w20545;
assign w29335 = ~w29333 & ~w29334;
assign w29336 = pi05156 & ~w20545;
assign w29337 = ~pi02707 & w20545;
assign w29338 = ~w29336 & ~w29337;
assign w29339 = pi05157 & ~w20545;
assign w29340 = w18234 & w18278;
assign w29341 = ~w29339 & ~w29340;
assign w29342 = pi05158 & ~w20545;
assign w29343 = ~pi02723 & w20545;
assign w29344 = ~w29342 & ~w29343;
assign w29345 = pi05159 & ~w20545;
assign w29346 = w18092 & w18278;
assign w29347 = ~w29345 & ~w29346;
assign w29348 = pi05160 & ~w20545;
assign w29349 = ~pi02710 & w20545;
assign w29350 = ~w29348 & ~w29349;
assign w29351 = pi05161 & ~w20538;
assign w29352 = ~pi02705 & w20538;
assign w29353 = ~w29351 & ~w29352;
assign w29354 = pi05162 & ~w20538;
assign w29355 = ~pi02707 & w20538;
assign w29356 = ~w29354 & ~w29355;
assign w29357 = pi05163 & ~w20538;
assign w29358 = ~pi02160 & w20538;
assign w29359 = ~w29357 & ~w29358;
assign w29360 = pi05164 & ~w20538;
assign w29361 = ~pi02723 & w20538;
assign w29362 = ~w29360 & ~w29361;
assign w29363 = pi05165 & ~w20538;
assign w29364 = ~pi02709 & w20538;
assign w29365 = ~w29363 & ~w29364;
assign w29366 = pi05166 & ~w20538;
assign w29367 = ~pi02710 & w20538;
assign w29368 = ~w29366 & ~w29367;
assign w29369 = pi05167 & ~w20478;
assign w29370 = ~pi02705 & w20478;
assign w29371 = ~w29369 & ~w29370;
assign w29372 = pi05168 & ~w20478;
assign w29373 = ~pi02706 & w20478;
assign w29374 = ~w29372 & ~w29373;
assign w29375 = pi05169 & ~w20478;
assign w29376 = ~pi02707 & w20478;
assign w29377 = ~w29375 & ~w29376;
assign w29378 = pi05170 & ~w20478;
assign w29379 = ~pi02160 & w20478;
assign w29380 = ~w29378 & ~w29379;
assign w29381 = pi05171 & ~w20478;
assign w29382 = ~pi02723 & w20478;
assign w29383 = ~w29381 & ~w29382;
assign w29384 = pi05172 & ~w20478;
assign w29385 = ~pi02709 & w20478;
assign w29386 = ~w29384 & ~w29385;
assign w29387 = pi05173 & ~w20478;
assign w29388 = w17837 & w18364;
assign w29389 = ~w29387 & ~w29388;
assign w29390 = pi05174 & ~w21270;
assign w29391 = ~pi02704 & w21270;
assign w29392 = ~w29390 & ~w29391;
assign w29393 = pi05175 & ~w20466;
assign w29394 = ~pi02706 & w20466;
assign w29395 = ~w29393 & ~w29394;
assign w29396 = pi05176 & ~w20466;
assign w29397 = ~pi02707 & w20466;
assign w29398 = ~w29396 & ~w29397;
assign w29399 = pi05177 & ~w20466;
assign w29400 = ~pi02160 & w20466;
assign w29401 = ~w29399 & ~w29400;
assign w29402 = pi05178 & ~w20466;
assign w29403 = ~pi02708 & w20466;
assign w29404 = ~w29402 & ~w29403;
assign w29405 = pi05179 & ~w20466;
assign w29406 = ~pi02709 & w20466;
assign w29407 = ~w29405 & ~w29406;
assign w29408 = pi05180 & ~w20466;
assign w29409 = ~pi02710 & w20466;
assign w29410 = ~w29408 & ~w29409;
assign w29411 = pi05181 & ~w20457;
assign w29412 = ~pi02705 & w20457;
assign w29413 = ~w29411 & ~w29412;
assign w29414 = pi05182 & ~w20457;
assign w29415 = ~pi02706 & w20457;
assign w29416 = ~w29414 & ~w29415;
assign w29417 = pi05183 & ~w20457;
assign w29418 = ~pi02707 & w20457;
assign w29419 = ~w29417 & ~w29418;
assign w29420 = pi05184 & ~w20457;
assign w29421 = ~pi02160 & w20457;
assign w29422 = ~w29420 & ~w29421;
assign w29423 = pi05185 & ~w20457;
assign w29424 = ~pi02708 & w20457;
assign w29425 = ~w29423 & ~w29424;
assign w29426 = pi05186 & ~w20457;
assign w29427 = ~pi02709 & w20457;
assign w29428 = ~w29426 & ~w29427;
assign w29429 = pi05187 & ~w20457;
assign w29430 = ~pi02710 & w20457;
assign w29431 = ~w29429 & ~w29430;
assign w29432 = pi05188 & ~w20415;
assign w29433 = ~pi02706 & w20415;
assign w29434 = ~w29432 & ~w29433;
assign w29435 = pi05189 & ~w20415;
assign w29436 = w17822 & w18067;
assign w29437 = ~w29435 & ~w29436;
assign w29438 = pi05190 & ~w20415;
assign w29439 = ~pi02160 & w20415;
assign w29440 = ~w29438 & ~w29439;
assign w29441 = pi05191 & ~w20415;
assign w29442 = ~pi02708 & w20415;
assign w29443 = ~w29441 & ~w29442;
assign w29444 = pi05192 & ~w20415;
assign w29445 = ~pi02709 & w20415;
assign w29446 = ~w29444 & ~w29445;
assign w29447 = pi05193 & ~w20415;
assign w29448 = ~pi02710 & w20415;
assign w29449 = ~w29447 & ~w29448;
assign w29450 = pi05194 & ~w18531;
assign w29451 = ~pi02705 & w18531;
assign w29452 = ~w29450 & ~w29451;
assign w29453 = pi05195 & ~w18531;
assign w29454 = w17775 & w17925;
assign w29455 = ~w29453 & ~w29454;
assign w29456 = pi05196 & ~w18531;
assign w29457 = w17775 & w18067;
assign w29458 = ~w29456 & ~w29457;
assign w29459 = pi05197 & ~w18531;
assign w29460 = ~pi02160 & w18531;
assign w29461 = ~w29459 & ~w29460;
assign w29462 = pi05198 & ~w18531;
assign w29463 = ~pi02708 & w18531;
assign w29464 = ~w29462 & ~w29463;
assign w29465 = pi05199 & ~w18531;
assign w29466 = ~pi02709 & w18531;
assign w29467 = ~w29465 & ~w29466;
assign w29468 = pi05200 & ~w18531;
assign w29469 = w17775 & w18364;
assign w29470 = ~w29468 & ~w29469;
assign w29471 = pi05201 & ~w20386;
assign w29472 = ~pi02706 & w20386;
assign w29473 = ~w29471 & ~w29472;
assign w29474 = pi05202 & ~w20386;
assign w29475 = ~pi02707 & w20386;
assign w29476 = ~w29474 & ~w29475;
assign w29477 = pi05203 & ~w20386;
assign w29478 = ~pi02160 & w20386;
assign w29479 = ~w29477 & ~w29478;
assign w29480 = pi05204 & ~w20386;
assign w29481 = ~pi02708 & w20386;
assign w29482 = ~w29480 & ~w29481;
assign w29483 = pi05205 & ~w20386;
assign w29484 = ~pi02709 & w20386;
assign w29485 = ~w29483 & ~w29484;
assign w29486 = pi05206 & ~w20386;
assign w29487 = w17573 & w18364;
assign w29488 = ~w29486 & ~w29487;
assign w29489 = pi05207 & ~w20147;
assign w29490 = w17028 & w18578;
assign w29491 = ~w29489 & ~w29490;
assign w29492 = pi05208 & ~w20147;
assign w29493 = w17028 & w17925;
assign w29494 = ~w29492 & ~w29493;
assign w29495 = pi05209 & ~w20147;
assign w29496 = w17028 & w18067;
assign w29497 = ~w29495 & ~w29496;
assign w29498 = pi05210 & ~w20147;
assign w29499 = w17028 & w18234;
assign w29500 = ~w29498 & ~w29499;
assign w29501 = pi05211 & ~w20147;
assign w29502 = w17028 & w18689;
assign w29503 = ~w29501 & ~w29502;
assign w29504 = pi05212 & ~w20147;
assign w29505 = w17028 & w18092;
assign w29506 = ~w29504 & ~w29505;
assign w29507 = pi05213 & ~w20147;
assign w29508 = w17028 & w18364;
assign w29509 = ~w29507 & ~w29508;
assign w29510 = pi05214 & ~w20111;
assign w29511 = w17053 & w17925;
assign w29512 = ~w29510 & ~w29511;
assign w29513 = pi05215 & ~w20111;
assign w29514 = ~pi02707 & w20111;
assign w29515 = ~w29513 & ~w29514;
assign w29516 = pi05216 & ~w20111;
assign w29517 = ~pi02160 & w20111;
assign w29518 = ~w29516 & ~w29517;
assign w29519 = pi05217 & ~w20111;
assign w29520 = ~pi02708 & w20111;
assign w29521 = ~w29519 & ~w29520;
assign w29522 = pi05218 & ~w20111;
assign w29523 = ~pi02709 & w20111;
assign w29524 = ~w29522 & ~w29523;
assign w29525 = pi05219 & ~w20111;
assign w29526 = ~pi02710 & w20111;
assign w29527 = ~w29525 & ~w29526;
assign w29528 = pi05220 & ~w19926;
assign w29529 = ~pi02705 & w19926;
assign w29530 = ~w29528 & ~w29529;
assign w29531 = pi05221 & ~w19926;
assign w29532 = ~pi02706 & w19926;
assign w29533 = ~w29531 & ~w29532;
assign w29534 = pi05222 & ~w19926;
assign w29535 = ~pi02707 & w19926;
assign w29536 = ~w29534 & ~w29535;
assign w29537 = pi05223 & ~w19926;
assign w29538 = ~pi02160 & w19926;
assign w29539 = ~w29537 & ~w29538;
assign w29540 = pi05224 & ~w19926;
assign w29541 = ~pi02708 & w19926;
assign w29542 = ~w29540 & ~w29541;
assign w29543 = pi05225 & ~w19926;
assign w29544 = ~pi02709 & w19926;
assign w29545 = ~w29543 & ~w29544;
assign w29546 = pi05226 & ~w19926;
assign w29547 = ~pi02710 & w19926;
assign w29548 = ~w29546 & ~w29547;
assign w29549 = pi05227 & ~w19787;
assign w29550 = ~pi02706 & w19787;
assign w29551 = ~w29549 & ~w29550;
assign w29552 = pi05228 & ~w19787;
assign w29553 = ~pi02707 & w19787;
assign w29554 = ~w29552 & ~w29553;
assign w29555 = pi05229 & ~w19787;
assign w29556 = ~pi02160 & w19787;
assign w29557 = ~w29555 & ~w29556;
assign w29558 = pi05230 & ~w19787;
assign w29559 = ~pi02708 & w19787;
assign w29560 = ~w29558 & ~w29559;
assign w29561 = pi05231 & ~w19787;
assign w29562 = ~pi02709 & w19787;
assign w29563 = ~w29561 & ~w29562;
assign w29564 = pi05232 & ~w19787;
assign w29565 = ~pi02710 & w19787;
assign w29566 = ~w29564 & ~w29565;
assign w29567 = pi05233 & ~w19876;
assign w29568 = ~pi02705 & w19876;
assign w29569 = ~w29567 & ~w29568;
assign w29570 = pi05234 & ~w19876;
assign w29571 = w17406 & w17925;
assign w29572 = ~w29570 & ~w29571;
assign w29573 = pi05235 & ~w19876;
assign w29574 = w17406 & w18067;
assign w29575 = ~w29573 & ~w29574;
assign w29576 = pi05236 & ~w19876;
assign w29577 = ~pi02160 & w19876;
assign w29578 = ~w29576 & ~w29577;
assign w29579 = pi05237 & ~w19876;
assign w29580 = ~pi02708 & w19876;
assign w29581 = ~w29579 & ~w29580;
assign w29582 = pi05238 & ~w19876;
assign w29583 = w17406 & w18092;
assign w29584 = ~w29582 & ~w29583;
assign w29585 = pi05239 & ~w19876;
assign w29586 = ~pi02710 & w19876;
assign w29587 = ~w29585 & ~w29586;
assign w29588 = pi05240 & ~w19630;
assign w29589 = ~pi02706 & w19630;
assign w29590 = ~w29588 & ~w29589;
assign w29591 = pi05241 & ~w19630;
assign w29592 = ~pi02707 & w19630;
assign w29593 = ~w29591 & ~w29592;
assign w29594 = pi05242 & ~w19630;
assign w29595 = w18234 & w19629;
assign w29596 = ~w29594 & ~w29595;
assign w29597 = pi05243 & ~w19630;
assign w29598 = ~pi02708 & w19630;
assign w29599 = ~w29597 & ~w29598;
assign w29600 = pi05244 & ~w19630;
assign w29601 = ~pi02709 & w19630;
assign w29602 = ~w29600 & ~w29601;
assign w29603 = pi05245 & ~w19630;
assign w29604 = ~pi02710 & w19630;
assign w29605 = ~w29603 & ~w29604;
assign w29606 = pi05246 & ~w19656;
assign w29607 = ~pi02705 & w19656;
assign w29608 = ~w29606 & ~w29607;
assign w29609 = pi05247 & ~w19656;
assign w29610 = ~pi02706 & w19656;
assign w29611 = ~w29609 & ~w29610;
assign w29612 = pi05248 & ~w19656;
assign w29613 = ~pi02707 & w19656;
assign w29614 = ~w29612 & ~w29613;
assign w29615 = pi05249 & ~w19656;
assign w29616 = ~pi02160 & w19656;
assign w29617 = ~w29615 & ~w29616;
assign w29618 = pi05250 & ~w19656;
assign w29619 = ~pi02708 & w19656;
assign w29620 = ~w29618 & ~w29619;
assign w29621 = pi05251 & ~w19656;
assign w29622 = ~pi02709 & w19656;
assign w29623 = ~w29621 & ~w29622;
assign w29624 = pi05252 & ~w19656;
assign w29625 = w18364 & w19655;
assign w29626 = ~w29624 & ~w29625;
assign w29627 = pi05253 & ~w19597;
assign w29628 = ~pi02706 & w19597;
assign w29629 = ~w29627 & ~w29628;
assign w29630 = pi05254 & ~w19597;
assign w29631 = ~pi02707 & w19597;
assign w29632 = ~w29630 & ~w29631;
assign w29633 = pi05255 & ~w19597;
assign w29634 = ~pi02160 & w19597;
assign w29635 = ~w29633 & ~w29634;
assign w29636 = pi05256 & ~w19597;
assign w29637 = ~pi02708 & w19597;
assign w29638 = ~w29636 & ~w29637;
assign w29639 = pi05257 & ~w19597;
assign w29640 = ~pi02709 & w19597;
assign w29641 = ~w29639 & ~w29640;
assign w29642 = pi05258 & ~w19597;
assign w29643 = ~pi02710 & w19597;
assign w29644 = ~w29642 & ~w29643;
assign w29645 = pi05259 & ~w19523;
assign w29646 = w17279 & w18578;
assign w29647 = ~w29645 & ~w29646;
assign w29648 = pi05260 & ~w19523;
assign w29649 = w17279 & w17925;
assign w29650 = ~w29648 & ~w29649;
assign w29651 = pi05261 & ~w19523;
assign w29652 = w17279 & w18067;
assign w29653 = ~w29651 & ~w29652;
assign w29654 = pi05262 & ~w19523;
assign w29655 = w17279 & w18234;
assign w29656 = ~w29654 & ~w29655;
assign w29657 = pi05263 & ~w19523;
assign w29658 = w17279 & w18689;
assign w29659 = ~w29657 & ~w29658;
assign w29660 = pi05264 & ~w19523;
assign w29661 = w17279 & w18092;
assign w29662 = ~w29660 & ~w29661;
assign w29663 = pi05265 & ~w19523;
assign w29664 = w17279 & w18364;
assign w29665 = ~w29663 & ~w29664;
assign w29666 = pi05266 & ~w19283;
assign w29667 = ~pi02706 & w19283;
assign w29668 = ~w29666 & ~w29667;
assign w29669 = pi05267 & ~w19283;
assign w29670 = ~pi02707 & w19283;
assign w29671 = ~w29669 & ~w29670;
assign w29672 = pi05268 & ~w19283;
assign w29673 = ~pi02160 & w19283;
assign w29674 = ~w29672 & ~w29673;
assign w29675 = pi05269 & ~w19283;
assign w29676 = ~pi02708 & w19283;
assign w29677 = ~w29675 & ~w29676;
assign w29678 = pi05270 & ~w19283;
assign w29679 = ~pi02709 & w19283;
assign w29680 = ~w29678 & ~w29679;
assign w29681 = pi05271 & ~w19283;
assign w29682 = ~pi02710 & w19283;
assign w29683 = ~w29681 & ~w29682;
assign w29684 = pi05272 & ~w19000;
assign w29685 = ~pi02705 & w19000;
assign w29686 = ~w29684 & ~w29685;
assign w29687 = pi05273 & ~w19000;
assign w29688 = ~pi02706 & w19000;
assign w29689 = ~w29687 & ~w29688;
assign w29690 = pi05274 & ~w19000;
assign w29691 = ~pi02707 & w19000;
assign w29692 = ~w29690 & ~w29691;
assign w29693 = pi05275 & ~w19000;
assign w29694 = w18234 & w18726;
assign w29695 = ~w29693 & ~w29694;
assign w29696 = pi05276 & ~w19000;
assign w29697 = ~pi02708 & w19000;
assign w29698 = ~w29696 & ~w29697;
assign w29699 = pi05277 & ~w19000;
assign w29700 = ~pi02709 & w19000;
assign w29701 = ~w29699 & ~w29700;
assign w29702 = pi05278 & ~w19000;
assign w29703 = w18364 & w18726;
assign w29704 = ~w29702 & ~w29703;
assign w29705 = pi05279 & ~w19210;
assign w29706 = ~pi02706 & w19210;
assign w29707 = ~w29705 & ~w29706;
assign w29708 = pi05280 & ~w19210;
assign w29709 = ~pi02707 & w19210;
assign w29710 = ~w29708 & ~w29709;
assign w29711 = pi05281 & ~w19210;
assign w29712 = ~pi02160 & w19210;
assign w29713 = ~w29711 & ~w29712;
assign w29714 = pi05282 & ~w19210;
assign w29715 = ~pi02708 & w19210;
assign w29716 = ~w29714 & ~w29715;
assign w29717 = pi05283 & ~w19210;
assign w29718 = ~pi02709 & w19210;
assign w29719 = ~w29717 & ~w29718;
assign w29720 = pi05284 & ~w19210;
assign w29721 = ~pi02710 & w19210;
assign w29722 = ~w29720 & ~w29721;
assign w29723 = pi05285 & ~w19138;
assign w29724 = ~pi02705 & w19138;
assign w29725 = ~w29723 & ~w29724;
assign w29726 = pi05286 & ~w19138;
assign w29727 = ~pi02706 & w19138;
assign w29728 = ~w29726 & ~w29727;
assign w29729 = pi05287 & ~w19138;
assign w29730 = ~pi02707 & w19138;
assign w29731 = ~w29729 & ~w29730;
assign w29732 = pi05288 & ~w19138;
assign w29733 = ~pi02160 & w19138;
assign w29734 = ~w29732 & ~w29733;
assign w29735 = pi05289 & ~w19138;
assign w29736 = ~pi02708 & w19138;
assign w29737 = ~w29735 & ~w29736;
assign w29738 = pi05290 & ~w19138;
assign w29739 = ~pi02709 & w19138;
assign w29740 = ~w29738 & ~w29739;
assign w29741 = pi05291 & ~w19138;
assign w29742 = ~pi02710 & w19138;
assign w29743 = ~w29741 & ~w29742;
assign w29744 = pi05292 & ~w21367;
assign w29745 = ~pi09812 & w21367;
assign w29746 = ~w29744 & ~w29745;
assign w29747 = pi05293 & ~w19111;
assign w29748 = ~pi02706 & w19111;
assign w29749 = ~w29747 & ~w29748;
assign w29750 = pi05294 & ~w19111;
assign w29751 = ~pi02707 & w19111;
assign w29752 = ~w29750 & ~w29751;
assign w29753 = pi05295 & ~w19111;
assign w29754 = ~pi02723 & w19111;
assign w29755 = ~w29753 & ~w29754;
assign w29756 = pi05296 & ~w19111;
assign w29757 = ~pi02708 & w19111;
assign w29758 = ~w29756 & ~w29757;
assign w29759 = pi05297 & ~w19111;
assign w29760 = ~pi02709 & w19111;
assign w29761 = ~w29759 & ~w29760;
assign w29762 = pi05298 & ~w19111;
assign w29763 = ~pi02710 & w19111;
assign w29764 = ~w29762 & ~w29763;
assign w29765 = pi05299 & ~w18794;
assign w29766 = ~pi02705 & w18794;
assign w29767 = ~w29765 & ~w29766;
assign w29768 = pi05300 & ~w18794;
assign w29769 = ~pi02706 & w18794;
assign w29770 = ~w29768 & ~w29769;
assign w29771 = pi05301 & ~w18794;
assign w29772 = ~pi02707 & w18794;
assign w29773 = ~w29771 & ~w29772;
assign w29774 = pi05302 & ~w18794;
assign w29775 = ~pi02723 & w18794;
assign w29776 = ~w29774 & ~w29775;
assign w29777 = pi05303 & ~w18794;
assign w29778 = ~pi02708 & w18794;
assign w29779 = ~w29777 & ~w29778;
assign w29780 = pi05304 & ~w18794;
assign w29781 = ~pi02709 & w18794;
assign w29782 = ~w29780 & ~w29781;
assign w29783 = pi05305 & ~w18971;
assign w29784 = w17084 & w18578;
assign w29785 = ~w29783 & ~w29784;
assign w29786 = pi05306 & ~w18971;
assign w29787 = w17084 & w17925;
assign w29788 = ~w29786 & ~w29787;
assign w29789 = pi05307 & ~w18971;
assign w29790 = w17084 & w18067;
assign w29791 = ~w29789 & ~w29790;
assign w29792 = pi05308 & ~w18971;
assign w29793 = w17084 & w17671;
assign w29794 = ~w29792 & ~w29793;
assign w29795 = pi05309 & ~w18971;
assign w29796 = w17084 & w18689;
assign w29797 = ~w29795 & ~w29796;
assign w29798 = pi05310 & ~w18971;
assign w29799 = w17084 & w18092;
assign w29800 = ~w29798 & ~w29799;
assign w29801 = pi05311 & ~w18971;
assign w29802 = w17084 & w18364;
assign w29803 = ~w29801 & ~w29802;
assign w29804 = pi05312 & ~w18893;
assign w29805 = ~pi02705 & w18893;
assign w29806 = ~w29804 & ~w29805;
assign w29807 = pi05313 & ~w18893;
assign w29808 = ~pi02706 & w18893;
assign w29809 = ~w29807 & ~w29808;
assign w29810 = pi05314 & ~w18893;
assign w29811 = ~pi02707 & w18893;
assign w29812 = ~w29810 & ~w29811;
assign w29813 = pi05315 & ~w18893;
assign w29814 = w16970 & w17671;
assign w29815 = ~w29813 & ~w29814;
assign w29816 = pi05316 & ~w18893;
assign w29817 = ~pi02708 & w18893;
assign w29818 = ~w29816 & ~w29817;
assign w29819 = pi05317 & ~w18893;
assign w29820 = ~pi02709 & w18893;
assign w29821 = ~w29819 & ~w29820;
assign w29822 = pi05318 & ~w18879;
assign w29823 = ~pi02705 & w18879;
assign w29824 = ~w29822 & ~w29823;
assign w29825 = pi05319 & ~w18879;
assign w29826 = ~pi02706 & w18879;
assign w29827 = ~w29825 & ~w29826;
assign w29828 = pi05320 & ~w18879;
assign w29829 = w17808 & w18067;
assign w29830 = ~w29828 & ~w29829;
assign w29831 = pi05321 & ~w18879;
assign w29832 = ~pi02723 & w18879;
assign w29833 = ~w29831 & ~w29832;
assign w29834 = pi05322 & ~w21356;
assign w29835 = ~pi02178 & w21356;
assign w29836 = ~w29834 & ~w29835;
assign w29837 = pi05323 & ~w18879;
assign w29838 = ~pi02708 & w18879;
assign w29839 = ~w29837 & ~w29838;
assign w29840 = pi05324 & ~w18879;
assign w29841 = ~pi02709 & w18879;
assign w29842 = ~w29840 & ~w29841;
assign w29843 = pi05325 & ~w18879;
assign w29844 = ~pi02710 & w18879;
assign w29845 = ~w29843 & ~w29844;
assign w29846 = pi05326 & ~w17280;
assign w29847 = ~pi02178 & w17280;
assign w29848 = ~w29846 & ~w29847;
assign w29849 = pi05327 & ~w18827;
assign w29850 = ~pi02705 & w18827;
assign w29851 = ~w29849 & ~w29850;
assign w29852 = pi05328 & ~w18827;
assign w29853 = ~pi02707 & w18827;
assign w29854 = ~w29852 & ~w29853;
assign w29855 = pi05329 & ~w18827;
assign w29856 = ~pi02160 & w18827;
assign w29857 = ~w29855 & ~w29856;
assign w29858 = pi05330 & ~w18827;
assign w29859 = ~pi02723 & w18827;
assign w29860 = ~w29858 & ~w29859;
assign w29861 = pi05331 & ~w18827;
assign w29862 = ~pi02709 & w18827;
assign w29863 = ~w29861 & ~w29862;
assign w29864 = pi05332 & ~w18827;
assign w29865 = ~pi02710 & w18827;
assign w29866 = ~w29864 & ~w29865;
assign w29867 = pi05333 & ~w18714;
assign w29868 = ~pi02705 & w18714;
assign w29869 = ~w29867 & ~w29868;
assign w29870 = pi05334 & ~w18714;
assign w29871 = w17495 & w18067;
assign w29872 = ~w29870 & ~w29871;
assign w29873 = pi05335 & ~w18714;
assign w29874 = ~pi02160 & w18714;
assign w29875 = ~w29873 & ~w29874;
assign w29876 = pi05336 & ~w18714;
assign w29877 = w17495 & w18689;
assign w29878 = ~w29876 & ~w29877;
assign w29879 = pi05337 & ~w18714;
assign w29880 = ~pi02709 & w18714;
assign w29881 = ~w29879 & ~w29880;
assign w29882 = pi05338 & ~w18714;
assign w29883 = ~pi02723 & w18714;
assign w29884 = ~w29882 & ~w29883;
assign w29885 = pi05339 & ~w18714;
assign w29886 = ~pi02710 & w18714;
assign w29887 = ~w29885 & ~w29886;
assign w29888 = pi05340 & ~w18014;
assign w29889 = w17450 & w18578;
assign w29890 = ~w29888 & ~w29889;
assign w29891 = pi05341 & ~w18014;
assign w29892 = w17450 & w18067;
assign w29893 = ~w29891 & ~w29892;
assign w29894 = pi05342 & ~w18014;
assign w29895 = w17450 & w18234;
assign w29896 = ~w29894 & ~w29895;
assign w29897 = pi05343 & ~w18014;
assign w29898 = w17450 & w17671;
assign w29899 = ~w29897 & ~w29898;
assign w29900 = pi05344 & ~w18014;
assign w29901 = w17450 & w18092;
assign w29902 = ~w29900 & ~w29901;
assign w29903 = pi05345 & ~w18014;
assign w29904 = w17450 & w18364;
assign w29905 = ~w29903 & ~w29904;
assign w29906 = pi05346 & ~w18496;
assign w29907 = ~pi02705 & w18496;
assign w29908 = ~w29906 & ~w29907;
assign w29909 = pi05347 & ~w18496;
assign w29910 = ~pi02707 & w18496;
assign w29911 = ~w29909 & ~w29910;
assign w29912 = pi05348 & ~w21162;
assign w29913 = ~pi02720 & w21162;
assign w29914 = ~w29912 & ~w29913;
assign w29915 = pi05349 & ~w18496;
assign w29916 = w17436 & w18234;
assign w29917 = ~w29915 & ~w29916;
assign w29918 = pi05350 & ~w18496;
assign w29919 = w17436 & w17671;
assign w29920 = ~w29918 & ~w29919;
assign w29921 = pi05351 & ~w18496;
assign w29922 = ~pi02708 & w18496;
assign w29923 = ~w29921 & ~w29922;
assign w29924 = pi05352 & ~w18496;
assign w29925 = w17436 & w18092;
assign w29926 = ~w29924 & ~w29925;
assign w29927 = pi05353 & ~w18496;
assign w29928 = ~pi02710 & w18496;
assign w29929 = ~w29927 & ~w29928;
assign w29930 = pi05354 & ~w18389;
assign w29931 = ~pi02706 & w18389;
assign w29932 = ~w29930 & ~w29931;
assign w29933 = pi05355 & ~w18389;
assign w29934 = ~pi02707 & w18389;
assign w29935 = ~w29933 & ~w29934;
assign w29936 = pi05356 & ~w18389;
assign w29937 = ~pi02160 & w18389;
assign w29938 = ~w29936 & ~w29937;
assign w29939 = pi05357 & ~w18389;
assign w29940 = ~pi02708 & w18389;
assign w29941 = ~w29939 & ~w29940;
assign w29942 = pi05358 & ~w18389;
assign w29943 = ~pi02709 & w18389;
assign w29944 = ~w29942 & ~w29943;
assign w29945 = pi05359 & ~w18389;
assign w29946 = ~pi02710 & w18389;
assign w29947 = ~w29945 & ~w29946;
assign w29948 = pi05360 & ~w18362;
assign w29949 = ~pi02706 & w18362;
assign w29950 = ~w29948 & ~w29949;
assign w29951 = pi05361 & ~w18362;
assign w29952 = ~pi02707 & w18362;
assign w29953 = ~w29951 & ~w29952;
assign w29954 = pi05362 & ~w18362;
assign w29955 = ~pi02160 & w18362;
assign w29956 = ~w29954 & ~w29955;
assign w29957 = pi05363 & ~w18362;
assign w29958 = w16912 & w17671;
assign w29959 = ~w29957 & ~w29958;
assign w29960 = pi05364 & ~w18362;
assign w29961 = ~pi02708 & w18362;
assign w29962 = ~w29960 & ~w29961;
assign w29963 = pi05365 & ~w18362;
assign w29964 = w16912 & w18092;
assign w29965 = ~w29963 & ~w29964;
assign w29966 = pi05366 & ~w21000;
assign w29967 = w17311 & w19655;
assign w29968 = ~w29966 & ~w29967;
assign w29969 = pi05367 & ~w18287;
assign w29970 = ~pi02705 & w18287;
assign w29971 = ~w29969 & ~w29970;
assign w29972 = pi05368 & ~w18287;
assign w29973 = ~pi02706 & w18287;
assign w29974 = ~w29972 & ~w29973;
assign w29975 = pi05369 & ~w18287;
assign w29976 = ~pi02707 & w18287;
assign w29977 = ~w29975 & ~w29976;
assign w29978 = pi05370 & ~w18287;
assign w29979 = ~pi02723 & w18287;
assign w29980 = ~w29978 & ~w29979;
assign w29981 = pi05371 & ~w18287;
assign w29982 = w17284 & w18689;
assign w29983 = ~w29981 & ~w29982;
assign w29984 = pi05372 & ~w18287;
assign w29985 = ~pi02709 & w18287;
assign w29986 = ~w29984 & ~w29985;
assign w29987 = ~w16928 & w17428;
assign w29988 = pi05373 & ~w29987;
assign w29989 = ~pi09812 & w29987;
assign w29990 = ~w29988 & ~w29989;
assign w29991 = pi05374 & ~w18142;
assign w29992 = w17177 & w18578;
assign w29993 = ~w29991 & ~w29992;
assign w29994 = pi05375 & ~w18142;
assign w29995 = ~pi02706 & w18142;
assign w29996 = ~w29994 & ~w29995;
assign w29997 = pi05376 & ~w18142;
assign w29998 = ~pi02707 & w18142;
assign w29999 = ~w29997 & ~w29998;
assign w30000 = pi05377 & ~w18142;
assign w30001 = ~pi02160 & w18142;
assign w30002 = ~w30000 & ~w30001;
assign w30003 = pi05378 & ~w18142;
assign w30004 = ~pi02723 & w18142;
assign w30005 = ~w30003 & ~w30004;
assign w30006 = pi05379 & ~w18142;
assign w30007 = ~pi02708 & w18142;
assign w30008 = ~w30006 & ~w30007;
assign w30009 = pi05380 & ~w18142;
assign w30010 = ~pi02709 & w18142;
assign w30011 = ~w30009 & ~w30010;
assign w30012 = pi05381 & ~w18178;
assign w30013 = ~pi02705 & w18178;
assign w30014 = ~w30012 & ~w30013;
assign w30015 = pi05382 & ~w18178;
assign w30016 = ~pi02706 & w18178;
assign w30017 = ~w30015 & ~w30016;
assign w30018 = pi05383 & ~w18178;
assign w30019 = ~pi02707 & w18178;
assign w30020 = ~w30018 & ~w30019;
assign w30021 = pi05384 & ~w18178;
assign w30022 = ~pi02723 & w18178;
assign w30023 = ~w30021 & ~w30022;
assign w30024 = pi05385 & ~w18178;
assign w30025 = w18177 & w18689;
assign w30026 = ~w30024 & ~w30025;
assign w30027 = pi05386 & ~w18178;
assign w30028 = w18092 & w18177;
assign w30029 = ~w30027 & ~w30028;
assign w30030 = pi05387 & ~w18112;
assign w30031 = ~pi02705 & w18112;
assign w30032 = ~w30030 & ~w30031;
assign w30033 = pi05388 & ~w18112;
assign w30034 = w17565 & w17925;
assign w30035 = ~w30033 & ~w30034;
assign w30036 = pi05389 & ~w18112;
assign w30037 = ~pi02707 & w18112;
assign w30038 = ~w30036 & ~w30037;
assign w30039 = pi05390 & ~w18112;
assign w30040 = ~pi02160 & w18112;
assign w30041 = ~w30039 & ~w30040;
assign w30042 = pi05391 & ~w18112;
assign w30043 = ~pi02723 & w18112;
assign w30044 = ~w30042 & ~w30043;
assign w30045 = pi05392 & ~w18112;
assign w30046 = ~pi02708 & w18112;
assign w30047 = ~w30045 & ~w30046;
assign w30048 = pi05393 & ~w18112;
assign w30049 = ~pi02709 & w18112;
assign w30050 = ~w30048 & ~w30049;
assign w30051 = pi05394 & ~w18041;
assign w30052 = ~pi02705 & w18041;
assign w30053 = ~w30051 & ~w30052;
assign w30054 = pi05395 & ~w18041;
assign w30055 = w17925 & w18040;
assign w30056 = ~w30054 & ~w30055;
assign w30057 = pi05396 & ~w24403;
assign w30058 = ~pi09954 & w24403;
assign w30059 = ~w30057 & ~w30058;
assign w30060 = pi05397 & ~w18041;
assign w30061 = ~pi02160 & w18041;
assign w30062 = ~w30060 & ~w30061;
assign w30063 = pi05398 & ~w18041;
assign w30064 = w17671 & w18040;
assign w30065 = ~w30063 & ~w30064;
assign w30066 = pi05399 & ~w18041;
assign w30067 = ~pi02708 & w18041;
assign w30068 = ~w30066 & ~w30067;
assign w30069 = pi05400 & ~w18041;
assign w30070 = ~pi02710 & w18041;
assign w30071 = ~w30069 & ~w30070;
assign w30072 = pi05401 & ~w17918;
assign w30073 = ~pi02705 & w17918;
assign w30074 = ~w30072 & ~w30073;
assign w30075 = pi05402 & ~w17918;
assign w30076 = ~pi02706 & w17918;
assign w30077 = ~w30075 & ~w30076;
assign w30078 = pi05403 & ~w17918;
assign w30079 = ~pi02707 & w17918;
assign w30080 = ~w30078 & ~w30079;
assign w30081 = pi05404 & ~w17918;
assign w30082 = ~pi02160 & w17918;
assign w30083 = ~w30081 & ~w30082;
assign w30084 = pi05405 & ~w17918;
assign w30085 = w17671 & w17917;
assign w30086 = ~w30084 & ~w30085;
assign w30087 = pi05406 & ~w17918;
assign w30088 = ~pi02708 & w17918;
assign w30089 = ~w30087 & ~w30088;
assign w30090 = pi05407 & ~w17918;
assign w30091 = ~pi02710 & w17918;
assign w30092 = ~w30090 & ~w30091;
assign w30093 = pi05408 & ~w17669;
assign w30094 = ~pi02705 & w17669;
assign w30095 = ~w30093 & ~w30094;
assign w30096 = pi05409 & ~w17669;
assign w30097 = ~pi02706 & w17669;
assign w30098 = ~w30096 & ~w30097;
assign w30099 = pi05410 & ~w17669;
assign w30100 = ~pi02160 & w17669;
assign w30101 = ~w30099 & ~w30100;
assign w30102 = pi05411 & ~w17669;
assign w30103 = ~pi02708 & w17669;
assign w30104 = ~w30102 & ~w30103;
assign w30105 = pi05412 & ~w17669;
assign w30106 = ~pi02709 & w17669;
assign w30107 = ~w30105 & ~w30106;
assign w30108 = pi05413 & ~w17669;
assign w30109 = ~pi02710 & w17669;
assign w30110 = ~w30108 & ~w30109;
assign w30111 = pi05414 & ~w17637;
assign w30112 = ~pi02705 & w17637;
assign w30113 = ~w30111 & ~w30112;
assign w30114 = pi05415 & ~w17637;
assign w30115 = ~pi02706 & w17637;
assign w30116 = ~w30114 & ~w30115;
assign w30117 = pi05416 & ~w17637;
assign w30118 = ~pi02707 & w17637;
assign w30119 = ~w30117 & ~w30118;
assign w30120 = pi05417 & ~w17637;
assign w30121 = ~pi02160 & w17637;
assign w30122 = ~w30120 & ~w30121;
assign w30123 = pi05418 & ~w17637;
assign w30124 = ~pi02723 & w17637;
assign w30125 = ~w30123 & ~w30124;
assign w30126 = pi05419 & ~w17637;
assign w30127 = ~pi02708 & w17637;
assign w30128 = ~w30126 & ~w30127;
assign w30129 = pi05420 & ~w17637;
assign w30130 = ~pi02710 & w17637;
assign w30131 = ~w30129 & ~w30130;
assign w30132 = pi05421 & ~w16962;
assign w30133 = ~pi02705 & w16962;
assign w30134 = ~w30132 & ~w30133;
assign w30135 = pi05422 & ~w16962;
assign w30136 = w16961 & w17925;
assign w30137 = ~w30135 & ~w30136;
assign w30138 = pi05423 & ~w16962;
assign w30139 = w16961 & w18234;
assign w30140 = ~w30138 & ~w30139;
assign w30141 = pi05424 & ~w16962;
assign w30142 = ~pi02723 & w16962;
assign w30143 = ~w30141 & ~w30142;
assign w30144 = pi05425 & ~w16962;
assign w30145 = w16961 & w18689;
assign w30146 = ~w30144 & ~w30145;
assign w30147 = pi05426 & ~w16962;
assign w30148 = ~pi02710 & w16962;
assign w30149 = ~w30147 & ~w30148;
assign w30150 = pi05427 & ~w20974;
assign w30151 = w17193 & w19596;
assign w30152 = ~w30150 & ~w30151;
assign w30153 = ~w16892 & w18009;
assign w30154 = pi05428 & ~w30153;
assign w30155 = ~pi02705 & w30153;
assign w30156 = ~w30154 & ~w30155;
assign w30157 = pi05429 & ~w30153;
assign w30158 = ~pi02706 & w30153;
assign w30159 = ~w30157 & ~w30158;
assign w30160 = pi05430 & ~w30153;
assign w30161 = ~pi02707 & w30153;
assign w30162 = ~w30160 & ~w30161;
assign w30163 = pi05431 & ~w21202;
assign w30164 = ~pi09812 & w21202;
assign w30165 = ~w30163 & ~w30164;
assign w30166 = pi05432 & ~w30153;
assign w30167 = ~pi02160 & w30153;
assign w30168 = ~w30166 & ~w30167;
assign w30169 = pi05433 & ~w30153;
assign w30170 = ~pi02708 & w30153;
assign w30171 = ~w30169 & ~w30170;
assign w30172 = pi05434 & ~w30153;
assign w30173 = ~pi02709 & w30153;
assign w30174 = ~w30172 & ~w30173;
assign w30175 = pi05435 & ~w30153;
assign w30176 = ~pi02710 & w30153;
assign w30177 = ~w30175 & ~w30176;
assign w30178 = ~w16892 & w17650;
assign w30179 = pi05436 & ~w30178;
assign w30180 = ~pi02705 & w30178;
assign w30181 = ~w30179 & ~w30180;
assign w30182 = pi05437 & ~w30178;
assign w30183 = ~pi02706 & w30178;
assign w30184 = ~w30182 & ~w30183;
assign w30185 = pi05438 & ~w30178;
assign w30186 = ~pi02707 & w30178;
assign w30187 = ~w30185 & ~w30186;
assign w30188 = pi05439 & ~w30178;
assign w30189 = ~pi02723 & w30178;
assign w30190 = ~w30188 & ~w30189;
assign w30191 = pi05440 & ~w30178;
assign w30192 = ~pi02708 & w30178;
assign w30193 = ~w30191 & ~w30192;
assign w30194 = pi05441 & ~w30178;
assign w30195 = ~pi02709 & w30178;
assign w30196 = ~w30194 & ~w30195;
assign w30197 = pi05442 & ~w30178;
assign w30198 = ~pi02710 & w30178;
assign w30199 = ~w30197 & ~w30198;
assign w30200 = ~w16892 & w18622;
assign w30201 = pi05443 & ~w30200;
assign w30202 = ~pi02705 & w30200;
assign w30203 = ~w30201 & ~w30202;
assign w30204 = pi05444 & ~w30200;
assign w30205 = ~pi02706 & w30200;
assign w30206 = ~w30204 & ~w30205;
assign w30207 = pi05445 & ~w30200;
assign w30208 = ~pi02707 & w30200;
assign w30209 = ~w30207 & ~w30208;
assign w30210 = pi05446 & ~w30200;
assign w30211 = ~pi02723 & w30200;
assign w30212 = ~w30210 & ~w30211;
assign w30213 = pi05447 & ~w30200;
assign w30214 = ~pi02708 & w30200;
assign w30215 = ~w30213 & ~w30214;
assign w30216 = pi05448 & ~w30200;
assign w30217 = ~pi02709 & w30200;
assign w30218 = ~w30216 & ~w30217;
assign w30219 = pi05449 & ~w21266;
assign w30220 = ~pi09961 & w21266;
assign w30221 = ~w30219 & ~w30220;
assign w30222 = ~w16892 & w17190;
assign w30223 = pi05450 & ~w30222;
assign w30224 = ~pi02705 & w30222;
assign w30225 = ~w30223 & ~w30224;
assign w30226 = pi05451 & ~w30222;
assign w30227 = ~pi02706 & w30222;
assign w30228 = ~w30226 & ~w30227;
assign w30229 = pi05452 & ~w30222;
assign w30230 = ~pi02160 & w30222;
assign w30231 = ~w30229 & ~w30230;
assign w30232 = pi05453 & ~w30222;
assign w30233 = ~pi02723 & w30222;
assign w30234 = ~w30232 & ~w30233;
assign w30235 = pi05454 & ~w30222;
assign w30236 = w17190 & w18689;
assign w30237 = ~w30235 & ~w30236;
assign w30238 = pi05455 & ~w30222;
assign w30239 = ~pi02709 & w30222;
assign w30240 = ~w30238 & ~w30239;
assign w30241 = pi05456 & ~w30222;
assign w30242 = ~pi02710 & w30222;
assign w30243 = ~w30241 & ~w30242;
assign w30244 = ~w16892 & w17600;
assign w30245 = pi05457 & ~w30244;
assign w30246 = ~pi02705 & w30244;
assign w30247 = ~w30245 & ~w30246;
assign w30248 = pi05458 & ~w30244;
assign w30249 = ~pi02706 & w30244;
assign w30250 = ~w30248 & ~w30249;
assign w30251 = pi05459 & ~w30244;
assign w30252 = ~pi02160 & w30244;
assign w30253 = ~w30251 & ~w30252;
assign w30254 = pi05460 & ~w30244;
assign w30255 = w17600 & w17671;
assign w30256 = ~w30254 & ~w30255;
assign w30257 = pi05461 & ~w30244;
assign w30258 = ~pi02708 & w30244;
assign w30259 = ~w30257 & ~w30258;
assign w30260 = pi05462 & ~w30244;
assign w30261 = w17600 & w18364;
assign w30262 = ~w30260 & ~w30261;
assign w30263 = ~w16892 & w17375;
assign w30264 = pi05463 & ~w30263;
assign w30265 = ~pi02705 & w30263;
assign w30266 = ~w30264 & ~w30265;
assign w30267 = pi05464 & ~w30263;
assign w30268 = ~pi02706 & w30263;
assign w30269 = ~w30267 & ~w30268;
assign w30270 = pi05465 & ~w30263;
assign w30271 = ~pi02160 & w30263;
assign w30272 = ~w30270 & ~w30271;
assign w30273 = pi05466 & ~w30263;
assign w30274 = ~pi02723 & w30263;
assign w30275 = ~w30273 & ~w30274;
assign w30276 = pi05467 & ~w30263;
assign w30277 = ~pi02708 & w30263;
assign w30278 = ~w30276 & ~w30277;
assign w30279 = pi05468 & ~w30263;
assign w30280 = ~pi02709 & w30263;
assign w30281 = ~w30279 & ~w30280;
assign w30282 = pi05469 & ~w30263;
assign w30283 = ~pi02710 & w30263;
assign w30284 = ~w30282 & ~w30283;
assign w30285 = ~w16892 & w18731;
assign w30286 = pi05470 & ~w30285;
assign w30287 = ~pi02705 & w30285;
assign w30288 = ~w30286 & ~w30287;
assign w30289 = pi05471 & ~w30285;
assign w30290 = ~pi02706 & w30285;
assign w30291 = ~w30289 & ~w30290;
assign w30292 = pi05472 & ~w18727;
assign w30293 = ~pi02704 & w18727;
assign w30294 = ~w30292 & ~w30293;
assign w30295 = pi05473 & ~w30285;
assign w30296 = ~pi02160 & w30285;
assign w30297 = ~w30295 & ~w30296;
assign w30298 = pi05474 & ~w30285;
assign w30299 = ~pi02723 & w30285;
assign w30300 = ~w30298 & ~w30299;
assign w30301 = pi05475 & ~w30285;
assign w30302 = ~pi02709 & w30285;
assign w30303 = ~w30301 & ~w30302;
assign w30304 = pi05476 & ~w30285;
assign w30305 = ~pi02710 & w30285;
assign w30306 = ~w30304 & ~w30305;
assign w30307 = ~w16892 & w18683;
assign w30308 = pi05477 & ~w30307;
assign w30309 = ~pi02705 & w30307;
assign w30310 = ~w30308 & ~w30309;
assign w30311 = pi05478 & ~w30307;
assign w30312 = ~pi02707 & w30307;
assign w30313 = ~w30311 & ~w30312;
assign w30314 = pi05479 & ~w30307;
assign w30315 = ~pi02160 & w30307;
assign w30316 = ~w30314 & ~w30315;
assign w30317 = pi05480 & ~w30307;
assign w30318 = ~pi02723 & w30307;
assign w30319 = ~w30317 & ~w30318;
assign w30320 = pi05481 & ~w30307;
assign w30321 = ~pi02708 & w30307;
assign w30322 = ~w30320 & ~w30321;
assign w30323 = pi05482 & ~w30307;
assign w30324 = ~pi02709 & w30307;
assign w30325 = ~w30323 & ~w30324;
assign w30326 = pi05483 & ~w30307;
assign w30327 = ~pi02710 & w30307;
assign w30328 = ~w30326 & ~w30327;
assign w30329 = ~w16892 & w18348;
assign w30330 = pi05484 & ~w30329;
assign w30331 = ~pi02705 & w30329;
assign w30332 = ~w30330 & ~w30331;
assign w30333 = pi05485 & ~w30329;
assign w30334 = ~pi02707 & w30329;
assign w30335 = ~w30333 & ~w30334;
assign w30336 = pi05486 & ~w30329;
assign w30337 = ~pi02160 & w30329;
assign w30338 = ~w30336 & ~w30337;
assign w30339 = pi05487 & ~w30329;
assign w30340 = ~pi02723 & w30329;
assign w30341 = ~w30339 & ~w30340;
assign w30342 = pi05488 & ~w30329;
assign w30343 = ~pi02709 & w30329;
assign w30344 = ~w30342 & ~w30343;
assign w30345 = pi05489 & ~w30329;
assign w30346 = ~pi02710 & w30329;
assign w30347 = ~w30345 & ~w30346;
assign w30348 = ~w16892 & w17521;
assign w30349 = pi05490 & ~w30348;
assign w30350 = ~pi02705 & w30348;
assign w30351 = ~w30349 & ~w30350;
assign w30352 = pi05491 & ~w30348;
assign w30353 = ~pi02707 & w30348;
assign w30354 = ~w30352 & ~w30353;
assign w30355 = pi05492 & ~w30348;
assign w30356 = ~pi02160 & w30348;
assign w30357 = ~w30355 & ~w30356;
assign w30358 = pi05493 & ~w30348;
assign w30359 = ~pi02723 & w30348;
assign w30360 = ~w30358 & ~w30359;
assign w30361 = pi05494 & ~w30348;
assign w30362 = ~pi02708 & w30348;
assign w30363 = ~w30361 & ~w30362;
assign w30364 = pi05495 & ~w30348;
assign w30365 = ~pi02709 & w30348;
assign w30366 = ~w30364 & ~w30365;
assign w30367 = pi05496 & ~w30348;
assign w30368 = ~pi02710 & w30348;
assign w30369 = ~w30367 & ~w30368;
assign w30370 = ~w16892 & w17325;
assign w30371 = pi05497 & ~w30370;
assign w30372 = w17325 & w18578;
assign w30373 = ~w30371 & ~w30372;
assign w30374 = pi05498 & ~w30370;
assign w30375 = ~pi02707 & w30370;
assign w30376 = ~w30374 & ~w30375;
assign w30377 = pi05499 & ~w30370;
assign w30378 = w17325 & w18234;
assign w30379 = ~w30377 & ~w30378;
assign w30380 = pi05500 & ~w30370;
assign w30381 = w17325 & w17671;
assign w30382 = ~w30380 & ~w30381;
assign w30383 = pi05501 & ~w30370;
assign w30384 = ~pi02709 & w30370;
assign w30385 = ~w30383 & ~w30384;
assign w30386 = pi05502 & ~w30370;
assign w30387 = w17325 & w18364;
assign w30388 = ~w30386 & ~w30387;
assign w30389 = ~w16892 & w17474;
assign w30390 = pi05503 & ~w30389;
assign w30391 = ~pi02705 & w30389;
assign w30392 = ~w30390 & ~w30391;
assign w30393 = pi05504 & ~w30389;
assign w30394 = ~pi02707 & w30389;
assign w30395 = ~w30393 & ~w30394;
assign w30396 = pi05505 & ~w30389;
assign w30397 = w17474 & w18234;
assign w30398 = ~w30396 & ~w30397;
assign w30399 = pi05506 & ~w30389;
assign w30400 = ~pi02723 & w30389;
assign w30401 = ~w30399 & ~w30400;
assign w30402 = pi05507 & ~w30389;
assign w30403 = ~pi02708 & w30389;
assign w30404 = ~w30402 & ~w30403;
assign w30405 = pi05508 & ~w30389;
assign w30406 = ~pi02709 & w30389;
assign w30407 = ~w30405 & ~w30406;
assign w30408 = pi05509 & ~w30389;
assign w30409 = ~pi02710 & w30389;
assign w30410 = ~w30408 & ~w30409;
assign w30411 = ~w16892 & w17320;
assign w30412 = pi05510 & ~w30411;
assign w30413 = ~pi02705 & w30411;
assign w30414 = ~w30412 & ~w30413;
assign w30415 = pi05511 & ~w30411;
assign w30416 = ~pi02707 & w30411;
assign w30417 = ~w30415 & ~w30416;
assign w30418 = pi05512 & ~w30411;
assign w30419 = ~pi02160 & w30411;
assign w30420 = ~w30418 & ~w30419;
assign w30421 = pi05513 & ~w30411;
assign w30422 = ~pi02723 & w30411;
assign w30423 = ~w30421 & ~w30422;
assign w30424 = pi05514 & ~w30411;
assign w30425 = ~pi02709 & w30411;
assign w30426 = ~w30424 & ~w30425;
assign w30427 = pi05515 & ~w30411;
assign w30428 = ~pi02710 & w30411;
assign w30429 = ~w30427 & ~w30428;
assign w30430 = ~w16892 & w17344;
assign w30431 = pi05516 & ~w30430;
assign w30432 = ~pi02705 & w30430;
assign w30433 = ~w30431 & ~w30432;
assign w30434 = pi05517 & ~w30430;
assign w30435 = w17344 & w18067;
assign w30436 = ~w30434 & ~w30435;
assign w30437 = pi05518 & ~w30430;
assign w30438 = ~pi02160 & w30430;
assign w30439 = ~w30437 & ~w30438;
assign w30440 = pi05519 & ~w30430;
assign w30441 = ~pi02723 & w30430;
assign w30442 = ~w30440 & ~w30441;
assign w30443 = pi05520 & ~w30430;
assign w30444 = ~pi02708 & w30430;
assign w30445 = ~w30443 & ~w30444;
assign w30446 = pi05521 & ~w30430;
assign w30447 = ~pi02709 & w30430;
assign w30448 = ~w30446 & ~w30447;
assign w30449 = pi05522 & ~w30430;
assign w30450 = ~pi02710 & w30430;
assign w30451 = ~w30449 & ~w30450;
assign w30452 = ~w16892 & w17162;
assign w30453 = pi05523 & ~w30452;
assign w30454 = ~pi02705 & w30452;
assign w30455 = ~w30453 & ~w30454;
assign w30456 = pi05524 & ~w30452;
assign w30457 = ~pi02707 & w30452;
assign w30458 = ~w30456 & ~w30457;
assign w30459 = pi05525 & ~w30452;
assign w30460 = ~pi02160 & w30452;
assign w30461 = ~w30459 & ~w30460;
assign w30462 = pi05526 & ~w30452;
assign w30463 = ~pi02723 & w30452;
assign w30464 = ~w30462 & ~w30463;
assign w30465 = pi05527 & ~w30452;
assign w30466 = ~pi02709 & w30452;
assign w30467 = ~w30465 & ~w30466;
assign w30468 = pi05528 & ~w30452;
assign w30469 = ~pi02710 & w30452;
assign w30470 = ~w30468 & ~w30469;
assign w30471 = ~w16892 & w17244;
assign w30472 = pi05529 & ~w30471;
assign w30473 = ~pi02705 & w30471;
assign w30474 = ~w30472 & ~w30473;
assign w30475 = pi05530 & ~w30471;
assign w30476 = ~pi02707 & w30471;
assign w30477 = ~w30475 & ~w30476;
assign w30478 = pi05531 & ~w30471;
assign w30479 = ~pi02160 & w30471;
assign w30480 = ~w30478 & ~w30479;
assign w30481 = pi05532 & ~w30471;
assign w30482 = ~pi02723 & w30471;
assign w30483 = ~w30481 & ~w30482;
assign w30484 = pi05533 & ~w30471;
assign w30485 = ~pi02708 & w30471;
assign w30486 = ~w30484 & ~w30485;
assign w30487 = pi05534 & ~w30471;
assign w30488 = ~pi02709 & w30471;
assign w30489 = ~w30487 & ~w30488;
assign w30490 = pi05535 & ~w30471;
assign w30491 = ~pi02710 & w30471;
assign w30492 = ~w30490 & ~w30491;
assign w30493 = ~w16892 & w19306;
assign w30494 = pi05536 & ~w30493;
assign w30495 = ~pi02705 & w30493;
assign w30496 = ~w30494 & ~w30495;
assign w30497 = pi05537 & ~w30493;
assign w30498 = w18067 & w19306;
assign w30499 = ~w30497 & ~w30498;
assign w30500 = pi05538 & ~w30493;
assign w30501 = w18234 & w19306;
assign w30502 = ~w30500 & ~w30501;
assign w30503 = pi05539 & ~w30493;
assign w30504 = w17671 & w19306;
assign w30505 = ~w30503 & ~w30504;
assign w30506 = pi05540 & ~w30493;
assign w30507 = w18092 & w19306;
assign w30508 = ~w30506 & ~w30507;
assign w30509 = pi05541 & ~w30493;
assign w30510 = w18364 & w19306;
assign w30511 = ~w30509 & ~w30510;
assign w30512 = ~w16892 & w18217;
assign w30513 = pi05542 & ~w30512;
assign w30514 = ~pi02705 & w30512;
assign w30515 = ~w30513 & ~w30514;
assign w30516 = pi05543 & ~w30512;
assign w30517 = ~pi02707 & w30512;
assign w30518 = ~w30516 & ~w30517;
assign w30519 = pi05544 & ~w30512;
assign w30520 = ~pi02160 & w30512;
assign w30521 = ~w30519 & ~w30520;
assign w30522 = pi05545 & ~w30512;
assign w30523 = w17671 & w18217;
assign w30524 = ~w30522 & ~w30523;
assign w30525 = pi05546 & ~w30512;
assign w30526 = ~pi02708 & w30512;
assign w30527 = ~w30525 & ~w30526;
assign w30528 = pi05547 & ~w30512;
assign w30529 = ~pi02709 & w30512;
assign w30530 = ~w30528 & ~w30529;
assign w30531 = pi05548 & ~w30512;
assign w30532 = w18217 & w18364;
assign w30533 = ~w30531 & ~w30532;
assign w30534 = ~w16892 & w17739;
assign w30535 = pi05549 & ~w30534;
assign w30536 = w17739 & w18578;
assign w30537 = ~w30535 & ~w30536;
assign w30538 = pi05550 & ~w30534;
assign w30539 = ~pi02707 & w30534;
assign w30540 = ~w30538 & ~w30539;
assign w30541 = pi05551 & ~w30534;
assign w30542 = ~pi02160 & w30534;
assign w30543 = ~w30541 & ~w30542;
assign w30544 = pi05552 & ~w30534;
assign w30545 = ~pi02723 & w30534;
assign w30546 = ~w30544 & ~w30545;
assign w30547 = pi05553 & ~w30534;
assign w30548 = ~pi02709 & w30534;
assign w30549 = ~w30547 & ~w30548;
assign w30550 = pi05554 & ~w30534;
assign w30551 = ~pi02710 & w30534;
assign w30552 = ~w30550 & ~w30551;
assign w30553 = ~w16892 & w16986;
assign w30554 = pi05555 & ~w30553;
assign w30555 = ~pi02705 & w30553;
assign w30556 = ~w30554 & ~w30555;
assign w30557 = pi05556 & ~w30553;
assign w30558 = ~pi02707 & w30553;
assign w30559 = ~w30557 & ~w30558;
assign w30560 = pi05557 & ~w30553;
assign w30561 = ~pi02160 & w30553;
assign w30562 = ~w30560 & ~w30561;
assign w30563 = pi05558 & ~w30553;
assign w30564 = ~pi02723 & w30553;
assign w30565 = ~w30563 & ~w30564;
assign w30566 = pi05559 & ~w30553;
assign w30567 = ~pi02708 & w30553;
assign w30568 = ~w30566 & ~w30567;
assign w30569 = pi05560 & ~w30553;
assign w30570 = ~pi02709 & w30553;
assign w30571 = ~w30569 & ~w30570;
assign w30572 = pi05561 & ~w30553;
assign w30573 = ~pi02710 & w30553;
assign w30574 = ~w30572 & ~w30573;
assign w30575 = ~w16892 & w17694;
assign w30576 = pi05562 & ~w30575;
assign w30577 = ~pi02705 & w30575;
assign w30578 = ~w30576 & ~w30577;
assign w30579 = pi05563 & ~w30575;
assign w30580 = ~pi02707 & w30575;
assign w30581 = ~w30579 & ~w30580;
assign w30582 = pi05564 & ~w30575;
assign w30583 = ~pi02160 & w30575;
assign w30584 = ~w30582 & ~w30583;
assign w30585 = pi05565 & ~w30575;
assign w30586 = ~pi02723 & w30575;
assign w30587 = ~w30585 & ~w30586;
assign w30588 = pi05566 & ~w30575;
assign w30589 = ~pi02709 & w30575;
assign w30590 = ~w30588 & ~w30589;
assign w30591 = pi05567 & ~w30575;
assign w30592 = ~pi02710 & w30575;
assign w30593 = ~w30591 & ~w30592;
assign w30594 = ~w16892 & w20923;
assign w30595 = pi05568 & ~w30594;
assign w30596 = ~pi02705 & w30594;
assign w30597 = ~w30595 & ~w30596;
assign w30598 = pi05569 & ~w30594;
assign w30599 = w18067 & w20923;
assign w30600 = ~w30598 & ~w30599;
assign w30601 = pi05570 & ~w30594;
assign w30602 = ~pi02160 & w30594;
assign w30603 = ~w30601 & ~w30602;
assign w30604 = pi05571 & ~w30594;
assign w30605 = ~pi02723 & w30594;
assign w30606 = ~w30604 & ~w30605;
assign w30607 = pi05572 & ~w30594;
assign w30608 = ~pi02708 & w30594;
assign w30609 = ~w30607 & ~w30608;
assign w30610 = pi05573 & ~w30594;
assign w30611 = ~pi02709 & w30594;
assign w30612 = ~w30610 & ~w30611;
assign w30613 = pi05574 & ~w30594;
assign w30614 = ~pi02710 & w30594;
assign w30615 = ~w30613 & ~w30614;
assign w30616 = ~w16892 & w17148;
assign w30617 = pi05575 & ~w30616;
assign w30618 = ~pi02705 & w30616;
assign w30619 = ~w30617 & ~w30618;
assign w30620 = pi05576 & ~w30616;
assign w30621 = ~pi02707 & w30616;
assign w30622 = ~w30620 & ~w30621;
assign w30623 = pi05577 & ~w30616;
assign w30624 = ~pi02160 & w30616;
assign w30625 = ~w30623 & ~w30624;
assign w30626 = pi05578 & ~w30616;
assign w30627 = ~pi02723 & w30616;
assign w30628 = ~w30626 & ~w30627;
assign w30629 = pi05579 & ~w30616;
assign w30630 = ~pi02709 & w30616;
assign w30631 = ~w30629 & ~w30630;
assign w30632 = pi05580 & ~w30616;
assign w30633 = w17148 & w18364;
assign w30634 = ~w30632 & ~w30633;
assign w30635 = ~w16892 & w18563;
assign w30636 = pi05581 & ~w30635;
assign w30637 = ~pi02705 & w30635;
assign w30638 = ~w30636 & ~w30637;
assign w30639 = pi05582 & ~w30635;
assign w30640 = ~pi02707 & w30635;
assign w30641 = ~w30639 & ~w30640;
assign w30642 = pi05583 & ~w30635;
assign w30643 = ~pi02160 & w30635;
assign w30644 = ~w30642 & ~w30643;
assign w30645 = pi05584 & ~w30635;
assign w30646 = ~pi02723 & w30635;
assign w30647 = ~w30645 & ~w30646;
assign w30648 = pi05585 & ~w30635;
assign w30649 = ~pi02708 & w30635;
assign w30650 = ~w30648 & ~w30649;
assign w30651 = pi05586 & ~w30635;
assign w30652 = w18092 & w18563;
assign w30653 = ~w30651 & ~w30652;
assign w30654 = pi05587 & ~w30635;
assign w30655 = ~pi02710 & w30635;
assign w30656 = ~w30654 & ~w30655;
assign w30657 = pi05588 & ~w21925;
assign w30658 = ~pi02705 & w21925;
assign w30659 = ~w30657 & ~w30658;
assign w30660 = pi05589 & ~w21925;
assign w30661 = ~pi02707 & w21925;
assign w30662 = ~w30660 & ~w30661;
assign w30663 = pi05590 & ~w21925;
assign w30664 = ~pi02160 & w21925;
assign w30665 = ~w30663 & ~w30664;
assign w30666 = pi05591 & ~w21925;
assign w30667 = w17671 & w18813;
assign w30668 = ~w30666 & ~w30667;
assign w30669 = pi05592 & ~w21925;
assign w30670 = ~pi02709 & w21925;
assign w30671 = ~w30669 & ~w30670;
assign w30672 = pi05593 & ~w21925;
assign w30673 = w18364 & w18813;
assign w30674 = ~w30672 & ~w30673;
assign w30675 = pi05594 & ~w21990;
assign w30676 = w18578 & w18781;
assign w30677 = ~w30675 & ~w30676;
assign w30678 = pi05595 & ~w21990;
assign w30679 = ~pi02707 & w21990;
assign w30680 = ~w30678 & ~w30679;
assign w30681 = pi05596 & ~w21990;
assign w30682 = ~pi02160 & w21990;
assign w30683 = ~w30681 & ~w30682;
assign w30684 = pi05597 & ~w21990;
assign w30685 = w17671 & w18781;
assign w30686 = ~w30684 & ~w30685;
assign w30687 = pi05598 & ~w21990;
assign w30688 = ~pi02708 & w21990;
assign w30689 = ~w30687 & ~w30688;
assign w30690 = pi05599 & ~w21990;
assign w30691 = ~pi02709 & w21990;
assign w30692 = ~w30690 & ~w30691;
assign w30693 = pi05600 & ~w21990;
assign w30694 = ~pi02710 & w21990;
assign w30695 = ~w30693 & ~w30694;
assign w30696 = pi05601 & ~w21972;
assign w30697 = ~pi02705 & w21972;
assign w30698 = ~w30696 & ~w30697;
assign w30699 = pi05602 & ~w21972;
assign w30700 = w17505 & w18067;
assign w30701 = ~w30699 & ~w30700;
assign w30702 = pi05603 & ~w21972;
assign w30703 = ~pi02160 & w21972;
assign w30704 = ~w30702 & ~w30703;
assign w30705 = pi05604 & ~w21972;
assign w30706 = ~pi02723 & w21972;
assign w30707 = ~w30705 & ~w30706;
assign w30708 = pi05605 & ~w21972;
assign w30709 = ~pi02709 & w21972;
assign w30710 = ~w30708 & ~w30709;
assign w30711 = pi05606 & ~w21972;
assign w30712 = ~pi02710 & w21972;
assign w30713 = ~w30711 & ~w30712;
assign w30714 = pi05607 & ~w21948;
assign w30715 = ~pi02705 & w21948;
assign w30716 = ~w30714 & ~w30715;
assign w30717 = pi05608 & ~w21948;
assign w30718 = ~pi02707 & w21948;
assign w30719 = ~w30717 & ~w30718;
assign w30720 = pi05609 & ~w21948;
assign w30721 = ~pi02160 & w21948;
assign w30722 = ~w30720 & ~w30721;
assign w30723 = pi05610 & ~w21948;
assign w30724 = ~pi02723 & w21948;
assign w30725 = ~w30723 & ~w30724;
assign w30726 = pi05611 & ~w21948;
assign w30727 = ~pi02708 & w21948;
assign w30728 = ~w30726 & ~w30727;
assign w30729 = pi05612 & ~w21948;
assign w30730 = ~pi02709 & w21948;
assign w30731 = ~w30729 & ~w30730;
assign w30732 = pi05613 & ~w21948;
assign w30733 = w18364 & w18449;
assign w30734 = ~w30732 & ~w30733;
assign w30735 = pi05614 & ~w21921;
assign w30736 = ~pi02705 & w21921;
assign w30737 = ~w30735 & ~w30736;
assign w30738 = pi05615 & ~w21921;
assign w30739 = ~pi02707 & w21921;
assign w30740 = ~w30738 & ~w30739;
assign w30741 = pi05616 & ~w21921;
assign w30742 = ~pi02160 & w21921;
assign w30743 = ~w30741 & ~w30742;
assign w30744 = pi05617 & ~w21921;
assign w30745 = ~pi02723 & w21921;
assign w30746 = ~w30744 & ~w30745;
assign w30747 = pi05618 & ~w21921;
assign w30748 = ~pi02709 & w21921;
assign w30749 = ~w30747 & ~w30748;
assign w30750 = pi05619 & ~w21921;
assign w30751 = ~pi02710 & w21921;
assign w30752 = ~w30750 & ~w30751;
assign w30753 = pi05620 & ~w21937;
assign w30754 = ~pi02705 & w21937;
assign w30755 = ~w30753 & ~w30754;
assign w30756 = pi05621 & ~w21937;
assign w30757 = ~pi02707 & w21937;
assign w30758 = ~w30756 & ~w30757;
assign w30759 = pi05622 & ~w21937;
assign w30760 = ~pi02160 & w21937;
assign w30761 = ~w30759 & ~w30760;
assign w30762 = pi05623 & ~w21937;
assign w30763 = ~pi02723 & w21937;
assign w30764 = ~w30762 & ~w30763;
assign w30765 = pi05624 & ~w21937;
assign w30766 = ~pi02708 & w21937;
assign w30767 = ~w30765 & ~w30766;
assign w30768 = pi05625 & ~w21937;
assign w30769 = ~pi02709 & w21937;
assign w30770 = ~w30768 & ~w30769;
assign w30771 = pi05626 & ~w21937;
assign w30772 = ~pi02710 & w21937;
assign w30773 = ~w30771 & ~w30772;
assign w30774 = pi05627 & ~w17340;
assign w30775 = ~pi02705 & w17340;
assign w30776 = ~w30774 & ~w30775;
assign w30777 = pi05628 & ~w17340;
assign w30778 = w17339 & w18067;
assign w30779 = ~w30777 & ~w30778;
assign w30780 = pi05629 & ~w17340;
assign w30781 = ~pi02160 & w17340;
assign w30782 = ~w30780 & ~w30781;
assign w30783 = pi05630 & ~w17340;
assign w30784 = w17339 & w17671;
assign w30785 = ~w30783 & ~w30784;
assign w30786 = pi05631 & ~w17340;
assign w30787 = ~pi02709 & w17340;
assign w30788 = ~w30786 & ~w30787;
assign w30789 = pi05632 & ~w17340;
assign w30790 = ~pi02710 & w17340;
assign w30791 = ~w30789 & ~w30790;
assign w30792 = pi05633 & ~w21477;
assign w30793 = w17300 & w18578;
assign w30794 = ~w30792 & ~w30793;
assign w30795 = pi05634 & ~w21477;
assign w30796 = ~pi02707 & w21477;
assign w30797 = ~w30795 & ~w30796;
assign w30798 = pi05635 & ~w21477;
assign w30799 = ~pi02160 & w21477;
assign w30800 = ~w30798 & ~w30799;
assign w30801 = pi05636 & ~w21477;
assign w30802 = ~pi02723 & w21477;
assign w30803 = ~w30801 & ~w30802;
assign w30804 = pi05637 & ~w21477;
assign w30805 = ~pi02708 & w21477;
assign w30806 = ~w30804 & ~w30805;
assign w30807 = pi05638 & ~w21477;
assign w30808 = ~pi02709 & w21477;
assign w30809 = ~w30807 & ~w30808;
assign w30810 = pi05639 & ~w21477;
assign w30811 = ~pi02710 & w21477;
assign w30812 = ~w30810 & ~w30811;
assign w30813 = pi05640 & ~w21056;
assign w30814 = ~pi02705 & w21056;
assign w30815 = ~w30813 & ~w30814;
assign w30816 = pi05641 & ~w21056;
assign w30817 = ~pi02707 & w21056;
assign w30818 = ~w30816 & ~w30817;
assign w30819 = pi05642 & ~w21056;
assign w30820 = ~pi02160 & w21056;
assign w30821 = ~w30819 & ~w30820;
assign w30822 = pi05643 & ~w21056;
assign w30823 = ~pi02723 & w21056;
assign w30824 = ~w30822 & ~w30823;
assign w30825 = pi05644 & ~w21056;
assign w30826 = ~pi02709 & w21056;
assign w30827 = ~w30825 & ~w30826;
assign w30828 = pi05645 & ~w21056;
assign w30829 = ~pi02710 & w21056;
assign w30830 = ~w30828 & ~w30829;
assign w30831 = pi05646 & ~w21011;
assign w30832 = ~pi02705 & w21011;
assign w30833 = ~w30831 & ~w30832;
assign w30834 = pi05647 & ~w21011;
assign w30835 = ~pi02707 & w21011;
assign w30836 = ~w30834 & ~w30835;
assign w30837 = pi05648 & ~w21011;
assign w30838 = ~pi02160 & w21011;
assign w30839 = ~w30837 & ~w30838;
assign w30840 = pi05649 & ~w21011;
assign w30841 = ~pi02723 & w21011;
assign w30842 = ~w30840 & ~w30841;
assign w30843 = pi05650 & ~w21011;
assign w30844 = ~pi02708 & w21011;
assign w30845 = ~w30843 & ~w30844;
assign w30846 = pi05651 & ~w21011;
assign w30847 = w17264 & w18092;
assign w30848 = ~w30846 & ~w30847;
assign w30849 = pi05652 & ~w21011;
assign w30850 = ~pi02710 & w21011;
assign w30851 = ~w30849 & ~w30850;
assign w30852 = pi05653 & ~w20731;
assign w30853 = ~pi02705 & w20731;
assign w30854 = ~w30852 & ~w30853;
assign w30855 = pi05654 & ~w20731;
assign w30856 = ~pi02707 & w20731;
assign w30857 = ~w30855 & ~w30856;
assign w30858 = pi05655 & ~w20731;
assign w30859 = ~pi02160 & w20731;
assign w30860 = ~w30858 & ~w30859;
assign w30861 = pi05656 & ~w20731;
assign w30862 = ~pi02723 & w20731;
assign w30863 = ~w30861 & ~w30862;
assign w30864 = pi05657 & ~w20731;
assign w30865 = ~pi02709 & w20731;
assign w30866 = ~w30864 & ~w30865;
assign w30867 = pi05658 & ~w20731;
assign w30868 = ~pi02710 & w20731;
assign w30869 = ~w30867 & ~w30868;
assign w30870 = pi05659 & ~w20664;
assign w30871 = w17681 & w18578;
assign w30872 = ~w30870 & ~w30871;
assign w30873 = pi05660 & ~w20664;
assign w30874 = ~pi02707 & w20664;
assign w30875 = ~w30873 & ~w30874;
assign w30876 = pi05661 & ~w20664;
assign w30877 = w17681 & w18234;
assign w30878 = ~w30876 & ~w30877;
assign w30879 = pi05662 & ~w20664;
assign w30880 = ~pi02723 & w20664;
assign w30881 = ~w30879 & ~w30880;
assign w30882 = pi05663 & ~w20664;
assign w30883 = ~pi02708 & w20664;
assign w30884 = ~w30882 & ~w30883;
assign w30885 = pi05664 & ~w20664;
assign w30886 = ~pi02709 & w20664;
assign w30887 = ~w30885 & ~w30886;
assign w30888 = pi05665 & ~w20664;
assign w30889 = ~pi02710 & w20664;
assign w30890 = ~w30888 & ~w30889;
assign w30891 = pi05666 & ~w20647;
assign w30892 = ~pi02705 & w20647;
assign w30893 = ~w30891 & ~w30892;
assign w30894 = pi05667 & ~w20647;
assign w30895 = ~pi02707 & w20647;
assign w30896 = ~w30894 & ~w30895;
assign w30897 = ~w16992 & w19379;
assign w30898 = pi05668 & ~w30897;
assign w30899 = ~pi02703 & w30897;
assign w30900 = ~w30898 & ~w30899;
assign w30901 = pi05669 & ~w20647;
assign w30902 = ~pi02160 & w20647;
assign w30903 = ~w30901 & ~w30902;
assign w30904 = pi05670 & ~w30897;
assign w30905 = w17811 & w19379;
assign w30906 = ~w30904 & ~w30905;
assign w30907 = pi05671 & ~w20647;
assign w30908 = ~pi02708 & w20647;
assign w30909 = ~w30907 & ~w30908;
assign w30910 = pi05672 & ~w20647;
assign w30911 = ~pi02709 & w20647;
assign w30912 = ~w30910 & ~w30911;
assign w30913 = pi05673 & ~w30897;
assign w30914 = w19379 & w19797;
assign w30915 = ~w30913 & ~w30914;
assign w30916 = pi05674 & ~w20519;
assign w30917 = ~pi02705 & w20519;
assign w30918 = ~w30916 & ~w30917;
assign w30919 = pi05675 & ~w20519;
assign w30920 = ~pi02706 & w20519;
assign w30921 = ~w30919 & ~w30920;
assign w30922 = pi05676 & ~w30897;
assign w30923 = ~pi02718 & w30897;
assign w30924 = ~w30922 & ~w30923;
assign w30925 = pi05677 & ~w20519;
assign w30926 = ~pi02707 & w20519;
assign w30927 = ~w30925 & ~w30926;
assign w30928 = pi05678 & ~w20519;
assign w30929 = ~pi02160 & w20519;
assign w30930 = ~w30928 & ~w30929;
assign w30931 = pi05679 & ~w30897;
assign w30932 = ~pi02167 & w30897;
assign w30933 = ~w30931 & ~w30932;
assign w30934 = pi05680 & ~w20519;
assign w30935 = ~pi02708 & w20519;
assign w30936 = ~w30934 & ~w30935;
assign w30937 = pi05681 & ~w20519;
assign w30938 = ~pi02709 & w20519;
assign w30939 = ~w30937 & ~w30938;
assign w30940 = pi05682 & ~w30897;
assign w30941 = ~pi02164 & w30897;
assign w30942 = ~w30940 & ~w30941;
assign w30943 = pi05683 & ~w20562;
assign w30944 = w18578 & w20561;
assign w30945 = ~w30943 & ~w30944;
assign w30946 = pi05684 & ~w30897;
assign w30947 = ~pi02722 & w30897;
assign w30948 = ~w30946 & ~w30947;
assign w30949 = pi05685 & ~w20562;
assign w30950 = ~pi02706 & w20562;
assign w30951 = ~w30949 & ~w30950;
assign w30952 = pi05686 & ~w30897;
assign w30953 = ~pi02719 & w30897;
assign w30954 = ~w30952 & ~w30953;
assign w30955 = pi05687 & ~w20562;
assign w30956 = ~pi02160 & w20562;
assign w30957 = ~w30955 & ~w30956;
assign w30958 = pi05688 & ~w20562;
assign w30959 = w17671 & w20561;
assign w30960 = ~w30958 & ~w30959;
assign w30961 = pi05689 & ~w20562;
assign w30962 = ~pi02708 & w20562;
assign w30963 = ~w30961 & ~w30962;
assign w30964 = pi05690 & ~w20562;
assign w30965 = ~pi02709 & w20562;
assign w30966 = ~w30964 & ~w30965;
assign w30967 = pi05691 & ~w20485;
assign w30968 = ~pi02703 & w20485;
assign w30969 = ~w30967 & ~w30968;
assign w30970 = pi05692 & ~w20562;
assign w30971 = ~pi02710 & w20562;
assign w30972 = ~w30970 & ~w30971;
assign w30973 = pi05693 & ~w20485;
assign w30974 = ~pi02169 & w20485;
assign w30975 = ~w30973 & ~w30974;
assign w30976 = pi05694 & ~w20485;
assign w30977 = ~pi02718 & w20485;
assign w30978 = ~w30976 & ~w30977;
assign w30979 = pi05695 & ~w20485;
assign w30980 = ~pi02167 & w20485;
assign w30981 = ~w30979 & ~w30980;
assign w30982 = pi05696 & ~w20485;
assign w30983 = ~pi02164 & w20485;
assign w30984 = ~w30982 & ~w30983;
assign w30985 = pi05697 & ~w20485;
assign w30986 = ~pi02719 & w20485;
assign w30987 = ~w30985 & ~w30986;
assign w30988 = pi05698 & ~w20471;
assign w30989 = w18578 & w20470;
assign w30990 = ~w30988 & ~w30989;
assign w30991 = pi05699 & ~w20471;
assign w30992 = ~pi02707 & w20471;
assign w30993 = ~w30991 & ~w30992;
assign w30994 = pi05700 & ~w20471;
assign w30995 = ~pi02160 & w20471;
assign w30996 = ~w30994 & ~w30995;
assign w30997 = pi05701 & ~w20471;
assign w30998 = ~pi02723 & w20471;
assign w30999 = ~w30997 & ~w30998;
assign w31000 = pi05702 & ~w20471;
assign w31001 = ~pi02708 & w20471;
assign w31002 = ~w31000 & ~w31001;
assign w31003 = pi05703 & ~w20471;
assign w31004 = ~pi02709 & w20471;
assign w31005 = ~w31003 & ~w31004;
assign w31006 = pi05704 & ~w20471;
assign w31007 = ~pi02710 & w20471;
assign w31008 = ~w31006 & ~w31007;
assign w31009 = pi05705 & ~w20237;
assign w31010 = ~pi02705 & w20237;
assign w31011 = ~w31009 & ~w31010;
assign w31012 = pi05706 & ~w20237;
assign w31013 = ~pi02707 & w20237;
assign w31014 = ~w31012 & ~w31013;
assign w31015 = pi05707 & ~w20237;
assign w31016 = ~pi02160 & w20237;
assign w31017 = ~w31015 & ~w31016;
assign w31018 = pi05708 & ~w20237;
assign w31019 = ~pi02723 & w20237;
assign w31020 = ~w31018 & ~w31019;
assign w31021 = pi05709 & ~w20237;
assign w31022 = w18032 & w18092;
assign w31023 = ~w31021 & ~w31022;
assign w31024 = pi05710 & ~w20237;
assign w31025 = ~pi02710 & w20237;
assign w31026 = ~w31024 & ~w31025;
assign w31027 = pi05711 & ~w20390;
assign w31028 = ~pi02705 & w20390;
assign w31029 = ~w31027 & ~w31028;
assign w31030 = ~w16928 & w17767;
assign w31031 = pi05712 & ~w31030;
assign w31032 = ~pi02720 & w31030;
assign w31033 = ~w31031 & ~w31032;
assign w31034 = pi05713 & ~w20390;
assign w31035 = ~pi02707 & w20390;
assign w31036 = ~w31034 & ~w31035;
assign w31037 = pi05714 & ~w20390;
assign w31038 = ~pi02160 & w20390;
assign w31039 = ~w31037 & ~w31038;
assign w31040 = pi05715 & ~w20390;
assign w31041 = ~pi02723 & w20390;
assign w31042 = ~w31040 & ~w31041;
assign w31043 = pi05716 & ~w20390;
assign w31044 = ~pi02708 & w20390;
assign w31045 = ~w31043 & ~w31044;
assign w31046 = pi05717 & ~w20390;
assign w31047 = ~pi02709 & w20390;
assign w31048 = ~w31046 & ~w31047;
assign w31049 = pi05718 & ~w20390;
assign w31050 = ~pi02710 & w20390;
assign w31051 = ~w31049 & ~w31050;
assign w31052 = pi05719 & ~w19974;
assign w31053 = ~pi02703 & w19974;
assign w31054 = ~w31052 & ~w31053;
assign w31055 = pi05720 & ~w19974;
assign w31056 = ~pi02169 & w19974;
assign w31057 = ~w31055 & ~w31056;
assign w31058 = pi05721 & ~w19974;
assign w31059 = ~pi02718 & w19974;
assign w31060 = ~w31058 & ~w31059;
assign w31061 = ~w16892 & w17540;
assign w31062 = pi05722 & ~w31061;
assign w31063 = ~pi02705 & w31061;
assign w31064 = ~w31062 & ~w31063;
assign w31065 = pi05723 & ~w31061;
assign w31066 = ~pi02706 & w31061;
assign w31067 = ~w31065 & ~w31066;
assign w31068 = pi05724 & ~w19974;
assign w31069 = ~pi02164 & w19974;
assign w31070 = ~w31068 & ~w31069;
assign w31071 = pi05725 & ~w31061;
assign w31072 = ~pi02707 & w31061;
assign w31073 = ~w31071 & ~w31072;
assign w31074 = pi05726 & ~w31061;
assign w31075 = ~pi02160 & w31061;
assign w31076 = ~w31074 & ~w31075;
assign w31077 = pi05727 & ~w31061;
assign w31078 = ~pi02723 & w31061;
assign w31079 = ~w31077 & ~w31078;
assign w31080 = pi05728 & ~w19974;
assign w31081 = ~pi02719 & w19974;
assign w31082 = ~w31080 & ~w31081;
assign w31083 = pi05729 & ~w31061;
assign w31084 = ~pi02708 & w31061;
assign w31085 = ~w31083 & ~w31084;
assign w31086 = pi05730 & ~w31061;
assign w31087 = ~pi02709 & w31061;
assign w31088 = ~w31086 & ~w31087;
assign w31089 = pi05731 & ~w31061;
assign w31090 = ~pi02710 & w31061;
assign w31091 = ~w31089 & ~w31090;
assign w31092 = pi05732 & ~w19039;
assign w31093 = ~pi02721 & w19039;
assign w31094 = ~w31092 & ~w31093;
assign w31095 = pi05733 & ~w19039;
assign w31096 = ~pi02169 & w19039;
assign w31097 = ~w31095 & ~w31096;
assign w31098 = pi05734 & ~w19039;
assign w31099 = w17586 & w18027;
assign w31100 = ~w31098 & ~w31099;
assign w31101 = pi05735 & ~w18982;
assign w31102 = ~pi02705 & w18982;
assign w31103 = ~w31101 & ~w31102;
assign w31104 = pi05736 & ~w19039;
assign w31105 = ~pi02164 & w19039;
assign w31106 = ~w31104 & ~w31105;
assign w31107 = pi05737 & ~w18982;
assign w31108 = ~pi02706 & w18982;
assign w31109 = ~w31107 & ~w31108;
assign w31110 = pi05738 & ~w18982;
assign w31111 = ~pi02707 & w18982;
assign w31112 = ~w31110 & ~w31111;
assign w31113 = pi05739 & ~w18982;
assign w31114 = ~pi02723 & w18982;
assign w31115 = ~w31113 & ~w31114;
assign w31116 = pi05740 & ~w19039;
assign w31117 = w18027 & w19312;
assign w31118 = ~w31116 & ~w31117;
assign w31119 = pi05741 & ~w18982;
assign w31120 = ~pi02708 & w18982;
assign w31121 = ~w31119 & ~w31120;
assign w31122 = pi05742 & ~w18982;
assign w31123 = ~pi02709 & w18982;
assign w31124 = ~w31122 & ~w31123;
assign w31125 = pi05743 & ~w18982;
assign w31126 = ~pi02710 & w18982;
assign w31127 = ~w31125 & ~w31126;
assign w31128 = pi05744 & ~w19039;
assign w31129 = ~pi02719 & w19039;
assign w31130 = ~w31128 & ~w31129;
assign w31131 = pi05745 & ~w18586;
assign w31132 = ~pi02705 & w18586;
assign w31133 = ~w31131 & ~w31132;
assign w31134 = pi05746 & ~w18586;
assign w31135 = ~pi02707 & w18586;
assign w31136 = ~w31134 & ~w31135;
assign w31137 = pi05747 & ~w18586;
assign w31138 = w18234 & w18585;
assign w31139 = ~w31137 & ~w31138;
assign w31140 = pi05748 & ~w18586;
assign w31141 = ~pi02723 & w18586;
assign w31142 = ~w31140 & ~w31141;
assign w31143 = pi05749 & ~w18586;
assign w31144 = ~pi02709 & w18586;
assign w31145 = ~w31143 & ~w31144;
assign w31146 = pi05750 & ~w18586;
assign w31147 = ~pi02710 & w18586;
assign w31148 = ~w31146 & ~w31147;
assign w31149 = pi05751 & ~w18679;
assign w31150 = ~pi02705 & w18679;
assign w31151 = ~w31149 & ~w31150;
assign w31152 = pi05752 & ~w18679;
assign w31153 = ~pi02707 & w18679;
assign w31154 = ~w31152 & ~w31153;
assign w31155 = pi05753 & ~w18679;
assign w31156 = ~pi02160 & w18679;
assign w31157 = ~w31155 & ~w31156;
assign w31158 = pi05754 & ~w18679;
assign w31159 = w17671 & w18526;
assign w31160 = ~w31158 & ~w31159;
assign w31161 = pi05755 & ~w18679;
assign w31162 = ~pi02708 & w18679;
assign w31163 = ~w31161 & ~w31162;
assign w31164 = pi05756 & ~w18679;
assign w31165 = w18092 & w18526;
assign w31166 = ~w31164 & ~w31165;
assign w31167 = pi05757 & ~w18679;
assign w31168 = ~pi02710 & w18679;
assign w31169 = ~w31167 & ~w31168;
assign w31170 = pi05758 & ~w18641;
assign w31171 = w18291 & w18578;
assign w31172 = ~w31170 & ~w31171;
assign w31173 = pi05759 & ~w18641;
assign w31174 = ~pi02707 & w18641;
assign w31175 = ~w31173 & ~w31174;
assign w31176 = pi05760 & ~w18641;
assign w31177 = ~pi02160 & w18641;
assign w31178 = ~w31176 & ~w31177;
assign w31179 = pi05761 & ~w18641;
assign w31180 = ~pi02723 & w18641;
assign w31181 = ~w31179 & ~w31180;
assign w31182 = pi05762 & ~w18641;
assign w31183 = ~pi02709 & w18641;
assign w31184 = ~w31182 & ~w31183;
assign w31185 = pi05763 & ~w18641;
assign w31186 = ~pi02710 & w18641;
assign w31187 = ~w31185 & ~w31186;
assign w31188 = pi05764 & ~w18605;
assign w31189 = w17411 & w18578;
assign w31190 = ~w31188 & ~w31189;
assign w31191 = pi05765 & ~w18605;
assign w31192 = w17411 & w18067;
assign w31193 = ~w31191 & ~w31192;
assign w31194 = pi05766 & ~w18605;
assign w31195 = w17411 & w18234;
assign w31196 = ~w31194 & ~w31195;
assign w31197 = pi05767 & ~w18605;
assign w31198 = w17411 & w17671;
assign w31199 = ~w31197 & ~w31198;
assign w31200 = pi05768 & ~w18605;
assign w31201 = w17411 & w18689;
assign w31202 = ~w31200 & ~w31201;
assign w31203 = pi05769 & ~w18605;
assign w31204 = w17411 & w18092;
assign w31205 = ~w31203 & ~w31204;
assign w31206 = pi05770 & ~w18605;
assign w31207 = w17411 & w18364;
assign w31208 = ~w31206 & ~w31207;
assign w31209 = pi05771 & ~w18547;
assign w31210 = ~pi02705 & w18547;
assign w31211 = ~w31209 & ~w31210;
assign w31212 = pi05772 & ~w17997;
assign w31213 = ~pi02703 & w17997;
assign w31214 = ~w31212 & ~w31213;
assign w31215 = pi05773 & ~w18547;
assign w31216 = ~pi02707 & w18547;
assign w31217 = ~w31215 & ~w31216;
assign w31218 = pi05774 & ~w18547;
assign w31219 = ~pi02160 & w18547;
assign w31220 = ~w31218 & ~w31219;
assign w31221 = pi05775 & ~w18547;
assign w31222 = ~pi02723 & w18547;
assign w31223 = ~w31221 & ~w31222;
assign w31224 = pi05776 & ~w18547;
assign w31225 = ~pi02708 & w18547;
assign w31226 = ~w31224 & ~w31225;
assign w31227 = pi05777 & ~w18547;
assign w31228 = w17305 & w18092;
assign w31229 = ~w31227 & ~w31228;
assign w31230 = pi05778 & ~w18547;
assign w31231 = ~pi02710 & w18547;
assign w31232 = ~w31230 & ~w31231;
assign w31233 = pi05779 & ~w18411;
assign w31234 = ~pi02705 & w18411;
assign w31235 = ~w31233 & ~w31234;
assign w31236 = pi05780 & ~w17997;
assign w31237 = ~pi02718 & w17997;
assign w31238 = ~w31236 & ~w31237;
assign w31239 = pi05781 & ~w18411;
assign w31240 = ~pi02706 & w18411;
assign w31241 = ~w31239 & ~w31240;
assign w31242 = pi05782 & ~w18411;
assign w31243 = ~pi02707 & w18411;
assign w31244 = ~w31242 & ~w31243;
assign w31245 = pi05783 & ~w17997;
assign w31246 = ~pi02167 & w17997;
assign w31247 = ~w31245 & ~w31246;
assign w31248 = pi05784 & ~w18411;
assign w31249 = ~pi02160 & w18411;
assign w31250 = ~w31248 & ~w31249;
assign w31251 = pi05785 & ~w17997;
assign w31252 = ~pi02164 & w17997;
assign w31253 = ~w31251 & ~w31252;
assign w31254 = pi05786 & ~w18411;
assign w31255 = ~pi02708 & w18411;
assign w31256 = ~w31254 & ~w31255;
assign w31257 = pi05787 & ~w18411;
assign w31258 = ~pi02709 & w18411;
assign w31259 = ~w31257 & ~w31258;
assign w31260 = pi05788 & ~w17997;
assign w31261 = ~pi02719 & w17997;
assign w31262 = ~w31260 & ~w31261;
assign w31263 = pi05789 & ~w17997;
assign w31264 = ~pi02722 & w17997;
assign w31265 = ~w31263 & ~w31264;
assign w31266 = pi05790 & ~w18393;
assign w31267 = ~pi02705 & w18393;
assign w31268 = ~w31266 & ~w31267;
assign w31269 = ~w16928 & w19306;
assign w31270 = pi05791 & ~w31269;
assign w31271 = ~pi02720 & w31269;
assign w31272 = ~w31270 & ~w31271;
assign w31273 = pi05792 & ~w18393;
assign w31274 = ~pi02707 & w18393;
assign w31275 = ~w31273 & ~w31274;
assign w31276 = pi05793 & ~w18393;
assign w31277 = w17767 & w18234;
assign w31278 = ~w31276 & ~w31277;
assign w31279 = pi05794 & ~w18182;
assign w31280 = ~pi02703 & w18182;
assign w31281 = ~w31279 & ~w31280;
assign w31282 = pi05795 & ~w18393;
assign w31283 = ~pi02723 & w18393;
assign w31284 = ~w31282 & ~w31283;
assign w31285 = pi05796 & ~w18182;
assign w31286 = ~pi02721 & w18182;
assign w31287 = ~w31285 & ~w31286;
assign w31288 = pi05797 & ~w18393;
assign w31289 = ~pi02708 & w18393;
assign w31290 = ~w31288 & ~w31289;
assign w31291 = pi05798 & ~w18393;
assign w31292 = w17767 & w18092;
assign w31293 = ~w31291 & ~w31292;
assign w31294 = pi05799 & ~w18393;
assign w31295 = ~pi02710 & w18393;
assign w31296 = ~w31294 & ~w31295;
assign w31297 = pi05800 & ~w18271;
assign w31298 = ~pi02705 & w18271;
assign w31299 = ~w31297 & ~w31298;
assign w31300 = pi05801 & ~w18182;
assign w31301 = ~pi02718 & w18182;
assign w31302 = ~w31300 & ~w31301;
assign w31303 = pi05802 & ~w18271;
assign w31304 = w17686 & w18067;
assign w31305 = ~w31303 & ~w31304;
assign w31306 = pi05803 & ~w18182;
assign w31307 = ~pi02167 & w18182;
assign w31308 = ~w31306 & ~w31307;
assign w31309 = pi05804 & ~w18271;
assign w31310 = w17686 & w18234;
assign w31311 = ~w31309 & ~w31310;
assign w31312 = pi05805 & ~w18182;
assign w31313 = ~pi02164 & w18182;
assign w31314 = ~w31312 & ~w31313;
assign w31315 = pi05806 & ~w18271;
assign w31316 = ~pi02708 & w18271;
assign w31317 = ~w31315 & ~w31316;
assign w31318 = pi05807 & ~w18271;
assign w31319 = w17686 & w18092;
assign w31320 = ~w31318 & ~w31319;
assign w31321 = pi05808 & ~w18271;
assign w31322 = ~pi02710 & w18271;
assign w31323 = ~w31321 & ~w31322;
assign w31324 = pi05809 & ~w18182;
assign w31325 = ~pi02722 & w18182;
assign w31326 = ~w31324 & ~w31325;
assign w31327 = pi05810 & ~w18243;
assign w31328 = w17614 & w18578;
assign w31329 = ~w31327 & ~w31328;
assign w31330 = pi05811 & ~w18243;
assign w31331 = ~pi02706 & w18243;
assign w31332 = ~w31330 & ~w31331;
assign w31333 = pi05812 & ~w18243;
assign w31334 = w17614 & w18067;
assign w31335 = ~w31333 & ~w31334;
assign w31336 = pi05813 & ~w18243;
assign w31337 = ~pi02160 & w18243;
assign w31338 = ~w31336 & ~w31337;
assign w31339 = pi05814 & ~w18134;
assign w31340 = ~pi02703 & w18134;
assign w31341 = ~w31339 & ~w31340;
assign w31342 = pi05815 & ~w18243;
assign w31343 = ~pi02708 & w18243;
assign w31344 = ~w31342 & ~w31343;
assign w31345 = pi05816 & ~w18243;
assign w31346 = ~pi02709 & w18243;
assign w31347 = ~w31345 & ~w31346;
assign w31348 = ~w16928 & w17996;
assign w31349 = pi05817 & ~w31348;
assign w31350 = w17193 & w17996;
assign w31351 = ~w31349 & ~w31350;
assign w31352 = pi05818 & ~w18243;
assign w31353 = ~pi02710 & w18243;
assign w31354 = ~w31352 & ~w31353;
assign w31355 = pi05819 & ~w17527;
assign w31356 = ~pi02705 & w17527;
assign w31357 = ~w31355 & ~w31356;
assign w31358 = pi05820 & ~w18134;
assign w31359 = ~pi02169 & w18134;
assign w31360 = ~w31358 & ~w31359;
assign w31361 = pi05821 & ~w17527;
assign w31362 = ~pi02706 & w17527;
assign w31363 = ~w31361 & ~w31362;
assign w31364 = pi05822 & ~w17527;
assign w31365 = ~pi02707 & w17527;
assign w31366 = ~w31364 & ~w31365;
assign w31367 = pi05823 & ~w18134;
assign w31368 = w17183 & w17586;
assign w31369 = ~w31367 & ~w31368;
assign w31370 = pi05824 & ~w17527;
assign w31371 = ~pi02160 & w17527;
assign w31372 = ~w31370 & ~w31371;
assign w31373 = pi05825 & ~w17527;
assign w31374 = w17526 & w17671;
assign w31375 = ~w31373 & ~w31374;
assign w31376 = pi05826 & ~w18134;
assign w31377 = ~pi02164 & w18134;
assign w31378 = ~w31376 & ~w31377;
assign w31379 = pi05827 & ~w17527;
assign w31380 = ~pi02708 & w17527;
assign w31381 = ~w31379 & ~w31380;
assign w31382 = pi05828 & ~w17527;
assign w31383 = w17526 & w18364;
assign w31384 = ~w31382 & ~w31383;
assign w31385 = pi05829 & ~w17923;
assign w31386 = w17922 & w18578;
assign w31387 = ~w31385 & ~w31386;
assign w31388 = pi05830 & ~w18134;
assign w31389 = ~pi02722 & w18134;
assign w31390 = ~w31388 & ~w31389;
assign w31391 = pi05831 & ~w18134;
assign w31392 = ~pi02719 & w18134;
assign w31393 = ~w31391 & ~w31392;
assign w31394 = pi05832 & ~w17923;
assign w31395 = w17922 & w18067;
assign w31396 = ~w31394 & ~w31395;
assign w31397 = pi05833 & ~w17923;
assign w31398 = w17922 & w18234;
assign w31399 = ~w31397 & ~w31398;
assign w31400 = pi05834 & ~w17726;
assign w31401 = ~pi02703 & w17726;
assign w31402 = ~w31400 & ~w31401;
assign w31403 = pi05835 & ~w17923;
assign w31404 = w17671 & w17922;
assign w31405 = ~w31403 & ~w31404;
assign w31406 = pi05836 & ~w17923;
assign w31407 = w17922 & w18689;
assign w31408 = ~w31406 & ~w31407;
assign w31409 = pi05837 & ~w17923;
assign w31410 = w17922 & w18092;
assign w31411 = ~w31409 & ~w31410;
assign w31412 = pi05838 & ~w17923;
assign w31413 = w17922 & w18364;
assign w31414 = ~w31412 & ~w31413;
assign w31415 = pi05839 & ~w17642;
assign w31416 = ~pi02705 & w17642;
assign w31417 = ~w31415 & ~w31416;
assign w31418 = pi05840 & ~w17726;
assign w31419 = ~pi02169 & w17726;
assign w31420 = ~w31418 & ~w31419;
assign w31421 = pi05841 & ~w17642;
assign w31422 = ~pi02707 & w17642;
assign w31423 = ~w31421 & ~w31422;
assign w31424 = pi05842 & ~w17726;
assign w31425 = ~pi02718 & w17726;
assign w31426 = ~w31424 & ~w31425;
assign w31427 = pi05843 & ~w17642;
assign w31428 = ~pi02160 & w17642;
assign w31429 = ~w31427 & ~w31428;
assign w31430 = pi05844 & ~w17726;
assign w31431 = ~pi02167 & w17726;
assign w31432 = ~w31430 & ~w31431;
assign w31433 = pi05845 & ~w17642;
assign w31434 = ~pi02708 & w17642;
assign w31435 = ~w31433 & ~w31434;
assign w31436 = pi05846 & ~w17642;
assign w31437 = ~pi02709 & w17642;
assign w31438 = ~w31436 & ~w31437;
assign w31439 = pi05847 & ~w17726;
assign w31440 = ~pi02164 & w17726;
assign w31441 = ~w31439 & ~w31440;
assign w31442 = pi05848 & ~w17642;
assign w31443 = w17641 & w18364;
assign w31444 = ~w31442 & ~w31443;
assign w31445 = pi05849 & ~w17726;
assign w31446 = ~pi02722 & w17726;
assign w31447 = ~w31445 & ~w31446;
assign w31448 = ~w16892 & w21154;
assign w31449 = pi05850 & ~w31448;
assign w31450 = ~pi02705 & w31448;
assign w31451 = ~w31449 & ~w31450;
assign w31452 = pi05851 & ~w17726;
assign w31453 = ~pi02719 & w17726;
assign w31454 = ~w31452 & ~w31453;
assign w31455 = pi05852 & ~w31448;
assign w31456 = ~pi02707 & w31448;
assign w31457 = ~w31455 & ~w31456;
assign w31458 = pi05853 & ~w31448;
assign w31459 = ~pi02160 & w31448;
assign w31460 = ~w31458 & ~w31459;
assign w31461 = pi05854 & ~w31448;
assign w31462 = ~pi02723 & w31448;
assign w31463 = ~w31461 & ~w31462;
assign w31464 = pi05855 & ~w31448;
assign w31465 = ~pi02708 & w31448;
assign w31466 = ~w31464 & ~w31465;
assign w31467 = pi05856 & ~w31448;
assign w31468 = ~pi02709 & w31448;
assign w31469 = ~w31467 & ~w31468;
assign w31470 = pi05857 & ~w31448;
assign w31471 = w18364 & w21154;
assign w31472 = ~w31470 & ~w31471;
assign w31473 = ~w16892 & w20720;
assign w31474 = pi05858 & ~w31473;
assign w31475 = ~pi02705 & w31473;
assign w31476 = ~w31474 & ~w31475;
assign w31477 = ~w16992 & w17349;
assign w31478 = pi05859 & ~w31477;
assign w31479 = ~pi02169 & w31477;
assign w31480 = ~w31478 & ~w31479;
assign w31481 = pi05860 & ~w31477;
assign w31482 = w17349 & w17586;
assign w31483 = ~w31481 & ~w31482;
assign w31484 = pi05861 & ~w31473;
assign w31485 = ~pi02706 & w31473;
assign w31486 = ~w31484 & ~w31485;
assign w31487 = pi05862 & ~w31473;
assign w31488 = ~pi02707 & w31473;
assign w31489 = ~w31487 & ~w31488;
assign w31490 = pi05863 & ~w31473;
assign w31491 = ~pi02160 & w31473;
assign w31492 = ~w31490 & ~w31491;
assign w31493 = pi05864 & ~w31477;
assign w31494 = w17349 & w19273;
assign w31495 = ~w31493 & ~w31494;
assign w31496 = pi05865 & ~w31473;
assign w31497 = ~pi02708 & w31473;
assign w31498 = ~w31496 & ~w31497;
assign w31499 = pi05866 & ~w31473;
assign w31500 = ~pi02709 & w31473;
assign w31501 = ~w31499 & ~w31500;
assign w31502 = pi05867 & ~w31477;
assign w31503 = ~pi02164 & w31477;
assign w31504 = ~w31502 & ~w31503;
assign w31505 = ~w16892 & w18631;
assign w31506 = pi05868 & ~w31505;
assign w31507 = ~pi02705 & w31505;
assign w31508 = ~w31506 & ~w31507;
assign w31509 = pi05869 & ~w31477;
assign w31510 = ~pi02722 & w31477;
assign w31511 = ~w31509 & ~w31510;
assign w31512 = pi05870 & ~w31477;
assign w31513 = w17349 & w17594;
assign w31514 = ~w31512 & ~w31513;
assign w31515 = pi05871 & ~w31505;
assign w31516 = ~pi02707 & w31505;
assign w31517 = ~w31515 & ~w31516;
assign w31518 = pi05872 & ~w31505;
assign w31519 = ~pi02160 & w31505;
assign w31520 = ~w31518 & ~w31519;
assign w31521 = pi05873 & ~w31505;
assign w31522 = ~pi02723 & w31505;
assign w31523 = ~w31521 & ~w31522;
assign w31524 = pi05874 & ~w31505;
assign w31525 = w18631 & w18689;
assign w31526 = ~w31524 & ~w31525;
assign w31527 = pi05875 & ~w31505;
assign w31528 = ~pi02709 & w31505;
assign w31529 = ~w31527 & ~w31528;
assign w31530 = ~w16992 & w17210;
assign w31531 = pi05876 & ~w31530;
assign w31532 = ~pi02703 & w31530;
assign w31533 = ~w31531 & ~w31532;
assign w31534 = pi05877 & ~w31530;
assign w31535 = ~pi02721 & w31530;
assign w31536 = ~w31534 & ~w31535;
assign w31537 = ~w16892 & w17334;
assign w31538 = pi05878 & ~w31537;
assign w31539 = w17334 & w18578;
assign w31540 = ~w31538 & ~w31539;
assign w31541 = pi05879 & ~w31530;
assign w31542 = ~pi02169 & w31530;
assign w31543 = ~w31541 & ~w31542;
assign w31544 = pi05880 & ~w31537;
assign w31545 = ~pi02707 & w31537;
assign w31546 = ~w31544 & ~w31545;
assign w31547 = pi05881 & ~w31530;
assign w31548 = w17210 & w17586;
assign w31549 = ~w31547 & ~w31548;
assign w31550 = pi05882 & ~w31530;
assign w31551 = w17210 & w19273;
assign w31552 = ~w31550 & ~w31551;
assign w31553 = pi05883 & ~w31537;
assign w31554 = w17334 & w17671;
assign w31555 = ~w31553 & ~w31554;
assign w31556 = pi05884 & ~w31537;
assign w31557 = ~pi02708 & w31537;
assign w31558 = ~w31556 & ~w31557;
assign w31559 = pi05885 & ~w31537;
assign w31560 = ~pi02709 & w31537;
assign w31561 = ~w31559 & ~w31560;
assign w31562 = pi05886 & ~w31537;
assign w31563 = w17334 & w18364;
assign w31564 = ~w31562 & ~w31563;
assign w31565 = pi05887 & ~w31530;
assign w31566 = ~pi02164 & w31530;
assign w31567 = ~w31565 & ~w31566;
assign w31568 = ~w16892 & w20775;
assign w31569 = pi05888 & ~w31568;
assign w31570 = ~pi02705 & w31568;
assign w31571 = ~w31569 & ~w31570;
assign w31572 = pi05889 & ~w31568;
assign w31573 = ~pi02706 & w31568;
assign w31574 = ~w31572 & ~w31573;
assign w31575 = pi05890 & ~w31568;
assign w31576 = ~pi02707 & w31568;
assign w31577 = ~w31575 & ~w31576;
assign w31578 = pi05891 & ~w31568;
assign w31579 = ~pi02160 & w31568;
assign w31580 = ~w31578 & ~w31579;
assign w31581 = pi05892 & ~w31530;
assign w31582 = ~pi02719 & w31530;
assign w31583 = ~w31581 & ~w31582;
assign w31584 = pi05893 & ~w31568;
assign w31585 = w18689 & w20775;
assign w31586 = ~w31584 & ~w31585;
assign w31587 = pi05894 & ~w31568;
assign w31588 = ~pi02709 & w31568;
assign w31589 = ~w31587 & ~w31588;
assign w31590 = pi05895 & ~w31568;
assign w31591 = ~pi02710 & w31568;
assign w31592 = ~w31590 & ~w31591;
assign w31593 = ~w16892 & w17583;
assign w31594 = pi05896 & ~w31593;
assign w31595 = ~pi02706 & w31593;
assign w31596 = ~w31594 & ~w31595;
assign w31597 = pi05897 & ~w31593;
assign w31598 = ~pi02707 & w31593;
assign w31599 = ~w31597 & ~w31598;
assign w31600 = pi05898 & ~w31593;
assign w31601 = ~pi02160 & w31593;
assign w31602 = ~w31600 & ~w31601;
assign w31603 = pi05899 & ~w31593;
assign w31604 = ~pi02723 & w31593;
assign w31605 = ~w31603 & ~w31604;
assign w31606 = pi05900 & ~w31593;
assign w31607 = ~pi02708 & w31593;
assign w31608 = ~w31606 & ~w31607;
assign w31609 = pi05901 & ~w31593;
assign w31610 = w17583 & w18092;
assign w31611 = ~w31609 & ~w31610;
assign w31612 = pi05902 & ~w31593;
assign w31613 = ~pi02710 & w31593;
assign w31614 = ~w31612 & ~w31613;
assign w31615 = ~w16892 & w20566;
assign w31616 = pi05903 & ~w31615;
assign w31617 = ~pi02706 & w31615;
assign w31618 = ~w31616 & ~w31617;
assign w31619 = pi05904 & ~w31615;
assign w31620 = ~pi02707 & w31615;
assign w31621 = ~w31619 & ~w31620;
assign w31622 = pi05905 & ~w31615;
assign w31623 = ~pi02160 & w31615;
assign w31624 = ~w31622 & ~w31623;
assign w31625 = pi05906 & ~w31615;
assign w31626 = ~pi02708 & w31615;
assign w31627 = ~w31625 & ~w31626;
assign w31628 = pi05907 & ~w31615;
assign w31629 = ~pi02709 & w31615;
assign w31630 = ~w31628 & ~w31629;
assign w31631 = pi05908 & ~w31615;
assign w31632 = ~pi02710 & w31615;
assign w31633 = ~w31631 & ~w31632;
assign w31634 = ~w16892 & w20170;
assign w31635 = pi05909 & ~w31634;
assign w31636 = w17925 & w20170;
assign w31637 = ~w31635 & ~w31636;
assign w31638 = pi05910 & ~w31634;
assign w31639 = ~pi02707 & w31634;
assign w31640 = ~w31638 & ~w31639;
assign w31641 = pi05911 & ~w31634;
assign w31642 = ~pi02160 & w31634;
assign w31643 = ~w31641 & ~w31642;
assign w31644 = pi05912 & ~w31634;
assign w31645 = ~pi02723 & w31634;
assign w31646 = ~w31644 & ~w31645;
assign w31647 = pi05913 & ~w31634;
assign w31648 = ~pi02708 & w31634;
assign w31649 = ~w31647 & ~w31648;
assign w31650 = pi05914 & ~w31634;
assign w31651 = ~pi02709 & w31634;
assign w31652 = ~w31650 & ~w31651;
assign w31653 = pi05915 & ~w31634;
assign w31654 = ~pi02710 & w31634;
assign w31655 = ~w31653 & ~w31654;
assign w31656 = ~w16892 & w16931;
assign w31657 = pi05916 & ~w31656;
assign w31658 = w16931 & w17925;
assign w31659 = ~w31657 & ~w31658;
assign w31660 = pi05917 & ~w31656;
assign w31661 = ~pi02707 & w31656;
assign w31662 = ~w31660 & ~w31661;
assign w31663 = pi05918 & ~w31656;
assign w31664 = ~pi02160 & w31656;
assign w31665 = ~w31663 & ~w31664;
assign w31666 = pi05919 & ~w31656;
assign w31667 = ~pi02708 & w31656;
assign w31668 = ~w31666 & ~w31667;
assign w31669 = pi05920 & ~w31656;
assign w31670 = ~pi02709 & w31656;
assign w31671 = ~w31669 & ~w31670;
assign w31672 = w16941 & ~w16992;
assign w31673 = pi05921 & ~w31672;
assign w31674 = ~pi02703 & w31672;
assign w31675 = ~w31673 & ~w31674;
assign w31676 = ~w16928 & w18278;
assign w31677 = pi05922 & ~w31676;
assign w31678 = ~pi02178 & w31676;
assign w31679 = ~w31677 & ~w31678;
assign w31680 = ~w16892 & w18772;
assign w31681 = pi05923 & ~w31680;
assign w31682 = ~pi02705 & w31680;
assign w31683 = ~w31681 & ~w31682;
assign w31684 = pi05924 & ~w31672;
assign w31685 = w16941 & w17811;
assign w31686 = ~w31684 & ~w31685;
assign w31687 = pi05925 & ~w31680;
assign w31688 = ~pi02706 & w31680;
assign w31689 = ~w31687 & ~w31688;
assign w31690 = pi05926 & ~w31680;
assign w31691 = ~pi02707 & w31680;
assign w31692 = ~w31690 & ~w31691;
assign w31693 = pi05927 & ~w31672;
assign w31694 = ~pi02169 & w31672;
assign w31695 = ~w31693 & ~w31694;
assign w31696 = pi05928 & ~w31680;
assign w31697 = ~pi02160 & w31680;
assign w31698 = ~w31696 & ~w31697;
assign w31699 = pi05929 & ~w31680;
assign w31700 = ~pi02723 & w31680;
assign w31701 = ~w31699 & ~w31700;
assign w31702 = pi05930 & ~w31680;
assign w31703 = ~pi02709 & w31680;
assign w31704 = ~w31702 & ~w31703;
assign w31705 = pi05931 & ~w31680;
assign w31706 = ~pi02710 & w31680;
assign w31707 = ~w31705 & ~w31706;
assign w31708 = pi05932 & ~w31672;
assign w31709 = ~pi02167 & w31672;
assign w31710 = ~w31708 & ~w31709;
assign w31711 = pi05933 & ~w31672;
assign w31712 = ~pi02164 & w31672;
assign w31713 = ~w31711 & ~w31712;
assign w31714 = pi05934 & ~w31672;
assign w31715 = ~pi02722 & w31672;
assign w31716 = ~w31714 & ~w31715;
assign w31717 = pi05935 & ~w31672;
assign w31718 = w16941 & w17594;
assign w31719 = ~w31717 & ~w31718;
assign w31720 = ~w16892 & w18300;
assign w31721 = pi05936 & ~w31720;
assign w31722 = w17925 & w18300;
assign w31723 = ~w31721 & ~w31722;
assign w31724 = pi05937 & ~w31720;
assign w31725 = ~pi02707 & w31720;
assign w31726 = ~w31724 & ~w31725;
assign w31727 = pi05938 & ~w31720;
assign w31728 = ~pi02160 & w31720;
assign w31729 = ~w31727 & ~w31728;
assign w31730 = pi05939 & ~w31720;
assign w31731 = w17671 & w18300;
assign w31732 = ~w31730 & ~w31731;
assign w31733 = pi05940 & ~w31720;
assign w31734 = ~pi02708 & w31720;
assign w31735 = ~w31733 & ~w31734;
assign w31736 = pi05941 & ~w31720;
assign w31737 = ~pi02709 & w31720;
assign w31738 = ~w31736 & ~w31737;
assign w31739 = pi05942 & ~w31720;
assign w31740 = ~pi02710 & w31720;
assign w31741 = ~w31739 & ~w31740;
assign w31742 = pi05943 & ~w21135;
assign w31743 = ~pi02705 & w21135;
assign w31744 = ~w31742 & ~w31743;
assign w31745 = pi05944 & ~w29203;
assign w31746 = ~pi02721 & w29203;
assign w31747 = ~w31745 & ~w31746;
assign w31748 = pi05945 & ~w21135;
assign w31749 = ~pi02706 & w21135;
assign w31750 = ~w31748 & ~w31749;
assign w31751 = pi05946 & ~w29203;
assign w31752 = w18278 & w19797;
assign w31753 = ~w31751 & ~w31752;
assign w31754 = pi05947 & ~w21135;
assign w31755 = ~pi02160 & w21135;
assign w31756 = ~w31754 & ~w31755;
assign w31757 = pi05948 & ~w21135;
assign w31758 = ~pi02723 & w21135;
assign w31759 = ~w31757 & ~w31758;
assign w31760 = pi05949 & ~w21135;
assign w31761 = ~pi02709 & w21135;
assign w31762 = ~w31760 & ~w31761;
assign w31763 = pi05950 & ~w21135;
assign w31764 = ~pi02710 & w21135;
assign w31765 = ~w31763 & ~w31764;
assign w31766 = pi05951 & ~w29203;
assign w31767 = ~pi02167 & w29203;
assign w31768 = ~w31766 & ~w31767;
assign w31769 = pi05952 & ~w29203;
assign w31770 = ~pi02718 & w29203;
assign w31771 = ~w31769 & ~w31770;
assign w31772 = pi05953 & ~w29203;
assign w31773 = ~pi02164 & w29203;
assign w31774 = ~w31772 & ~w31773;
assign w31775 = pi05954 & ~w29203;
assign w31776 = ~pi02722 & w29203;
assign w31777 = ~w31775 & ~w31776;
assign w31778 = pi05955 & ~w29203;
assign w31779 = ~pi02719 & w29203;
assign w31780 = ~w31778 & ~w31779;
assign w31781 = pi05956 & ~w21030;
assign w31782 = ~pi02705 & w21030;
assign w31783 = ~w31781 & ~w31782;
assign w31784 = pi05957 & ~w20953;
assign w31785 = ~pi02721 & w20953;
assign w31786 = ~w31784 & ~w31785;
assign w31787 = pi05958 & ~w21030;
assign w31788 = ~pi02706 & w21030;
assign w31789 = ~w31787 & ~w31788;
assign w31790 = pi05959 & ~w20953;
assign w31791 = ~pi02169 & w20953;
assign w31792 = ~w31790 & ~w31791;
assign w31793 = pi05960 & ~w21030;
assign w31794 = ~pi02160 & w21030;
assign w31795 = ~w31793 & ~w31794;
assign w31796 = pi05961 & ~w21030;
assign w31797 = ~pi02723 & w21030;
assign w31798 = ~w31796 & ~w31797;
assign w31799 = pi05962 & ~w21030;
assign w31800 = w17754 & w18689;
assign w31801 = ~w31799 & ~w31800;
assign w31802 = pi05963 & ~w21030;
assign w31803 = ~pi02709 & w21030;
assign w31804 = ~w31802 & ~w31803;
assign w31805 = pi05964 & ~w21030;
assign w31806 = w17754 & w18364;
assign w31807 = ~w31805 & ~w31806;
assign w31808 = pi05965 & ~w20953;
assign w31809 = ~pi02167 & w20953;
assign w31810 = ~w31808 & ~w31809;
assign w31811 = pi05966 & ~w20953;
assign w31812 = ~pi02164 & w20953;
assign w31813 = ~w31811 & ~w31812;
assign w31814 = pi05967 & ~w20953;
assign w31815 = w18001 & w19312;
assign w31816 = ~w31814 & ~w31815;
assign w31817 = pi05968 & ~w20953;
assign w31818 = ~pi02719 & w20953;
assign w31819 = ~w31817 & ~w31818;
assign w31820 = pi05969 & ~w20698;
assign w31821 = ~pi02703 & w20698;
assign w31822 = ~w31820 & ~w31821;
assign w31823 = pi05970 & ~w20698;
assign w31824 = w17811 & w17837;
assign w31825 = ~w31823 & ~w31824;
assign w31826 = pi05971 & ~w20596;
assign w31827 = ~pi02706 & w20596;
assign w31828 = ~w31826 & ~w31827;
assign w31829 = pi05972 & ~w20698;
assign w31830 = w17837 & w19797;
assign w31831 = ~w31829 & ~w31830;
assign w31832 = pi05973 & ~w20596;
assign w31833 = ~pi02160 & w20596;
assign w31834 = ~w31832 & ~w31833;
assign w31835 = pi05974 & ~w20596;
assign w31836 = ~pi02723 & w20596;
assign w31837 = ~w31835 & ~w31836;
assign w31838 = pi05975 & ~w20596;
assign w31839 = ~pi02708 & w20596;
assign w31840 = ~w31838 & ~w31839;
assign w31841 = pi05976 & ~w20596;
assign w31842 = ~pi02709 & w20596;
assign w31843 = ~w31841 & ~w31842;
assign w31844 = pi05977 & ~w20596;
assign w31845 = ~pi02710 & w20596;
assign w31846 = ~w31844 & ~w31845;
assign w31847 = pi05978 & ~w20698;
assign w31848 = ~pi02167 & w20698;
assign w31849 = ~w31847 & ~w31848;
assign w31850 = pi05979 & ~w20600;
assign w31851 = ~pi02705 & w20600;
assign w31852 = ~w31850 & ~w31851;
assign w31853 = pi05980 & ~w20600;
assign w31854 = ~pi02706 & w20600;
assign w31855 = ~w31853 & ~w31854;
assign w31856 = pi05981 & ~w20698;
assign w31857 = ~pi02164 & w20698;
assign w31858 = ~w31856 & ~w31857;
assign w31859 = pi05982 & ~w20600;
assign w31860 = ~pi02160 & w20600;
assign w31861 = ~w31859 & ~w31860;
assign w31862 = pi05983 & ~w20698;
assign w31863 = ~pi02722 & w20698;
assign w31864 = ~w31862 & ~w31863;
assign w31865 = pi05984 & ~w20600;
assign w31866 = ~pi02723 & w20600;
assign w31867 = ~w31865 & ~w31866;
assign w31868 = pi05985 & ~w20600;
assign w31869 = w17289 & w18092;
assign w31870 = ~w31868 & ~w31869;
assign w31871 = pi05986 & ~w20698;
assign w31872 = ~pi02719 & w20698;
assign w31873 = ~w31871 & ~w31872;
assign w31874 = pi05987 & ~w20600;
assign w31875 = ~pi02710 & w20600;
assign w31876 = ~w31874 & ~w31875;
assign w31877 = ~w16992 & w20465;
assign w31878 = pi05988 & ~w31877;
assign w31879 = w17532 & w20465;
assign w31880 = ~w31878 & ~w31879;
assign w31881 = pi05989 & ~w20574;
assign w31882 = w17925 & w17938;
assign w31883 = ~w31881 & ~w31882;
assign w31884 = pi05990 & ~w20574;
assign w31885 = w17938 & w18067;
assign w31886 = ~w31884 & ~w31885;
assign w31887 = pi05991 & ~w31877;
assign w31888 = w17811 & w20465;
assign w31889 = ~w31887 & ~w31888;
assign w31890 = pi05992 & ~w20574;
assign w31891 = w17938 & w18234;
assign w31892 = ~w31890 & ~w31891;
assign w31893 = pi05993 & ~w20574;
assign w31894 = w17671 & w17938;
assign w31895 = ~w31893 & ~w31894;
assign w31896 = pi05994 & ~w31877;
assign w31897 = w19797 & w20465;
assign w31898 = ~w31896 & ~w31897;
assign w31899 = pi05995 & ~w20574;
assign w31900 = w17938 & w18092;
assign w31901 = ~w31899 & ~w31900;
assign w31902 = pi05996 & ~w20574;
assign w31903 = w17938 & w18364;
assign w31904 = ~w31902 & ~w31903;
assign w31905 = pi05997 & ~w31877;
assign w31906 = w17586 & w20465;
assign w31907 = ~w31905 & ~w31906;
assign w31908 = pi05998 & ~w31877;
assign w31909 = w19273 & w20465;
assign w31910 = ~w31908 & ~w31909;
assign w31911 = pi05999 & ~w20489;
assign w31912 = ~pi02706 & w20489;
assign w31913 = ~w31911 & ~w31912;
assign w31914 = pi06000 & ~w31877;
assign w31915 = w17620 & w20465;
assign w31916 = ~w31914 & ~w31915;
assign w31917 = pi06001 & ~w30635;
assign w31918 = ~pi02706 & w30635;
assign w31919 = ~w31917 & ~w31918;
assign w31920 = pi06002 & ~w20489;
assign w31921 = ~pi02160 & w20489;
assign w31922 = ~w31920 & ~w31921;
assign w31923 = pi06003 & ~w31877;
assign w31924 = w19312 & w20465;
assign w31925 = ~w31923 & ~w31924;
assign w31926 = pi06004 & ~w20489;
assign w31927 = ~pi02723 & w20489;
assign w31928 = ~w31926 & ~w31927;
assign w31929 = pi06005 & ~w20489;
assign w31930 = ~pi02708 & w20489;
assign w31931 = ~w31929 & ~w31930;
assign w31932 = pi06006 & ~w20489;
assign w31933 = ~pi02709 & w20489;
assign w31934 = ~w31932 & ~w31933;
assign w31935 = pi06007 & ~w20489;
assign w31936 = ~pi02710 & w20489;
assign w31937 = ~w31935 & ~w31936;
assign w31938 = pi06008 & ~w31877;
assign w31939 = w17594 & w20465;
assign w31940 = ~w31938 & ~w31939;
assign w31941 = pi06009 & ~w20446;
assign w31942 = ~pi02706 & w20446;
assign w31943 = ~w31941 & ~w31942;
assign w31944 = pi06010 & ~w20446;
assign w31945 = ~pi02707 & w20446;
assign w31946 = ~w31944 & ~w31945;
assign w31947 = pi06011 & ~w20446;
assign w31948 = ~pi02160 & w20446;
assign w31949 = ~w31947 & ~w31948;
assign w31950 = pi06012 & ~w20446;
assign w31951 = ~pi02708 & w20446;
assign w31952 = ~w31950 & ~w31951;
assign w31953 = pi06013 & ~w20446;
assign w31954 = w17108 & w18092;
assign w31955 = ~w31953 & ~w31954;
assign w31956 = pi06014 & ~w20446;
assign w31957 = ~pi02710 & w20446;
assign w31958 = ~w31956 & ~w31957;
assign w31959 = pi06015 & ~w17099;
assign w31960 = ~pi02706 & w17099;
assign w31961 = ~w31959 & ~w31960;
assign w31962 = pi06016 & ~w17099;
assign w31963 = ~pi02707 & w17099;
assign w31964 = ~w31962 & ~w31963;
assign w31965 = pi06017 & ~w17099;
assign w31966 = ~pi02160 & w17099;
assign w31967 = ~w31965 & ~w31966;
assign w31968 = pi06018 & ~w17099;
assign w31969 = w17098 & w17671;
assign w31970 = ~w31968 & ~w31969;
assign w31971 = pi06019 & ~w17099;
assign w31972 = w17098 & w18689;
assign w31973 = ~w31971 & ~w31972;
assign w31974 = pi06020 & ~w17099;
assign w31975 = w17098 & w18092;
assign w31976 = ~w31974 & ~w31975;
assign w31977 = pi06021 & ~w17099;
assign w31978 = w17098 & w18364;
assign w31979 = ~w31977 & ~w31978;
assign w31980 = pi06022 & ~w20245;
assign w31981 = ~pi02706 & w20245;
assign w31982 = ~w31980 & ~w31981;
assign w31983 = pi06023 & ~w20245;
assign w31984 = ~pi02707 & w20245;
assign w31985 = ~w31983 & ~w31984;
assign w31986 = pi06024 & ~w20245;
assign w31987 = ~pi02160 & w20245;
assign w31988 = ~w31986 & ~w31987;
assign w31989 = pi06025 & ~w20245;
assign w31990 = ~pi02708 & w20245;
assign w31991 = ~w31989 & ~w31990;
assign w31992 = pi06026 & ~w20245;
assign w31993 = ~pi02709 & w20245;
assign w31994 = ~w31992 & ~w31993;
assign w31995 = pi06027 & ~w20245;
assign w31996 = ~pi02710 & w20245;
assign w31997 = ~w31995 & ~w31996;
assign w31998 = pi06028 & ~w18703;
assign w31999 = w17811 & w17814;
assign w32000 = ~w31998 & ~w31999;
assign w32001 = pi06029 & ~w18703;
assign w32002 = w17814 & w19797;
assign w32003 = ~w32001 & ~w32002;
assign w32004 = pi06030 & ~w18543;
assign w32005 = ~pi02705 & w18543;
assign w32006 = ~w32004 & ~w32005;
assign w32007 = pi06031 & ~w18703;
assign w32008 = w17586 & w17814;
assign w32009 = ~w32007 & ~w32008;
assign w32010 = pi06032 & ~w18543;
assign w32011 = ~pi02706 & w18543;
assign w32012 = ~w32010 & ~w32011;
assign w32013 = pi06033 & ~w18703;
assign w32014 = w17814 & w19273;
assign w32015 = ~w32013 & ~w32014;
assign w32016 = pi06034 & ~w18543;
assign w32017 = ~pi02707 & w18543;
assign w32018 = ~w32016 & ~w32017;
assign w32019 = pi06035 & ~w18703;
assign w32020 = w17620 & w17814;
assign w32021 = ~w32019 & ~w32020;
assign w32022 = pi06036 & ~w18543;
assign w32023 = ~pi02723 & w18543;
assign w32024 = ~w32022 & ~w32023;
assign w32025 = pi06037 & ~w18543;
assign w32026 = w18542 & w18689;
assign w32027 = ~w32025 & ~w32026;
assign w32028 = pi06038 & ~w18703;
assign w32029 = w17814 & w19312;
assign w32030 = ~w32028 & ~w32029;
assign w32031 = pi06039 & ~w18543;
assign w32032 = w18364 & w18542;
assign w32033 = ~w32031 & ~w32032;
assign w32034 = pi06040 & ~w18663;
assign w32035 = w18578 & w18662;
assign w32036 = ~w32034 & ~w32035;
assign w32037 = pi06041 & ~w18663;
assign w32038 = w17925 & w18662;
assign w32039 = ~w32037 & ~w32038;
assign w32040 = pi06042 & ~w18663;
assign w32041 = w18067 & w18662;
assign w32042 = ~w32040 & ~w32041;
assign w32043 = pi06043 & ~w18590;
assign w32044 = ~pi02703 & w18590;
assign w32045 = ~w32043 & ~w32044;
assign w32046 = pi06044 & ~w18663;
assign w32047 = w18234 & w18662;
assign w32048 = ~w32046 & ~w32047;
assign w32049 = pi06045 & ~w18663;
assign w32050 = w17671 & w18662;
assign w32051 = ~w32049 & ~w32050;
assign w32052 = pi06046 & ~w18590;
assign w32053 = ~pi02721 & w18590;
assign w32054 = ~w32052 & ~w32053;
assign w32055 = pi06047 & ~w18663;
assign w32056 = w18662 & w18689;
assign w32057 = ~w32055 & ~w32056;
assign w32058 = pi06048 & ~w18663;
assign w32059 = w18364 & w18662;
assign w32060 = ~w32058 & ~w32059;
assign w32061 = pi06049 & ~w18590;
assign w32062 = ~pi02169 & w18590;
assign w32063 = ~w32061 & ~w32062;
assign w32064 = pi06050 & ~w18590;
assign w32065 = ~pi02718 & w18590;
assign w32066 = ~w32064 & ~w32065;
assign w32067 = pi06051 & ~w18618;
assign w32068 = ~pi02706 & w18618;
assign w32069 = ~w32067 & ~w32068;
assign w32070 = pi06052 & ~w18590;
assign w32071 = ~pi02167 & w18590;
assign w32072 = ~w32070 & ~w32071;
assign w32073 = pi06053 & ~w18618;
assign w32074 = ~pi02707 & w18618;
assign w32075 = ~w32073 & ~w32074;
assign w32076 = pi06054 & ~w22189;
assign w32077 = ~pi02160 & w22189;
assign w32078 = ~w32076 & ~w32077;
assign w32079 = pi06055 & ~w18590;
assign w32080 = ~pi02164 & w18590;
assign w32081 = ~w32079 & ~w32080;
assign w32082 = pi06056 & ~w18618;
assign w32083 = ~pi02723 & w18618;
assign w32084 = ~w32082 & ~w32083;
assign w32085 = pi06057 & ~w18618;
assign w32086 = ~pi02708 & w18618;
assign w32087 = ~w32085 & ~w32086;
assign w32088 = pi06058 & ~w18618;
assign w32089 = ~pi02709 & w18618;
assign w32090 = ~w32088 & ~w32089;
assign w32091 = pi06059 & ~w18590;
assign w32092 = ~pi02722 & w18590;
assign w32093 = ~w32091 & ~w32092;
assign w32094 = pi06060 & ~w18618;
assign w32095 = w18364 & w18617;
assign w32096 = ~w32094 & ~w32095;
assign w32097 = pi06061 & ~w18601;
assign w32098 = ~pi02705 & w18601;
assign w32099 = ~w32097 & ~w32098;
assign w32100 = pi06062 & ~w18601;
assign w32101 = ~pi02706 & w18601;
assign w32102 = ~w32100 & ~w32101;
assign w32103 = pi06063 & ~w18601;
assign w32104 = ~pi02707 & w18601;
assign w32105 = ~w32103 & ~w32104;
assign w32106 = pi06064 & ~w18559;
assign w32107 = w17532 & w17775;
assign w32108 = ~w32106 & ~w32107;
assign w32109 = pi06065 & ~w18601;
assign w32110 = ~pi02723 & w18601;
assign w32111 = ~w32109 & ~w32110;
assign w32112 = pi06066 & ~w18601;
assign w32113 = ~pi02708 & w18601;
assign w32114 = ~w32112 & ~w32113;
assign w32115 = pi06067 & ~w18601;
assign w32116 = w18092 & w18554;
assign w32117 = ~w32115 & ~w32116;
assign w32118 = pi06068 & ~w18559;
assign w32119 = w17775 & w19797;
assign w32120 = ~w32118 & ~w32119;
assign w32121 = pi06069 & ~w18559;
assign w32122 = w17775 & w17811;
assign w32123 = ~w32121 & ~w32122;
assign w32124 = pi06070 & ~w18559;
assign w32125 = w17775 & w19273;
assign w32126 = ~w32124 & ~w32125;
assign w32127 = pi06071 & ~w18559;
assign w32128 = w17586 & w17775;
assign w32129 = ~w32127 & ~w32128;
assign w32130 = pi06072 & ~w18559;
assign w32131 = w17620 & w17775;
assign w32132 = ~w32130 & ~w32131;
assign w32133 = pi06073 & ~w18559;
assign w32134 = w17775 & w19312;
assign w32135 = ~w32133 & ~w32134;
assign w32136 = pi06074 & ~w17040;
assign w32137 = ~pi02705 & w17040;
assign w32138 = ~w32136 & ~w32137;
assign w32139 = pi06075 & ~w17040;
assign w32140 = ~pi02706 & w17040;
assign w32141 = ~w32139 & ~w32140;
assign w32142 = pi06076 & ~w17040;
assign w32143 = ~pi02707 & w17040;
assign w32144 = ~w32142 & ~w32143;
assign w32145 = ~w16992 & w17573;
assign w32146 = pi06077 & ~w32145;
assign w32147 = ~pi02703 & w32145;
assign w32148 = ~w32146 & ~w32147;
assign w32149 = pi06078 & ~w17040;
assign w32150 = ~pi02723 & w17040;
assign w32151 = ~w32149 & ~w32150;
assign w32152 = pi06079 & ~w32145;
assign w32153 = ~pi02721 & w32145;
assign w32154 = ~w32152 & ~w32153;
assign w32155 = pi06080 & ~w17040;
assign w32156 = ~pi02708 & w17040;
assign w32157 = ~w32155 & ~w32156;
assign w32158 = pi06081 & ~w17040;
assign w32159 = ~pi02710 & w17040;
assign w32160 = ~w32158 & ~w32159;
assign w32161 = pi06082 & ~w32145;
assign w32162 = ~pi02169 & w32145;
assign w32163 = ~w32161 & ~w32162;
assign w32164 = pi06083 & ~w32145;
assign w32165 = ~pi02718 & w32145;
assign w32166 = ~w32164 & ~w32165;
assign w32167 = pi06084 & ~w32145;
assign w32168 = ~pi02164 & w32145;
assign w32169 = ~w32167 & ~w32168;
assign w32170 = pi06085 & ~w32145;
assign w32171 = ~pi02167 & w32145;
assign w32172 = ~w32170 & ~w32171;
assign w32173 = pi06086 & ~w32145;
assign w32174 = w17573 & w19312;
assign w32175 = ~w32173 & ~w32174;
assign w32176 = pi06087 & ~w32145;
assign w32177 = w17573 & w17594;
assign w32178 = ~w32176 & ~w32177;
assign w32179 = pi06088 & ~w18400;
assign w32180 = ~pi02721 & w18400;
assign w32181 = ~w32179 & ~w32180;
assign w32182 = pi06089 & ~w18400;
assign w32183 = ~pi02169 & w18400;
assign w32184 = ~w32182 & ~w32183;
assign w32185 = pi06090 & ~w18455;
assign w32186 = w18454 & w18578;
assign w32187 = ~w32185 & ~w32186;
assign w32188 = pi06091 & ~w18400;
assign w32189 = w17028 & w17586;
assign w32190 = ~w32188 & ~w32189;
assign w32191 = pi06092 & ~w18455;
assign w32192 = w18067 & w18454;
assign w32193 = ~w32191 & ~w32192;
assign w32194 = pi06093 & ~w18455;
assign w32195 = w18234 & w18454;
assign w32196 = ~w32194 & ~w32195;
assign w32197 = pi06094 & ~w18455;
assign w32198 = w17671 & w18454;
assign w32199 = ~w32197 & ~w32198;
assign w32200 = pi06095 & ~w18455;
assign w32201 = w18454 & w18689;
assign w32202 = ~w32200 & ~w32201;
assign w32203 = pi06096 & ~w18455;
assign w32204 = w18092 & w18454;
assign w32205 = ~w32203 & ~w32204;
assign w32206 = pi06097 & ~w18400;
assign w32207 = w17028 & w17620;
assign w32208 = ~w32206 & ~w32207;
assign w32209 = pi06098 & ~w18455;
assign w32210 = w18364 & w18454;
assign w32211 = ~w32209 & ~w32210;
assign w32212 = pi06099 & ~w18400;
assign w32213 = ~pi02722 & w18400;
assign w32214 = ~w32212 & ~w32213;
assign w32215 = pi06100 & ~w18378;
assign w32216 = ~pi02705 & w18378;
assign w32217 = ~w32215 & ~w32216;
assign w32218 = pi06101 & ~w18378;
assign w32219 = ~pi02707 & w18378;
assign w32220 = ~w32218 & ~w32219;
assign w32221 = pi06102 & ~w18400;
assign w32222 = ~pi02719 & w18400;
assign w32223 = ~w32221 & ~w32222;
assign w32224 = pi06103 & ~w18378;
assign w32225 = w17710 & w18234;
assign w32226 = ~w32224 & ~w32225;
assign w32227 = pi06104 & ~w18378;
assign w32228 = ~pi02723 & w18378;
assign w32229 = ~w32227 & ~w32228;
assign w32230 = pi06105 & ~w18378;
assign w32231 = ~pi02708 & w18378;
assign w32232 = ~w32230 & ~w32231;
assign w32233 = pi06106 & ~w18378;
assign w32234 = ~pi02709 & w18378;
assign w32235 = ~w32233 & ~w32234;
assign w32236 = pi06107 & ~w18378;
assign w32237 = ~pi02710 & w18378;
assign w32238 = ~w32236 & ~w32237;
assign w32239 = ~w16892 & w18468;
assign w32240 = pi06108 & ~w32239;
assign w32241 = ~pi02705 & w32239;
assign w32242 = ~w32240 & ~w32241;
assign w32243 = pi06109 & ~w18151;
assign w32244 = ~pi02169 & w18151;
assign w32245 = ~w32243 & ~w32244;
assign w32246 = pi06110 & ~w32239;
assign w32247 = ~pi02706 & w32239;
assign w32248 = ~w32246 & ~w32247;
assign w32249 = pi06111 & ~w18151;
assign w32250 = ~pi02718 & w18151;
assign w32251 = ~w32249 & ~w32250;
assign w32252 = pi06112 & ~w32239;
assign w32253 = w18067 & w18468;
assign w32254 = ~w32252 & ~w32253;
assign w32255 = pi06113 & ~w32239;
assign w32256 = ~pi02160 & w32239;
assign w32257 = ~w32255 & ~w32256;
assign w32258 = pi06114 & ~w32239;
assign w32259 = ~pi02723 & w32239;
assign w32260 = ~w32258 & ~w32259;
assign w32261 = pi06115 & ~w32239;
assign w32262 = ~pi02708 & w32239;
assign w32263 = ~w32261 & ~w32262;
assign w32264 = pi06116 & ~w32239;
assign w32265 = w18092 & w18468;
assign w32266 = ~w32264 & ~w32265;
assign w32267 = pi06117 & ~w32239;
assign w32268 = ~pi02710 & w32239;
assign w32269 = ~w32267 & ~w32268;
assign w32270 = pi06118 & ~w18164;
assign w32271 = ~pi02705 & w18164;
assign w32272 = ~w32270 & ~w32271;
assign w32273 = pi06119 & ~w18151;
assign w32274 = ~pi02722 & w18151;
assign w32275 = ~w32273 & ~w32274;
assign w32276 = pi06120 & ~w18151;
assign w32277 = ~pi02719 & w18151;
assign w32278 = ~w32276 & ~w32277;
assign w32279 = pi06121 & ~w18164;
assign w32280 = ~pi02707 & w18164;
assign w32281 = ~w32279 & ~w32280;
assign w32282 = pi06122 & ~w18164;
assign w32283 = ~pi02160 & w18164;
assign w32284 = ~w32282 & ~w32283;
assign w32285 = pi06123 & ~w18164;
assign w32286 = ~pi02723 & w18164;
assign w32287 = ~w32285 & ~w32286;
assign w32288 = ~w16992 & w17006;
assign w32289 = pi06124 & ~w32288;
assign w32290 = w17006 & w17532;
assign w32291 = ~w32289 & ~w32290;
assign w32292 = pi06125 & ~w18164;
assign w32293 = ~pi02708 & w18164;
assign w32294 = ~w32292 & ~w32293;
assign w32295 = pi06126 & ~w18164;
assign w32296 = ~pi02709 & w18164;
assign w32297 = ~w32295 & ~w32296;
assign w32298 = pi06127 & ~w32288;
assign w32299 = ~pi02721 & w32288;
assign w32300 = ~w32298 & ~w32299;
assign w32301 = pi06128 & ~w17973;
assign w32302 = ~pi02705 & w17973;
assign w32303 = ~w32301 & ~w32302;
assign w32304 = pi06129 & ~w32288;
assign w32305 = ~pi02169 & w32288;
assign w32306 = ~w32304 & ~w32305;
assign w32307 = pi06130 & ~w32288;
assign w32308 = ~pi02718 & w32288;
assign w32309 = ~w32307 & ~w32308;
assign w32310 = pi06131 & ~w17973;
assign w32311 = ~pi02707 & w17973;
assign w32312 = ~w32310 & ~w32311;
assign w32313 = pi06132 & ~w17973;
assign w32314 = w17631 & w18234;
assign w32315 = ~w32313 & ~w32314;
assign w32316 = pi06133 & ~w32288;
assign w32317 = ~pi02167 & w32288;
assign w32318 = ~w32316 & ~w32317;
assign w32319 = pi06134 & ~w17973;
assign w32320 = ~pi02708 & w17973;
assign w32321 = ~w32319 & ~w32320;
assign w32322 = pi06135 & ~w17973;
assign w32323 = ~pi02709 & w17973;
assign w32324 = ~w32322 & ~w32323;
assign w32325 = pi06136 & ~w17973;
assign w32326 = ~pi02710 & w17973;
assign w32327 = ~w32325 & ~w32326;
assign w32328 = pi06137 & ~w32288;
assign w32329 = ~pi02164 & w32288;
assign w32330 = ~w32328 & ~w32329;
assign w32331 = pi06138 & ~w32288;
assign w32332 = ~pi02722 & w32288;
assign w32333 = ~w32331 & ~w32332;
assign w32334 = pi06139 & ~w32288;
assign w32335 = ~pi02719 & w32288;
assign w32336 = ~w32334 & ~w32335;
assign w32337 = pi06140 & ~w17735;
assign w32338 = ~pi02721 & w17735;
assign w32339 = ~w32337 & ~w32338;
assign w32340 = pi06141 & ~w17780;
assign w32341 = w17416 & w18578;
assign w32342 = ~w32340 & ~w32341;
assign w32343 = pi06142 & ~w17780;
assign w32344 = w17416 & w17925;
assign w32345 = ~w32343 & ~w32344;
assign w32346 = pi06143 & ~w17780;
assign w32347 = w17416 & w18067;
assign w32348 = ~w32346 & ~w32347;
assign w32349 = pi06144 & ~w17780;
assign w32350 = w17416 & w18234;
assign w32351 = ~w32349 & ~w32350;
assign w32352 = pi06145 & ~w17735;
assign w32353 = ~pi02718 & w17735;
assign w32354 = ~w32352 & ~w32353;
assign w32355 = pi06146 & ~w17735;
assign w32356 = ~pi02167 & w17735;
assign w32357 = ~w32355 & ~w32356;
assign w32358 = pi06147 & ~w17780;
assign w32359 = w17416 & w18689;
assign w32360 = ~w32358 & ~w32359;
assign w32361 = pi06148 & ~w17780;
assign w32362 = w17416 & w18092;
assign w32363 = ~w32361 & ~w32362;
assign w32364 = pi06149 & ~w17780;
assign w32365 = w17416 & w18364;
assign w32366 = ~w32364 & ~w32365;
assign w32367 = pi06150 & ~w17735;
assign w32368 = ~pi02164 & w17735;
assign w32369 = ~w32367 & ~w32368;
assign w32370 = pi06151 & ~w17735;
assign w32371 = w17734 & w19312;
assign w32372 = ~w32370 & ~w32371;
assign w32373 = pi06152 & ~w17735;
assign w32374 = ~pi02719 & w17735;
assign w32375 = ~w32373 & ~w32374;
assign w32376 = pi06153 & ~w17407;
assign w32377 = ~pi02721 & w17407;
assign w32378 = ~w32376 & ~w32377;
assign w32379 = pi06154 & ~w17407;
assign w32380 = ~pi02169 & w17407;
assign w32381 = ~w32379 & ~w32380;
assign w32382 = pi06155 & ~w17407;
assign w32383 = ~pi02718 & w17407;
assign w32384 = ~w32382 & ~w32383;
assign w32385 = pi06156 & ~w21281;
assign w32386 = ~pi02705 & w21281;
assign w32387 = ~w32385 & ~w32386;
assign w32388 = pi06157 & ~w17407;
assign w32389 = ~pi02164 & w17407;
assign w32390 = ~w32388 & ~w32389;
assign w32391 = pi06158 & ~w21281;
assign w32392 = ~pi02706 & w21281;
assign w32393 = ~w32391 & ~w32392;
assign w32394 = pi06159 & ~w17407;
assign w32395 = ~pi02722 & w17407;
assign w32396 = ~w32394 & ~w32395;
assign w32397 = pi06160 & ~w17407;
assign w32398 = ~pi02719 & w17407;
assign w32399 = ~w32397 & ~w32398;
assign w32400 = pi06161 & ~w21281;
assign w32401 = ~pi02160 & w21281;
assign w32402 = ~w32400 & ~w32401;
assign w32403 = pi06162 & ~w21281;
assign w32404 = ~pi02723 & w21281;
assign w32405 = ~w32403 & ~w32404;
assign w32406 = pi06163 & ~w21281;
assign w32407 = ~pi02708 & w21281;
assign w32408 = ~w32406 & ~w32407;
assign w32409 = pi06164 & ~w21281;
assign w32410 = ~pi02709 & w21281;
assign w32411 = ~w32409 & ~w32410;
assign w32412 = pi06165 & ~w21281;
assign w32413 = ~pi02710 & w21281;
assign w32414 = ~w32412 & ~w32413;
assign w32415 = ~w16892 & w17125;
assign w32416 = pi06166 & ~w32415;
assign w32417 = ~pi02705 & w32415;
assign w32418 = ~w32416 & ~w32417;
assign w32419 = pi06167 & ~w32415;
assign w32420 = ~pi02706 & w32415;
assign w32421 = ~w32419 & ~w32420;
assign w32422 = ~w16992 & w19629;
assign w32423 = pi06168 & ~w32422;
assign w32424 = ~pi02721 & w32422;
assign w32425 = ~w32423 & ~w32424;
assign w32426 = pi06169 & ~w32422;
assign w32427 = w19629 & w19797;
assign w32428 = ~w32426 & ~w32427;
assign w32429 = pi06170 & ~w32415;
assign w32430 = ~pi02160 & w32415;
assign w32431 = ~w32429 & ~w32430;
assign w32432 = pi06171 & ~w32415;
assign w32433 = ~pi02723 & w32415;
assign w32434 = ~w32432 & ~w32433;
assign w32435 = pi06172 & ~w32415;
assign w32436 = ~pi02708 & w32415;
assign w32437 = ~w32435 & ~w32436;
assign w32438 = pi06173 & ~w32415;
assign w32439 = ~pi02709 & w32415;
assign w32440 = ~w32438 & ~w32439;
assign w32441 = pi06174 & ~w32415;
assign w32442 = ~pi02710 & w32415;
assign w32443 = ~w32441 & ~w32442;
assign w32444 = pi06175 & ~w32422;
assign w32445 = ~pi02167 & w32422;
assign w32446 = ~w32444 & ~w32445;
assign w32447 = pi06176 & ~w32422;
assign w32448 = ~pi02164 & w32422;
assign w32449 = ~w32447 & ~w32448;
assign w32450 = pi06177 & ~w32422;
assign w32451 = ~pi02722 & w32422;
assign w32452 = ~w32450 & ~w32451;
assign w32453 = pi06178 & ~w32422;
assign w32454 = ~pi02719 & w32422;
assign w32455 = ~w32453 & ~w32454;
assign w32456 = ~w16992 & w19655;
assign w32457 = pi06179 & ~w32456;
assign w32458 = ~pi02721 & w32456;
assign w32459 = ~w32457 & ~w32458;
assign w32460 = pi06180 & ~w32456;
assign w32461 = ~pi02169 & w32456;
assign w32462 = ~w32460 & ~w32461;
assign w32463 = pi06181 & ~w32456;
assign w32464 = ~pi02718 & w32456;
assign w32465 = ~w32463 & ~w32464;
assign w32466 = ~w16892 & w17239;
assign w32467 = pi06182 & ~w32466;
assign w32468 = w17239 & w18578;
assign w32469 = ~w32467 & ~w32468;
assign w32470 = pi06183 & ~w32456;
assign w32471 = ~pi02164 & w32456;
assign w32472 = ~w32470 & ~w32471;
assign w32473 = pi06184 & ~w32466;
assign w32474 = ~pi02706 & w32466;
assign w32475 = ~w32473 & ~w32474;
assign w32476 = pi06185 & ~w32456;
assign w32477 = ~pi02722 & w32456;
assign w32478 = ~w32476 & ~w32477;
assign w32479 = pi06186 & ~w32466;
assign w32480 = ~pi02160 & w32466;
assign w32481 = ~w32479 & ~w32480;
assign w32482 = pi06187 & ~w32466;
assign w32483 = ~pi02723 & w32466;
assign w32484 = ~w32482 & ~w32483;
assign w32485 = pi06188 & ~w32456;
assign w32486 = ~pi02719 & w32456;
assign w32487 = ~w32485 & ~w32486;
assign w32488 = pi06189 & ~w32466;
assign w32489 = ~pi02708 & w32466;
assign w32490 = ~w32488 & ~w32489;
assign w32491 = pi06190 & ~w32466;
assign w32492 = ~pi02709 & w32466;
assign w32493 = ~w32491 & ~w32492;
assign w32494 = pi06191 & ~w32466;
assign w32495 = ~pi02710 & w32466;
assign w32496 = ~w32494 & ~w32495;
assign w32497 = ~w16892 & w17167;
assign w32498 = pi06192 & ~w32497;
assign w32499 = ~pi02705 & w32497;
assign w32500 = ~w32498 & ~w32499;
assign w32501 = pi06193 & ~w32497;
assign w32502 = ~pi02706 & w32497;
assign w32503 = ~w32501 & ~w32502;
assign w32504 = ~w16992 & w19596;
assign w32505 = pi06194 & ~w32504;
assign w32506 = ~pi02721 & w32504;
assign w32507 = ~w32505 & ~w32506;
assign w32508 = pi06195 & ~w32497;
assign w32509 = ~pi02160 & w32497;
assign w32510 = ~w32508 & ~w32509;
assign w32511 = pi06196 & ~w32504;
assign w32512 = ~pi02169 & w32504;
assign w32513 = ~w32511 & ~w32512;
assign w32514 = pi06197 & ~w32497;
assign w32515 = ~pi02723 & w32497;
assign w32516 = ~w32514 & ~w32515;
assign w32517 = pi06198 & ~w32497;
assign w32518 = ~pi02709 & w32497;
assign w32519 = ~w32517 & ~w32518;
assign w32520 = pi06199 & ~w32497;
assign w32521 = ~pi02710 & w32497;
assign w32522 = ~w32520 & ~w32521;
assign w32523 = pi06200 & ~w32504;
assign w32524 = ~pi02718 & w32504;
assign w32525 = ~w32523 & ~w32524;
assign w32526 = pi06201 & ~w32504;
assign w32527 = ~pi02167 & w32504;
assign w32528 = ~w32526 & ~w32527;
assign w32529 = pi06202 & ~w32504;
assign w32530 = ~pi02164 & w32504;
assign w32531 = ~w32529 & ~w32530;
assign w32532 = pi06203 & ~w32504;
assign w32533 = ~pi02722 & w32504;
assign w32534 = ~w32532 & ~w32533;
assign w32535 = pi06204 & ~w32504;
assign w32536 = ~pi02719 & w32504;
assign w32537 = ~w32535 & ~w32536;
assign w32538 = ~w16892 & w17205;
assign w32539 = pi06205 & ~w32538;
assign w32540 = w17205 & w18578;
assign w32541 = ~w32539 & ~w32540;
assign w32542 = pi06206 & ~w32538;
assign w32543 = w17205 & w17925;
assign w32544 = ~w32542 & ~w32543;
assign w32545 = pi06207 & ~w20425;
assign w32546 = ~pi02721 & w20425;
assign w32547 = ~w32545 & ~w32546;
assign w32548 = pi06208 & ~w32538;
assign w32549 = ~pi02160 & w32538;
assign w32550 = ~w32548 & ~w32549;
assign w32551 = pi06209 & ~w20425;
assign w32552 = ~pi02169 & w20425;
assign w32553 = ~w32551 & ~w32552;
assign w32554 = pi06210 & ~w32538;
assign w32555 = ~pi02723 & w32538;
assign w32556 = ~w32554 & ~w32555;
assign w32557 = pi06211 & ~w32538;
assign w32558 = ~pi02709 & w32538;
assign w32559 = ~w32557 & ~w32558;
assign w32560 = pi06212 & ~w20425;
assign w32561 = ~pi02718 & w20425;
assign w32562 = ~w32560 & ~w32561;
assign w32563 = pi06213 & ~w32538;
assign w32564 = ~pi02710 & w32538;
assign w32565 = ~w32563 & ~w32564;
assign w32566 = ~w16892 & w17366;
assign w32567 = pi06214 & ~w32566;
assign w32568 = ~pi02705 & w32566;
assign w32569 = ~w32567 & ~w32568;
assign w32570 = pi06215 & ~w20425;
assign w32571 = ~pi02167 & w20425;
assign w32572 = ~w32570 & ~w32571;
assign w32573 = pi06216 & ~w32566;
assign w32574 = ~pi02706 & w32566;
assign w32575 = ~w32573 & ~w32574;
assign w32576 = pi06217 & ~w32566;
assign w32577 = w17366 & w18067;
assign w32578 = ~w32576 & ~w32577;
assign w32579 = pi06218 & ~w32566;
assign w32580 = ~pi02160 & w32566;
assign w32581 = ~w32579 & ~w32580;
assign w32582 = pi06219 & ~w20425;
assign w32583 = ~pi02722 & w20425;
assign w32584 = ~w32582 & ~w32583;
assign w32585 = pi06220 & ~w32566;
assign w32586 = ~pi02723 & w32566;
assign w32587 = ~w32585 & ~w32586;
assign w32588 = pi06221 & ~w32566;
assign w32589 = ~pi02708 & w32566;
assign w32590 = ~w32588 & ~w32589;
assign w32591 = pi06222 & ~w32566;
assign w32592 = ~pi02709 & w32566;
assign w32593 = ~w32591 & ~w32592;
assign w32594 = pi06223 & ~w32566;
assign w32595 = ~pi02710 & w32566;
assign w32596 = ~w32594 & ~w32595;
assign w32597 = pi06224 & ~w21045;
assign w32598 = ~pi02706 & w21045;
assign w32599 = ~w32597 & ~w32598;
assign w32600 = pi06225 & ~w21045;
assign w32601 = ~pi02707 & w21045;
assign w32602 = ~w32600 & ~w32601;
assign w32603 = pi06226 & ~w21045;
assign w32604 = ~pi02160 & w21045;
assign w32605 = ~w32603 & ~w32604;
assign w32606 = pi06227 & ~w21045;
assign w32607 = ~pi02723 & w21045;
assign w32608 = ~w32606 & ~w32607;
assign w32609 = pi06228 & ~w21045;
assign w32610 = ~pi02708 & w21045;
assign w32611 = ~w32609 & ~w32610;
assign w32612 = pi06229 & ~w21045;
assign w32613 = ~pi02709 & w21045;
assign w32614 = ~w32612 & ~w32613;
assign w32615 = pi06230 & ~w21045;
assign w32616 = ~pi02710 & w21045;
assign w32617 = ~w32615 & ~w32616;
assign w32618 = pi06231 & ~w20806;
assign w32619 = ~pi02706 & w20806;
assign w32620 = ~w32618 & ~w32619;
assign w32621 = pi06232 & ~w20806;
assign w32622 = ~pi02707 & w20806;
assign w32623 = ~w32621 & ~w32622;
assign w32624 = pi06233 & ~w20806;
assign w32625 = ~pi02160 & w20806;
assign w32626 = ~w32624 & ~w32625;
assign w32627 = pi06234 & ~w20806;
assign w32628 = ~pi02708 & w20806;
assign w32629 = ~w32627 & ~w32628;
assign w32630 = pi06235 & ~w20806;
assign w32631 = ~pi02709 & w20806;
assign w32632 = ~w32630 & ~w32631;
assign w32633 = pi06236 & ~w20806;
assign w32634 = ~pi02710 & w20806;
assign w32635 = ~w32633 & ~w32634;
assign w32636 = pi06237 & ~w20860;
assign w32637 = ~pi02706 & w20860;
assign w32638 = ~w32636 & ~w32637;
assign w32639 = pi06238 & ~w20860;
assign w32640 = ~pi02707 & w20860;
assign w32641 = ~w32639 & ~w32640;
assign w32642 = pi06239 & ~w20860;
assign w32643 = ~pi02160 & w20860;
assign w32644 = ~w32642 & ~w32643;
assign w32645 = pi06240 & ~w20860;
assign w32646 = w17023 & w17671;
assign w32647 = ~w32645 & ~w32646;
assign w32648 = pi06241 & ~w20860;
assign w32649 = ~pi02708 & w20860;
assign w32650 = ~w32648 & ~w32649;
assign w32651 = pi06242 & ~w20860;
assign w32652 = w17023 & w18092;
assign w32653 = ~w32651 & ~w32652;
assign w32654 = pi06243 & ~w20860;
assign w32655 = ~pi02710 & w20860;
assign w32656 = ~w32654 & ~w32655;
assign w32657 = pi06244 & ~w20625;
assign w32658 = ~pi02706 & w20625;
assign w32659 = ~w32657 & ~w32658;
assign w32660 = pi06245 & ~w20625;
assign w32661 = ~pi02707 & w20625;
assign w32662 = ~w32660 & ~w32661;
assign w32663 = pi06246 & ~w20625;
assign w32664 = ~pi02160 & w20625;
assign w32665 = ~w32663 & ~w32664;
assign w32666 = pi06247 & ~w20625;
assign w32667 = ~pi02708 & w20625;
assign w32668 = ~w32666 & ~w32667;
assign w32669 = pi06248 & ~w20625;
assign w32670 = ~pi02709 & w20625;
assign w32671 = ~w32669 & ~w32670;
assign w32672 = pi06249 & ~w20625;
assign w32673 = ~pi02710 & w20625;
assign w32674 = ~w32672 & ~w32673;
assign w32675 = pi06250 & ~w20523;
assign w32676 = ~pi02706 & w20523;
assign w32677 = ~w32675 & ~w32676;
assign w32678 = pi06251 & ~w20249;
assign w32679 = ~pi02703 & w20249;
assign w32680 = ~w32678 & ~w32679;
assign w32681 = pi06252 & ~w20523;
assign w32682 = ~pi02707 & w20523;
assign w32683 = ~w32681 & ~w32682;
assign w32684 = pi06253 & ~w20523;
assign w32685 = ~pi02160 & w20523;
assign w32686 = ~w32684 & ~w32685;
assign w32687 = pi06254 & ~w20249;
assign w32688 = ~pi02721 & w20249;
assign w32689 = ~w32687 & ~w32688;
assign w32690 = pi06255 & ~w20249;
assign w32691 = ~pi02169 & w20249;
assign w32692 = ~w32690 & ~w32691;
assign w32693 = pi06256 & ~w20523;
assign w32694 = ~pi02723 & w20523;
assign w32695 = ~w32693 & ~w32694;
assign w32696 = pi06257 & ~w20523;
assign w32697 = ~pi02709 & w20523;
assign w32698 = ~w32696 & ~w32697;
assign w32699 = pi06258 & ~w20249;
assign w32700 = ~pi02718 & w20249;
assign w32701 = ~w32699 & ~w32700;
assign w32702 = pi06259 & ~w20523;
assign w32703 = ~pi02710 & w20523;
assign w32704 = ~w32702 & ~w32703;
assign w32705 = pi06260 & ~w20249;
assign w32706 = ~pi02167 & w20249;
assign w32707 = ~w32705 & ~w32706;
assign w32708 = pi06261 & ~w20527;
assign w32709 = ~pi02706 & w20527;
assign w32710 = ~w32708 & ~w32709;
assign w32711 = pi06262 & ~w20527;
assign w32712 = ~pi02707 & w20527;
assign w32713 = ~w32711 & ~w32712;
assign w32714 = pi06263 & ~w26184;
assign w32715 = ~pi02715 & w26184;
assign w32716 = ~w32714 & ~w32715;
assign w32717 = pi06264 & ~w20527;
assign w32718 = ~pi02160 & w20527;
assign w32719 = ~w32717 & ~w32718;
assign w32720 = pi06265 & ~w20527;
assign w32721 = ~pi02723 & w20527;
assign w32722 = ~w32720 & ~w32721;
assign w32723 = pi06266 & ~w20249;
assign w32724 = ~pi02722 & w20249;
assign w32725 = ~w32723 & ~w32724;
assign w32726 = pi06267 & ~w20527;
assign w32727 = ~pi02708 & w20527;
assign w32728 = ~w32726 & ~w32727;
assign w32729 = pi06268 & ~w20527;
assign w32730 = ~pi02709 & w20527;
assign w32731 = ~w32729 & ~w32730;
assign w32732 = pi06269 & ~w20527;
assign w32733 = ~pi02710 & w20527;
assign w32734 = ~w32732 & ~w32733;
assign w32735 = pi06270 & ~w20249;
assign w32736 = ~pi02719 & w20249;
assign w32737 = ~w32735 & ~w32736;
assign w32738 = pi06271 & ~w20318;
assign w32739 = w17114 & w17925;
assign w32740 = ~w32738 & ~w32739;
assign w32741 = pi06272 & ~w20299;
assign w32742 = ~pi02703 & w20299;
assign w32743 = ~w32741 & ~w32742;
assign w32744 = pi06273 & ~w20318;
assign w32745 = ~pi02707 & w20318;
assign w32746 = ~w32744 & ~w32745;
assign w32747 = pi06274 & ~w20299;
assign w32748 = ~pi02721 & w20299;
assign w32749 = ~w32747 & ~w32748;
assign w32750 = pi06275 & ~w20318;
assign w32751 = ~pi02723 & w20318;
assign w32752 = ~w32750 & ~w32751;
assign w32753 = pi06276 & ~w20318;
assign w32754 = ~pi02708 & w20318;
assign w32755 = ~w32753 & ~w32754;
assign w32756 = pi06277 & ~w20299;
assign w32757 = ~pi02169 & w20299;
assign w32758 = ~w32756 & ~w32757;
assign w32759 = pi06278 & ~w20318;
assign w32760 = w17114 & w18364;
assign w32761 = ~w32759 & ~w32760;
assign w32762 = pi06279 & ~w20299;
assign w32763 = ~pi02718 & w20299;
assign w32764 = ~w32762 & ~w32763;
assign w32765 = pi06280 & ~w20273;
assign w32766 = ~pi02705 & w20273;
assign w32767 = ~w32765 & ~w32766;
assign w32768 = pi06281 & ~w20299;
assign w32769 = ~pi02167 & w20299;
assign w32770 = ~w32768 & ~w32769;
assign w32771 = pi06282 & ~w20273;
assign w32772 = ~pi02706 & w20273;
assign w32773 = ~w32771 & ~w32772;
assign w32774 = pi06283 & ~w20273;
assign w32775 = ~pi02707 & w20273;
assign w32776 = ~w32774 & ~w32775;
assign w32777 = pi06284 & ~w20273;
assign w32778 = w17249 & w18234;
assign w32779 = ~w32777 & ~w32778;
assign w32780 = pi06285 & ~w20273;
assign w32781 = ~pi02723 & w20273;
assign w32782 = ~w32780 & ~w32781;
assign w32783 = pi06286 & ~w20299;
assign w32784 = ~pi02722 & w20299;
assign w32785 = ~w32783 & ~w32784;
assign w32786 = pi06287 & ~w20273;
assign w32787 = w17249 & w18092;
assign w32788 = ~w32786 & ~w32787;
assign w32789 = pi06288 & ~w20273;
assign w32790 = ~pi02710 & w20273;
assign w32791 = ~w32789 & ~w32790;
assign w32792 = pi06289 & ~w20299;
assign w32793 = ~pi02719 & w20299;
assign w32794 = ~w32792 & ~w32793;
assign w32795 = pi06290 & ~w18535;
assign w32796 = ~pi02706 & w18535;
assign w32797 = ~w32795 & ~w32796;
assign w32798 = pi06291 & ~w18637;
assign w32799 = ~pi02703 & w18637;
assign w32800 = ~w32798 & ~w32799;
assign w32801 = pi06292 & ~w18535;
assign w32802 = ~pi02707 & w18535;
assign w32803 = ~w32801 & ~w32802;
assign w32804 = pi06293 & ~w18535;
assign w32805 = ~pi02160 & w18535;
assign w32806 = ~w32804 & ~w32805;
assign w32807 = pi06294 & ~w18637;
assign w32808 = ~pi02721 & w18637;
assign w32809 = ~w32807 & ~w32808;
assign w32810 = pi06295 & ~w18535;
assign w32811 = ~pi02723 & w18535;
assign w32812 = ~w32810 & ~w32811;
assign w32813 = pi06296 & ~w18535;
assign w32814 = ~pi02708 & w18535;
assign w32815 = ~w32813 & ~w32814;
assign w32816 = pi06297 & ~w18535;
assign w32817 = ~pi02710 & w18535;
assign w32818 = ~w32816 & ~w32817;
assign w32819 = pi06298 & ~w18637;
assign w32820 = ~pi02169 & w18637;
assign w32821 = ~w32819 & ~w32820;
assign w32822 = pi06299 & ~w18637;
assign w32823 = w18636 & w19273;
assign w32824 = ~w32822 & ~w32823;
assign w32825 = pi06300 & ~w18637;
assign w32826 = ~pi02164 & w18637;
assign w32827 = ~w32825 & ~w32826;
assign w32828 = pi06301 & ~w18637;
assign w32829 = w17594 & w18636;
assign w32830 = ~w32828 & ~w32829;
assign w32831 = pi06302 & ~w18692;
assign w32832 = w17490 & w18578;
assign w32833 = ~w32831 & ~w32832;
assign w32834 = pi06303 & ~w18692;
assign w32835 = ~pi02707 & w18692;
assign w32836 = ~w32834 & ~w32835;
assign w32837 = pi06304 & ~w18692;
assign w32838 = ~pi02160 & w18692;
assign w32839 = ~w32837 & ~w32838;
assign w32840 = pi06305 & ~w18637;
assign w32841 = ~pi02722 & w18637;
assign w32842 = ~w32840 & ~w32841;
assign w32843 = pi06306 & ~w18692;
assign w32844 = ~pi02723 & w18692;
assign w32845 = ~w32843 & ~w32844;
assign w32846 = pi06307 & ~w18692;
assign w32847 = ~pi02708 & w18692;
assign w32848 = ~w32846 & ~w32847;
assign w32849 = pi06308 & ~w18692;
assign w32850 = w17490 & w18092;
assign w32851 = ~w32849 & ~w32850;
assign w32852 = pi06309 & ~w18692;
assign w32853 = w17490 & w18364;
assign w32854 = ~w32852 & ~w32853;
assign w32855 = pi06310 & ~w18646;
assign w32856 = ~pi02706 & w18646;
assign w32857 = ~w32855 & ~w32856;
assign w32858 = pi06311 & ~w18573;
assign w32859 = ~pi02703 & w18573;
assign w32860 = ~w32858 & ~w32859;
assign w32861 = pi06312 & ~w18646;
assign w32862 = ~pi02707 & w18646;
assign w32863 = ~w32861 & ~w32862;
assign w32864 = pi06313 & ~w18646;
assign w32865 = w17671 & w18645;
assign w32866 = ~w32864 & ~w32865;
assign w32867 = pi06314 & ~w18646;
assign w32868 = ~pi02708 & w18646;
assign w32869 = ~w32867 & ~w32868;
assign w32870 = pi06315 & ~w18646;
assign w32871 = ~pi02709 & w18646;
assign w32872 = ~w32870 & ~w32871;
assign w32873 = pi06316 & ~w21555;
assign w32874 = ~pi02703 & w21555;
assign w32875 = ~w32873 & ~w32874;
assign w32876 = pi06317 & ~w18646;
assign w32877 = ~pi02710 & w18646;
assign w32878 = ~w32876 & ~w32877;
assign w32879 = pi06318 & ~w18573;
assign w32880 = ~pi02169 & w18573;
assign w32881 = ~w32879 & ~w32880;
assign w32882 = pi06319 & ~w18573;
assign w32883 = w17586 & w18572;
assign w32884 = ~w32882 & ~w32883;
assign w32885 = pi06320 & ~w18573;
assign w32886 = ~pi02167 & w18573;
assign w32887 = ~w32885 & ~w32886;
assign w32888 = pi06321 & ~w18573;
assign w32889 = ~pi02164 & w18573;
assign w32890 = ~w32888 & ~w32889;
assign w32891 = pi06322 & ~w18573;
assign w32892 = w18572 & w19312;
assign w32893 = ~w32891 & ~w32892;
assign w32894 = pi06323 & ~w18573;
assign w32895 = ~pi02719 & w18573;
assign w32896 = ~w32894 & ~w32895;
assign w32897 = pi06324 & ~w18090;
assign w32898 = w17500 & w17925;
assign w32899 = ~w32897 & ~w32898;
assign w32900 = ~w16992 & w18808;
assign w32901 = pi06325 & ~w32900;
assign w32902 = ~pi02703 & w32900;
assign w32903 = ~w32901 & ~w32902;
assign w32904 = pi06326 & ~w18090;
assign w32905 = w17500 & w18067;
assign w32906 = ~w32904 & ~w32905;
assign w32907 = pi06327 & ~w32900;
assign w32908 = ~pi02721 & w32900;
assign w32909 = ~w32907 & ~w32908;
assign w32910 = pi06328 & ~w18090;
assign w32911 = w17500 & w17671;
assign w32912 = ~w32910 & ~w32911;
assign w32913 = pi06329 & ~w18090;
assign w32914 = w17500 & w18689;
assign w32915 = ~w32913 & ~w32914;
assign w32916 = pi06330 & ~w18090;
assign w32917 = w17500 & w18364;
assign w32918 = ~w32916 & ~w32917;
assign w32919 = pi06331 & ~w32900;
assign w32920 = ~pi02169 & w32900;
assign w32921 = ~w32919 & ~w32920;
assign w32922 = pi06332 & ~w32900;
assign w32923 = w17586 & w18808;
assign w32924 = ~w32922 & ~w32923;
assign w32925 = pi06333 & ~w32900;
assign w32926 = ~pi02167 & w32900;
assign w32927 = ~w32925 & ~w32926;
assign w32928 = pi06334 & ~w32900;
assign w32929 = ~pi02164 & w32900;
assign w32930 = ~w32928 & ~w32929;
assign w32931 = pi06335 & ~w32900;
assign w32932 = ~pi02719 & w32900;
assign w32933 = ~w32931 & ~w32932;
assign w32934 = pi06336 & ~w32900;
assign w32935 = ~pi02722 & w32900;
assign w32936 = ~w32934 & ~w32935;
assign w32937 = pi06337 & ~w18423;
assign w32938 = ~pi02706 & w18423;
assign w32939 = ~w32937 & ~w32938;
assign w32940 = pi06338 & ~w18423;
assign w32941 = ~pi02707 & w18423;
assign w32942 = ~w32940 & ~w32941;
assign w32943 = pi06339 & ~w18423;
assign w32944 = ~pi02160 & w18423;
assign w32945 = ~w32943 & ~w32944;
assign w32946 = pi06340 & ~w18423;
assign w32947 = ~pi02708 & w18423;
assign w32948 = ~w32946 & ~w32947;
assign w32949 = pi06341 & ~w18423;
assign w32950 = ~pi02709 & w18423;
assign w32951 = ~w32949 & ~w32950;
assign w32952 = pi06342 & ~w18423;
assign w32953 = ~pi02710 & w18423;
assign w32954 = ~w32952 & ~w32953;
assign w32955 = pi06343 & ~w18371;
assign w32956 = ~pi02706 & w18371;
assign w32957 = ~w32955 & ~w32956;
assign w32958 = pi06344 & ~w18371;
assign w32959 = ~pi02707 & w18371;
assign w32960 = ~w32958 & ~w32959;
assign w32961 = pi06345 & ~w18371;
assign w32962 = ~pi02160 & w18371;
assign w32963 = ~w32961 & ~w32962;
assign w32964 = pi06346 & ~w18371;
assign w32965 = ~pi02723 & w18371;
assign w32966 = ~w32964 & ~w32965;
assign w32967 = pi06347 & ~w18371;
assign w32968 = ~pi02708 & w18371;
assign w32969 = ~w32967 & ~w32968;
assign w32970 = pi06348 & ~w18371;
assign w32971 = ~pi02709 & w18371;
assign w32972 = ~w32970 & ~w32971;
assign w32973 = pi06349 & ~w18371;
assign w32974 = ~pi02710 & w18371;
assign w32975 = ~w32973 & ~w32974;
assign w32976 = pi06350 & ~w18222;
assign w32977 = w16999 & w17925;
assign w32978 = ~w32976 & ~w32977;
assign w32979 = pi06351 & ~w18222;
assign w32980 = ~pi02707 & w18222;
assign w32981 = ~w32979 & ~w32980;
assign w32982 = pi06352 & ~w18222;
assign w32983 = ~pi02160 & w18222;
assign w32984 = ~w32982 & ~w32983;
assign w32985 = pi06353 & ~w18222;
assign w32986 = ~pi02708 & w18222;
assign w32987 = ~w32985 & ~w32986;
assign w32988 = pi06354 & ~w18222;
assign w32989 = ~pi02709 & w18222;
assign w32990 = ~w32988 & ~w32989;
assign w32991 = pi06355 & ~w18222;
assign w32992 = ~pi02710 & w18222;
assign w32993 = ~w32991 & ~w32992;
assign w32994 = pi06356 & ~w18187;
assign w32995 = ~pi02721 & w18187;
assign w32996 = ~w32994 & ~w32995;
assign w32997 = pi06357 & ~w18187;
assign w32998 = ~pi02169 & w18187;
assign w32999 = ~w32997 & ~w32998;
assign w33000 = pi06358 & ~w17557;
assign w33001 = ~pi02705 & w17557;
assign w33002 = ~w33000 & ~w33001;
assign w33003 = pi06359 & ~w18187;
assign w33004 = ~pi02718 & w18187;
assign w33005 = ~w33003 & ~w33004;
assign w33006 = pi06360 & ~w17557;
assign w33007 = ~pi02706 & w17557;
assign w33008 = ~w33006 & ~w33007;
assign w33009 = pi06361 & ~w17557;
assign w33010 = ~pi02707 & w17557;
assign w33011 = ~w33009 & ~w33010;
assign w33012 = pi06362 & ~w18187;
assign w33013 = ~pi02167 & w18187;
assign w33014 = ~w33012 & ~w33013;
assign w33015 = pi06363 & ~w17557;
assign w33016 = w17556 & w17671;
assign w33017 = ~w33015 & ~w33016;
assign w33018 = pi06364 & ~w17557;
assign w33019 = ~pi02708 & w17557;
assign w33020 = ~w33018 & ~w33019;
assign w33021 = pi06365 & ~w17557;
assign w33022 = ~pi02709 & w17557;
assign w33023 = ~w33021 & ~w33022;
assign w33024 = pi06366 & ~w18187;
assign w33025 = ~pi02722 & w18187;
assign w33026 = ~w33024 & ~w33025;
assign w33027 = pi06367 & ~w18187;
assign w33028 = ~pi02164 & w18187;
assign w33029 = ~w33027 & ~w33028;
assign w33030 = pi06368 & ~w18187;
assign w33031 = ~pi02719 & w18187;
assign w33032 = ~w33030 & ~w33031;
assign w33033 = pi06369 & ~w17900;
assign w33034 = ~pi02721 & w17900;
assign w33035 = ~w33033 & ~w33034;
assign w33036 = pi06370 & ~w17856;
assign w33037 = w17855 & w18578;
assign w33038 = ~w33036 & ~w33037;
assign w33039 = pi06371 & ~w17900;
assign w33040 = ~pi02169 & w17900;
assign w33041 = ~w33039 & ~w33040;
assign w33042 = pi06372 & ~w17856;
assign w33043 = ~pi02706 & w17856;
assign w33044 = ~w33042 & ~w33043;
assign w33045 = pi06373 & ~w17856;
assign w33046 = ~pi02707 & w17856;
assign w33047 = ~w33045 & ~w33046;
assign w33048 = pi06374 & ~w17900;
assign w33049 = ~pi02718 & w17900;
assign w33050 = ~w33048 & ~w33049;
assign w33051 = pi06375 & ~w17900;
assign w33052 = w17084 & w19273;
assign w33053 = ~w33051 & ~w33052;
assign w33054 = pi06376 & ~w17856;
assign w33055 = ~pi02723 & w17856;
assign w33056 = ~w33054 & ~w33055;
assign w33057 = pi06377 & ~w17900;
assign w33058 = w17084 & w17620;
assign w33059 = ~w33057 & ~w33058;
assign w33060 = pi06378 & ~w17856;
assign w33061 = ~pi02708 & w17856;
assign w33062 = ~w33060 & ~w33061;
assign w33063 = pi06379 & ~w17856;
assign w33064 = ~pi02710 & w17856;
assign w33065 = ~w33063 & ~w33064;
assign w33066 = pi06380 & ~w17900;
assign w33067 = ~pi02722 & w17900;
assign w33068 = ~w33066 & ~w33067;
assign w33069 = pi06381 & ~w17900;
assign w33070 = ~pi02719 & w17900;
assign w33071 = ~w33069 & ~w33070;
assign w33072 = pi06382 & ~w17848;
assign w33073 = ~pi02721 & w17848;
assign w33074 = ~w33072 & ~w33073;
assign w33075 = pi06383 & ~w17848;
assign w33076 = ~pi02169 & w17848;
assign w33077 = ~w33075 & ~w33076;
assign w33078 = pi06384 & ~w17848;
assign w33079 = w16970 & w17586;
assign w33080 = ~w33078 & ~w33079;
assign w33081 = pi06385 & ~w17848;
assign w33082 = ~pi02164 & w17848;
assign w33083 = ~w33081 & ~w33082;
assign w33084 = pi06386 & ~w17848;
assign w33085 = ~pi02167 & w17848;
assign w33086 = ~w33084 & ~w33085;
assign w33087 = pi06387 & ~w17848;
assign w33088 = ~pi02722 & w17848;
assign w33089 = ~w33087 & ~w33088;
assign w33090 = pi06388 & ~w17827;
assign w33091 = ~pi02705 & w17827;
assign w33092 = ~w33090 & ~w33091;
assign w33093 = pi06389 & ~w17848;
assign w33094 = ~pi02719 & w17848;
assign w33095 = ~w33093 & ~w33094;
assign w33096 = pi06390 & ~w17827;
assign w33097 = ~pi02707 & w17827;
assign w33098 = ~w33096 & ~w33097;
assign w33099 = pi06391 & ~w17827;
assign w33100 = ~pi02160 & w17827;
assign w33101 = ~w33099 & ~w33100;
assign w33102 = pi06392 & ~w17827;
assign w33103 = w17461 & w17671;
assign w33104 = ~w33102 & ~w33103;
assign w33105 = pi06393 & ~w17827;
assign w33106 = ~pi02708 & w17827;
assign w33107 = ~w33105 & ~w33106;
assign w33108 = pi06394 & ~w17827;
assign w33109 = ~pi02709 & w17827;
assign w33110 = ~w33108 & ~w33109;
assign w33111 = pi06395 & ~w17827;
assign w33112 = ~pi02710 & w17827;
assign w33113 = ~w33111 & ~w33112;
assign w33114 = pi06396 & ~w17809;
assign w33115 = ~pi02169 & w17809;
assign w33116 = ~w33114 & ~w33115;
assign w33117 = pi06397 & ~w17809;
assign w33118 = ~pi02718 & w17809;
assign w33119 = ~w33117 & ~w33118;
assign w33120 = pi06398 & ~w17809;
assign w33121 = ~pi02167 & w17809;
assign w33122 = ~w33120 & ~w33121;
assign w33123 = pi06399 & ~w17809;
assign w33124 = w17620 & w17808;
assign w33125 = ~w33123 & ~w33124;
assign w33126 = pi06400 & ~w17809;
assign w33127 = ~pi02722 & w17809;
assign w33128 = ~w33126 & ~w33127;
assign w33129 = pi06401 & ~w17809;
assign w33130 = ~pi02719 & w17809;
assign w33131 = ~w33129 & ~w33130;
assign w33132 = pi06402 & ~w17706;
assign w33133 = w17119 & w17925;
assign w33134 = ~w33132 & ~w33133;
assign w33135 = pi06403 & ~w17706;
assign w33136 = ~pi02707 & w17706;
assign w33137 = ~w33135 & ~w33136;
assign w33138 = pi06404 & ~w17706;
assign w33139 = w17119 & w18234;
assign w33140 = ~w33138 & ~w33139;
assign w33141 = pi06405 & ~w17706;
assign w33142 = ~pi02708 & w17706;
assign w33143 = ~w33141 & ~w33142;
assign w33144 = pi06406 & ~w17706;
assign w33145 = ~pi02709 & w17706;
assign w33146 = ~w33144 & ~w33145;
assign w33147 = pi06407 & ~w17706;
assign w33148 = w17119 & w18364;
assign w33149 = ~w33147 & ~w33148;
assign w33150 = pi06408 & ~w17391;
assign w33151 = ~pi02703 & w17391;
assign w33152 = ~w33150 & ~w33151;
assign w33153 = pi06409 & ~w17391;
assign w33154 = ~pi02169 & w17391;
assign w33155 = ~w33153 & ~w33154;
assign w33156 = pi06410 & ~w17391;
assign w33157 = ~pi02718 & w17391;
assign w33158 = ~w33156 & ~w33157;
assign w33159 = pi06411 & ~w17391;
assign w33160 = ~pi02167 & w17391;
assign w33161 = ~w33159 & ~w33160;
assign w33162 = pi06412 & ~w17391;
assign w33163 = ~pi02164 & w17391;
assign w33164 = ~w33162 & ~w33163;
assign w33165 = pi06413 & ~w17391;
assign w33166 = ~pi02722 & w17391;
assign w33167 = ~w33165 & ~w33166;
assign w33168 = pi06414 & ~w17391;
assign w33169 = w17390 & w17594;
assign w33170 = ~w33168 & ~w33169;
assign w33171 = pi06415 & ~w16923;
assign w33172 = ~pi02706 & w16923;
assign w33173 = ~w33171 & ~w33172;
assign w33174 = pi06416 & ~w16923;
assign w33175 = ~pi02707 & w16923;
assign w33176 = ~w33174 & ~w33175;
assign w33177 = pi06417 & ~w16923;
assign w33178 = ~pi02160 & w16923;
assign w33179 = ~w33177 & ~w33178;
assign w33180 = pi06418 & ~w16923;
assign w33181 = ~pi02708 & w16923;
assign w33182 = ~w33180 & ~w33181;
assign w33183 = pi06419 & ~w16923;
assign w33184 = w16922 & w18092;
assign w33185 = ~w33183 & ~w33184;
assign w33186 = ~w16992 & w17495;
assign w33187 = pi06420 & ~w33186;
assign w33188 = ~pi02703 & w33186;
assign w33189 = ~w33187 & ~w33188;
assign w33190 = ~w16905 & w17239;
assign w33191 = pi06421 & ~w33190;
assign w33192 = ~pi02716 & w33190;
assign w33193 = ~w33191 & ~w33192;
assign w33194 = ~w16892 & w17226;
assign w33195 = pi06422 & ~w33194;
assign w33196 = ~pi02705 & w33194;
assign w33197 = ~w33195 & ~w33196;
assign w33198 = pi06423 & ~w33186;
assign w33199 = ~pi02721 & w33186;
assign w33200 = ~w33198 & ~w33199;
assign w33201 = pi06424 & ~w33194;
assign w33202 = ~pi02706 & w33194;
assign w33203 = ~w33201 & ~w33202;
assign w33204 = pi06425 & ~w33194;
assign w33205 = ~pi02707 & w33194;
assign w33206 = ~w33204 & ~w33205;
assign w33207 = pi06426 & ~w33186;
assign w33208 = ~pi02169 & w33186;
assign w33209 = ~w33207 & ~w33208;
assign w33210 = pi06427 & ~w33194;
assign w33211 = ~pi02160 & w33194;
assign w33212 = ~w33210 & ~w33211;
assign w33213 = pi06428 & ~w33194;
assign w33214 = ~pi02723 & w33194;
assign w33215 = ~w33213 & ~w33214;
assign w33216 = pi06429 & ~w33194;
assign w33217 = ~pi02708 & w33194;
assign w33218 = ~w33216 & ~w33217;
assign w33219 = pi06430 & ~w33194;
assign w33220 = ~pi02709 & w33194;
assign w33221 = ~w33219 & ~w33220;
assign w33222 = pi06431 & ~w33186;
assign w33223 = ~pi02167 & w33186;
assign w33224 = ~w33222 & ~w33223;
assign w33225 = pi06432 & ~w33186;
assign w33226 = w17495 & w17620;
assign w33227 = ~w33225 & ~w33226;
assign w33228 = ~w16892 & w17259;
assign w33229 = pi06433 & ~w33228;
assign w33230 = ~pi02705 & w33228;
assign w33231 = ~w33229 & ~w33230;
assign w33232 = pi06434 & ~w33228;
assign w33233 = ~pi02706 & w33228;
assign w33234 = ~w33232 & ~w33233;
assign w33235 = pi06435 & ~w33228;
assign w33236 = ~pi02707 & w33228;
assign w33237 = ~w33235 & ~w33236;
assign w33238 = pi06436 & ~w33228;
assign w33239 = ~pi02160 & w33228;
assign w33240 = ~w33238 & ~w33239;
assign w33241 = pi06437 & ~w33186;
assign w33242 = ~pi02719 & w33186;
assign w33243 = ~w33241 & ~w33242;
assign w33244 = pi06438 & ~w33228;
assign w33245 = ~pi02723 & w33228;
assign w33246 = ~w33244 & ~w33245;
assign w33247 = pi06439 & ~w33228;
assign w33248 = ~pi02708 & w33228;
assign w33249 = ~w33247 & ~w33248;
assign w33250 = pi06440 & ~w33228;
assign w33251 = ~pi02709 & w33228;
assign w33252 = ~w33250 & ~w33251;
assign w33253 = pi06441 & ~w33228;
assign w33254 = ~pi02710 & w33228;
assign w33255 = ~w33253 & ~w33254;
assign w33256 = ~w16892 & w17762;
assign w33257 = pi06442 & ~w33256;
assign w33258 = w17762 & w17925;
assign w33259 = ~w33257 & ~w33258;
assign w33260 = pi06443 & ~w33256;
assign w33261 = ~pi02707 & w33256;
assign w33262 = ~w33260 & ~w33261;
assign w33263 = pi06444 & ~w33256;
assign w33264 = ~pi02160 & w33256;
assign w33265 = ~w33263 & ~w33264;
assign w33266 = pi06445 & ~w33256;
assign w33267 = w17762 & w18689;
assign w33268 = ~w33266 & ~w33267;
assign w33269 = pi06446 & ~w33256;
assign w33270 = ~pi02709 & w33256;
assign w33271 = ~w33269 & ~w33270;
assign w33272 = pi06447 & ~w33256;
assign w33273 = ~pi02710 & w33256;
assign w33274 = ~w33272 & ~w33273;
assign w33275 = ~w16892 & w17535;
assign w33276 = pi06448 & ~w33275;
assign w33277 = ~pi02706 & w33275;
assign w33278 = ~w33276 & ~w33277;
assign w33279 = pi06449 & ~w33275;
assign w33280 = ~pi02707 & w33275;
assign w33281 = ~w33279 & ~w33280;
assign w33282 = pi06450 & ~w33275;
assign w33283 = ~pi02160 & w33275;
assign w33284 = ~w33282 & ~w33283;
assign w33285 = pi06451 & ~w33275;
assign w33286 = w17535 & w17671;
assign w33287 = ~w33285 & ~w33286;
assign w33288 = pi06452 & ~w33275;
assign w33289 = ~pi02708 & w33275;
assign w33290 = ~w33288 & ~w33289;
assign w33291 = pi06453 & ~w33275;
assign w33292 = w17535 & w18092;
assign w33293 = ~w33291 & ~w33292;
assign w33294 = pi06454 & ~w33275;
assign w33295 = ~pi02710 & w33275;
assign w33296 = ~w33294 & ~w33295;
assign w33297 = ~w16992 & w17450;
assign w33298 = pi06455 & ~w33297;
assign w33299 = ~pi02721 & w33297;
assign w33300 = ~w33298 & ~w33299;
assign w33301 = pi06456 & ~w33297;
assign w33302 = ~pi02169 & w33297;
assign w33303 = ~w33301 & ~w33302;
assign w33304 = pi06457 & ~w33297;
assign w33305 = w17450 & w17586;
assign w33306 = ~w33304 & ~w33305;
assign w33307 = pi06458 & ~w21500;
assign w33308 = ~pi02705 & w21500;
assign w33309 = ~w33307 & ~w33308;
assign w33310 = pi06459 & ~w21500;
assign w33311 = ~pi02706 & w21500;
assign w33312 = ~w33310 & ~w33311;
assign w33313 = pi06460 & ~w33297;
assign w33314 = ~pi02164 & w33297;
assign w33315 = ~w33313 & ~w33314;
assign w33316 = pi06461 & ~w33297;
assign w33317 = ~pi02722 & w33297;
assign w33318 = ~w33316 & ~w33317;
assign w33319 = pi06462 & ~w21500;
assign w33320 = ~pi02160 & w21500;
assign w33321 = ~w33319 & ~w33320;
assign w33322 = pi06463 & ~w33297;
assign w33323 = ~pi02719 & w33297;
assign w33324 = ~w33322 & ~w33323;
assign w33325 = pi06464 & ~w21500;
assign w33326 = ~pi02723 & w21500;
assign w33327 = ~w33325 & ~w33326;
assign w33328 = pi06465 & ~w21500;
assign w33329 = ~pi02708 & w21500;
assign w33330 = ~w33328 & ~w33329;
assign w33331 = pi06466 & ~w21500;
assign w33332 = ~pi02709 & w21500;
assign w33333 = ~w33331 & ~w33332;
assign w33334 = ~w16992 & w17436;
assign w33335 = pi06467 & ~w33334;
assign w33336 = ~pi02703 & w33334;
assign w33337 = ~w33335 & ~w33336;
assign w33338 = pi06468 & ~w33334;
assign w33339 = ~pi02721 & w33334;
assign w33340 = ~w33338 & ~w33339;
assign w33341 = pi06469 & ~w21407;
assign w33342 = ~pi02711 & w21407;
assign w33343 = ~w33341 & ~w33342;
assign w33344 = pi06470 & ~w21407;
assign w33345 = ~pi02712 & w21407;
assign w33346 = ~w33344 & ~w33345;
assign w33347 = pi06471 & ~w33334;
assign w33348 = ~pi02169 & w33334;
assign w33349 = ~w33347 & ~w33348;
assign w33350 = pi06472 & ~w21407;
assign w33351 = ~pi02713 & w21407;
assign w33352 = ~w33350 & ~w33351;
assign w33353 = pi06473 & ~w33334;
assign w33354 = ~pi02718 & w33334;
assign w33355 = ~w33353 & ~w33354;
assign w33356 = pi06474 & ~w21929;
assign w33357 = w17375 & w19273;
assign w33358 = ~w33356 & ~w33357;
assign w33359 = pi06475 & ~w21407;
assign w33360 = ~pi02715 & w21407;
assign w33361 = ~w33359 & ~w33360;
assign w33362 = pi06476 & ~w33334;
assign w33363 = ~pi02167 & w33334;
assign w33364 = ~w33362 & ~w33363;
assign w33365 = pi06477 & ~w21407;
assign w33366 = ~pi02716 & w21407;
assign w33367 = ~w33365 & ~w33366;
assign w33368 = pi06478 & ~w21407;
assign w33369 = ~pi02717 & w21407;
assign w33370 = ~w33368 & ~w33369;
assign w33371 = pi06479 & ~w20895;
assign w33372 = w17603 & w18745;
assign w33373 = ~w33371 & ~w33372;
assign w33374 = pi06480 & ~w33334;
assign w33375 = ~pi02164 & w33334;
assign w33376 = ~w33374 & ~w33375;
assign w33377 = pi06481 & ~w20895;
assign w33378 = ~pi02712 & w20895;
assign w33379 = ~w33377 & ~w33378;
assign w33380 = pi06482 & ~w33334;
assign w33381 = ~pi02722 & w33334;
assign w33382 = ~w33380 & ~w33381;
assign w33383 = pi06483 & ~w20895;
assign w33384 = ~pi02713 & w20895;
assign w33385 = ~w33383 & ~w33384;
assign w33386 = pi06484 & ~w20895;
assign w33387 = w17742 & w18745;
assign w33388 = ~w33386 & ~w33387;
assign w33389 = pi06485 & ~w20895;
assign w33390 = w17317 & w18745;
assign w33391 = ~w33389 & ~w33390;
assign w33392 = pi06486 & ~w33334;
assign w33393 = w17436 & w17594;
assign w33394 = ~w33392 & ~w33393;
assign w33395 = pi06487 & ~w20895;
assign w33396 = w16973 & w18745;
assign w33397 = ~w33395 & ~w33396;
assign w33398 = pi06488 & ~w20871;
assign w33399 = ~pi02712 & w20871;
assign w33400 = ~w33398 & ~w33399;
assign w33401 = pi06489 & ~w20871;
assign w33402 = ~pi02170 & w20871;
assign w33403 = ~w33401 & ~w33402;
assign w33404 = pi06490 & ~w20871;
assign w33405 = ~pi02713 & w20871;
assign w33406 = ~w33404 & ~w33405;
assign w33407 = pi06491 & ~w20871;
assign w33408 = ~pi02714 & w20871;
assign w33409 = ~w33407 & ~w33408;
assign w33410 = pi06492 & ~w20871;
assign w33411 = ~pi02715 & w20871;
assign w33412 = ~w33410 & ~w33411;
assign w33413 = pi06493 & ~w20871;
assign w33414 = ~pi02716 & w20871;
assign w33415 = ~w33413 & ~w33414;
assign w33416 = pi06494 & ~w20871;
assign w33417 = w16973 & w17977;
assign w33418 = ~w33416 & ~w33417;
assign w33419 = pi06495 & ~w20493;
assign w33420 = w17020 & w18027;
assign w33421 = ~w33419 & ~w33420;
assign w33422 = pi06496 & ~w20493;
assign w33423 = ~pi02170 & w20493;
assign w33424 = ~w33422 & ~w33423;
assign w33425 = pi06497 & ~w20493;
assign w33426 = ~pi02713 & w20493;
assign w33427 = ~w33425 & ~w33426;
assign w33428 = pi06498 & ~w20493;
assign w33429 = ~pi02715 & w20493;
assign w33430 = ~w33428 & ~w33429;
assign w33431 = pi06499 & ~w20493;
assign w33432 = w17317 & w18027;
assign w33433 = ~w33431 & ~w33432;
assign w33434 = w16978 & ~w16992;
assign w33435 = pi06500 & ~w33434;
assign w33436 = ~pi02703 & w33434;
assign w33437 = ~w33435 & ~w33436;
assign w33438 = pi06501 & ~w33434;
assign w33439 = ~pi02721 & w33434;
assign w33440 = ~w33438 & ~w33439;
assign w33441 = pi06502 & ~w33434;
assign w33442 = w16978 & w19797;
assign w33443 = ~w33441 & ~w33442;
assign w33444 = pi06503 & ~w33434;
assign w33445 = ~pi02718 & w33434;
assign w33446 = ~w33444 & ~w33445;
assign w33447 = pi06504 & ~w33434;
assign w33448 = ~pi02167 & w33434;
assign w33449 = ~w33447 & ~w33448;
assign w33450 = pi06505 & ~w33434;
assign w33451 = ~pi02164 & w33434;
assign w33452 = ~w33450 & ~w33451;
assign w33453 = pi06506 & ~w33434;
assign w33454 = ~pi02722 & w33434;
assign w33455 = ~w33453 & ~w33454;
assign w33456 = pi06507 & ~w33434;
assign w33457 = ~pi02719 & w33434;
assign w33458 = ~w33456 & ~w33457;
assign w33459 = pi06508 & ~w20306;
assign w33460 = ~pi02712 & w20306;
assign w33461 = ~w33459 & ~w33460;
assign w33462 = pi06509 & ~w20306;
assign w33463 = w17996 & w20209;
assign w33464 = ~w33462 & ~w33463;
assign w33465 = pi06510 & ~w20306;
assign w33466 = w17929 & w17996;
assign w33467 = ~w33465 & ~w33466;
assign w33468 = pi06511 & ~w20306;
assign w33469 = ~pi02715 & w20306;
assign w33470 = ~w33468 & ~w33469;
assign w33471 = pi06512 & ~w20306;
assign w33472 = w17317 & w17996;
assign w33473 = ~w33471 & ~w33472;
assign w33474 = pi06513 & ~w20306;
assign w33475 = w16973 & w17996;
assign w33476 = ~w33474 & ~w33475;
assign w33477 = pi06514 & ~w20230;
assign w33478 = w17231 & w17603;
assign w33479 = ~w33477 & ~w33478;
assign w33480 = pi06515 & ~w20230;
assign w33481 = ~pi02712 & w20230;
assign w33482 = ~w33480 & ~w33481;
assign w33483 = pi06516 & ~w20257;
assign w33484 = ~pi02721 & w20257;
assign w33485 = ~w33483 & ~w33484;
assign w33486 = pi06517 & ~w20230;
assign w33487 = w17231 & w20209;
assign w33488 = ~w33486 & ~w33487;
assign w33489 = pi06518 & ~w20230;
assign w33490 = ~pi02713 & w20230;
assign w33491 = ~w33489 & ~w33490;
assign w33492 = pi06519 & ~w20257;
assign w33493 = ~pi02169 & w20257;
assign w33494 = ~w33492 & ~w33493;
assign w33495 = pi06520 & ~w20230;
assign w33496 = w17231 & w17742;
assign w33497 = ~w33495 & ~w33496;
assign w33498 = pi06521 & ~w20257;
assign w33499 = ~pi02718 & w20257;
assign w33500 = ~w33498 & ~w33499;
assign w33501 = pi06522 & ~w20230;
assign w33502 = ~pi02716 & w20230;
assign w33503 = ~w33501 & ~w33502;
assign w33504 = pi06523 & ~w20230;
assign w33505 = w16973 & w17231;
assign w33506 = ~w33504 & ~w33505;
assign w33507 = pi06524 & ~w20257;
assign w33508 = ~pi02167 & w20257;
assign w33509 = ~w33507 & ~w33508;
assign w33510 = pi06525 & ~w20068;
assign w33511 = ~pi02712 & w20068;
assign w33512 = ~w33510 & ~w33511;
assign w33513 = pi06526 & ~w20068;
assign w33514 = ~pi02170 & w20068;
assign w33515 = ~w33513 & ~w33514;
assign w33516 = pi06527 & ~w20068;
assign w33517 = ~pi02713 & w20068;
assign w33518 = ~w33516 & ~w33517;
assign w33519 = pi06528 & ~w20257;
assign w33520 = ~pi02722 & w20257;
assign w33521 = ~w33519 & ~w33520;
assign w33522 = pi06529 & ~w20068;
assign w33523 = ~pi02714 & w20068;
assign w33524 = ~w33522 & ~w33523;
assign w33525 = pi06530 & ~w20257;
assign w33526 = ~pi02719 & w20257;
assign w33527 = ~w33525 & ~w33526;
assign w33528 = pi06531 & ~w20068;
assign w33529 = ~pi02715 & w20068;
assign w33530 = ~w33528 & ~w33529;
assign w33531 = pi06532 & ~w20068;
assign w33532 = ~pi02716 & w20068;
assign w33533 = ~w33531 & ~w33532;
assign w33534 = pi06533 & ~w18675;
assign w33535 = w17284 & w17532;
assign w33536 = ~w33534 & ~w33535;
assign w33537 = pi06534 & ~w18918;
assign w33538 = w17385 & w17603;
assign w33539 = ~w33537 & ~w33538;
assign w33540 = pi06535 & ~w18918;
assign w33541 = ~pi02712 & w18918;
assign w33542 = ~w33540 & ~w33541;
assign w33543 = pi06536 & ~w18675;
assign w33544 = ~pi02721 & w18675;
assign w33545 = ~w33543 & ~w33544;
assign w33546 = pi06537 & ~w18918;
assign w33547 = w17385 & w17929;
assign w33548 = ~w33546 & ~w33547;
assign w33549 = pi06538 & ~w18675;
assign w33550 = ~pi02169 & w18675;
assign w33551 = ~w33549 & ~w33550;
assign w33552 = pi06539 & ~w18918;
assign w33553 = ~pi02714 & w18918;
assign w33554 = ~w33552 & ~w33553;
assign w33555 = pi06540 & ~w18675;
assign w33556 = ~pi02718 & w18675;
assign w33557 = ~w33555 & ~w33556;
assign w33558 = pi06541 & ~w18918;
assign w33559 = ~pi02716 & w18918;
assign w33560 = ~w33558 & ~w33559;
assign w33561 = pi06542 & ~w18918;
assign w33562 = ~pi02717 & w18918;
assign w33563 = ~w33561 & ~w33562;
assign w33564 = pi06543 & ~w18671;
assign w33565 = ~pi02711 & w18671;
assign w33566 = ~w33564 & ~w33565;
assign w33567 = pi06544 & ~w18675;
assign w33568 = ~pi02167 & w18675;
assign w33569 = ~w33567 & ~w33568;
assign w33570 = pi06545 & ~w18671;
assign w33571 = w17020 & w17349;
assign w33572 = ~w33570 & ~w33571;
assign w33573 = pi06546 & ~w18671;
assign w33574 = ~pi02170 & w18671;
assign w33575 = ~w33573 & ~w33574;
assign w33576 = pi06547 & ~w18671;
assign w33577 = ~pi02713 & w18671;
assign w33578 = ~w33576 & ~w33577;
assign w33579 = pi06548 & ~w18671;
assign w33580 = ~pi02714 & w18671;
assign w33581 = ~w33579 & ~w33580;
assign w33582 = pi06549 & ~w18675;
assign w33583 = ~pi02722 & w18675;
assign w33584 = ~w33582 & ~w33583;
assign w33585 = pi06550 & ~w18675;
assign w33586 = ~pi02719 & w18675;
assign w33587 = ~w33585 & ~w33586;
assign w33588 = pi06551 & ~w18671;
assign w33589 = ~pi02716 & w18671;
assign w33590 = ~w33588 & ~w33589;
assign w33591 = pi06552 & ~w18671;
assign w33592 = ~pi02717 & w18671;
assign w33593 = ~w33591 & ~w33592;
assign w33594 = pi06553 & ~w18581;
assign w33595 = ~pi02703 & w18581;
assign w33596 = ~w33594 & ~w33595;
assign w33597 = pi06554 & ~w18597;
assign w33598 = ~pi02712 & w18597;
assign w33599 = ~w33597 & ~w33598;
assign w33600 = pi06555 & ~w18581;
assign w33601 = ~pi02721 & w18581;
assign w33602 = ~w33600 & ~w33601;
assign w33603 = pi06556 & ~w18597;
assign w33604 = ~pi02170 & w18597;
assign w33605 = ~w33603 & ~w33604;
assign w33606 = pi06557 & ~w18597;
assign w33607 = ~pi02713 & w18597;
assign w33608 = ~w33606 & ~w33607;
assign w33609 = pi06558 & ~w18581;
assign w33610 = ~pi02169 & w18581;
assign w33611 = ~w33609 & ~w33610;
assign w33612 = pi06559 & ~w18597;
assign w33613 = w17210 & w17742;
assign w33614 = ~w33612 & ~w33613;
assign w33615 = pi06560 & ~w18597;
assign w33616 = w17210 & w17317;
assign w33617 = ~w33615 & ~w33616;
assign w33618 = pi06561 & ~w18581;
assign w33619 = ~pi02718 & w18581;
assign w33620 = ~w33618 & ~w33619;
assign w33621 = pi06562 & ~w18597;
assign w33622 = ~pi02717 & w18597;
assign w33623 = ~w33621 & ~w33622;
assign w33624 = pi06563 & ~w18581;
assign w33625 = w17177 & w17620;
assign w33626 = ~w33624 & ~w33625;
assign w33627 = pi06564 & ~w18581;
assign w33628 = ~pi02722 & w18581;
assign w33629 = ~w33627 & ~w33628;
assign w33630 = pi06565 & ~w18581;
assign w33631 = ~pi02719 & w18581;
assign w33632 = ~w33630 & ~w33631;
assign w33633 = pi06566 & ~w16942;
assign w33634 = ~pi02712 & w16942;
assign w33635 = ~w33633 & ~w33634;
assign w33636 = pi06567 & ~w16942;
assign w33637 = w16941 & w20209;
assign w33638 = ~w33636 & ~w33637;
assign w33639 = pi06568 & ~w16942;
assign w33640 = ~pi02713 & w16942;
assign w33641 = ~w33639 & ~w33640;
assign w33642 = pi06569 & ~w16942;
assign w33643 = ~pi02714 & w16942;
assign w33644 = ~w33642 & ~w33643;
assign w33645 = pi06570 & ~w16942;
assign w33646 = ~pi02715 & w16942;
assign w33647 = ~w33645 & ~w33646;
assign w33648 = pi06571 & ~w16942;
assign w33649 = w16941 & w17317;
assign w33650 = ~w33648 & ~w33649;
assign w33651 = pi06572 & ~w16942;
assign w33652 = ~pi02717 & w16942;
assign w33653 = ~w33651 & ~w33652;
assign w33654 = pi06573 & ~w18330;
assign w33655 = w17811 & w18177;
assign w33656 = ~w33654 & ~w33655;
assign w33657 = pi06574 & ~w18330;
assign w33658 = ~pi02169 & w18330;
assign w33659 = ~w33657 & ~w33658;
assign w33660 = pi06575 & ~w18330;
assign w33661 = ~pi02718 & w18330;
assign w33662 = ~w33660 & ~w33661;
assign w33663 = pi06576 & ~w18330;
assign w33664 = ~pi02167 & w18330;
assign w33665 = ~w33663 & ~w33664;
assign w33666 = pi06577 & ~w18279;
assign w33667 = ~pi02712 & w18279;
assign w33668 = ~w33666 & ~w33667;
assign w33669 = pi06578 & ~w18279;
assign w33670 = ~pi02170 & w18279;
assign w33671 = ~w33669 & ~w33670;
assign w33672 = pi06579 & ~w18279;
assign w33673 = w17929 & w18278;
assign w33674 = ~w33672 & ~w33673;
assign w33675 = pi06580 & ~w18279;
assign w33676 = ~pi02714 & w18279;
assign w33677 = ~w33675 & ~w33676;
assign w33678 = pi06581 & ~w18330;
assign w33679 = ~pi02722 & w18330;
assign w33680 = ~w33678 & ~w33679;
assign w33681 = pi06582 & ~w18279;
assign w33682 = w18059 & w18278;
assign w33683 = ~w33681 & ~w33682;
assign w33684 = pi06583 & ~w18279;
assign w33685 = ~pi02716 & w18279;
assign w33686 = ~w33684 & ~w33685;
assign w33687 = pi06584 & ~w18330;
assign w33688 = w17594 & w18177;
assign w33689 = ~w33687 & ~w33688;
assign w33690 = pi06585 & ~w18279;
assign w33691 = ~pi02717 & w18279;
assign w33692 = ~w33690 & ~w33691;
assign w33693 = pi06586 & ~w18002;
assign w33694 = ~pi02712 & w18002;
assign w33695 = ~w33693 & ~w33694;
assign w33696 = pi06587 & ~w17566;
assign w33697 = ~pi02703 & w17566;
assign w33698 = ~w33696 & ~w33697;
assign w33699 = pi06588 & ~w18002;
assign w33700 = ~pi02170 & w18002;
assign w33701 = ~w33699 & ~w33700;
assign w33702 = pi06589 & ~w17566;
assign w33703 = ~pi02721 & w17566;
assign w33704 = ~w33702 & ~w33703;
assign w33705 = pi06590 & ~w18002;
assign w33706 = ~pi02714 & w18002;
assign w33707 = ~w33705 & ~w33706;
assign w33708 = pi06591 & ~w18002;
assign w33709 = ~pi02715 & w18002;
assign w33710 = ~w33708 & ~w33709;
assign w33711 = pi06592 & ~w18002;
assign w33712 = ~pi02716 & w18002;
assign w33713 = ~w33711 & ~w33712;
assign w33714 = pi06593 & ~w18002;
assign w33715 = ~pi02717 & w18002;
assign w33716 = ~w33714 & ~w33715;
assign w33717 = pi06594 & ~w17838;
assign w33718 = ~pi02711 & w17838;
assign w33719 = ~w33717 & ~w33718;
assign w33720 = pi06595 & ~w17566;
assign w33721 = ~pi02718 & w17566;
assign w33722 = ~w33720 & ~w33721;
assign w33723 = pi06596 & ~w17838;
assign w33724 = ~pi02712 & w17838;
assign w33725 = ~w33723 & ~w33724;
assign w33726 = pi06597 & ~w17566;
assign w33727 = ~pi02167 & w17566;
assign w33728 = ~w33726 & ~w33727;
assign w33729 = pi06598 & ~w17838;
assign w33730 = w17837 & w20209;
assign w33731 = ~w33729 & ~w33730;
assign w33732 = pi06599 & ~w17838;
assign w33733 = ~pi02713 & w17838;
assign w33734 = ~w33732 & ~w33733;
assign w33735 = pi06600 & ~w17838;
assign w33736 = ~pi02714 & w17838;
assign w33737 = ~w33735 & ~w33736;
assign w33738 = pi06601 & ~w17566;
assign w33739 = ~pi02722 & w17566;
assign w33740 = ~w33738 & ~w33739;
assign w33741 = pi06602 & ~w17838;
assign w33742 = ~pi02716 & w17838;
assign w33743 = ~w33741 & ~w33742;
assign w33744 = pi06603 & ~w17838;
assign w33745 = ~pi02717 & w17838;
assign w33746 = ~w33744 & ~w33745;
assign w33747 = ~w16905 & w20465;
assign w33748 = pi06604 & ~w33747;
assign w33749 = ~pi02711 & w33747;
assign w33750 = ~w33748 & ~w33749;
assign w33751 = pi06605 & ~w33747;
assign w33752 = ~pi02712 & w33747;
assign w33753 = ~w33751 & ~w33752;
assign w33754 = pi06606 & ~w33747;
assign w33755 = ~pi02170 & w33747;
assign w33756 = ~w33754 & ~w33755;
assign w33757 = pi06607 & ~w33747;
assign w33758 = ~pi02713 & w33747;
assign w33759 = ~w33757 & ~w33758;
assign w33760 = pi06608 & ~w33747;
assign w33761 = ~pi02714 & w33747;
assign w33762 = ~w33760 & ~w33761;
assign w33763 = pi06609 & ~w33747;
assign w33764 = ~pi02715 & w33747;
assign w33765 = ~w33763 & ~w33764;
assign w33766 = pi06610 & ~w33747;
assign w33767 = ~pi02716 & w33747;
assign w33768 = ~w33766 & ~w33767;
assign w33769 = pi06611 & ~w33747;
assign w33770 = ~pi02717 & w33747;
assign w33771 = ~w33769 & ~w33770;
assign w33772 = pi06612 & ~w17815;
assign w33773 = ~pi02712 & w17815;
assign w33774 = ~w33772 & ~w33773;
assign w33775 = pi06613 & ~w17815;
assign w33776 = ~pi02170 & w17815;
assign w33777 = ~w33775 & ~w33776;
assign w33778 = pi06614 & ~w17815;
assign w33779 = w17814 & w17929;
assign w33780 = ~w33778 & ~w33779;
assign w33781 = pi06615 & ~w17815;
assign w33782 = w17814 & w18059;
assign w33783 = ~w33781 & ~w33782;
assign w33784 = pi06616 & ~w17815;
assign w33785 = ~pi02716 & w17815;
assign w33786 = ~w33784 & ~w33785;
assign w33787 = pi06617 & ~w17815;
assign w33788 = ~pi02717 & w17815;
assign w33789 = ~w33787 & ~w33788;
assign w33790 = pi06618 & ~w17823;
assign w33791 = w17020 & w17822;
assign w33792 = ~w33790 & ~w33791;
assign w33793 = pi06619 & ~w17823;
assign w33794 = ~pi02170 & w17823;
assign w33795 = ~w33793 & ~w33794;
assign w33796 = pi06620 & ~w17823;
assign w33797 = ~pi02713 & w17823;
assign w33798 = ~w33796 & ~w33797;
assign w33799 = pi06621 & ~w17823;
assign w33800 = ~pi02714 & w17823;
assign w33801 = ~w33799 & ~w33800;
assign w33802 = pi06622 & ~w17823;
assign w33803 = ~pi02715 & w17823;
assign w33804 = ~w33802 & ~w33803;
assign w33805 = pi06623 & ~w17823;
assign w33806 = w17317 & w17822;
assign w33807 = ~w33805 & ~w33806;
assign w33808 = pi06624 & ~w17823;
assign w33809 = ~pi02717 & w17823;
assign w33810 = ~w33808 & ~w33809;
assign w33811 = pi06625 & ~w17776;
assign w33812 = ~pi02712 & w17776;
assign w33813 = ~w33811 & ~w33812;
assign w33814 = pi06626 & ~w17776;
assign w33815 = ~pi02170 & w17776;
assign w33816 = ~w33814 & ~w33815;
assign w33817 = pi06627 & ~w17776;
assign w33818 = ~pi02713 & w17776;
assign w33819 = ~w33817 & ~w33818;
assign w33820 = pi06628 & ~w17776;
assign w33821 = ~pi02715 & w17776;
assign w33822 = ~w33820 & ~w33821;
assign w33823 = pi06629 & ~w17776;
assign w33824 = ~pi02716 & w17776;
assign w33825 = ~w33823 & ~w33824;
assign w33826 = pi06630 & ~w17776;
assign w33827 = ~pi02717 & w17776;
assign w33828 = ~w33826 & ~w33827;
assign w33829 = ~w16992 & w17466;
assign w33830 = pi06631 & ~w33829;
assign w33831 = ~pi02164 & w33829;
assign w33832 = ~w33830 & ~w33831;
assign w33833 = pi06632 & ~w17574;
assign w33834 = w17020 & w17573;
assign w33835 = ~w33833 & ~w33834;
assign w33836 = pi06633 & ~w17574;
assign w33837 = w17573 & w20209;
assign w33838 = ~w33836 & ~w33837;
assign w33839 = pi06634 & ~w17574;
assign w33840 = ~pi02713 & w17574;
assign w33841 = ~w33839 & ~w33840;
assign w33842 = pi06635 & ~w17574;
assign w33843 = ~pi02714 & w17574;
assign w33844 = ~w33842 & ~w33843;
assign w33845 = pi06636 & ~w17574;
assign w33846 = ~pi02715 & w17574;
assign w33847 = ~w33845 & ~w33846;
assign w33848 = pi06637 & ~w17574;
assign w33849 = w17317 & w17573;
assign w33850 = ~w33848 & ~w33849;
assign w33851 = pi06638 & ~w17574;
assign w33852 = ~pi02717 & w17574;
assign w33853 = ~w33851 & ~w33852;
assign w33854 = pi06639 & ~w17029;
assign w33855 = ~pi02712 & w17029;
assign w33856 = ~w33854 & ~w33855;
assign w33857 = pi06640 & ~w17029;
assign w33858 = ~pi02170 & w17029;
assign w33859 = ~w33857 & ~w33858;
assign w33860 = pi06641 & ~w17029;
assign w33861 = ~pi02713 & w17029;
assign w33862 = ~w33860 & ~w33861;
assign w33863 = pi06642 & ~w17029;
assign w33864 = ~pi02715 & w17029;
assign w33865 = ~w33863 & ~w33864;
assign w33866 = pi06643 & ~w17029;
assign w33867 = ~pi02716 & w17029;
assign w33868 = ~w33866 & ~w33867;
assign w33869 = pi06644 & ~w17029;
assign w33870 = ~pi02717 & w17029;
assign w33871 = ~w33869 & ~w33870;
assign w33872 = pi06645 & ~w17054;
assign w33873 = ~pi02712 & w17054;
assign w33874 = ~w33872 & ~w33873;
assign w33875 = pi06646 & ~w17054;
assign w33876 = ~pi02170 & w17054;
assign w33877 = ~w33875 & ~w33876;
assign w33878 = pi06647 & ~w17054;
assign w33879 = ~pi02713 & w17054;
assign w33880 = ~w33878 & ~w33879;
assign w33881 = pi06648 & ~w17054;
assign w33882 = ~pi02714 & w17054;
assign w33883 = ~w33881 & ~w33882;
assign w33884 = pi06649 & ~w17054;
assign w33885 = ~pi02715 & w17054;
assign w33886 = ~w33884 & ~w33885;
assign w33887 = pi06650 & ~w17054;
assign w33888 = w17053 & w17317;
assign w33889 = ~w33887 & ~w33888;
assign w33890 = pi06651 & ~w17054;
assign w33891 = ~pi02717 & w17054;
assign w33892 = ~w33890 & ~w33891;
assign w33893 = pi06652 & ~w17007;
assign w33894 = ~pi02712 & w17007;
assign w33895 = ~w33893 & ~w33894;
assign w33896 = pi06653 & ~w17007;
assign w33897 = ~pi02170 & w17007;
assign w33898 = ~w33896 & ~w33897;
assign w33899 = pi06654 & ~w17007;
assign w33900 = ~pi02713 & w17007;
assign w33901 = ~w33899 & ~w33900;
assign w33902 = pi06655 & ~w17007;
assign w33903 = ~pi02715 & w17007;
assign w33904 = ~w33902 & ~w33903;
assign w33905 = pi06656 & ~w17007;
assign w33906 = ~pi02716 & w17007;
assign w33907 = ~w33905 & ~w33906;
assign w33908 = pi06657 & ~w17007;
assign w33909 = ~pi02717 & w17007;
assign w33910 = ~w33908 & ~w33909;
assign w33911 = pi06658 & ~w21070;
assign w33912 = ~pi02703 & w21070;
assign w33913 = ~w33911 & ~w33912;
assign w33914 = ~w16905 & w17734;
assign w33915 = pi06659 & ~w33914;
assign w33916 = ~pi02712 & w33914;
assign w33917 = ~w33915 & ~w33916;
assign w33918 = pi06660 & ~w33914;
assign w33919 = ~pi02170 & w33914;
assign w33920 = ~w33918 & ~w33919;
assign w33921 = pi06661 & ~w33914;
assign w33922 = ~pi02713 & w33914;
assign w33923 = ~w33921 & ~w33922;
assign w33924 = pi06662 & ~w33914;
assign w33925 = ~pi02714 & w33914;
assign w33926 = ~w33924 & ~w33925;
assign w33927 = pi06663 & ~w33914;
assign w33928 = ~pi02715 & w33914;
assign w33929 = ~w33927 & ~w33928;
assign w33930 = pi06664 & ~w33914;
assign w33931 = ~pi02716 & w33914;
assign w33932 = ~w33930 & ~w33931;
assign w33933 = pi06665 & ~w33914;
assign w33934 = ~pi02717 & w33914;
assign w33935 = ~w33933 & ~w33934;
assign w33936 = ~w16905 & w17406;
assign w33937 = pi06666 & ~w33936;
assign w33938 = ~pi02712 & w33936;
assign w33939 = ~w33937 & ~w33938;
assign w33940 = pi06667 & ~w33936;
assign w33941 = ~pi02170 & w33936;
assign w33942 = ~w33940 & ~w33941;
assign w33943 = pi06668 & ~w33936;
assign w33944 = ~pi02713 & w33936;
assign w33945 = ~w33943 & ~w33944;
assign w33946 = pi06669 & ~w33936;
assign w33947 = ~pi02715 & w33936;
assign w33948 = ~w33946 & ~w33947;
assign w33949 = pi06670 & ~w33936;
assign w33950 = ~pi02716 & w33936;
assign w33951 = ~w33949 & ~w33950;
assign w33952 = pi06671 & ~w33936;
assign w33953 = ~pi02717 & w33936;
assign w33954 = ~w33952 & ~w33953;
assign w33955 = ~w16905 & w19629;
assign w33956 = pi06672 & ~w33955;
assign w33957 = ~pi02712 & w33955;
assign w33958 = ~w33956 & ~w33957;
assign w33959 = pi06673 & ~w33955;
assign w33960 = ~pi02170 & w33955;
assign w33961 = ~w33959 & ~w33960;
assign w33962 = pi06674 & ~w33955;
assign w33963 = ~pi02713 & w33955;
assign w33964 = ~w33962 & ~w33963;
assign w33965 = pi06675 & ~w33955;
assign w33966 = ~pi02714 & w33955;
assign w33967 = ~w33965 & ~w33966;
assign w33968 = ~w16992 & w18040;
assign w33969 = pi06676 & ~w33968;
assign w33970 = ~pi02703 & w33968;
assign w33971 = ~w33969 & ~w33970;
assign w33972 = pi06677 & ~w33955;
assign w33973 = ~pi02715 & w33955;
assign w33974 = ~w33972 & ~w33973;
assign w33975 = pi06678 & ~w33968;
assign w33976 = ~pi02721 & w33968;
assign w33977 = ~w33975 & ~w33976;
assign w33978 = pi06679 & ~w33955;
assign w33979 = ~pi02716 & w33955;
assign w33980 = ~w33978 & ~w33979;
assign w33981 = pi06680 & ~w33955;
assign w33982 = ~pi02717 & w33955;
assign w33983 = ~w33981 & ~w33982;
assign w33984 = ~w16905 & w19655;
assign w33985 = pi06681 & ~w33984;
assign w33986 = w17603 & w19655;
assign w33987 = ~w33985 & ~w33986;
assign w33988 = pi06682 & ~w33984;
assign w33989 = ~pi02170 & w33984;
assign w33990 = ~w33988 & ~w33989;
assign w33991 = pi06683 & ~w33968;
assign w33992 = ~pi02718 & w33968;
assign w33993 = ~w33991 & ~w33992;
assign w33994 = pi06684 & ~w33984;
assign w33995 = ~pi02713 & w33984;
assign w33996 = ~w33994 & ~w33995;
assign w33997 = pi06685 & ~w33968;
assign w33998 = ~pi02167 & w33968;
assign w33999 = ~w33997 & ~w33998;
assign w34000 = pi06686 & ~w33984;
assign w34001 = w18059 & w19655;
assign w34002 = ~w34000 & ~w34001;
assign w34003 = pi06687 & ~w33984;
assign w34004 = ~pi02716 & w33984;
assign w34005 = ~w34003 & ~w34004;
assign w34006 = pi06688 & ~w33968;
assign w34007 = ~pi02722 & w33968;
assign w34008 = ~w34006 & ~w34007;
assign w34009 = pi06689 & ~w33984;
assign w34010 = ~pi02717 & w33984;
assign w34011 = ~w34009 & ~w34010;
assign w34012 = ~w16905 & w19596;
assign w34013 = pi06690 & ~w34012;
assign w34014 = ~pi02711 & w34012;
assign w34015 = ~w34013 & ~w34014;
assign w34016 = pi06691 & ~w34012;
assign w34017 = ~pi02712 & w34012;
assign w34018 = ~w34016 & ~w34017;
assign w34019 = pi06692 & ~w34012;
assign w34020 = ~pi02170 & w34012;
assign w34021 = ~w34019 & ~w34020;
assign w34022 = pi06693 & ~w34012;
assign w34023 = ~pi02713 & w34012;
assign w34024 = ~w34022 & ~w34023;
assign w34025 = pi06694 & ~w34012;
assign w34026 = w17742 & w19596;
assign w34027 = ~w34025 & ~w34026;
assign w34028 = pi06695 & ~w33968;
assign w34029 = ~pi02164 & w33968;
assign w34030 = ~w34028 & ~w34029;
assign w34031 = pi06696 & ~w34012;
assign w34032 = ~pi02716 & w34012;
assign w34033 = ~w34031 & ~w34032;
assign w34034 = pi06697 & ~w34012;
assign w34035 = ~pi02717 & w34012;
assign w34036 = ~w34034 & ~w34035;
assign w34037 = pi06698 & ~w21232;
assign w34038 = ~pi02712 & w21232;
assign w34039 = ~w34037 & ~w34038;
assign w34040 = pi06699 & ~w21232;
assign w34041 = ~pi02170 & w21232;
assign w34042 = ~w34040 & ~w34041;
assign w34043 = pi06700 & ~w21232;
assign w34044 = w17279 & w17929;
assign w34045 = ~w34043 & ~w34044;
assign w34046 = pi06701 & ~w21232;
assign w34047 = w17279 & w17742;
assign w34048 = ~w34046 & ~w34047;
assign w34049 = pi06702 & ~w21232;
assign w34050 = ~pi02715 & w21232;
assign w34051 = ~w34049 & ~w34050;
assign w34052 = pi06703 & ~w21232;
assign w34053 = ~pi02716 & w21232;
assign w34054 = ~w34052 & ~w34053;
assign w34055 = pi06704 & ~w21232;
assign w34056 = ~pi02717 & w21232;
assign w34057 = ~w34055 & ~w34056;
assign w34058 = pi06705 & ~w20531;
assign w34059 = w17811 & w17917;
assign w34060 = ~w34058 & ~w34059;
assign w34061 = pi06706 & ~w20531;
assign w34062 = w17917 & w19797;
assign w34063 = ~w34061 & ~w34062;
assign w34064 = pi06707 & ~w20531;
assign w34065 = w17586 & w17917;
assign w34066 = ~w34064 & ~w34065;
assign w34067 = pi06708 & ~w20531;
assign w34068 = w17620 & w17917;
assign w34069 = ~w34067 & ~w34068;
assign w34070 = ~w16905 & w19282;
assign w34071 = pi06709 & ~w34070;
assign w34072 = ~pi02711 & w34070;
assign w34073 = ~w34071 & ~w34072;
assign w34074 = pi06710 & ~w34070;
assign w34075 = ~pi02712 & w34070;
assign w34076 = ~w34074 & ~w34075;
assign w34077 = pi06711 & ~w34070;
assign w34078 = ~pi02170 & w34070;
assign w34079 = ~w34077 & ~w34078;
assign w34080 = pi06712 & ~w34070;
assign w34081 = ~pi02713 & w34070;
assign w34082 = ~w34080 & ~w34081;
assign w34083 = pi06713 & ~w34070;
assign w34084 = ~pi02714 & w34070;
assign w34085 = ~w34083 & ~w34084;
assign w34086 = pi06714 & ~w34070;
assign w34087 = ~pi02715 & w34070;
assign w34088 = ~w34086 & ~w34087;
assign w34089 = pi06715 & ~w34070;
assign w34090 = ~pi02716 & w34070;
assign w34091 = ~w34089 & ~w34090;
assign w34092 = pi06716 & ~w20531;
assign w34093 = w17594 & w17917;
assign w34094 = ~w34092 & ~w34093;
assign w34095 = pi06717 & ~w34070;
assign w34096 = w16973 & w19282;
assign w34097 = ~w34095 & ~w34096;
assign w34098 = pi06718 & ~w20322;
assign w34099 = ~pi02712 & w20322;
assign w34100 = ~w34098 & ~w34099;
assign w34101 = pi06719 & ~w20322;
assign w34102 = ~pi02170 & w20322;
assign w34103 = ~w34101 & ~w34102;
assign w34104 = pi06720 & ~w20322;
assign w34105 = ~pi02713 & w20322;
assign w34106 = ~w34104 & ~w34105;
assign w34107 = pi06721 & ~w20322;
assign w34108 = ~pi02715 & w20322;
assign w34109 = ~w34107 & ~w34108;
assign w34110 = pi06722 & ~w20322;
assign w34111 = ~pi02716 & w20322;
assign w34112 = ~w34110 & ~w34111;
assign w34113 = pi06723 & ~w20322;
assign w34114 = ~pi02717 & w20322;
assign w34115 = ~w34113 & ~w34114;
assign w34116 = pi06724 & ~w20310;
assign w34117 = ~pi02712 & w20310;
assign w34118 = ~w34116 & ~w34117;
assign w34119 = pi06725 & ~w20310;
assign w34120 = ~pi02170 & w20310;
assign w34121 = ~w34119 & ~w34120;
assign w34122 = pi06726 & ~w20310;
assign w34123 = ~pi02713 & w20310;
assign w34124 = ~w34122 & ~w34123;
assign w34125 = pi06727 & ~w20310;
assign w34126 = w17742 & w18636;
assign w34127 = ~w34125 & ~w34126;
assign w34128 = pi06728 & ~w20310;
assign w34129 = ~pi02715 & w20310;
assign w34130 = ~w34128 & ~w34129;
assign w34131 = pi06729 & ~w20310;
assign w34132 = ~pi02716 & w20310;
assign w34133 = ~w34131 & ~w34132;
assign w34134 = pi06730 & ~w20292;
assign w34135 = w17532 & w17668;
assign w34136 = ~w34134 & ~w34135;
assign w34137 = pi06731 & ~w20292;
assign w34138 = w17668 & w17811;
assign w34139 = ~w34137 & ~w34138;
assign w34140 = pi06732 & ~w20292;
assign w34141 = w17668 & w19797;
assign w34142 = ~w34140 & ~w34141;
assign w34143 = pi06733 & ~w20292;
assign w34144 = w17586 & w17668;
assign w34145 = ~w34143 & ~w34144;
assign w34146 = pi06734 & ~w20292;
assign w34147 = w17620 & w17668;
assign w34148 = ~w34146 & ~w34147;
assign w34149 = pi06735 & ~w20285;
assign w34150 = ~pi02711 & w20285;
assign w34151 = ~w34149 & ~w34150;
assign w34152 = pi06736 & ~w20285;
assign w34153 = w17020 & w18572;
assign w34154 = ~w34152 & ~w34153;
assign w34155 = pi06737 & ~w20285;
assign w34156 = w17929 & w18572;
assign w34157 = ~w34155 & ~w34156;
assign w34158 = pi06738 & ~w20292;
assign w34159 = w17668 & w19312;
assign w34160 = ~w34158 & ~w34159;
assign w34161 = pi06739 & ~w20285;
assign w34162 = ~pi02714 & w20285;
assign w34163 = ~w34161 & ~w34162;
assign w34164 = pi06740 & ~w20285;
assign w34165 = ~pi02715 & w20285;
assign w34166 = ~w34164 & ~w34165;
assign w34167 = pi06741 & ~w20292;
assign w34168 = w17594 & w17668;
assign w34169 = ~w34167 & ~w34168;
assign w34170 = pi06742 & ~w20285;
assign w34171 = ~pi02716 & w20285;
assign w34172 = ~w34170 & ~w34171;
assign w34173 = pi06743 & ~w20285;
assign w34174 = ~pi02717 & w20285;
assign w34175 = ~w34173 & ~w34174;
assign w34176 = pi06744 & ~w19402;
assign w34177 = ~pi02712 & w19402;
assign w34178 = ~w34176 & ~w34177;
assign w34179 = pi06745 & ~w19402;
assign w34180 = ~pi02170 & w19402;
assign w34181 = ~w34179 & ~w34180;
assign w34182 = pi06746 & ~w19402;
assign w34183 = ~pi02713 & w19402;
assign w34184 = ~w34182 & ~w34183;
assign w34185 = pi06747 & ~w19402;
assign w34186 = ~pi02715 & w19402;
assign w34187 = ~w34185 & ~w34186;
assign w34188 = pi06748 & ~w19402;
assign w34189 = ~pi02716 & w19402;
assign w34190 = ~w34188 & ~w34189;
assign w34191 = pi06749 & ~w19402;
assign w34192 = ~pi02717 & w19402;
assign w34193 = ~w34191 & ~w34192;
assign w34194 = pi06750 & ~w18518;
assign w34195 = ~pi02721 & w18518;
assign w34196 = ~w34194 & ~w34195;
assign w34197 = pi06751 & ~w18518;
assign w34198 = w17636 & w19797;
assign w34199 = ~w34197 & ~w34198;
assign w34200 = pi06752 & ~w18518;
assign w34201 = ~pi02718 & w18518;
assign w34202 = ~w34200 & ~w34201;
assign w34203 = pi06753 & ~w18518;
assign w34204 = ~pi02167 & w18518;
assign w34205 = ~w34203 & ~w34204;
assign w34206 = pi06754 & ~w18518;
assign w34207 = ~pi02164 & w18518;
assign w34208 = ~w34206 & ~w34207;
assign w34209 = pi06755 & ~w18696;
assign w34210 = w17603 & w18186;
assign w34211 = ~w34209 & ~w34210;
assign w34212 = pi06756 & ~w18696;
assign w34213 = ~pi02712 & w18696;
assign w34214 = ~w34212 & ~w34213;
assign w34215 = pi06757 & ~w18696;
assign w34216 = ~pi02170 & w18696;
assign w34217 = ~w34215 & ~w34216;
assign w34218 = pi06758 & ~w18696;
assign w34219 = ~pi02713 & w18696;
assign w34220 = ~w34218 & ~w34219;
assign w34221 = pi06759 & ~w18696;
assign w34222 = ~pi02714 & w18696;
assign w34223 = ~w34221 & ~w34222;
assign w34224 = pi06760 & ~w18518;
assign w34225 = ~pi02719 & w18518;
assign w34226 = ~w34224 & ~w34225;
assign w34227 = pi06761 & ~w18696;
assign w34228 = ~pi02716 & w18696;
assign w34229 = ~w34227 & ~w34228;
assign w34230 = pi06762 & ~w18696;
assign w34231 = ~pi02717 & w18696;
assign w34232 = ~w34230 & ~w34231;
assign w34233 = pi06763 & ~w18667;
assign w34234 = w17020 & w17084;
assign w34235 = ~w34233 & ~w34234;
assign w34236 = pi06764 & ~w18667;
assign w34237 = ~pi02170 & w18667;
assign w34238 = ~w34236 & ~w34237;
assign w34239 = pi06765 & ~w18667;
assign w34240 = w17084 & w17929;
assign w34241 = ~w34239 & ~w34240;
assign w34242 = pi06766 & ~w18667;
assign w34243 = ~pi02714 & w18667;
assign w34244 = ~w34242 & ~w34243;
assign w34245 = pi06767 & ~w18667;
assign w34246 = ~pi02715 & w18667;
assign w34247 = ~w34245 & ~w34246;
assign w34248 = pi06768 & ~w18667;
assign w34249 = w17084 & w17317;
assign w34250 = ~w34248 & ~w34249;
assign w34251 = pi06769 & ~w18667;
assign w34252 = ~pi02717 & w18667;
assign w34253 = ~w34251 & ~w34252;
assign w34254 = pi06770 & ~w16971;
assign w34255 = ~pi02712 & w16971;
assign w34256 = ~w34254 & ~w34255;
assign w34257 = pi06771 & ~w16971;
assign w34258 = ~pi02170 & w16971;
assign w34259 = ~w34257 & ~w34258;
assign w34260 = pi06772 & ~w16971;
assign w34261 = ~pi02713 & w16971;
assign w34262 = ~w34260 & ~w34261;
assign w34263 = pi06773 & ~w16971;
assign w34264 = w16970 & w18059;
assign w34265 = ~w34263 & ~w34264;
assign w34266 = pi06774 & ~w18256;
assign w34267 = ~pi02703 & w18256;
assign w34268 = ~w34266 & ~w34267;
assign w34269 = pi06775 & ~w16971;
assign w34270 = ~pi02716 & w16971;
assign w34271 = ~w34269 & ~w34270;
assign w34272 = ~w16905 & w17808;
assign w34273 = pi06776 & ~w34272;
assign w34274 = ~pi02711 & w34272;
assign w34275 = ~w34273 & ~w34274;
assign w34276 = pi06777 & ~w18256;
assign w34277 = w16961 & w17811;
assign w34278 = ~w34276 & ~w34277;
assign w34279 = pi06778 & ~w34272;
assign w34280 = ~pi02712 & w34272;
assign w34281 = ~w34279 & ~w34280;
assign w34282 = pi06779 & ~w34272;
assign w34283 = ~pi02170 & w34272;
assign w34284 = ~w34282 & ~w34283;
assign w34285 = pi06780 & ~w18256;
assign w34286 = ~pi02169 & w18256;
assign w34287 = ~w34285 & ~w34286;
assign w34288 = pi06781 & ~w34272;
assign w34289 = ~pi02713 & w34272;
assign w34290 = ~w34288 & ~w34289;
assign w34291 = pi06782 & ~w34272;
assign w34292 = ~pi02714 & w34272;
assign w34293 = ~w34291 & ~w34292;
assign w34294 = pi06783 & ~w34272;
assign w34295 = ~pi02715 & w34272;
assign w34296 = ~w34294 & ~w34295;
assign w34297 = pi06784 & ~w34272;
assign w34298 = ~pi02716 & w34272;
assign w34299 = ~w34297 & ~w34298;
assign w34300 = pi06785 & ~w34272;
assign w34301 = ~pi02717 & w34272;
assign w34302 = ~w34300 & ~w34301;
assign w34303 = pi06786 & ~w18256;
assign w34304 = w16961 & w17620;
assign w34305 = ~w34303 & ~w34304;
assign w34306 = pi06787 & ~w18256;
assign w34307 = ~pi02722 & w18256;
assign w34308 = ~w34306 & ~w34307;
assign w34309 = pi06788 & ~w18256;
assign w34310 = w16961 & w17594;
assign w34311 = ~w34309 & ~w34310;
assign w34312 = ~w16905 & w17390;
assign w34313 = pi06789 & ~w34312;
assign w34314 = ~pi02711 & w34312;
assign w34315 = ~w34313 & ~w34314;
assign w34316 = pi06790 & ~w18010;
assign w34317 = ~pi02721 & w18010;
assign w34318 = ~w34316 & ~w34317;
assign w34319 = pi06791 & ~w34312;
assign w34320 = ~pi02712 & w34312;
assign w34321 = ~w34319 & ~w34320;
assign w34322 = pi06792 & ~w34312;
assign w34323 = ~pi02170 & w34312;
assign w34324 = ~w34322 & ~w34323;
assign w34325 = pi06793 & ~w18010;
assign w34326 = ~pi02169 & w18010;
assign w34327 = ~w34325 & ~w34326;
assign w34328 = pi06794 & ~w34312;
assign w34329 = ~pi02713 & w34312;
assign w34330 = ~w34328 & ~w34329;
assign w34331 = pi06795 & ~w34312;
assign w34332 = ~pi02714 & w34312;
assign w34333 = ~w34331 & ~w34332;
assign w34334 = pi06796 & ~w34312;
assign w34335 = ~pi02715 & w34312;
assign w34336 = ~w34334 & ~w34335;
assign w34337 = pi06797 & ~w34312;
assign w34338 = ~pi02716 & w34312;
assign w34339 = ~w34337 & ~w34338;
assign w34340 = pi06798 & ~w34312;
assign w34341 = w16973 & w17390;
assign w34342 = ~w34340 & ~w34341;
assign w34343 = pi06799 & ~w18010;
assign w34344 = ~pi02164 & w18010;
assign w34345 = ~w34343 & ~w34344;
assign w34346 = pi06800 & ~w18010;
assign w34347 = ~pi02722 & w18010;
assign w34348 = ~w34346 & ~w34347;
assign w34349 = pi06801 & ~w18010;
assign w34350 = ~pi02719 & w18010;
assign w34351 = ~w34349 & ~w34350;
assign w34352 = pi06802 & ~w18101;
assign w34353 = ~pi02712 & w18101;
assign w34354 = ~w34352 & ~w34353;
assign w34355 = pi06803 & ~w18101;
assign w34356 = ~pi02170 & w18101;
assign w34357 = ~w34355 & ~w34356;
assign w34358 = pi06804 & ~w18101;
assign w34359 = ~pi02713 & w18101;
assign w34360 = ~w34358 & ~w34359;
assign w34361 = pi06805 & ~w18101;
assign w34362 = ~pi02714 & w18101;
assign w34363 = ~w34361 & ~w34362;
assign w34364 = pi06806 & ~w18101;
assign w34365 = w17495 & w18059;
assign w34366 = ~w34364 & ~w34365;
assign w34367 = pi06807 & ~w18101;
assign w34368 = ~pi02716 & w18101;
assign w34369 = ~w34367 & ~w34368;
assign w34370 = pi06808 & ~w18101;
assign w34371 = ~pi02717 & w18101;
assign w34372 = ~w34370 & ~w34371;
assign w34373 = pi06809 & ~w17798;
assign w34374 = ~pi02712 & w17798;
assign w34375 = ~w34373 & ~w34374;
assign w34376 = pi06810 & ~w17798;
assign w34377 = ~pi02170 & w17798;
assign w34378 = ~w34376 & ~w34377;
assign w34379 = pi06811 & ~w17798;
assign w34380 = ~pi02713 & w17798;
assign w34381 = ~w34379 & ~w34380;
assign w34382 = pi06812 & ~w17798;
assign w34383 = ~pi02715 & w17798;
assign w34384 = ~w34382 & ~w34383;
assign w34385 = pi06813 & ~w17798;
assign w34386 = ~pi02716 & w17798;
assign w34387 = ~w34385 & ~w34386;
assign w34388 = pi06814 & ~w17798;
assign w34389 = ~pi02717 & w17798;
assign w34390 = ~w34388 & ~w34389;
assign w34391 = pi06815 & ~w17745;
assign w34392 = ~pi02712 & w17745;
assign w34393 = ~w34391 & ~w34392;
assign w34394 = pi06816 & ~w17745;
assign w34395 = ~pi02170 & w17745;
assign w34396 = ~w34394 & ~w34395;
assign w34397 = pi06817 & ~w17745;
assign w34398 = ~pi02713 & w17745;
assign w34399 = ~w34397 & ~w34398;
assign w34400 = pi06818 & ~w17745;
assign w34401 = ~pi02714 & w17745;
assign w34402 = ~w34400 & ~w34401;
assign w34403 = pi06819 & ~w17745;
assign w34404 = ~pi02715 & w17745;
assign w34405 = ~w34403 & ~w34404;
assign w34406 = pi06820 & ~w17745;
assign w34407 = ~pi02716 & w17745;
assign w34408 = ~w34406 & ~w34407;
assign w34409 = pi06821 & ~w17745;
assign w34410 = ~pi02717 & w17745;
assign w34411 = ~w34409 & ~w34410;
assign w34412 = pi06822 & ~w17651;
assign w34413 = ~pi02721 & w17651;
assign w34414 = ~w34412 & ~w34413;
assign w34415 = pi06823 & ~w17651;
assign w34416 = ~pi02169 & w17651;
assign w34417 = ~w34415 & ~w34416;
assign w34418 = pi06824 & ~w17651;
assign w34419 = ~pi02718 & w17651;
assign w34420 = ~w34418 & ~w34419;
assign w34421 = pi06825 & ~w17651;
assign w34422 = ~pi02167 & w17651;
assign w34423 = ~w34421 & ~w34422;
assign w34424 = pi06826 & ~w17651;
assign w34425 = ~pi02722 & w17651;
assign w34426 = ~w34424 & ~w34425;
assign w34427 = pi06827 & ~w17651;
assign w34428 = ~pi02719 & w17651;
assign w34429 = ~w34427 & ~w34428;
assign w34430 = ~w16992 & w18622;
assign w34431 = pi06828 & ~w34430;
assign w34432 = ~pi02703 & w34430;
assign w34433 = ~w34431 & ~w34432;
assign w34434 = pi06829 & ~w16979;
assign w34435 = ~pi02712 & w16979;
assign w34436 = ~w34434 & ~w34435;
assign w34437 = pi06830 & ~w16979;
assign w34438 = ~pi02170 & w16979;
assign w34439 = ~w34437 & ~w34438;
assign w34440 = pi06831 & ~w34430;
assign w34441 = ~pi02721 & w34430;
assign w34442 = ~w34440 & ~w34441;
assign w34443 = pi06832 & ~w16979;
assign w34444 = ~pi02713 & w16979;
assign w34445 = ~w34443 & ~w34444;
assign w34446 = pi06833 & ~w16979;
assign w34447 = w16978 & w17742;
assign w34448 = ~w34446 & ~w34447;
assign w34449 = pi06834 & ~w34430;
assign w34450 = ~pi02169 & w34430;
assign w34451 = ~w34449 & ~w34450;
assign w34452 = pi06835 & ~w34430;
assign w34453 = ~pi02718 & w34430;
assign w34454 = ~w34452 & ~w34453;
assign w34455 = pi06836 & ~w16979;
assign w34456 = w16978 & w17317;
assign w34457 = ~w34455 & ~w34456;
assign w34458 = pi06837 & ~w34430;
assign w34459 = ~pi02167 & w34430;
assign w34460 = ~w34458 & ~w34459;
assign w34461 = pi06838 & ~w34430;
assign w34462 = w17620 & w18622;
assign w34463 = ~w34461 & ~w34462;
assign w34464 = pi06839 & ~w34430;
assign w34465 = ~pi02722 & w34430;
assign w34466 = ~w34464 & ~w34465;
assign w34467 = pi06840 & ~w34430;
assign w34468 = ~pi02719 & w34430;
assign w34469 = ~w34467 & ~w34468;
assign w34470 = pi06841 & ~w16913;
assign w34471 = w16912 & w17020;
assign w34472 = ~w34470 & ~w34471;
assign w34473 = pi06842 & ~w16913;
assign w34474 = ~pi02170 & w16913;
assign w34475 = ~w34473 & ~w34474;
assign w34476 = pi06843 & ~w16913;
assign w34477 = ~pi02713 & w16913;
assign w34478 = ~w34476 & ~w34477;
assign w34479 = pi06844 & ~w16913;
assign w34480 = ~pi02714 & w16913;
assign w34481 = ~w34479 & ~w34480;
assign w34482 = pi06845 & ~w16913;
assign w34483 = w16912 & w18059;
assign w34484 = ~w34482 & ~w34483;
assign w34485 = pi06846 & ~w16913;
assign w34486 = ~pi02716 & w16913;
assign w34487 = ~w34485 & ~w34486;
assign w34488 = pi06847 & ~w16913;
assign w34489 = ~pi02717 & w16913;
assign w34490 = ~w34488 & ~w34489;
assign w34491 = ~w16905 & w17284;
assign w34492 = pi06848 & ~w34491;
assign w34493 = ~pi02712 & w34491;
assign w34494 = ~w34492 & ~w34493;
assign w34495 = pi06849 & ~w34491;
assign w34496 = ~pi02170 & w34491;
assign w34497 = ~w34495 & ~w34496;
assign w34498 = pi06850 & ~w34491;
assign w34499 = ~pi02713 & w34491;
assign w34500 = ~w34498 & ~w34499;
assign w34501 = pi06851 & ~w34491;
assign w34502 = ~pi02715 & w34491;
assign w34503 = ~w34501 & ~w34502;
assign w34504 = pi06852 & ~w34491;
assign w34505 = ~pi02716 & w34491;
assign w34506 = ~w34504 & ~w34505;
assign w34507 = pi06853 & ~w34491;
assign w34508 = w16973 & w17284;
assign w34509 = ~w34507 & ~w34508;
assign w34510 = ~w16992 & w17190;
assign w34511 = pi06854 & ~w34510;
assign w34512 = w17190 & w17532;
assign w34513 = ~w34511 & ~w34512;
assign w34514 = ~w16905 & w17177;
assign w34515 = pi06855 & ~w34514;
assign w34516 = ~pi02712 & w34514;
assign w34517 = ~w34515 & ~w34516;
assign w34518 = pi06856 & ~w34514;
assign w34519 = ~pi02170 & w34514;
assign w34520 = ~w34518 & ~w34519;
assign w34521 = pi06857 & ~w34510;
assign w34522 = w17190 & w17811;
assign w34523 = ~w34521 & ~w34522;
assign w34524 = pi06858 & ~w34514;
assign w34525 = ~pi02713 & w34514;
assign w34526 = ~w34524 & ~w34525;
assign w34527 = pi06859 & ~w34514;
assign w34528 = ~pi02714 & w34514;
assign w34529 = ~w34527 & ~w34528;
assign w34530 = pi06860 & ~w34514;
assign w34531 = w17177 & w18059;
assign w34532 = ~w34530 & ~w34531;
assign w34533 = pi06861 & ~w34510;
assign w34534 = ~pi02718 & w34510;
assign w34535 = ~w34533 & ~w34534;
assign w34536 = pi06862 & ~w34514;
assign w34537 = w16973 & w17177;
assign w34538 = ~w34536 & ~w34537;
assign w34539 = pi06863 & ~w34510;
assign w34540 = ~pi02169 & w34510;
assign w34541 = ~w34539 & ~w34540;
assign w34542 = pi06864 & ~w34510;
assign w34543 = ~pi02164 & w34510;
assign w34544 = ~w34542 & ~w34543;
assign w34545 = pi06865 & ~w34510;
assign w34546 = ~pi02722 & w34510;
assign w34547 = ~w34545 & ~w34546;
assign w34548 = pi06866 & ~w34510;
assign w34549 = ~pi02719 & w34510;
assign w34550 = ~w34548 & ~w34549;
assign w34551 = ~w16905 & w18177;
assign w34552 = pi06867 & ~w34551;
assign w34553 = ~pi02712 & w34551;
assign w34554 = ~w34552 & ~w34553;
assign w34555 = pi06868 & ~w34551;
assign w34556 = ~pi02170 & w34551;
assign w34557 = ~w34555 & ~w34556;
assign w34558 = pi06869 & ~w34551;
assign w34559 = w17929 & w18177;
assign w34560 = ~w34558 & ~w34559;
assign w34561 = pi06870 & ~w34551;
assign w34562 = ~pi02714 & w34551;
assign w34563 = ~w34561 & ~w34562;
assign w34564 = pi06871 & ~w34551;
assign w34565 = ~pi02715 & w34551;
assign w34566 = ~w34564 & ~w34565;
assign w34567 = pi06872 & ~w34551;
assign w34568 = ~pi02716 & w34551;
assign w34569 = ~w34567 & ~w34568;
assign w34570 = pi06873 & ~w34551;
assign w34571 = w16973 & w18177;
assign w34572 = ~w34570 & ~w34571;
assign w34573 = ~w16905 & w17565;
assign w34574 = pi06874 & ~w34573;
assign w34575 = ~pi02712 & w34573;
assign w34576 = ~w34574 & ~w34575;
assign w34577 = pi06875 & ~w34573;
assign w34578 = ~pi02170 & w34573;
assign w34579 = ~w34577 & ~w34578;
assign w34580 = pi06876 & ~w34573;
assign w34581 = ~pi02713 & w34573;
assign w34582 = ~w34580 & ~w34581;
assign w34583 = pi06877 & ~w34573;
assign w34584 = ~pi02715 & w34573;
assign w34585 = ~w34583 & ~w34584;
assign w34586 = pi06878 & ~w34573;
assign w34587 = w17317 & w17565;
assign w34588 = ~w34586 & ~w34587;
assign w34589 = pi06879 & ~w34573;
assign w34590 = w16973 & w17565;
assign w34591 = ~w34589 & ~w34590;
assign w34592 = ~w16992 & w17600;
assign w34593 = pi06880 & ~w34592;
assign w34594 = w17600 & w17811;
assign w34595 = ~w34593 & ~w34594;
assign w34596 = pi06881 & ~w34592;
assign w34597 = ~pi02169 & w34592;
assign w34598 = ~w34596 & ~w34597;
assign w34599 = pi06882 & ~w34592;
assign w34600 = ~pi02718 & w34592;
assign w34601 = ~w34599 & ~w34600;
assign w34602 = pi06883 & ~w34592;
assign w34603 = w17600 & w19273;
assign w34604 = ~w34602 & ~w34603;
assign w34605 = pi06884 & ~w34592;
assign w34606 = ~pi02164 & w34592;
assign w34607 = ~w34605 & ~w34606;
assign w34608 = pi06885 & ~w34592;
assign w34609 = ~pi02722 & w34592;
assign w34610 = ~w34608 & ~w34609;
assign w34611 = pi06886 & ~w34592;
assign w34612 = ~pi02719 & w34592;
assign w34613 = ~w34611 & ~w34612;
assign w34614 = pi06887 & ~w21929;
assign w34615 = ~pi02721 & w21929;
assign w34616 = ~w34614 & ~w34615;
assign w34617 = pi06888 & ~w21929;
assign w34618 = w17375 & w19797;
assign w34619 = ~w34617 & ~w34618;
assign w34620 = pi06889 & ~w21929;
assign w34621 = ~pi02718 & w21929;
assign w34622 = ~w34620 & ~w34621;
assign w34623 = pi06890 & ~w21929;
assign w34624 = ~pi02164 & w21929;
assign w34625 = ~w34623 & ~w34624;
assign w34626 = pi06891 & ~w21929;
assign w34627 = ~pi02722 & w21929;
assign w34628 = ~w34626 & ~w34627;
assign w34629 = ~w16905 & w18040;
assign w34630 = pi06892 & ~w34629;
assign w34631 = ~pi02711 & w34629;
assign w34632 = ~w34630 & ~w34631;
assign w34633 = pi06893 & ~w34629;
assign w34634 = ~pi02712 & w34629;
assign w34635 = ~w34633 & ~w34634;
assign w34636 = pi06894 & ~w34629;
assign w34637 = ~pi02170 & w34629;
assign w34638 = ~w34636 & ~w34637;
assign w34639 = pi06895 & ~w21293;
assign w34640 = ~pi02703 & w21293;
assign w34641 = ~w34639 & ~w34640;
assign w34642 = pi06896 & ~w34629;
assign w34643 = ~pi02713 & w34629;
assign w34644 = ~w34642 & ~w34643;
assign w34645 = pi06897 & ~w34629;
assign w34646 = ~pi02714 & w34629;
assign w34647 = ~w34645 & ~w34646;
assign w34648 = pi06898 & ~w21293;
assign w34649 = w17811 & w18731;
assign w34650 = ~w34648 & ~w34649;
assign w34651 = pi06899 & ~w34629;
assign w34652 = ~pi02715 & w34629;
assign w34653 = ~w34651 & ~w34652;
assign w34654 = pi06900 & ~w34629;
assign w34655 = w17317 & w18040;
assign w34656 = ~w34654 & ~w34655;
assign w34657 = pi06901 & ~w21293;
assign w34658 = ~pi02718 & w21293;
assign w34659 = ~w34657 & ~w34658;
assign w34660 = pi06902 & ~w34629;
assign w34661 = ~pi02717 & w34629;
assign w34662 = ~w34660 & ~w34661;
assign w34663 = pi06903 & ~w21293;
assign w34664 = w17620 & w18731;
assign w34665 = ~w34663 & ~w34664;
assign w34666 = pi06904 & ~w21293;
assign w34667 = ~pi02722 & w21293;
assign w34668 = ~w34666 & ~w34667;
assign w34669 = pi06905 & ~w21467;
assign w34670 = w17603 & w17917;
assign w34671 = ~w34669 & ~w34670;
assign w34672 = pi06906 & ~w21467;
assign w34673 = ~pi02712 & w21467;
assign w34674 = ~w34672 & ~w34673;
assign w34675 = pi06907 & ~w21467;
assign w34676 = ~pi02170 & w21467;
assign w34677 = ~w34675 & ~w34676;
assign w34678 = pi06908 & ~w21460;
assign w34679 = ~pi02703 & w21460;
assign w34680 = ~w34678 & ~w34679;
assign w34681 = pi06909 & ~w21467;
assign w34682 = ~pi02713 & w21467;
assign w34683 = ~w34681 & ~w34682;
assign w34684 = pi06910 & ~w21467;
assign w34685 = ~pi02714 & w21467;
assign w34686 = ~w34684 & ~w34685;
assign w34687 = pi06911 & ~w21460;
assign w34688 = ~pi02721 & w21460;
assign w34689 = ~w34687 & ~w34688;
assign w34690 = pi06912 & ~w21467;
assign w34691 = ~pi02715 & w21467;
assign w34692 = ~w34690 & ~w34691;
assign w34693 = pi06913 & ~w21467;
assign w34694 = ~pi02717 & w21467;
assign w34695 = ~w34693 & ~w34694;
assign w34696 = pi06914 & ~w21460;
assign w34697 = ~pi02169 & w21460;
assign w34698 = ~w34696 & ~w34697;
assign w34699 = pi06915 & ~w21460;
assign w34700 = ~pi02718 & w21460;
assign w34701 = ~w34699 & ~w34700;
assign w34702 = pi06916 & ~w21460;
assign w34703 = ~pi02164 & w21460;
assign w34704 = ~w34702 & ~w34703;
assign w34705 = pi06917 & ~w21460;
assign w34706 = ~pi02722 & w21460;
assign w34707 = ~w34705 & ~w34706;
assign w34708 = pi06918 & ~w18507;
assign w34709 = ~pi02711 & w18507;
assign w34710 = ~w34708 & ~w34709;
assign w34711 = pi06919 & ~w18507;
assign w34712 = ~pi02712 & w18507;
assign w34713 = ~w34711 & ~w34712;
assign w34714 = pi06920 & ~w18507;
assign w34715 = w17668 & w20209;
assign w34716 = ~w34714 & ~w34715;
assign w34717 = pi06921 & ~w20326;
assign w34718 = ~pi02703 & w20326;
assign w34719 = ~w34717 & ~w34718;
assign w34720 = pi06922 & ~w18507;
assign w34721 = w17668 & w17929;
assign w34722 = ~w34720 & ~w34721;
assign w34723 = pi06923 & ~w18507;
assign w34724 = ~pi02714 & w18507;
assign w34725 = ~w34723 & ~w34724;
assign w34726 = pi06924 & ~w20326;
assign w34727 = ~pi02721 & w20326;
assign w34728 = ~w34726 & ~w34727;
assign w34729 = pi06925 & ~w18507;
assign w34730 = ~pi02715 & w18507;
assign w34731 = ~w34729 & ~w34730;
assign w34732 = pi06926 & ~w20326;
assign w34733 = ~pi02169 & w20326;
assign w34734 = ~w34732 & ~w34733;
assign w34735 = pi06927 & ~w18507;
assign w34736 = ~pi02717 & w18507;
assign w34737 = ~w34735 & ~w34736;
assign w34738 = pi06928 & ~w20326;
assign w34739 = w17586 & w18348;
assign w34740 = ~w34738 & ~w34739;
assign w34741 = pi06929 & ~w20326;
assign w34742 = ~pi02164 & w20326;
assign w34743 = ~w34741 & ~w34742;
assign w34744 = pi06930 & ~w20326;
assign w34745 = ~pi02722 & w20326;
assign w34746 = ~w34744 & ~w34745;
assign w34747 = pi06931 & ~w20314;
assign w34748 = ~pi02711 & w20314;
assign w34749 = ~w34747 & ~w34748;
assign w34750 = pi06932 & ~w20326;
assign w34751 = ~pi02719 & w20326;
assign w34752 = ~w34750 & ~w34751;
assign w34753 = pi06933 & ~w20314;
assign w34754 = w17636 & w20209;
assign w34755 = ~w34753 & ~w34754;
assign w34756 = pi06934 & ~w20314;
assign w34757 = ~pi02713 & w20314;
assign w34758 = ~w34756 & ~w34757;
assign w34759 = pi06935 & ~w20265;
assign w34760 = ~pi02703 & w20265;
assign w34761 = ~w34759 & ~w34760;
assign w34762 = pi06936 & ~w20314;
assign w34763 = ~pi02714 & w20314;
assign w34764 = ~w34762 & ~w34763;
assign w34765 = pi06937 & ~w20265;
assign w34766 = ~pi02721 & w20265;
assign w34767 = ~w34765 & ~w34766;
assign w34768 = pi06938 & ~w20314;
assign w34769 = ~pi02715 & w20314;
assign w34770 = ~w34768 & ~w34769;
assign w34771 = pi06939 & ~w20265;
assign w34772 = ~pi02169 & w20265;
assign w34773 = ~w34771 & ~w34772;
assign w34774 = pi06940 & ~w20314;
assign w34775 = ~pi02717 & w20314;
assign w34776 = ~w34774 & ~w34775;
assign w34777 = pi06941 & ~w20265;
assign w34778 = ~pi02718 & w20265;
assign w34779 = ~w34777 & ~w34778;
assign w34780 = pi06942 & ~w20265;
assign w34781 = ~pi02164 & w20265;
assign w34782 = ~w34780 & ~w34781;
assign w34783 = pi06943 & ~w20265;
assign w34784 = ~pi02722 & w20265;
assign w34785 = ~w34783 & ~w34784;
assign w34786 = pi06944 & ~w20151;
assign w34787 = ~pi02711 & w20151;
assign w34788 = ~w34786 & ~w34787;
assign w34789 = pi06945 & ~w20151;
assign w34790 = ~pi02712 & w20151;
assign w34791 = ~w34789 & ~w34790;
assign w34792 = pi06946 & ~w20151;
assign w34793 = ~pi02170 & w20151;
assign w34794 = ~w34792 & ~w34793;
assign w34795 = pi06947 & ~w19154;
assign w34796 = ~pi02703 & w19154;
assign w34797 = ~w34795 & ~w34796;
assign w34798 = pi06948 & ~w20151;
assign w34799 = ~pi02713 & w20151;
assign w34800 = ~w34798 & ~w34799;
assign w34801 = pi06949 & ~w20151;
assign w34802 = ~pi02714 & w20151;
assign w34803 = ~w34801 & ~w34802;
assign w34804 = pi06950 & ~w19154;
assign w34805 = ~pi02721 & w19154;
assign w34806 = ~w34804 & ~w34805;
assign w34807 = pi06951 & ~w20151;
assign w34808 = ~pi02715 & w20151;
assign w34809 = ~w34807 & ~w34808;
assign w34810 = pi06952 & ~w19154;
assign w34811 = ~pi02169 & w19154;
assign w34812 = ~w34810 & ~w34811;
assign w34813 = pi06953 & ~w20151;
assign w34814 = ~pi02717 & w20151;
assign w34815 = ~w34813 & ~w34814;
assign w34816 = pi06954 & ~w19963;
assign w34817 = ~pi02711 & w19963;
assign w34818 = ~w34816 & ~w34817;
assign w34819 = pi06955 & ~w19154;
assign w34820 = w17325 & w17586;
assign w34821 = ~w34819 & ~w34820;
assign w34822 = pi06956 & ~w19963;
assign w34823 = ~pi02170 & w19963;
assign w34824 = ~w34822 & ~w34823;
assign w34825 = pi06957 & ~w19963;
assign w34826 = ~pi02713 & w19963;
assign w34827 = ~w34825 & ~w34826;
assign w34828 = pi06958 & ~w19963;
assign w34829 = ~pi02714 & w19963;
assign w34830 = ~w34828 & ~w34829;
assign w34831 = pi06959 & ~w19963;
assign w34832 = ~pi02715 & w19963;
assign w34833 = ~w34831 & ~w34832;
assign w34834 = pi06960 & ~w19963;
assign w34835 = ~pi02716 & w19963;
assign w34836 = ~w34834 & ~w34835;
assign w34837 = pi06961 & ~w19154;
assign w34838 = w17325 & w17620;
assign w34839 = ~w34837 & ~w34838;
assign w34840 = pi06962 & ~w19963;
assign w34841 = ~pi02717 & w19963;
assign w34842 = ~w34840 & ~w34841;
assign w34843 = pi06963 & ~w19154;
assign w34844 = ~pi02722 & w19154;
assign w34845 = ~w34843 & ~w34844;
assign w34846 = pi06964 & ~w19154;
assign w34847 = ~pi02719 & w19154;
assign w34848 = ~w34846 & ~w34847;
assign w34849 = pi06965 & ~w19455;
assign w34850 = ~pi02721 & w19455;
assign w34851 = ~w34849 & ~w34850;
assign w34852 = pi06966 & ~w19455;
assign w34853 = ~pi02169 & w19455;
assign w34854 = ~w34852 & ~w34853;
assign w34855 = pi06967 & ~w19455;
assign w34856 = ~pi02718 & w19455;
assign w34857 = ~w34855 & ~w34856;
assign w34858 = pi06968 & ~w19455;
assign w34859 = ~pi02164 & w19455;
assign w34860 = ~w34858 & ~w34859;
assign w34861 = pi06969 & ~w18522;
assign w34862 = w17603 & w17650;
assign w34863 = ~w34861 & ~w34862;
assign w34864 = pi06970 & ~w19455;
assign w34865 = ~pi02722 & w19455;
assign w34866 = ~w34864 & ~w34865;
assign w34867 = pi06971 & ~w19455;
assign w34868 = ~pi02719 & w19455;
assign w34869 = ~w34867 & ~w34868;
assign w34870 = pi06972 & ~w18522;
assign w34871 = ~pi02170 & w18522;
assign w34872 = ~w34870 & ~w34871;
assign w34873 = pi06973 & ~w18568;
assign w34874 = ~pi02703 & w18568;
assign w34875 = ~w34873 & ~w34874;
assign w34876 = pi06974 & ~w18522;
assign w34877 = w17650 & w17929;
assign w34878 = ~w34876 & ~w34877;
assign w34879 = pi06975 & ~w18522;
assign w34880 = ~pi02714 & w18522;
assign w34881 = ~w34879 & ~w34880;
assign w34882 = pi06976 & ~w18568;
assign w34883 = ~pi02721 & w18568;
assign w34884 = ~w34882 & ~w34883;
assign w34885 = pi06977 & ~w18522;
assign w34886 = ~pi02715 & w18522;
assign w34887 = ~w34885 & ~w34886;
assign w34888 = pi06978 & ~w18568;
assign w34889 = ~pi02169 & w18568;
assign w34890 = ~w34888 & ~w34889;
assign w34891 = pi06979 & ~w18522;
assign w34892 = ~pi02717 & w18522;
assign w34893 = ~w34891 & ~w34892;
assign w34894 = pi06980 & ~w18623;
assign w34895 = ~pi02711 & w18623;
assign w34896 = ~w34894 & ~w34895;
assign w34897 = pi06981 & ~w18568;
assign w34898 = ~pi02718 & w18568;
assign w34899 = ~w34897 & ~w34898;
assign w34900 = pi06982 & ~w18623;
assign w34901 = w18622 & w20209;
assign w34902 = ~w34900 & ~w34901;
assign w34903 = pi06983 & ~w18623;
assign w34904 = w17929 & w18622;
assign w34905 = ~w34903 & ~w34904;
assign w34906 = pi06984 & ~w18623;
assign w34907 = w17742 & w18622;
assign w34908 = ~w34906 & ~w34907;
assign w34909 = pi06985 & ~w18623;
assign w34910 = w18059 & w18622;
assign w34911 = ~w34909 & ~w34910;
assign w34912 = pi06986 & ~w18623;
assign w34913 = w17317 & w18622;
assign w34914 = ~w34912 & ~w34913;
assign w34915 = pi06987 & ~w18568;
assign w34916 = ~pi02164 & w18568;
assign w34917 = ~w34915 & ~w34916;
assign w34918 = pi06988 & ~w18623;
assign w34919 = ~pi02717 & w18623;
assign w34920 = ~w34918 & ~w34919;
assign w34921 = pi06989 & ~w18568;
assign w34922 = ~pi02722 & w18568;
assign w34923 = ~w34921 & ~w34922;
assign w34924 = pi06990 & ~w18568;
assign w34925 = ~pi02719 & w18568;
assign w34926 = ~w34924 & ~w34925;
assign w34927 = pi06991 & ~w18283;
assign w34928 = ~pi02721 & w18283;
assign w34929 = ~w34927 & ~w34928;
assign w34930 = pi06992 & ~w18283;
assign w34931 = ~pi02169 & w18283;
assign w34932 = ~w34930 & ~w34931;
assign w34933 = pi06993 & ~w18127;
assign w34934 = ~pi02711 & w18127;
assign w34935 = ~w34933 & ~w34934;
assign w34936 = pi06994 & ~w18283;
assign w34937 = ~pi02718 & w18283;
assign w34938 = ~w34936 & ~w34937;
assign w34939 = pi06995 & ~w18127;
assign w34940 = ~pi02170 & w18127;
assign w34941 = ~w34939 & ~w34940;
assign w34942 = pi06996 & ~w18127;
assign w34943 = ~pi02713 & w18127;
assign w34944 = ~w34942 & ~w34943;
assign w34945 = pi06997 & ~w18283;
assign w34946 = w17344 & w19273;
assign w34947 = ~w34945 & ~w34946;
assign w34948 = pi06998 & ~w18127;
assign w34949 = ~pi02715 & w18127;
assign w34950 = ~w34948 & ~w34949;
assign w34951 = pi06999 & ~w18127;
assign w34952 = ~pi02716 & w18127;
assign w34953 = ~w34951 & ~w34952;
assign w34954 = pi07000 & ~w18283;
assign w34955 = ~pi02164 & w18283;
assign w34956 = ~w34954 & ~w34955;
assign w34957 = pi07001 & ~w18127;
assign w34958 = ~pi02717 & w18127;
assign w34959 = ~w34957 & ~w34958;
assign w34960 = pi07002 & ~w18283;
assign w34961 = ~pi02722 & w18283;
assign w34962 = ~w34960 & ~w34961;
assign w34963 = pi07003 & ~w18283;
assign w34964 = ~pi02719 & w18283;
assign w34965 = ~w34963 & ~w34964;
assign w34966 = pi07004 & ~w17702;
assign w34967 = ~pi02703 & w17702;
assign w34968 = ~w34966 & ~w34967;
assign w34969 = pi07005 & ~w17702;
assign w34970 = ~pi02721 & w17702;
assign w34971 = ~w34969 & ~w34970;
assign w34972 = pi07006 & ~w17702;
assign w34973 = ~pi02169 & w17702;
assign w34974 = ~w34972 & ~w34973;
assign w34975 = pi07007 & ~w17601;
assign w34976 = ~pi02712 & w17601;
assign w34977 = ~w34975 & ~w34976;
assign w34978 = pi07008 & ~w17702;
assign w34979 = ~pi02718 & w17702;
assign w34980 = ~w34978 & ~w34979;
assign w34981 = pi07009 & ~w17601;
assign w34982 = ~pi02170 & w17601;
assign w34983 = ~w34981 & ~w34982;
assign w34984 = pi07010 & ~w17702;
assign w34985 = ~pi02167 & w17702;
assign w34986 = ~w34984 & ~w34985;
assign w34987 = pi07011 & ~w17601;
assign w34988 = ~pi02714 & w17601;
assign w34989 = ~w34987 & ~w34988;
assign w34990 = pi07012 & ~w17601;
assign w34991 = ~pi02715 & w17601;
assign w34992 = ~w34990 & ~w34991;
assign w34993 = pi07013 & ~w17601;
assign w34994 = ~pi02716 & w17601;
assign w34995 = ~w34993 & ~w34994;
assign w34996 = pi07014 & ~w17601;
assign w34997 = ~pi02717 & w17601;
assign w34998 = ~w34996 & ~w34997;
assign w34999 = pi07015 & ~w17702;
assign w35000 = ~pi02164 & w17702;
assign w35001 = ~w34999 & ~w35000;
assign w35002 = pi07016 & ~w17702;
assign w35003 = ~pi02722 & w17702;
assign w35004 = ~w35002 & ~w35003;
assign w35005 = ~w16992 & w17244;
assign w35006 = pi07017 & ~w35005;
assign w35007 = ~pi02703 & w35005;
assign w35008 = ~w35006 & ~w35007;
assign w35009 = pi07018 & ~w35005;
assign w35010 = ~pi02721 & w35005;
assign w35011 = ~w35009 & ~w35010;
assign w35012 = pi07019 & ~w17376;
assign w35013 = ~pi02711 & w17376;
assign w35014 = ~w35012 & ~w35013;
assign w35015 = pi07020 & ~w35005;
assign w35016 = ~pi02169 & w35005;
assign w35017 = ~w35015 & ~w35016;
assign w35018 = pi07021 & ~w35005;
assign w35019 = ~pi02718 & w35005;
assign w35020 = ~w35018 & ~w35019;
assign w35021 = pi07022 & ~w17376;
assign w35022 = ~pi02170 & w17376;
assign w35023 = ~w35021 & ~w35022;
assign w35024 = pi07023 & ~w35005;
assign w35025 = w17244 & w19273;
assign w35026 = ~w35024 & ~w35025;
assign w35027 = pi07024 & ~w17376;
assign w35028 = ~pi02714 & w17376;
assign w35029 = ~w35027 & ~w35028;
assign w35030 = pi07025 & ~w17376;
assign w35031 = ~pi02715 & w17376;
assign w35032 = ~w35030 & ~w35031;
assign w35033 = pi07026 & ~w35005;
assign w35034 = ~pi02164 & w35005;
assign w35035 = ~w35033 & ~w35034;
assign w35036 = pi07027 & ~w17376;
assign w35037 = ~pi02716 & w17376;
assign w35038 = ~w35036 & ~w35037;
assign w35039 = pi07028 & ~w17376;
assign w35040 = ~pi02717 & w17376;
assign w35041 = ~w35039 & ~w35040;
assign w35042 = ~w16905 & w18731;
assign w35043 = pi07029 & ~w35042;
assign w35044 = ~pi02711 & w35042;
assign w35045 = ~w35043 & ~w35044;
assign w35046 = pi07030 & ~w35042;
assign w35047 = ~pi02712 & w35042;
assign w35048 = ~w35046 & ~w35047;
assign w35049 = pi07031 & ~w35042;
assign w35050 = ~pi02170 & w35042;
assign w35051 = ~w35049 & ~w35050;
assign w35052 = pi07032 & ~w35005;
assign w35053 = ~pi02719 & w35005;
assign w35054 = ~w35052 & ~w35053;
assign w35055 = pi07033 & ~w35042;
assign w35056 = ~pi02714 & w35042;
assign w35057 = ~w35055 & ~w35056;
assign w35058 = pi07034 & ~w35042;
assign w35059 = ~pi02715 & w35042;
assign w35060 = ~w35058 & ~w35059;
assign w35061 = pi07035 & ~w35042;
assign w35062 = ~pi02716 & w35042;
assign w35063 = ~w35061 & ~w35062;
assign w35064 = ~w16905 & w18683;
assign w35065 = pi07036 & ~w35064;
assign w35066 = w17603 & w18683;
assign w35067 = ~w35065 & ~w35066;
assign w35068 = pi07037 & ~w35064;
assign w35069 = w17020 & w18683;
assign w35070 = ~w35068 & ~w35069;
assign w35071 = pi07038 & ~w35064;
assign w35072 = ~pi02170 & w35064;
assign w35073 = ~w35071 & ~w35072;
assign w35074 = pi07039 & ~w35064;
assign w35075 = ~pi02713 & w35064;
assign w35076 = ~w35074 & ~w35075;
assign w35077 = pi07040 & ~w35064;
assign w35078 = ~pi02714 & w35064;
assign w35079 = ~w35077 & ~w35078;
assign w35080 = pi07041 & ~w35064;
assign w35081 = ~pi02715 & w35064;
assign w35082 = ~w35080 & ~w35081;
assign w35083 = pi07042 & ~w35064;
assign w35084 = ~pi02716 & w35064;
assign w35085 = ~w35083 & ~w35084;
assign w35086 = ~w16905 & w18348;
assign w35087 = pi07043 & ~w35086;
assign w35088 = w17603 & w18348;
assign w35089 = ~w35087 & ~w35088;
assign w35090 = pi07044 & ~w35086;
assign w35091 = ~pi02712 & w35086;
assign w35092 = ~w35090 & ~w35091;
assign w35093 = pi07045 & ~w35086;
assign w35094 = ~pi02170 & w35086;
assign w35095 = ~w35093 & ~w35094;
assign w35096 = pi07046 & ~w35086;
assign w35097 = ~pi02714 & w35086;
assign w35098 = ~w35096 & ~w35097;
assign w35099 = pi07047 & ~w35086;
assign w35100 = ~pi02715 & w35086;
assign w35101 = ~w35099 & ~w35100;
assign w35102 = ~w16992 & w19306;
assign w35103 = pi07048 & ~w35102;
assign w35104 = ~pi02703 & w35102;
assign w35105 = ~w35103 & ~w35104;
assign w35106 = pi07049 & ~w35086;
assign w35107 = ~pi02717 & w35086;
assign w35108 = ~w35106 & ~w35107;
assign w35109 = pi07050 & ~w35102;
assign w35110 = ~pi02721 & w35102;
assign w35111 = ~w35109 & ~w35110;
assign w35112 = ~w16905 & w17521;
assign w35113 = pi07051 & ~w35112;
assign w35114 = ~pi02711 & w35112;
assign w35115 = ~w35113 & ~w35114;
assign w35116 = pi07052 & ~w35112;
assign w35117 = ~pi02712 & w35112;
assign w35118 = ~w35116 & ~w35117;
assign w35119 = pi07053 & ~w35102;
assign w35120 = ~pi02169 & w35102;
assign w35121 = ~w35119 & ~w35120;
assign w35122 = pi07054 & ~w35112;
assign w35123 = ~pi02170 & w35112;
assign w35124 = ~w35122 & ~w35123;
assign w35125 = pi07055 & ~w35112;
assign w35126 = ~pi02713 & w35112;
assign w35127 = ~w35125 & ~w35126;
assign w35128 = pi07056 & ~w35112;
assign w35129 = w17521 & w17742;
assign w35130 = ~w35128 & ~w35129;
assign w35131 = pi07057 & ~w35112;
assign w35132 = ~pi02715 & w35112;
assign w35133 = ~w35131 & ~w35132;
assign w35134 = pi07058 & ~w35102;
assign w35135 = ~pi02167 & w35102;
assign w35136 = ~w35134 & ~w35135;
assign w35137 = pi07059 & ~w35112;
assign w35138 = ~pi02716 & w35112;
assign w35139 = ~w35137 & ~w35138;
assign w35140 = pi07060 & ~w35112;
assign w35141 = ~pi02717 & w35112;
assign w35142 = ~w35140 & ~w35141;
assign w35143 = pi07061 & ~w21456;
assign w35144 = ~pi02711 & w21456;
assign w35145 = ~w35143 & ~w35144;
assign w35146 = pi07062 & ~w21456;
assign w35147 = ~pi02712 & w21456;
assign w35148 = ~w35146 & ~w35147;
assign w35149 = pi07063 & ~w21456;
assign w35150 = ~pi02170 & w21456;
assign w35151 = ~w35149 & ~w35150;
assign w35152 = pi07064 & ~w35102;
assign w35153 = ~pi02719 & w35102;
assign w35154 = ~w35152 & ~w35153;
assign w35155 = pi07065 & ~w21456;
assign w35156 = w17325 & w17929;
assign w35157 = ~w35155 & ~w35156;
assign w35158 = pi07066 & ~w21456;
assign w35159 = ~pi02714 & w21456;
assign w35160 = ~w35158 & ~w35159;
assign w35161 = pi07067 & ~w21456;
assign w35162 = ~pi02715 & w21456;
assign w35163 = ~w35161 & ~w35162;
assign w35164 = pi07068 & ~w21456;
assign w35165 = ~pi02716 & w21456;
assign w35166 = ~w35164 & ~w35165;
assign w35167 = pi07069 & ~w21080;
assign w35168 = ~pi02711 & w21080;
assign w35169 = ~w35167 & ~w35168;
assign w35170 = pi07070 & ~w21080;
assign w35171 = ~pi02712 & w21080;
assign w35172 = ~w35170 & ~w35171;
assign w35173 = pi07071 & ~w21080;
assign w35174 = ~pi02170 & w21080;
assign w35175 = ~w35173 & ~w35174;
assign w35176 = pi07072 & ~w21080;
assign w35177 = w17474 & w17742;
assign w35178 = ~w35176 & ~w35177;
assign w35179 = pi07073 & ~w21080;
assign w35180 = ~pi02715 & w21080;
assign w35181 = ~w35179 & ~w35180;
assign w35182 = pi07074 & ~w21080;
assign w35183 = ~pi02716 & w21080;
assign w35184 = ~w35182 & ~w35183;
assign w35185 = pi07075 & ~w20442;
assign w35186 = ~pi02711 & w20442;
assign w35187 = ~w35185 & ~w35186;
assign w35188 = pi07076 & ~w20442;
assign w35189 = ~pi02712 & w20442;
assign w35190 = ~w35188 & ~w35189;
assign w35191 = pi07077 & ~w20442;
assign w35192 = ~pi02170 & w20442;
assign w35193 = ~w35191 & ~w35192;
assign w35194 = pi07078 & ~w20442;
assign w35195 = ~pi02713 & w20442;
assign w35196 = ~w35194 & ~w35195;
assign w35197 = pi07079 & ~w20442;
assign w35198 = ~pi02714 & w20442;
assign w35199 = ~w35197 & ~w35198;
assign w35200 = pi07080 & ~w20442;
assign w35201 = ~pi02715 & w20442;
assign w35202 = ~w35200 & ~w35201;
assign w35203 = pi07081 & ~w20442;
assign w35204 = ~pi02716 & w20442;
assign w35205 = ~w35203 & ~w35204;
assign w35206 = pi07082 & ~w20261;
assign w35207 = ~pi02711 & w20261;
assign w35208 = ~w35206 & ~w35207;
assign w35209 = pi07083 & ~w20261;
assign w35210 = w17020 & w17344;
assign w35211 = ~w35209 & ~w35210;
assign w35212 = pi07084 & ~w20261;
assign w35213 = w17344 & w20209;
assign w35214 = ~w35212 & ~w35213;
assign w35215 = pi07085 & ~w20261;
assign w35216 = ~pi02714 & w20261;
assign w35217 = ~w35215 & ~w35216;
assign w35218 = pi07086 & ~w20261;
assign w35219 = ~pi02715 & w20261;
assign w35220 = ~w35218 & ~w35219;
assign w35221 = pi07087 & ~w20261;
assign w35222 = w17317 & w17344;
assign w35223 = ~w35221 & ~w35222;
assign w35224 = pi07088 & ~w20337;
assign w35225 = ~pi02711 & w20337;
assign w35226 = ~w35224 & ~w35225;
assign w35227 = pi07089 & ~w20337;
assign w35228 = ~pi02712 & w20337;
assign w35229 = ~w35227 & ~w35228;
assign w35230 = pi07090 & ~w20337;
assign w35231 = ~pi02170 & w20337;
assign w35232 = ~w35230 & ~w35231;
assign w35233 = pi07091 & ~w20337;
assign w35234 = ~pi02713 & w20337;
assign w35235 = ~w35233 & ~w35234;
assign w35236 = pi07092 & ~w20337;
assign w35237 = ~pi02714 & w20337;
assign w35238 = ~w35236 & ~w35237;
assign w35239 = pi07093 & ~w20200;
assign w35240 = ~pi02703 & w20200;
assign w35241 = ~w35239 & ~w35240;
assign w35242 = pi07094 & ~w20337;
assign w35243 = w17162 & w18059;
assign w35244 = ~w35242 & ~w35243;
assign w35245 = pi07095 & ~w20200;
assign w35246 = ~pi02721 & w20200;
assign w35247 = ~w35245 & ~w35246;
assign w35248 = pi07096 & ~w20337;
assign w35249 = ~pi02717 & w20337;
assign w35250 = ~w35248 & ~w35249;
assign w35251 = pi07097 & ~w20330;
assign w35252 = w17244 & w17603;
assign w35253 = ~w35251 & ~w35252;
assign w35254 = pi07098 & ~w20330;
assign w35255 = ~pi02170 & w20330;
assign w35256 = ~w35254 & ~w35255;
assign w35257 = pi07099 & ~w20200;
assign w35258 = ~pi02169 & w20200;
assign w35259 = ~w35257 & ~w35258;
assign w35260 = pi07100 & ~w20330;
assign w35261 = ~pi02713 & w20330;
assign w35262 = ~w35260 & ~w35261;
assign w35263 = pi07101 & ~w20330;
assign w35264 = w17244 & w17742;
assign w35265 = ~w35263 & ~w35264;
assign w35266 = pi07102 & ~w20330;
assign w35267 = ~pi02715 & w20330;
assign w35268 = ~w35266 & ~w35267;
assign w35269 = pi07103 & ~w20200;
assign w35270 = ~pi02167 & w20200;
assign w35271 = ~w35269 & ~w35270;
assign w35272 = pi07104 & ~w20330;
assign w35273 = ~pi02716 & w20330;
assign w35274 = ~w35272 & ~w35273;
assign w35275 = pi07105 & ~w20330;
assign w35276 = ~pi02717 & w20330;
assign w35277 = ~w35275 & ~w35276;
assign w35278 = pi07106 & ~w20200;
assign w35279 = ~pi02164 & w20200;
assign w35280 = ~w35278 & ~w35279;
assign w35281 = pi07107 & ~w20200;
assign w35282 = ~pi02722 & w20200;
assign w35283 = ~w35281 & ~w35282;
assign w35284 = pi07108 & ~w18086;
assign w35285 = ~pi02703 & w18086;
assign w35286 = ~w35284 & ~w35285;
assign w35287 = pi07109 & ~w19307;
assign w35288 = ~pi02711 & w19307;
assign w35289 = ~w35287 & ~w35288;
assign w35290 = pi07110 & ~w18086;
assign w35291 = ~pi02721 & w18086;
assign w35292 = ~w35290 & ~w35291;
assign w35293 = pi07111 & ~w18086;
assign w35294 = w17739 & w19797;
assign w35295 = ~w35293 & ~w35294;
assign w35296 = pi07112 & ~w19307;
assign w35297 = ~pi02170 & w19307;
assign w35298 = ~w35296 & ~w35297;
assign w35299 = pi07113 & ~w19307;
assign w35300 = ~pi02713 & w19307;
assign w35301 = ~w35299 & ~w35300;
assign w35302 = pi07114 & ~w18086;
assign w35303 = ~pi02718 & w18086;
assign w35304 = ~w35302 & ~w35303;
assign w35305 = pi07115 & ~w19307;
assign w35306 = ~pi02715 & w19307;
assign w35307 = ~w35305 & ~w35306;
assign w35308 = pi07116 & ~w19307;
assign w35309 = ~pi02716 & w19307;
assign w35310 = ~w35308 & ~w35309;
assign w35311 = pi07117 & ~w18086;
assign w35312 = ~pi02167 & w18086;
assign w35313 = ~w35311 & ~w35312;
assign w35314 = pi07118 & ~w19307;
assign w35315 = ~pi02717 & w19307;
assign w35316 = ~w35314 & ~w35315;
assign w35317 = pi07119 & ~w18086;
assign w35318 = ~pi02164 & w18086;
assign w35319 = ~w35317 & ~w35318;
assign w35320 = pi07120 & ~w18086;
assign w35321 = ~pi02722 & w18086;
assign w35322 = ~w35320 & ~w35321;
assign w35323 = pi07121 & ~w18492;
assign w35324 = ~pi02703 & w18492;
assign w35325 = ~w35323 & ~w35324;
assign w35326 = pi07122 & ~w18492;
assign w35327 = ~pi02721 & w18492;
assign w35328 = ~w35326 & ~w35327;
assign w35329 = pi07123 & ~w18492;
assign w35330 = ~pi02169 & w18492;
assign w35331 = ~w35329 & ~w35330;
assign w35332 = pi07124 & ~w18492;
assign w35333 = w16986 & w19273;
assign w35334 = ~w35332 & ~w35333;
assign w35335 = pi07125 & ~w18218;
assign w35336 = ~pi02711 & w18218;
assign w35337 = ~w35335 & ~w35336;
assign w35338 = pi07126 & ~w18492;
assign w35339 = ~pi02164 & w18492;
assign w35340 = ~w35338 & ~w35339;
assign w35341 = pi07127 & ~w18218;
assign w35342 = ~pi02170 & w18218;
assign w35343 = ~w35341 & ~w35342;
assign w35344 = pi07128 & ~w18492;
assign w35345 = ~pi02722 & w18492;
assign w35346 = ~w35344 & ~w35345;
assign w35347 = pi07129 & ~w18218;
assign w35348 = w17929 & w18217;
assign w35349 = ~w35347 & ~w35348;
assign w35350 = pi07130 & ~w18218;
assign w35351 = ~pi02714 & w18218;
assign w35352 = ~w35350 & ~w35351;
assign w35353 = pi07131 & ~w18492;
assign w35354 = ~pi02719 & w18492;
assign w35355 = ~w35353 & ~w35354;
assign w35356 = pi07132 & ~w18218;
assign w35357 = ~pi02715 & w18218;
assign w35358 = ~w35356 & ~w35357;
assign w35359 = pi07133 & ~w18218;
assign w35360 = ~pi02716 & w18218;
assign w35361 = ~w35359 & ~w35360;
assign w35362 = pi07134 & ~w18218;
assign w35363 = ~pi02717 & w18218;
assign w35364 = ~w35362 & ~w35363;
assign w35365 = pi07135 & ~w17740;
assign w35366 = ~pi02711 & w17740;
assign w35367 = ~w35365 & ~w35366;
assign w35368 = pi07136 & ~w17740;
assign w35369 = ~pi02712 & w17740;
assign w35370 = ~w35368 & ~w35369;
assign w35371 = pi07137 & ~w17740;
assign w35372 = ~pi02170 & w17740;
assign w35373 = ~w35371 & ~w35372;
assign w35374 = pi07138 & ~w17740;
assign w35375 = ~pi02713 & w17740;
assign w35376 = ~w35374 & ~w35375;
assign w35377 = pi07139 & ~w17695;
assign w35378 = w17694 & w19797;
assign w35379 = ~w35377 & ~w35378;
assign w35380 = pi07140 & ~w17695;
assign w35381 = ~pi02718 & w17695;
assign w35382 = ~w35380 & ~w35381;
assign w35383 = pi07141 & ~w17740;
assign w35384 = ~pi02715 & w17740;
assign w35385 = ~w35383 & ~w35384;
assign w35386 = pi07142 & ~w17695;
assign w35387 = ~pi02167 & w17695;
assign w35388 = ~w35386 & ~w35387;
assign w35389 = pi07143 & ~w17740;
assign w35390 = ~pi02716 & w17740;
assign w35391 = ~w35389 & ~w35390;
assign w35392 = pi07144 & ~w17740;
assign w35393 = ~pi02717 & w17740;
assign w35394 = ~w35392 & ~w35393;
assign w35395 = pi07145 & ~w16987;
assign w35396 = ~pi02711 & w16987;
assign w35397 = ~w35395 & ~w35396;
assign w35398 = pi07146 & ~w16987;
assign w35399 = ~pi02712 & w16987;
assign w35400 = ~w35398 & ~w35399;
assign w35401 = pi07147 & ~w16987;
assign w35402 = ~pi02170 & w16987;
assign w35403 = ~w35401 & ~w35402;
assign w35404 = pi07148 & ~w17695;
assign w35405 = ~pi02722 & w17695;
assign w35406 = ~w35404 & ~w35405;
assign w35407 = pi07149 & ~w16987;
assign w35408 = ~pi02713 & w16987;
assign w35409 = ~w35407 & ~w35408;
assign w35410 = pi07150 & ~w16987;
assign w35411 = ~pi02715 & w16987;
assign w35412 = ~w35410 & ~w35411;
assign w35413 = pi07151 & ~w17695;
assign w35414 = ~pi02719 & w17695;
assign w35415 = ~w35413 & ~w35414;
assign w35416 = pi07152 & ~w16987;
assign w35417 = ~pi02716 & w16987;
assign w35418 = ~w35416 & ~w35417;
assign w35419 = ~w16905 & w17694;
assign w35420 = pi07153 & ~w35419;
assign w35421 = ~pi02711 & w35419;
assign w35422 = ~w35420 & ~w35421;
assign w35423 = pi07154 & ~w35419;
assign w35424 = ~pi02712 & w35419;
assign w35425 = ~w35423 & ~w35424;
assign w35426 = pi07155 & ~w35419;
assign w35427 = ~pi02170 & w35419;
assign w35428 = ~w35426 & ~w35427;
assign w35429 = pi07156 & ~w35419;
assign w35430 = ~pi02713 & w35419;
assign w35431 = ~w35429 & ~w35430;
assign w35432 = pi07157 & ~w35419;
assign w35433 = ~pi02714 & w35419;
assign w35434 = ~w35432 & ~w35433;
assign w35435 = pi07158 & ~w35419;
assign w35436 = ~pi02715 & w35419;
assign w35437 = ~w35435 & ~w35436;
assign w35438 = pi07159 & ~w35419;
assign w35439 = w17317 & w17694;
assign w35440 = ~w35438 & ~w35439;
assign w35441 = ~w16905 & w20923;
assign w35442 = pi07160 & ~w35441;
assign w35443 = ~pi02711 & w35441;
assign w35444 = ~w35442 & ~w35443;
assign w35445 = pi07161 & ~w35441;
assign w35446 = w17020 & w20923;
assign w35447 = ~w35445 & ~w35446;
assign w35448 = pi07162 & ~w35441;
assign w35449 = w20209 & w20923;
assign w35450 = ~w35448 & ~w35449;
assign w35451 = pi07163 & ~w35441;
assign w35452 = ~pi02714 & w35441;
assign w35453 = ~w35451 & ~w35452;
assign w35454 = pi07164 & ~w35441;
assign w35455 = ~pi02715 & w35441;
assign w35456 = ~w35454 & ~w35455;
assign w35457 = pi07165 & ~w35441;
assign w35458 = ~pi02716 & w35441;
assign w35459 = ~w35457 & ~w35458;
assign w35460 = pi07166 & ~w35441;
assign w35461 = ~pi02717 & w35441;
assign w35462 = ~w35460 & ~w35461;
assign w35463 = ~w16992 & w20923;
assign w35464 = pi07167 & ~w35463;
assign w35465 = ~pi02721 & w35463;
assign w35466 = ~w35464 & ~w35465;
assign w35467 = pi07168 & ~w35463;
assign w35468 = w19797 & w20923;
assign w35469 = ~w35467 & ~w35468;
assign w35470 = pi07169 & ~w35463;
assign w35471 = w17586 & w20923;
assign w35472 = ~w35470 & ~w35471;
assign w35473 = ~w16905 & w17148;
assign w35474 = pi07170 & ~w35473;
assign w35475 = ~pi02711 & w35473;
assign w35476 = ~w35474 & ~w35475;
assign w35477 = pi07171 & ~w35463;
assign w35478 = ~pi02167 & w35463;
assign w35479 = ~w35477 & ~w35478;
assign w35480 = pi07172 & ~w35473;
assign w35481 = ~pi02712 & w35473;
assign w35482 = ~w35480 & ~w35481;
assign w35483 = pi07173 & ~w35463;
assign w35484 = ~pi02164 & w35463;
assign w35485 = ~w35483 & ~w35484;
assign w35486 = pi07174 & ~w35473;
assign w35487 = ~pi02713 & w35473;
assign w35488 = ~w35486 & ~w35487;
assign w35489 = pi07175 & ~w35463;
assign w35490 = ~pi02722 & w35463;
assign w35491 = ~w35489 & ~w35490;
assign w35492 = pi07176 & ~w35463;
assign w35493 = ~pi02719 & w35463;
assign w35494 = ~w35492 & ~w35493;
assign w35495 = pi07177 & ~w35473;
assign w35496 = ~pi02715 & w35473;
assign w35497 = ~w35495 & ~w35496;
assign w35498 = pi07178 & ~w35473;
assign w35499 = ~pi02716 & w35473;
assign w35500 = ~w35498 & ~w35499;
assign w35501 = ~w16905 & w18563;
assign w35502 = pi07179 & ~w35501;
assign w35503 = w17603 & w18563;
assign w35504 = ~w35502 & ~w35503;
assign w35505 = pi07180 & ~w35501;
assign w35506 = ~pi02712 & w35501;
assign w35507 = ~w35505 & ~w35506;
assign w35508 = pi07181 & ~w35501;
assign w35509 = ~pi02170 & w35501;
assign w35510 = ~w35508 & ~w35509;
assign w35511 = pi07182 & ~w35501;
assign w35512 = ~pi02713 & w35501;
assign w35513 = ~w35511 & ~w35512;
assign w35514 = pi07183 & ~w35501;
assign w35515 = w17742 & w18563;
assign w35516 = ~w35514 & ~w35515;
assign w35517 = pi07184 & ~w35501;
assign w35518 = ~pi02715 & w35501;
assign w35519 = ~w35517 & ~w35518;
assign w35520 = pi07185 & ~w35501;
assign w35521 = w17317 & w18563;
assign w35522 = ~w35520 & ~w35521;
assign w35523 = pi07186 & ~w21285;
assign w35524 = ~pi02711 & w21285;
assign w35525 = ~w35523 & ~w35524;
assign w35526 = pi07187 & ~w21285;
assign w35527 = ~pi02712 & w21285;
assign w35528 = ~w35526 & ~w35527;
assign w35529 = pi07188 & ~w21285;
assign w35530 = ~pi02170 & w21285;
assign w35531 = ~w35529 & ~w35530;
assign w35532 = pi07189 & ~w21285;
assign w35533 = ~pi02714 & w21285;
assign w35534 = ~w35532 & ~w35533;
assign w35535 = pi07190 & ~w21285;
assign w35536 = ~pi02715 & w21285;
assign w35537 = ~w35535 & ~w35536;
assign w35538 = pi07191 & ~w21285;
assign w35539 = ~pi02716 & w21285;
assign w35540 = ~w35538 & ~w35539;
assign w35541 = pi07192 & ~w21285;
assign w35542 = ~pi02717 & w21285;
assign w35543 = ~w35541 & ~w35542;
assign w35544 = pi07193 & ~w21277;
assign w35545 = ~pi02711 & w21277;
assign w35546 = ~w35544 & ~w35545;
assign w35547 = pi07194 & ~w21277;
assign w35548 = ~pi02712 & w21277;
assign w35549 = ~w35547 & ~w35548;
assign w35550 = pi07195 & ~w21277;
assign w35551 = ~pi02170 & w21277;
assign w35552 = ~w35550 & ~w35551;
assign w35553 = pi07196 & ~w21555;
assign w35554 = ~pi02721 & w21555;
assign w35555 = ~w35553 & ~w35554;
assign w35556 = pi07197 & ~w21277;
assign w35557 = ~pi02713 & w21277;
assign w35558 = ~w35556 & ~w35557;
assign w35559 = pi07198 & ~w21555;
assign w35560 = w17148 & w19797;
assign w35561 = ~w35559 & ~w35560;
assign w35562 = pi07199 & ~w21277;
assign w35563 = w18059 & w18781;
assign w35564 = ~w35562 & ~w35563;
assign w35565 = pi07200 & ~w21277;
assign w35566 = ~pi02716 & w21277;
assign w35567 = ~w35565 & ~w35566;
assign w35568 = pi07201 & ~w21555;
assign w35569 = ~pi02718 & w21555;
assign w35570 = ~w35568 & ~w35569;
assign w35571 = pi07202 & ~w21555;
assign w35572 = ~pi02167 & w21555;
assign w35573 = ~w35571 & ~w35572;
assign w35574 = pi07203 & ~w21555;
assign w35575 = ~pi02164 & w21555;
assign w35576 = ~w35574 & ~w35575;
assign w35577 = pi07204 & ~w21555;
assign w35578 = ~pi02722 & w21555;
assign w35579 = ~w35577 & ~w35578;
assign w35580 = pi07205 & ~w21548;
assign w35581 = ~pi02711 & w21548;
assign w35582 = ~w35580 & ~w35581;
assign w35583 = pi07206 & ~w21548;
assign w35584 = ~pi02712 & w21548;
assign w35585 = ~w35583 & ~w35584;
assign w35586 = pi07207 & ~w21544;
assign w35587 = ~pi02703 & w21544;
assign w35588 = ~w35586 & ~w35587;
assign w35589 = pi07208 & ~w21548;
assign w35590 = ~pi02170 & w21548;
assign w35591 = ~w35589 & ~w35590;
assign w35592 = pi07209 & ~w21544;
assign w35593 = ~pi02721 & w21544;
assign w35594 = ~w35592 & ~w35593;
assign w35595 = pi07210 & ~w21548;
assign w35596 = ~pi02713 & w21548;
assign w35597 = ~w35595 & ~w35596;
assign w35598 = pi07211 & ~w21544;
assign w35599 = ~pi02169 & w21544;
assign w35600 = ~w35598 & ~w35599;
assign w35601 = pi07212 & ~w21548;
assign w35602 = ~pi02715 & w21548;
assign w35603 = ~w35601 & ~w35602;
assign w35604 = pi07213 & ~w21548;
assign w35605 = ~pi02716 & w21548;
assign w35606 = ~w35604 & ~w35605;
assign w35607 = pi07214 & ~w21544;
assign w35608 = ~pi02718 & w21544;
assign w35609 = ~w35607 & ~w35608;
assign w35610 = pi07215 & ~w21544;
assign w35611 = ~pi02167 & w21544;
assign w35612 = ~w35610 & ~w35611;
assign w35613 = pi07216 & ~w21544;
assign w35614 = ~pi02164 & w21544;
assign w35615 = ~w35613 & ~w35614;
assign w35616 = pi07217 & ~w21544;
assign w35617 = ~pi02722 & w21544;
assign w35618 = ~w35616 & ~w35617;
assign w35619 = ~w16905 & w18449;
assign w35620 = pi07218 & ~w35619;
assign w35621 = ~pi02711 & w35619;
assign w35622 = ~w35620 & ~w35621;
assign w35623 = pi07219 & ~w35619;
assign w35624 = ~pi02712 & w35619;
assign w35625 = ~w35623 & ~w35624;
assign w35626 = pi07220 & ~w21041;
assign w35627 = ~pi02703 & w21041;
assign w35628 = ~w35626 & ~w35627;
assign w35629 = pi07221 & ~w35619;
assign w35630 = ~pi02170 & w35619;
assign w35631 = ~w35629 & ~w35630;
assign w35632 = pi07222 & ~w35619;
assign w35633 = ~pi02713 & w35619;
assign w35634 = ~w35632 & ~w35633;
assign w35635 = pi07223 & ~w21041;
assign w35636 = ~pi02721 & w21041;
assign w35637 = ~w35635 & ~w35636;
assign w35638 = pi07224 & ~w35619;
assign w35639 = ~pi02714 & w35619;
assign w35640 = ~w35638 & ~w35639;
assign w35641 = pi07225 & ~w35619;
assign w35642 = ~pi02715 & w35619;
assign w35643 = ~w35641 & ~w35642;
assign w35644 = pi07226 & ~w35619;
assign w35645 = ~pi02716 & w35619;
assign w35646 = ~w35644 & ~w35645;
assign w35647 = pi07227 & ~w35619;
assign w35648 = ~pi02717 & w35619;
assign w35649 = ~w35647 & ~w35648;
assign w35650 = pi07228 & ~w21041;
assign w35651 = ~pi02167 & w21041;
assign w35652 = ~w35650 & ~w35651;
assign w35653 = pi07229 & ~w21041;
assign w35654 = ~pi02164 & w21041;
assign w35655 = ~w35653 & ~w35654;
assign w35656 = pi07230 & ~w21041;
assign w35657 = w18813 & w19312;
assign w35658 = ~w35656 & ~w35657;
assign w35659 = pi07231 & ~w19541;
assign w35660 = w17153 & w17603;
assign w35661 = ~w35659 & ~w35660;
assign w35662 = pi07232 & ~w19541;
assign w35663 = ~pi02712 & w19541;
assign w35664 = ~w35662 & ~w35663;
assign w35665 = ~w16992 & w18781;
assign w35666 = pi07233 & ~w35665;
assign w35667 = ~pi02703 & w35665;
assign w35668 = ~w35666 & ~w35667;
assign w35669 = pi07234 & ~w35665;
assign w35670 = w17811 & w18781;
assign w35671 = ~w35669 & ~w35670;
assign w35672 = pi07235 & ~w19541;
assign w35673 = ~pi02170 & w19541;
assign w35674 = ~w35672 & ~w35673;
assign w35675 = pi07236 & ~w19541;
assign w35676 = ~pi02713 & w19541;
assign w35677 = ~w35675 & ~w35676;
assign w35678 = pi07237 & ~w19541;
assign w35679 = ~pi02714 & w19541;
assign w35680 = ~w35678 & ~w35679;
assign w35681 = pi07238 & ~w35665;
assign w35682 = ~pi02169 & w35665;
assign w35683 = ~w35681 & ~w35682;
assign w35684 = pi07239 & ~w35665;
assign w35685 = ~pi02718 & w35665;
assign w35686 = ~w35684 & ~w35685;
assign w35687 = pi07240 & ~w19541;
assign w35688 = ~pi02716 & w19541;
assign w35689 = ~w35687 & ~w35688;
assign w35690 = pi07241 & ~w20222;
assign w35691 = ~pi02711 & w20222;
assign w35692 = ~w35690 & ~w35691;
assign w35693 = pi07242 & ~w35665;
assign w35694 = ~pi02167 & w35665;
assign w35695 = ~w35693 & ~w35694;
assign w35696 = pi07243 & ~w20222;
assign w35697 = ~pi02712 & w20222;
assign w35698 = ~w35696 & ~w35697;
assign w35699 = pi07244 & ~w35665;
assign w35700 = ~pi02722 & w35665;
assign w35701 = ~w35699 & ~w35700;
assign w35702 = pi07245 & ~w20222;
assign w35703 = ~pi02713 & w20222;
assign w35704 = ~w35702 & ~w35703;
assign w35705 = pi07246 & ~w20222;
assign w35706 = ~pi02714 & w20222;
assign w35707 = ~w35705 & ~w35706;
assign w35708 = pi07247 & ~w20222;
assign w35709 = ~pi02715 & w20222;
assign w35710 = ~w35708 & ~w35709;
assign w35711 = pi07248 & ~w20222;
assign w35712 = ~pi02716 & w20222;
assign w35713 = ~w35711 & ~w35712;
assign w35714 = pi07249 & ~w35665;
assign w35715 = ~pi02164 & w35665;
assign w35716 = ~w35714 & ~w35715;
assign w35717 = pi07250 & ~w20222;
assign w35718 = ~pi02717 & w20222;
assign w35719 = ~w35717 & ~w35718;
assign w35720 = pi07251 & ~w19485;
assign w35721 = ~pi02712 & w19485;
assign w35722 = ~w35720 & ~w35721;
assign w35723 = pi07252 & ~w35665;
assign w35724 = ~pi02719 & w35665;
assign w35725 = ~w35723 & ~w35724;
assign w35726 = pi07253 & ~w19485;
assign w35727 = ~pi02170 & w19485;
assign w35728 = ~w35726 & ~w35727;
assign w35729 = pi07254 & ~w19485;
assign w35730 = ~pi02714 & w19485;
assign w35731 = ~w35729 & ~w35730;
assign w35732 = pi07255 & ~w19485;
assign w35733 = ~pi02715 & w19485;
assign w35734 = ~w35732 & ~w35733;
assign w35735 = pi07256 & ~w19485;
assign w35736 = w17317 & w17339;
assign w35737 = ~w35735 & ~w35736;
assign w35738 = pi07257 & ~w17646;
assign w35739 = ~pi02703 & w17646;
assign w35740 = ~w35738 & ~w35739;
assign w35741 = pi07258 & ~w17646;
assign w35742 = ~pi02721 & w17646;
assign w35743 = ~w35741 & ~w35742;
assign w35744 = pi07259 & ~w17646;
assign w35745 = ~pi02169 & w17646;
assign w35746 = ~w35744 & ~w35745;
assign w35747 = pi07260 & ~w18418;
assign w35748 = ~pi02711 & w18418;
assign w35749 = ~w35747 & ~w35748;
assign w35750 = pi07261 & ~w17646;
assign w35751 = ~pi02718 & w17646;
assign w35752 = ~w35750 & ~w35751;
assign w35753 = pi07262 & ~w18418;
assign w35754 = ~pi02712 & w18418;
assign w35755 = ~w35753 & ~w35754;
assign w35756 = pi07263 & ~w18418;
assign w35757 = w17300 & w20209;
assign w35758 = ~w35756 & ~w35757;
assign w35759 = pi07264 & ~w17646;
assign w35760 = ~pi02164 & w17646;
assign w35761 = ~w35759 & ~w35760;
assign w35762 = pi07265 & ~w18418;
assign w35763 = ~pi02713 & w18418;
assign w35764 = ~w35762 & ~w35763;
assign w35765 = pi07266 & ~w18418;
assign w35766 = ~pi02714 & w18418;
assign w35767 = ~w35765 & ~w35766;
assign w35768 = pi07267 & ~w18418;
assign w35769 = ~pi02715 & w18418;
assign w35770 = ~w35768 & ~w35769;
assign w35771 = pi07268 & ~w18418;
assign w35772 = ~pi02716 & w18418;
assign w35773 = ~w35771 & ~w35772;
assign w35774 = pi07269 & ~w21488;
assign w35775 = ~pi02704 & w21488;
assign w35776 = ~w35774 & ~w35775;
assign w35777 = pi07270 & ~w18229;
assign w35778 = ~pi02711 & w18229;
assign w35779 = ~w35777 & ~w35778;
assign w35780 = pi07271 & ~w17646;
assign w35781 = ~pi02719 & w17646;
assign w35782 = ~w35780 & ~w35781;
assign w35783 = pi07272 & ~w18229;
assign w35784 = ~pi02712 & w18229;
assign w35785 = ~w35783 & ~w35784;
assign w35786 = pi07273 & ~w18229;
assign w35787 = ~pi02170 & w18229;
assign w35788 = ~w35786 & ~w35787;
assign w35789 = pi07274 & ~w18229;
assign w35790 = ~pi02713 & w18229;
assign w35791 = ~w35789 & ~w35790;
assign w35792 = pi07275 & ~w18229;
assign w35793 = ~pi02714 & w18229;
assign w35794 = ~w35792 & ~w35793;
assign w35795 = pi07276 & ~w18229;
assign w35796 = ~pi02715 & w18229;
assign w35797 = ~w35795 & ~w35796;
assign w35798 = pi07277 & ~w18229;
assign w35799 = ~pi02717 & w18229;
assign w35800 = ~w35798 & ~w35799;
assign w35801 = pi07278 & ~w18079;
assign w35802 = ~pi02711 & w18079;
assign w35803 = ~w35801 & ~w35802;
assign w35804 = pi07279 & ~w18079;
assign w35805 = ~pi02712 & w18079;
assign w35806 = ~w35804 & ~w35805;
assign w35807 = pi07280 & ~w18079;
assign w35808 = ~pi02713 & w18079;
assign w35809 = ~w35807 & ~w35808;
assign w35810 = pi07281 & ~w18079;
assign w35811 = ~pi02714 & w18079;
assign w35812 = ~w35810 & ~w35811;
assign w35813 = pi07282 & ~w18079;
assign w35814 = ~pi02715 & w18079;
assign w35815 = ~w35813 & ~w35814;
assign w35816 = pi07283 & ~w18079;
assign w35817 = ~pi02717 & w18079;
assign w35818 = ~w35816 & ~w35817;
assign w35819 = pi07284 & ~w17961;
assign w35820 = ~pi02711 & w17961;
assign w35821 = ~w35819 & ~w35820;
assign w35822 = pi07285 & ~w17961;
assign w35823 = w17020 & w17663;
assign w35824 = ~w35822 & ~w35823;
assign w35825 = ~w16992 & w18449;
assign w35826 = pi07286 & ~w35825;
assign w35827 = ~pi02703 & w35825;
assign w35828 = ~w35826 & ~w35827;
assign w35829 = pi07287 & ~w35825;
assign w35830 = ~pi02721 & w35825;
assign w35831 = ~w35829 & ~w35830;
assign w35832 = pi07288 & ~w17961;
assign w35833 = ~pi02170 & w17961;
assign w35834 = ~w35832 & ~w35833;
assign w35835 = pi07289 & ~w17961;
assign w35836 = w17663 & w17929;
assign w35837 = ~w35835 & ~w35836;
assign w35838 = pi07290 & ~w17961;
assign w35839 = ~pi02715 & w17961;
assign w35840 = ~w35838 & ~w35839;
assign w35841 = pi07291 & ~w35825;
assign w35842 = ~pi02169 & w35825;
assign w35843 = ~w35841 & ~w35842;
assign w35844 = pi07292 & ~w17961;
assign w35845 = ~pi02716 & w17961;
assign w35846 = ~w35844 & ~w35845;
assign w35847 = pi07293 & ~w17682;
assign w35848 = ~pi02711 & w17682;
assign w35849 = ~w35847 & ~w35848;
assign w35850 = pi07294 & ~w35825;
assign w35851 = ~pi02718 & w35825;
assign w35852 = ~w35850 & ~w35851;
assign w35853 = pi07295 & ~w17682;
assign w35854 = ~pi02712 & w17682;
assign w35855 = ~w35853 & ~w35854;
assign w35856 = pi07296 & ~w35825;
assign w35857 = ~pi02164 & w35825;
assign w35858 = ~w35856 & ~w35857;
assign w35859 = pi07297 & ~w17682;
assign w35860 = ~pi02713 & w17682;
assign w35861 = ~w35859 & ~w35860;
assign w35862 = pi07298 & ~w17682;
assign w35863 = ~pi02714 & w17682;
assign w35864 = ~w35862 & ~w35863;
assign w35865 = pi07299 & ~w17682;
assign w35866 = ~pi02715 & w17682;
assign w35867 = ~w35865 & ~w35866;
assign w35868 = pi07300 & ~w17682;
assign w35869 = ~pi02716 & w17682;
assign w35870 = ~w35868 & ~w35869;
assign w35871 = pi07301 & ~w35825;
assign w35872 = ~pi02167 & w35825;
assign w35873 = ~w35871 & ~w35872;
assign w35874 = pi07302 & ~w35825;
assign w35875 = ~pi02719 & w35825;
assign w35876 = ~w35874 & ~w35875;
assign w35877 = pi07303 & ~w17750;
assign w35878 = ~pi02711 & w17750;
assign w35879 = ~w35877 & ~w35878;
assign w35880 = pi07304 & ~w17750;
assign w35881 = ~pi02712 & w17750;
assign w35882 = ~w35880 & ~w35881;
assign w35883 = pi07305 & ~w35825;
assign w35884 = ~pi02722 & w35825;
assign w35885 = ~w35883 & ~w35884;
assign w35886 = pi07306 & ~w17750;
assign w35887 = ~pi02713 & w17750;
assign w35888 = ~w35886 & ~w35887;
assign w35889 = pi07307 & ~w17750;
assign w35890 = ~pi02714 & w17750;
assign w35891 = ~w35889 & ~w35890;
assign w35892 = pi07308 & ~w17750;
assign w35893 = ~pi02715 & w17750;
assign w35894 = ~w35892 & ~w35893;
assign w35895 = pi07309 & ~w17750;
assign w35896 = ~pi02717 & w17750;
assign w35897 = ~w35895 & ~w35896;
assign w35898 = pi07310 & ~w17659;
assign w35899 = w17603 & w17658;
assign w35900 = ~w35898 & ~w35899;
assign w35901 = pi07311 & ~w17659;
assign w35902 = w17020 & w17658;
assign w35903 = ~w35901 & ~w35902;
assign w35904 = pi07312 & ~w17659;
assign w35905 = ~pi02170 & w17659;
assign w35906 = ~w35904 & ~w35905;
assign w35907 = pi07313 & ~w17659;
assign w35908 = ~pi02713 & w17659;
assign w35909 = ~w35907 & ~w35908;
assign w35910 = pi07314 & ~w17659;
assign w35911 = ~pi02714 & w17659;
assign w35912 = ~w35910 & ~w35911;
assign w35913 = pi07315 & ~w17659;
assign w35914 = ~pi02715 & w17659;
assign w35915 = ~w35913 & ~w35914;
assign w35916 = pi07316 & ~w17659;
assign w35917 = ~pi02717 & w17659;
assign w35918 = ~w35916 & ~w35917;
assign w35919 = ~w16905 & w20561;
assign w35920 = pi07317 & ~w35919;
assign w35921 = w17603 & w20561;
assign w35922 = ~w35920 & ~w35921;
assign w35923 = pi07318 & ~w35919;
assign w35924 = ~pi02712 & w35919;
assign w35925 = ~w35923 & ~w35924;
assign w35926 = pi07319 & ~w35919;
assign w35927 = ~pi02713 & w35919;
assign w35928 = ~w35926 & ~w35927;
assign w35929 = ~w16992 & w17153;
assign w35930 = pi07320 & ~w35929;
assign w35931 = ~pi02703 & w35929;
assign w35932 = ~w35930 & ~w35931;
assign w35933 = pi07321 & ~w35919;
assign w35934 = ~pi02714 & w35919;
assign w35935 = ~w35933 & ~w35934;
assign w35936 = pi07322 & ~w35919;
assign w35937 = ~pi02715 & w35919;
assign w35938 = ~w35936 & ~w35937;
assign w35939 = pi07323 & ~w35919;
assign w35940 = ~pi02716 & w35919;
assign w35941 = ~w35939 & ~w35940;
assign w35942 = pi07324 & ~w35929;
assign w35943 = ~pi02169 & w35929;
assign w35944 = ~w35942 & ~w35943;
assign w35945 = pi07325 & ~w35919;
assign w35946 = ~pi02717 & w35919;
assign w35947 = ~w35945 & ~w35946;
assign w35948 = pi07326 & ~w35929;
assign w35949 = ~pi02718 & w35929;
assign w35950 = ~w35948 & ~w35949;
assign w35951 = pi07327 & ~w35929;
assign w35952 = ~pi02167 & w35929;
assign w35953 = ~w35951 & ~w35952;
assign w35954 = pi07328 & ~w35929;
assign w35955 = ~pi02164 & w35929;
assign w35956 = ~w35954 & ~w35955;
assign w35957 = pi07329 & ~w35929;
assign w35958 = ~pi02719 & w35929;
assign w35959 = ~w35957 & ~w35958;
assign w35960 = pi07330 & ~w33829;
assign w35961 = ~pi02703 & w33829;
assign w35962 = ~w35960 & ~w35961;
assign w35963 = pi07331 & ~w33829;
assign w35964 = w17466 & w17811;
assign w35965 = ~w35963 & ~w35964;
assign w35966 = ~w16905 & w20470;
assign w35967 = pi07332 & ~w35966;
assign w35968 = ~pi02711 & w35966;
assign w35969 = ~w35967 & ~w35968;
assign w35970 = pi07333 & ~w33829;
assign w35971 = ~pi02167 & w33829;
assign w35972 = ~w35970 & ~w35971;
assign w35973 = pi07334 & ~w35966;
assign w35974 = ~pi02712 & w35966;
assign w35975 = ~w35973 & ~w35974;
assign w35976 = pi07335 & ~w35966;
assign w35977 = ~pi02713 & w35966;
assign w35978 = ~w35976 & ~w35977;
assign w35979 = pi07336 & ~w35966;
assign w35980 = ~pi02714 & w35966;
assign w35981 = ~w35979 & ~w35980;
assign w35982 = pi07337 & ~w35966;
assign w35983 = ~pi02715 & w35966;
assign w35984 = ~w35982 & ~w35983;
assign w35985 = pi07338 & ~w35966;
assign w35986 = ~pi02716 & w35966;
assign w35987 = ~w35985 & ~w35986;
assign w35988 = pi07339 & ~w33829;
assign w35989 = ~pi02718 & w33829;
assign w35990 = ~w35988 & ~w35989;
assign w35991 = pi07340 & ~w33829;
assign w35992 = ~pi02722 & w33829;
assign w35993 = ~w35991 & ~w35992;
assign w35994 = pi07341 & ~w35966;
assign w35995 = ~pi02717 & w35966;
assign w35996 = ~w35994 & ~w35995;
assign w35997 = ~w16992 & w17339;
assign w35998 = pi07342 & ~w35997;
assign w35999 = ~pi02703 & w35997;
assign w36000 = ~w35998 & ~w35999;
assign w36001 = pi07343 & ~w33829;
assign w36002 = ~pi02719 & w33829;
assign w36003 = ~w36001 & ~w36002;
assign w36004 = pi07344 & ~w35997;
assign w36005 = ~pi02721 & w35997;
assign w36006 = ~w36004 & ~w36005;
assign w36007 = pi07345 & ~w35997;
assign w36008 = ~pi02169 & w35997;
assign w36009 = ~w36007 & ~w36008;
assign w36010 = pi07346 & ~w27595;
assign w36011 = ~pi02712 & w27595;
assign w36012 = ~w36010 & ~w36011;
assign w36013 = pi07347 & ~w35997;
assign w36014 = w17339 & w17586;
assign w36015 = ~w36013 & ~w36014;
assign w36016 = pi07348 & ~w35997;
assign w36017 = ~pi02167 & w35997;
assign w36018 = ~w36016 & ~w36017;
assign w36019 = pi07349 & ~w35997;
assign w36020 = ~pi02164 & w35997;
assign w36021 = ~w36019 & ~w36020;
assign w36022 = pi07350 & ~w27595;
assign w36023 = ~pi02713 & w27595;
assign w36024 = ~w36022 & ~w36023;
assign w36025 = pi07351 & ~w27595;
assign w36026 = ~pi02714 & w27595;
assign w36027 = ~w36025 & ~w36026;
assign w36028 = pi07352 & ~w27595;
assign w36029 = ~pi02715 & w27595;
assign w36030 = ~w36028 & ~w36029;
assign w36031 = pi07353 & ~w27595;
assign w36032 = ~pi02716 & w27595;
assign w36033 = ~w36031 & ~w36032;
assign w36034 = pi07354 & ~w35997;
assign w36035 = ~pi02722 & w35997;
assign w36036 = ~w36034 & ~w36035;
assign w36037 = pi07355 & ~w21318;
assign w36038 = w17603 & w17609;
assign w36039 = ~w36037 & ~w36038;
assign w36040 = pi07356 & ~w21318;
assign w36041 = w17020 & w17609;
assign w36042 = ~w36040 & ~w36041;
assign w36043 = pi07357 & ~w35997;
assign w36044 = ~pi02719 & w35997;
assign w36045 = ~w36043 & ~w36044;
assign w36046 = pi07358 & ~w21318;
assign w36047 = w17609 & w17929;
assign w36048 = ~w36046 & ~w36047;
assign w36049 = pi07359 & ~w21318;
assign w36050 = ~pi02714 & w21318;
assign w36051 = ~w36049 & ~w36050;
assign w36052 = pi07360 & ~w21318;
assign w36053 = w17609 & w18059;
assign w36054 = ~w36052 & ~w36053;
assign w36055 = pi07361 & ~w21318;
assign w36056 = w16973 & w17609;
assign w36057 = ~w36055 & ~w36056;
assign w36058 = pi07362 & ~w21105;
assign w36059 = w17540 & w17603;
assign w36060 = ~w36058 & ~w36059;
assign w36061 = pi07363 & ~w21105;
assign w36062 = w17020 & w17540;
assign w36063 = ~w36061 & ~w36062;
assign w36064 = pi07364 & ~w21105;
assign w36065 = ~pi02170 & w21105;
assign w36066 = ~w36064 & ~w36065;
assign w36067 = pi07365 & ~w21105;
assign w36068 = ~pi02713 & w21105;
assign w36069 = ~w36067 & ~w36068;
assign w36070 = pi07366 & ~w21105;
assign w36071 = w17540 & w17742;
assign w36072 = ~w36070 & ~w36071;
assign w36073 = pi07367 & ~w21105;
assign w36074 = ~pi02715 & w21105;
assign w36075 = ~w36073 & ~w36074;
assign w36076 = pi07368 & ~w21105;
assign w36077 = ~pi02717 & w21105;
assign w36078 = ~w36076 & ~w36077;
assign w36079 = pi07369 & ~w20946;
assign w36080 = ~pi02711 & w20946;
assign w36081 = ~w36079 & ~w36080;
assign w36082 = pi07370 & ~w20946;
assign w36083 = ~pi02712 & w20946;
assign w36084 = ~w36082 & ~w36083;
assign w36085 = pi07371 & ~w20946;
assign w36086 = ~pi02713 & w20946;
assign w36087 = ~w36085 & ~w36086;
assign w36088 = ~w16992 & w17300;
assign w36089 = pi07372 & ~w36088;
assign w36090 = ~pi02703 & w36088;
assign w36091 = ~w36089 & ~w36090;
assign w36092 = pi07373 & ~w20946;
assign w36093 = ~pi02714 & w20946;
assign w36094 = ~w36092 & ~w36093;
assign w36095 = pi07374 & ~w36088;
assign w36096 = ~pi02721 & w36088;
assign w36097 = ~w36095 & ~w36096;
assign w36098 = pi07375 & ~w20946;
assign w36099 = ~pi02716 & w20946;
assign w36100 = ~w36098 & ~w36099;
assign w36101 = pi07376 & ~w20946;
assign w36102 = ~pi02717 & w20946;
assign w36103 = ~w36101 & ~w36102;
assign w36104 = pi07377 & ~w20758;
assign w36105 = ~pi02711 & w20758;
assign w36106 = ~w36104 & ~w36105;
assign w36107 = pi07378 & ~w36088;
assign w36108 = ~pi02169 & w36088;
assign w36109 = ~w36107 & ~w36108;
assign w36110 = pi07379 & ~w36088;
assign w36111 = ~pi02718 & w36088;
assign w36112 = ~w36110 & ~w36111;
assign w36113 = pi07380 & ~w20758;
assign w36114 = w17020 & w18585;
assign w36115 = ~w36113 & ~w36114;
assign w36116 = pi07381 & ~w20758;
assign w36117 = ~pi02713 & w20758;
assign w36118 = ~w36116 & ~w36117;
assign w36119 = pi07382 & ~w20758;
assign w36120 = ~pi02714 & w20758;
assign w36121 = ~w36119 & ~w36120;
assign w36122 = pi07383 & ~w36088;
assign w36123 = w17300 & w19273;
assign w36124 = ~w36122 & ~w36123;
assign w36125 = pi07384 & ~w20758;
assign w36126 = ~pi02716 & w20758;
assign w36127 = ~w36125 & ~w36126;
assign w36128 = pi07385 & ~w36088;
assign w36129 = ~pi02164 & w36088;
assign w36130 = ~w36128 & ~w36129;
assign w36131 = pi07386 & ~w20758;
assign w36132 = w16973 & w18585;
assign w36133 = ~w36131 & ~w36132;
assign w36134 = pi07387 & ~w36088;
assign w36135 = ~pi02722 & w36088;
assign w36136 = ~w36134 & ~w36135;
assign w36137 = pi07388 & ~w18527;
assign w36138 = ~pi02712 & w18527;
assign w36139 = ~w36137 & ~w36138;
assign w36140 = pi07389 & ~w36088;
assign w36141 = ~pi02719 & w36088;
assign w36142 = ~w36140 & ~w36141;
assign w36143 = pi07390 & ~w19171;
assign w36144 = ~pi02703 & w19171;
assign w36145 = ~w36143 & ~w36144;
assign w36146 = pi07391 & ~w18527;
assign w36147 = w18526 & w20209;
assign w36148 = ~w36146 & ~w36147;
assign w36149 = pi07392 & ~w18527;
assign w36150 = w17929 & w18526;
assign w36151 = ~w36149 & ~w36150;
assign w36152 = pi07393 & ~w18527;
assign w36153 = w17742 & w18526;
assign w36154 = ~w36152 & ~w36153;
assign w36155 = pi07394 & ~w19171;
assign w36156 = ~pi02721 & w19171;
assign w36157 = ~w36155 & ~w36156;
assign w36158 = pi07395 & ~w18527;
assign w36159 = ~pi02716 & w18527;
assign w36160 = ~w36158 & ~w36159;
assign w36161 = pi07396 & ~w18527;
assign w36162 = w16973 & w18526;
assign w36163 = ~w36161 & ~w36162;
assign w36164 = pi07397 & ~w19171;
assign w36165 = ~pi02169 & w19171;
assign w36166 = ~w36164 & ~w36165;
assign w36167 = pi07398 & ~w19880;
assign w36168 = ~pi02712 & w19880;
assign w36169 = ~w36167 & ~w36168;
assign w36170 = pi07399 & ~w19880;
assign w36171 = ~pi02170 & w19880;
assign w36172 = ~w36170 & ~w36171;
assign w36173 = pi07400 & ~w19171;
assign w36174 = ~pi02167 & w19171;
assign w36175 = ~w36173 & ~w36174;
assign w36176 = pi07401 & ~w19880;
assign w36177 = ~pi02713 & w19880;
assign w36178 = ~w36176 & ~w36177;
assign w36179 = pi07402 & ~w19880;
assign w36180 = ~pi02714 & w19880;
assign w36181 = ~w36179 & ~w36180;
assign w36182 = pi07403 & ~w19880;
assign w36183 = ~pi02715 & w19880;
assign w36184 = ~w36182 & ~w36183;
assign w36185 = pi07404 & ~w19880;
assign w36186 = ~pi02716 & w19880;
assign w36187 = ~w36185 & ~w36186;
assign w36188 = pi07405 & ~w19171;
assign w36189 = ~pi02164 & w19171;
assign w36190 = ~w36188 & ~w36189;
assign w36191 = pi07406 & ~w19880;
assign w36192 = ~pi02717 & w19880;
assign w36193 = ~w36191 & ~w36192;
assign w36194 = pi07407 & ~w17954;
assign w36195 = ~pi02712 & w17954;
assign w36196 = ~w36194 & ~w36195;
assign w36197 = pi07408 & ~w19171;
assign w36198 = ~pi02722 & w19171;
assign w36199 = ~w36197 & ~w36198;
assign w36200 = pi07409 & ~w17954;
assign w36201 = ~pi02170 & w17954;
assign w36202 = ~w36200 & ~w36201;
assign w36203 = pi07410 & ~w17954;
assign w36204 = w17411 & w17929;
assign w36205 = ~w36203 & ~w36204;
assign w36206 = ~w16992 & w17264;
assign w36207 = pi07411 & ~w36206;
assign w36208 = ~pi02703 & w36206;
assign w36209 = ~w36207 & ~w36208;
assign w36210 = pi07412 & ~w17954;
assign w36211 = ~pi02714 & w17954;
assign w36212 = ~w36210 & ~w36211;
assign w36213 = pi07413 & ~w36206;
assign w36214 = ~pi02721 & w36206;
assign w36215 = ~w36213 & ~w36214;
assign w36216 = pi07414 & ~w17954;
assign w36217 = ~pi02716 & w17954;
assign w36218 = ~w36216 & ~w36217;
assign w36219 = pi07415 & ~w17954;
assign w36220 = ~pi02717 & w17954;
assign w36221 = ~w36219 & ~w36220;
assign w36222 = pi07416 & ~w18075;
assign w36223 = ~pi02711 & w18075;
assign w36224 = ~w36222 & ~w36223;
assign w36225 = pi07417 & ~w36206;
assign w36226 = ~pi02169 & w36206;
assign w36227 = ~w36225 & ~w36226;
assign w36228 = pi07418 & ~w18075;
assign w36229 = ~pi02712 & w18075;
assign w36230 = ~w36228 & ~w36229;
assign w36231 = pi07419 & ~w18075;
assign w36232 = ~pi02170 & w18075;
assign w36233 = ~w36231 & ~w36232;
assign w36234 = pi07420 & ~w36206;
assign w36235 = ~pi02718 & w36206;
assign w36236 = ~w36234 & ~w36235;
assign w36237 = pi07421 & ~w18075;
assign w36238 = ~pi02714 & w18075;
assign w36239 = ~w36237 & ~w36238;
assign w36240 = pi07422 & ~w36206;
assign w36241 = ~pi02167 & w36206;
assign w36242 = ~w36240 & ~w36241;
assign w36243 = pi07423 & ~w18075;
assign w36244 = ~pi02716 & w18075;
assign w36245 = ~w36243 & ~w36244;
assign w36246 = pi07424 & ~w36206;
assign w36247 = ~pi02164 & w36206;
assign w36248 = ~w36246 & ~w36247;
assign w36249 = pi07425 & ~w18075;
assign w36250 = ~pi02717 & w18075;
assign w36251 = ~w36249 & ~w36250;
assign w36252 = pi07426 & ~w18023;
assign w36253 = w17020 & w18022;
assign w36254 = ~w36252 & ~w36253;
assign w36255 = pi07427 & ~w36206;
assign w36256 = ~pi02722 & w36206;
assign w36257 = ~w36255 & ~w36256;
assign w36258 = pi07428 & ~w18023;
assign w36259 = ~pi02170 & w18023;
assign w36260 = ~w36258 & ~w36259;
assign w36261 = pi07429 & ~w18023;
assign w36262 = w17929 & w18022;
assign w36263 = ~w36261 & ~w36262;
assign w36264 = pi07430 & ~w36206;
assign w36265 = ~pi02719 & w36206;
assign w36266 = ~w36264 & ~w36265;
assign w36267 = pi07431 & ~w18023;
assign w36268 = w17742 & w18022;
assign w36269 = ~w36267 & ~w36268;
assign w36270 = pi07432 & ~w18023;
assign w36271 = ~pi02715 & w18023;
assign w36272 = ~w36270 & ~w36271;
assign w36273 = pi07433 & ~w18023;
assign w36274 = w17317 & w18022;
assign w36275 = ~w36273 & ~w36274;
assign w36276 = pi07434 & ~w18023;
assign w36277 = ~pi02717 & w18023;
assign w36278 = ~w36276 & ~w36277;
assign w36279 = pi07435 & ~w17664;
assign w36280 = ~pi02169 & w17664;
assign w36281 = ~w36279 & ~w36280;
assign w36282 = pi07436 & ~w17664;
assign w36283 = ~pi02718 & w17664;
assign w36284 = ~w36282 & ~w36283;
assign w36285 = pi07437 & ~w17664;
assign w36286 = w17663 & w19273;
assign w36287 = ~w36285 & ~w36286;
assign w36288 = pi07438 & ~w17664;
assign w36289 = w17663 & w19312;
assign w36290 = ~w36288 & ~w36289;
assign w36291 = pi07439 & ~w17664;
assign w36292 = ~pi02719 & w17664;
assign w36293 = ~w36291 & ~w36292;
assign w36294 = pi07440 & ~w17866;
assign w36295 = ~pi02703 & w17866;
assign w36296 = ~w36294 & ~w36295;
assign w36297 = pi07441 & ~w17768;
assign w36298 = ~pi02711 & w17768;
assign w36299 = ~w36297 & ~w36298;
assign w36300 = pi07442 & ~w17866;
assign w36301 = ~pi02721 & w17866;
assign w36302 = ~w36300 & ~w36301;
assign w36303 = pi07443 & ~w17866;
assign w36304 = ~pi02169 & w17866;
assign w36305 = ~w36303 & ~w36304;
assign w36306 = pi07444 & ~w17768;
assign w36307 = ~pi02712 & w17768;
assign w36308 = ~w36306 & ~w36307;
assign w36309 = pi07445 & ~w17768;
assign w36310 = ~pi02170 & w17768;
assign w36311 = ~w36309 & ~w36310;
assign w36312 = pi07446 & ~w17768;
assign w36313 = ~pi02713 & w17768;
assign w36314 = ~w36312 & ~w36313;
assign w36315 = pi07447 & ~w17768;
assign w36316 = ~pi02714 & w17768;
assign w36317 = ~w36315 & ~w36316;
assign w36318 = pi07448 & ~w17866;
assign w36319 = ~pi02167 & w17866;
assign w36320 = ~w36318 & ~w36319;
assign w36321 = pi07449 & ~w17768;
assign w36322 = ~pi02716 & w17768;
assign w36323 = ~w36321 & ~w36322;
assign w36324 = pi07450 & ~w17866;
assign w36325 = ~pi02164 & w17866;
assign w36326 = ~w36324 & ~w36325;
assign w36327 = pi07451 & ~w17768;
assign w36328 = ~pi02717 & w17768;
assign w36329 = ~w36327 & ~w36328;
assign w36330 = pi07452 & ~w17687;
assign w36331 = w17020 & w17686;
assign w36332 = ~w36330 & ~w36331;
assign w36333 = pi07453 & ~w17866;
assign w36334 = ~pi02722 & w17866;
assign w36335 = ~w36333 & ~w36334;
assign w36336 = pi07454 & ~w17687;
assign w36337 = ~pi02170 & w17687;
assign w36338 = ~w36336 & ~w36337;
assign w36339 = pi07455 & ~w17687;
assign w36340 = w17686 & w17929;
assign w36341 = ~w36339 & ~w36340;
assign w36342 = pi07456 & ~w17866;
assign w36343 = ~pi02719 & w17866;
assign w36344 = ~w36342 & ~w36343;
assign w36345 = pi07457 & ~w17687;
assign w36346 = w17686 & w17742;
assign w36347 = ~w36345 & ~w36346;
assign w36348 = pi07458 & ~w17687;
assign w36349 = ~pi02715 & w17687;
assign w36350 = ~w36348 & ~w36349;
assign w36351 = pi07459 & ~w17687;
assign w36352 = w17317 & w17686;
assign w36353 = ~w36351 & ~w36352;
assign w36354 = pi07460 & ~w17687;
assign w36355 = ~pi02717 & w17687;
assign w36356 = ~w36354 & ~w36355;
assign w36357 = ~w16905 & w17614;
assign w36358 = pi07461 & ~w36357;
assign w36359 = ~pi02711 & w36357;
assign w36360 = ~w36358 & ~w36359;
assign w36361 = pi07462 & ~w36357;
assign w36362 = w17020 & w17614;
assign w36363 = ~w36361 & ~w36362;
assign w36364 = pi07463 & ~w36357;
assign w36365 = ~pi02170 & w36357;
assign w36366 = ~w36364 & ~w36365;
assign w36367 = pi07464 & ~w20713;
assign w36368 = ~pi02169 & w20713;
assign w36369 = ~w36367 & ~w36368;
assign w36370 = pi07465 & ~w36357;
assign w36371 = ~pi02713 & w36357;
assign w36372 = ~w36370 & ~w36371;
assign w36373 = pi07466 & ~w36357;
assign w36374 = ~pi02714 & w36357;
assign w36375 = ~w36373 & ~w36374;
assign w36376 = pi07467 & ~w20713;
assign w36377 = ~pi02167 & w20713;
assign w36378 = ~w36376 & ~w36377;
assign w36379 = pi07468 & ~w36357;
assign w36380 = ~pi02715 & w36357;
assign w36381 = ~w36379 & ~w36380;
assign w36382 = pi07469 & ~w36357;
assign w36383 = ~pi02716 & w36357;
assign w36384 = ~w36382 & ~w36383;
assign w36385 = pi07470 & ~w20713;
assign w36386 = ~pi02164 & w20713;
assign w36387 = ~w36385 & ~w36386;
assign w36388 = pi07471 & ~w36357;
assign w36389 = ~pi02717 & w36357;
assign w36390 = ~w36388 & ~w36389;
assign w36391 = ~w16905 & w17526;
assign w36392 = pi07472 & ~w36391;
assign w36393 = ~pi02712 & w36391;
assign w36394 = ~w36392 & ~w36393;
assign w36395 = pi07473 & ~w20713;
assign w36396 = ~pi02722 & w20713;
assign w36397 = ~w36395 & ~w36396;
assign w36398 = pi07474 & ~w36391;
assign w36399 = ~pi02170 & w36391;
assign w36400 = ~w36398 & ~w36399;
assign w36401 = pi07475 & ~w20713;
assign w36402 = ~pi02719 & w20713;
assign w36403 = ~w36401 & ~w36402;
assign w36404 = pi07476 & ~w36391;
assign w36405 = ~pi02714 & w36391;
assign w36406 = ~w36404 & ~w36405;
assign w36407 = pi07477 & ~w36391;
assign w36408 = ~pi02715 & w36391;
assign w36409 = ~w36407 & ~w36408;
assign w36410 = pi07478 & ~w36391;
assign w36411 = ~pi02716 & w36391;
assign w36412 = ~w36410 & ~w36411;
assign w36413 = pi07479 & ~w36391;
assign w36414 = ~pi02717 & w36391;
assign w36415 = ~w36413 & ~w36414;
assign w36416 = ~w16905 & w17922;
assign w36417 = pi07480 & ~w36416;
assign w36418 = ~pi02711 & w36416;
assign w36419 = ~w36417 & ~w36418;
assign w36420 = pi07481 & ~w21600;
assign w36421 = ~pi02721 & w21600;
assign w36422 = ~w36420 & ~w36421;
assign w36423 = pi07482 & ~w36416;
assign w36424 = w17020 & w17922;
assign w36425 = ~w36423 & ~w36424;
assign w36426 = pi07483 & ~w36416;
assign w36427 = w17922 & w20209;
assign w36428 = ~w36426 & ~w36427;
assign w36429 = pi07484 & ~w21600;
assign w36430 = ~pi02169 & w21600;
assign w36431 = ~w36429 & ~w36430;
assign w36432 = pi07485 & ~w36416;
assign w36433 = ~pi02714 & w36416;
assign w36434 = ~w36432 & ~w36433;
assign w36435 = pi07486 & ~w21600;
assign w36436 = ~pi02718 & w21600;
assign w36437 = ~w36435 & ~w36436;
assign w36438 = pi07487 & ~w21600;
assign w36439 = ~pi02167 & w21600;
assign w36440 = ~w36438 & ~w36439;
assign w36441 = pi07488 & ~w36416;
assign w36442 = ~pi02716 & w36416;
assign w36443 = ~w36441 & ~w36442;
assign w36444 = pi07489 & ~w21600;
assign w36445 = ~pi02164 & w21600;
assign w36446 = ~w36444 & ~w36445;
assign w36447 = pi07490 & ~w36416;
assign w36448 = ~pi02717 & w36416;
assign w36449 = ~w36447 & ~w36448;
assign w36450 = ~w16905 & w17641;
assign w36451 = pi07491 & ~w36450;
assign w36452 = ~pi02712 & w36450;
assign w36453 = ~w36451 & ~w36452;
assign w36454 = pi07492 & ~w21600;
assign w36455 = ~pi02722 & w21600;
assign w36456 = ~w36454 & ~w36455;
assign w36457 = pi07493 & ~w36450;
assign w36458 = ~pi02170 & w36450;
assign w36459 = ~w36457 & ~w36458;
assign w36460 = pi07494 & ~w36450;
assign w36461 = ~pi02713 & w36450;
assign w36462 = ~w36460 & ~w36461;
assign w36463 = pi07495 & ~w21600;
assign w36464 = ~pi02719 & w21600;
assign w36465 = ~w36463 & ~w36464;
assign w36466 = pi07496 & ~w36450;
assign w36467 = ~pi02714 & w36450;
assign w36468 = ~w36466 & ~w36467;
assign w36469 = pi07497 & ~w36450;
assign w36470 = ~pi02715 & w36450;
assign w36471 = ~w36469 & ~w36470;
assign w36472 = ~w16992 & w20561;
assign w36473 = pi07498 & ~w36472;
assign w36474 = w17811 & w20561;
assign w36475 = ~w36473 & ~w36474;
assign w36476 = pi07499 & ~w36450;
assign w36477 = ~pi02716 & w36450;
assign w36478 = ~w36476 & ~w36477;
assign w36479 = pi07500 & ~w36450;
assign w36480 = ~pi02717 & w36450;
assign w36481 = ~w36479 & ~w36480;
assign w36482 = pi07501 & ~w21563;
assign w36483 = ~pi02712 & w21563;
assign w36484 = ~w36482 & ~w36483;
assign w36485 = pi07502 & ~w21563;
assign w36486 = ~pi02170 & w21563;
assign w36487 = ~w36485 & ~w36486;
assign w36488 = pi07503 & ~w36472;
assign w36489 = w19797 & w20561;
assign w36490 = ~w36488 & ~w36489;
assign w36491 = pi07504 & ~w21563;
assign w36492 = ~pi02714 & w21563;
assign w36493 = ~w36491 & ~w36492;
assign w36494 = pi07505 & ~w36472;
assign w36495 = w17586 & w20561;
assign w36496 = ~w36494 & ~w36495;
assign w36497 = pi07506 & ~w21563;
assign w36498 = ~pi02715 & w21563;
assign w36499 = ~w36497 & ~w36498;
assign w36500 = pi07507 & ~w21563;
assign w36501 = ~pi02716 & w21563;
assign w36502 = ~w36500 & ~w36501;
assign w36503 = pi07508 & ~w36472;
assign w36504 = w19273 & w20561;
assign w36505 = ~w36503 & ~w36504;
assign w36506 = pi07509 & ~w36472;
assign w36507 = w17620 & w20561;
assign w36508 = ~w36506 & ~w36507;
assign w36509 = pi07510 & ~w21563;
assign w36510 = ~pi02717 & w21563;
assign w36511 = ~w36509 & ~w36510;
assign w36512 = pi07511 & ~w21037;
assign w36513 = ~pi02712 & w21037;
assign w36514 = ~w36512 & ~w36513;
assign w36515 = pi07512 & ~w36472;
assign w36516 = w19312 & w20561;
assign w36517 = ~w36515 & ~w36516;
assign w36518 = pi07513 & ~w21037;
assign w36519 = ~pi02170 & w21037;
assign w36520 = ~w36518 & ~w36519;
assign w36521 = pi07514 & ~w21037;
assign w36522 = ~pi02714 & w21037;
assign w36523 = ~w36521 & ~w36522;
assign w36524 = pi07515 & ~w36472;
assign w36525 = w17594 & w20561;
assign w36526 = ~w36524 & ~w36525;
assign w36527 = pi07516 & ~w21037;
assign w36528 = w18059 & w20720;
assign w36529 = ~w36527 & ~w36528;
assign w36530 = pi07517 & ~w21037;
assign w36531 = ~pi02717 & w21037;
assign w36532 = ~w36530 & ~w36531;
assign w36533 = pi07518 & ~w20981;
assign w36534 = ~pi02711 & w20981;
assign w36535 = ~w36533 & ~w36534;
assign w36536 = pi07519 & ~w20981;
assign w36537 = ~pi02712 & w20981;
assign w36538 = ~w36536 & ~w36537;
assign w36539 = pi07520 & ~w20981;
assign w36540 = ~pi02170 & w20981;
assign w36541 = ~w36539 & ~w36540;
assign w36542 = pi07521 & ~w20981;
assign w36543 = ~pi02713 & w20981;
assign w36544 = ~w36542 & ~w36543;
assign w36545 = pi07522 & ~w20981;
assign w36546 = ~pi02714 & w20981;
assign w36547 = ~w36545 & ~w36546;
assign w36548 = pi07523 & ~w20981;
assign w36549 = ~pi02715 & w20981;
assign w36550 = ~w36548 & ~w36549;
assign w36551 = pi07524 & ~w20981;
assign w36552 = w16973 & w18631;
assign w36553 = ~w36551 & ~w36552;
assign w36554 = pi07525 & ~w20928;
assign w36555 = ~pi02711 & w20928;
assign w36556 = ~w36554 & ~w36555;
assign w36557 = pi07526 & ~w20928;
assign w36558 = ~pi02712 & w20928;
assign w36559 = ~w36557 & ~w36558;
assign w36560 = pi07527 & ~w20928;
assign w36561 = ~pi02713 & w20928;
assign w36562 = ~w36560 & ~w36561;
assign w36563 = pi07528 & ~w20928;
assign w36564 = ~pi02714 & w20928;
assign w36565 = ~w36563 & ~w36564;
assign w36566 = pi07529 & ~w20928;
assign w36567 = ~pi02715 & w20928;
assign w36568 = ~w36566 & ~w36567;
assign w36569 = pi07530 & ~w20928;
assign w36570 = ~pi02717 & w20928;
assign w36571 = ~w36569 & ~w36570;
assign w36572 = pi07531 & ~w20776;
assign w36573 = ~pi02711 & w20776;
assign w36574 = ~w36572 & ~w36573;
assign w36575 = pi07532 & ~w20776;
assign w36576 = w17020 & w20775;
assign w36577 = ~w36575 & ~w36576;
assign w36578 = pi07533 & ~w20776;
assign w36579 = ~pi02170 & w20776;
assign w36580 = ~w36578 & ~w36579;
assign w36581 = pi07534 & ~w20776;
assign w36582 = w17929 & w20775;
assign w36583 = ~w36581 & ~w36582;
assign w36584 = pi07535 & ~w20776;
assign w36585 = ~pi02714 & w20776;
assign w36586 = ~w36584 & ~w36585;
assign w36587 = pi07536 & ~w20776;
assign w36588 = ~pi02715 & w20776;
assign w36589 = ~w36587 & ~w36588;
assign w36590 = pi07537 & ~w20776;
assign w36591 = w16973 & w20775;
assign w36592 = ~w36590 & ~w36591;
assign w36593 = pi07538 & ~w20810;
assign w36594 = ~pi02711 & w20810;
assign w36595 = ~w36593 & ~w36594;
assign w36596 = pi07539 & ~w20810;
assign w36597 = w17020 & w17583;
assign w36598 = ~w36596 & ~w36597;
assign w36599 = pi07540 & ~w20810;
assign w36600 = w17583 & w17929;
assign w36601 = ~w36599 & ~w36600;
assign w36602 = pi07541 & ~w20810;
assign w36603 = w17583 & w17742;
assign w36604 = ~w36602 & ~w36603;
assign w36605 = pi07542 & ~w20810;
assign w36606 = ~pi02715 & w20810;
assign w36607 = ~w36605 & ~w36606;
assign w36608 = pi07543 & ~w20810;
assign w36609 = w17317 & w17583;
assign w36610 = ~w36608 & ~w36609;
assign w36611 = pi07544 & ~w20810;
assign w36612 = ~pi02717 & w20810;
assign w36613 = ~w36611 & ~w36612;
assign w36614 = pi07545 & ~w20567;
assign w36615 = ~pi02711 & w20567;
assign w36616 = ~w36614 & ~w36615;
assign w36617 = pi07546 & ~w20747;
assign w36618 = ~pi02721 & w20747;
assign w36619 = ~w36617 & ~w36618;
assign w36620 = pi07547 & ~w20567;
assign w36621 = ~pi02712 & w20567;
assign w36622 = ~w36620 & ~w36621;
assign w36623 = pi07548 & ~w20567;
assign w36624 = ~pi02170 & w20567;
assign w36625 = ~w36623 & ~w36624;
assign w36626 = pi07549 & ~w20747;
assign w36627 = ~pi02169 & w20747;
assign w36628 = ~w36626 & ~w36627;
assign w36629 = pi07550 & ~w20567;
assign w36630 = ~pi02714 & w20567;
assign w36631 = ~w36629 & ~w36630;
assign w36632 = pi07551 & ~w20747;
assign w36633 = ~pi02718 & w20747;
assign w36634 = ~w36632 & ~w36633;
assign w36635 = pi07552 & ~w20747;
assign w36636 = ~pi02167 & w20747;
assign w36637 = ~w36635 & ~w36636;
assign w36638 = pi07553 & ~w20567;
assign w36639 = ~pi02716 & w20567;
assign w36640 = ~w36638 & ~w36639;
assign w36641 = pi07554 & ~w20567;
assign w36642 = ~pi02717 & w20567;
assign w36643 = ~w36641 & ~w36642;
assign w36644 = pi07555 & ~w20171;
assign w36645 = ~pi02711 & w20171;
assign w36646 = ~w36644 & ~w36645;
assign w36647 = pi07556 & ~w20747;
assign w36648 = ~pi02164 & w20747;
assign w36649 = ~w36647 & ~w36648;
assign w36650 = pi07557 & ~w20171;
assign w36651 = w20170 & w20209;
assign w36652 = ~w36650 & ~w36651;
assign w36653 = pi07558 & ~w20171;
assign w36654 = w17929 & w20170;
assign w36655 = ~w36653 & ~w36654;
assign w36656 = pi07559 & ~w20747;
assign w36657 = ~pi02722 & w20747;
assign w36658 = ~w36656 & ~w36657;
assign w36659 = pi07560 & ~w20171;
assign w36660 = ~pi02714 & w20171;
assign w36661 = ~w36659 & ~w36660;
assign w36662 = pi07561 & ~w20171;
assign w36663 = ~pi02715 & w20171;
assign w36664 = ~w36662 & ~w36663;
assign w36665 = pi07562 & ~w20171;
assign w36666 = ~pi02716 & w20171;
assign w36667 = ~w36665 & ~w36666;
assign w36668 = pi07563 & ~w20185;
assign w36669 = ~pi02711 & w20185;
assign w36670 = ~w36668 & ~w36669;
assign w36671 = pi07564 & ~w20747;
assign w36672 = ~pi02719 & w20747;
assign w36673 = ~w36671 & ~w36672;
assign w36674 = pi07565 & ~w20185;
assign w36675 = ~pi02712 & w20185;
assign w36676 = ~w36674 & ~w36675;
assign w36677 = pi07566 & ~w20185;
assign w36678 = ~pi02713 & w20185;
assign w36679 = ~w36677 & ~w36678;
assign w36680 = pi07567 & ~w20185;
assign w36681 = ~pi02714 & w20185;
assign w36682 = ~w36680 & ~w36681;
assign w36683 = pi07568 & ~w20185;
assign w36684 = ~pi02715 & w20185;
assign w36685 = ~w36683 & ~w36684;
assign w36686 = ~w16928 & w17289;
assign w36687 = pi07569 & ~w36686;
assign w36688 = ~pi02720 & w36686;
assign w36689 = ~w36687 & ~w36688;
assign w36690 = pi07570 & ~w20185;
assign w36691 = ~pi02717 & w20185;
assign w36692 = ~w36690 & ~w36691;
assign w36693 = pi07571 & ~w18773;
assign w36694 = ~pi02711 & w18773;
assign w36695 = ~w36693 & ~w36694;
assign w36696 = pi07572 & ~w18773;
assign w36697 = ~pi02712 & w18773;
assign w36698 = ~w36696 & ~w36697;
assign w36699 = pi07573 & ~w18773;
assign w36700 = ~pi02170 & w18773;
assign w36701 = ~w36699 & ~w36700;
assign w36702 = pi07574 & ~w18773;
assign w36703 = w17929 & w18772;
assign w36704 = ~w36702 & ~w36703;
assign w36705 = pi07575 & ~w18773;
assign w36706 = ~pi02714 & w18773;
assign w36707 = ~w36705 & ~w36706;
assign w36708 = pi07576 & ~w18773;
assign w36709 = ~pi02715 & w18773;
assign w36710 = ~w36708 & ~w36709;
assign w36711 = pi07577 & ~w18773;
assign w36712 = ~pi02717 & w18773;
assign w36713 = ~w36711 & ~w36712;
assign w36714 = pi07578 & ~w18033;
assign w36715 = w17532 & w18032;
assign w36716 = ~w36714 & ~w36715;
assign w36717 = pi07579 & ~w18033;
assign w36718 = ~pi02721 & w18033;
assign w36719 = ~w36717 & ~w36718;
assign w36720 = pi07580 & ~w18033;
assign w36721 = w17586 & w18032;
assign w36722 = ~w36720 & ~w36721;
assign w36723 = pi07581 & ~w18033;
assign w36724 = ~pi02167 & w18033;
assign w36725 = ~w36723 & ~w36724;
assign w36726 = pi07582 & ~w18301;
assign w36727 = ~pi02711 & w18301;
assign w36728 = ~w36726 & ~w36727;
assign w36729 = pi07583 & ~w18301;
assign w36730 = ~pi02170 & w18301;
assign w36731 = ~w36729 & ~w36730;
assign w36732 = pi07584 & ~w18301;
assign w36733 = ~pi02713 & w18301;
assign w36734 = ~w36732 & ~w36733;
assign w36735 = pi07585 & ~w18301;
assign w36736 = ~pi02714 & w18301;
assign w36737 = ~w36735 & ~w36736;
assign w36738 = pi07586 & ~w18301;
assign w36739 = ~pi02715 & w18301;
assign w36740 = ~w36738 & ~w36739;
assign w36741 = pi07587 & ~w18033;
assign w36742 = ~pi02719 & w18033;
assign w36743 = ~w36741 & ~w36742;
assign w36744 = pi07588 & ~w18301;
assign w36745 = ~pi02716 & w18301;
assign w36746 = ~w36744 & ~w36745;
assign w36747 = pi07589 & ~w18301;
assign w36748 = ~pi02717 & w18301;
assign w36749 = ~w36747 & ~w36748;
assign w36750 = pi07590 & ~w17610;
assign w36751 = ~pi02703 & w17610;
assign w36752 = ~w36750 & ~w36751;
assign w36753 = pi07591 & ~w18033;
assign w36754 = ~pi02722 & w18033;
assign w36755 = ~w36753 & ~w36754;
assign w36756 = pi07592 & ~w17610;
assign w36757 = ~pi02721 & w17610;
assign w36758 = ~w36756 & ~w36757;
assign w36759 = pi07593 & ~w17610;
assign w36760 = ~pi02718 & w17610;
assign w36761 = ~w36759 & ~w36760;
assign w36762 = pi07594 & ~w17610;
assign w36763 = w17609 & w19273;
assign w36764 = ~w36762 & ~w36763;
assign w36765 = pi07595 & ~w17908;
assign w36766 = ~pi02711 & w17908;
assign w36767 = ~w36765 & ~w36766;
assign w36768 = pi07596 & ~w17610;
assign w36769 = w17609 & w17620;
assign w36770 = ~w36768 & ~w36769;
assign w36771 = pi07597 & ~w17908;
assign w36772 = ~pi02170 & w17908;
assign w36773 = ~w36771 & ~w36772;
assign w36774 = pi07598 & ~w17908;
assign w36775 = ~pi02713 & w17908;
assign w36776 = ~w36774 & ~w36775;
assign w36777 = pi07599 & ~w17908;
assign w36778 = ~pi02715 & w17908;
assign w36779 = ~w36777 & ~w36778;
assign w36780 = pi07600 & ~w17908;
assign w36781 = ~pi02714 & w17908;
assign w36782 = ~w36780 & ~w36781;
assign w36783 = pi07601 & ~w17908;
assign w36784 = w17317 & w17907;
assign w36785 = ~w36783 & ~w36784;
assign w36786 = pi07602 & ~w17908;
assign w36787 = ~pi02717 & w17908;
assign w36788 = ~w36786 & ~w36787;
assign w36789 = pi07603 & ~w17610;
assign w36790 = ~pi02719 & w17610;
assign w36791 = ~w36789 & ~w36790;
assign w36792 = pi07604 & ~w17755;
assign w36793 = ~pi02711 & w17755;
assign w36794 = ~w36792 & ~w36793;
assign w36795 = pi07605 & ~w17755;
assign w36796 = ~pi02712 & w17755;
assign w36797 = ~w36795 & ~w36796;
assign w36798 = pi07606 & ~w17755;
assign w36799 = ~pi02713 & w17755;
assign w36800 = ~w36798 & ~w36799;
assign w36801 = pi07607 & ~w17755;
assign w36802 = ~pi02714 & w17755;
assign w36803 = ~w36801 & ~w36802;
assign w36804 = pi07608 & ~w17755;
assign w36805 = w17754 & w18059;
assign w36806 = ~w36804 & ~w36805;
assign w36807 = pi07609 & ~w17755;
assign w36808 = ~pi02716 & w17755;
assign w36809 = ~w36807 & ~w36808;
assign w36810 = pi07610 & ~w17755;
assign w36811 = w16973 & w17754;
assign w36812 = ~w36810 & ~w36811;
assign w36813 = pi07611 & ~w17541;
assign w36814 = ~pi02721 & w17541;
assign w36815 = ~w36813 & ~w36814;
assign w36816 = pi07612 & ~w17541;
assign w36817 = w17540 & w19797;
assign w36818 = ~w36816 & ~w36817;
assign w36819 = pi07613 & ~w17541;
assign w36820 = ~pi02718 & w17541;
assign w36821 = ~w36819 & ~w36820;
assign w36822 = pi07614 & ~w17541;
assign w36823 = ~pi02167 & w17541;
assign w36824 = ~w36822 & ~w36823;
assign w36825 = pi07615 & ~w17429;
assign w36826 = ~pi02711 & w17429;
assign w36827 = ~w36825 & ~w36826;
assign w36828 = pi07616 & ~w17541;
assign w36829 = ~pi02164 & w17541;
assign w36830 = ~w36828 & ~w36829;
assign w36831 = pi07617 & ~w17429;
assign w36832 = ~pi02170 & w17429;
assign w36833 = ~w36831 & ~w36832;
assign w36834 = pi07618 & ~w17429;
assign w36835 = ~pi02713 & w17429;
assign w36836 = ~w36834 & ~w36835;
assign w36837 = pi07619 & ~w17429;
assign w36838 = ~pi02714 & w17429;
assign w36839 = ~w36837 & ~w36838;
assign w36840 = pi07620 & ~w17429;
assign w36841 = w17428 & w18059;
assign w36842 = ~w36840 & ~w36841;
assign w36843 = pi07621 & ~w17541;
assign w36844 = ~pi02719 & w17541;
assign w36845 = ~w36843 & ~w36844;
assign w36846 = pi07622 & ~w17429;
assign w36847 = ~pi02717 & w17429;
assign w36848 = ~w36846 & ~w36847;
assign w36849 = pi07623 & ~w17290;
assign w36850 = ~pi02711 & w17290;
assign w36851 = ~w36849 & ~w36850;
assign w36852 = pi07624 & ~w17290;
assign w36853 = w17020 & w17289;
assign w36854 = ~w36852 & ~w36853;
assign w36855 = pi07625 & ~w17290;
assign w36856 = ~pi02170 & w17290;
assign w36857 = ~w36855 & ~w36856;
assign w36858 = pi07626 & ~w17290;
assign w36859 = ~pi02713 & w17290;
assign w36860 = ~w36858 & ~w36859;
assign w36861 = pi07627 & ~w17290;
assign w36862 = ~pi02714 & w17290;
assign w36863 = ~w36861 & ~w36862;
assign w36864 = pi07628 & ~w17290;
assign w36865 = ~pi02715 & w17290;
assign w36866 = ~w36864 & ~w36865;
assign w36867 = pi07629 & ~w17290;
assign w36868 = ~pi02717 & w17290;
assign w36869 = ~w36867 & ~w36868;
assign w36870 = pi07630 & ~w21540;
assign w36871 = ~pi02711 & w21540;
assign w36872 = ~w36870 & ~w36871;
assign w36873 = pi07631 & ~w21540;
assign w36874 = w17020 & w17938;
assign w36875 = ~w36873 & ~w36874;
assign w36876 = pi07632 & ~w21540;
assign w36877 = ~pi02713 & w21540;
assign w36878 = ~w36876 & ~w36877;
assign w36879 = pi07633 & ~w21540;
assign w36880 = ~pi02714 & w21540;
assign w36881 = ~w36879 & ~w36880;
assign w36882 = pi07634 & ~w21540;
assign w36883 = ~pi02715 & w21540;
assign w36884 = ~w36882 & ~w36883;
assign w36885 = pi07635 & ~w21540;
assign w36886 = ~pi02717 & w21540;
assign w36887 = ~w36885 & ~w36886;
assign w36888 = ~w16905 & w17011;
assign w36889 = pi07636 & ~w36888;
assign w36890 = ~pi02711 & w36888;
assign w36891 = ~w36889 & ~w36890;
assign w36892 = ~w16992 & w18949;
assign w36893 = pi07637 & ~w36892;
assign w36894 = ~pi02703 & w36892;
assign w36895 = ~w36893 & ~w36894;
assign w36896 = pi07638 & ~w36888;
assign w36897 = ~pi02712 & w36888;
assign w36898 = ~w36896 & ~w36897;
assign w36899 = pi07639 & ~w36888;
assign w36900 = ~pi02170 & w36888;
assign w36901 = ~w36899 & ~w36900;
assign w36902 = pi07640 & ~w36892;
assign w36903 = ~pi02721 & w36892;
assign w36904 = ~w36902 & ~w36903;
assign w36905 = pi07641 & ~w36888;
assign w36906 = ~pi02713 & w36888;
assign w36907 = ~w36905 & ~w36906;
assign w36908 = pi07642 & ~w36892;
assign w36909 = ~pi02169 & w36892;
assign w36910 = ~w36908 & ~w36909;
assign w36911 = pi07643 & ~w36888;
assign w36912 = ~pi02715 & w36888;
assign w36913 = ~w36911 & ~w36912;
assign w36914 = pi07644 & ~w36888;
assign w36915 = ~pi02716 & w36888;
assign w36916 = ~w36914 & ~w36915;
assign w36917 = pi07645 & ~w36888;
assign w36918 = ~pi02717 & w36888;
assign w36919 = ~w36917 & ~w36918;
assign w36920 = ~w16905 & w17108;
assign w36921 = pi07646 & ~w36920;
assign w36922 = w17108 & w17603;
assign w36923 = ~w36921 & ~w36922;
assign w36924 = pi07647 & ~w36920;
assign w36925 = ~pi02712 & w36920;
assign w36926 = ~w36924 & ~w36925;
assign w36927 = pi07648 & ~w36920;
assign w36928 = ~pi02170 & w36920;
assign w36929 = ~w36927 & ~w36928;
assign w36930 = pi07649 & ~w36920;
assign w36931 = ~pi02713 & w36920;
assign w36932 = ~w36930 & ~w36931;
assign w36933 = pi07650 & ~w21202;
assign w36934 = w17128 & w17734;
assign w36935 = ~w36933 & ~w36934;
assign w36936 = pi07651 & ~w36892;
assign w36937 = ~pi02164 & w36892;
assign w36938 = ~w36936 & ~w36937;
assign w36939 = pi07652 & ~w36920;
assign w36940 = ~pi02714 & w36920;
assign w36941 = ~w36939 & ~w36940;
assign w36942 = pi07653 & ~w36920;
assign w36943 = ~pi02715 & w36920;
assign w36944 = ~w36942 & ~w36943;
assign w36945 = pi07654 & ~w36892;
assign w36946 = ~pi02722 & w36892;
assign w36947 = ~w36945 & ~w36946;
assign w36948 = pi07655 & ~w36892;
assign w36949 = ~pi02719 & w36892;
assign w36950 = ~w36948 & ~w36949;
assign w36951 = pi07656 & ~w36920;
assign w36952 = w16973 & w17108;
assign w36953 = ~w36951 & ~w36952;
assign w36954 = ~w16905 & w17098;
assign w36955 = pi07657 & ~w36954;
assign w36956 = ~pi02711 & w36954;
assign w36957 = ~w36955 & ~w36956;
assign w36958 = pi07658 & ~w36954;
assign w36959 = ~pi02712 & w36954;
assign w36960 = ~w36958 & ~w36959;
assign w36961 = pi07659 & ~w36954;
assign w36962 = ~pi02170 & w36954;
assign w36963 = ~w36961 & ~w36962;
assign w36964 = pi07660 & ~w36954;
assign w36965 = ~pi02713 & w36954;
assign w36966 = ~w36964 & ~w36965;
assign w36967 = pi07661 & ~w36954;
assign w36968 = ~pi02714 & w36954;
assign w36969 = ~w36967 & ~w36968;
assign w36970 = pi07662 & ~w21070;
assign w36971 = ~pi02169 & w21070;
assign w36972 = ~w36970 & ~w36971;
assign w36973 = pi07663 & ~w36954;
assign w36974 = ~pi02715 & w36954;
assign w36975 = ~w36973 & ~w36974;
assign w36976 = pi07664 & ~w36954;
assign w36977 = ~pi02716 & w36954;
assign w36978 = ~w36976 & ~w36977;
assign w36979 = pi07665 & ~w21070;
assign w36980 = ~pi02718 & w21070;
assign w36981 = ~w36979 & ~w36980;
assign w36982 = pi07666 & ~w36954;
assign w36983 = w16973 & w17098;
assign w36984 = ~w36982 & ~w36983;
assign w36985 = pi07667 & ~w21170;
assign w36986 = ~pi02711 & w21170;
assign w36987 = ~w36985 & ~w36986;
assign w36988 = pi07668 & ~w21070;
assign w36989 = ~pi02167 & w21070;
assign w36990 = ~w36988 & ~w36989;
assign w36991 = pi07669 & ~w21170;
assign w36992 = ~pi02170 & w21170;
assign w36993 = ~w36991 & ~w36992;
assign w36994 = pi07670 & ~w21170;
assign w36995 = w17929 & w20244;
assign w36996 = ~w36994 & ~w36995;
assign w36997 = pi07671 & ~w21170;
assign w36998 = w17742 & w20244;
assign w36999 = ~w36997 & ~w36998;
assign w37000 = pi07672 & ~w21170;
assign w37001 = ~pi02715 & w21170;
assign w37002 = ~w37000 & ~w37001;
assign w37003 = pi07673 & ~w21070;
assign w37004 = ~pi02722 & w21070;
assign w37005 = ~w37003 & ~w37004;
assign w37006 = pi07674 & ~w21220;
assign w37007 = ~pi02169 & w21220;
assign w37008 = ~w37006 & ~w37007;
assign w37009 = pi07675 & ~w21170;
assign w37010 = ~pi02717 & w21170;
assign w37011 = ~w37009 & ~w37010;
assign w37012 = pi07676 & ~w21070;
assign w37013 = w17594 & w18585;
assign w37014 = ~w37012 & ~w37013;
assign w37015 = pi07677 & ~w21115;
assign w37016 = ~pi02703 & w21115;
assign w37017 = ~w37015 & ~w37016;
assign w37018 = pi07678 & ~w21115;
assign w37019 = w17811 & w18526;
assign w37020 = ~w37018 & ~w37019;
assign w37021 = pi07679 & ~w21367;
assign w37022 = ~pi02178 & w21367;
assign w37023 = ~w37021 & ~w37022;
assign w37024 = pi07680 & ~w21115;
assign w37025 = ~pi02169 & w21115;
assign w37026 = ~w37024 & ~w37025;
assign w37027 = pi07681 & ~w21115;
assign w37028 = ~pi02167 & w21115;
assign w37029 = ~w37027 & ~w37028;
assign w37030 = pi07682 & ~w21115;
assign w37031 = ~pi02164 & w21115;
assign w37032 = ~w37030 & ~w37031;
assign w37033 = pi07683 & ~w21115;
assign w37034 = ~pi02722 & w21115;
assign w37035 = ~w37033 & ~w37034;
assign w37036 = pi07684 & ~w21088;
assign w37037 = ~pi02711 & w21088;
assign w37038 = ~w37036 & ~w37037;
assign w37039 = pi07685 & ~w21088;
assign w37040 = ~pi02712 & w21088;
assign w37041 = ~w37039 & ~w37040;
assign w37042 = pi07686 & ~w21088;
assign w37043 = ~pi02170 & w21088;
assign w37044 = ~w37042 & ~w37043;
assign w37045 = pi07687 & ~w20966;
assign w37046 = ~pi02703 & w20966;
assign w37047 = ~w37045 & ~w37046;
assign w37048 = pi07688 & ~w21088;
assign w37049 = ~pi02714 & w21088;
assign w37050 = ~w37048 & ~w37049;
assign w37051 = pi07689 & ~w20966;
assign w37052 = ~pi02721 & w20966;
assign w37053 = ~w37051 & ~w37052;
assign w37054 = pi07690 & ~w20966;
assign w37055 = ~pi02169 & w20966;
assign w37056 = ~w37054 & ~w37055;
assign w37057 = pi07691 & ~w21088;
assign w37058 = ~pi02715 & w21088;
assign w37059 = ~w37057 & ~w37058;
assign w37060 = pi07692 & ~w21088;
assign w37061 = ~pi02716 & w21088;
assign w37062 = ~w37060 & ~w37061;
assign w37063 = pi07693 & ~w20966;
assign w37064 = ~pi02718 & w20966;
assign w37065 = ~w37063 & ~w37064;
assign w37066 = pi07694 & ~w21088;
assign w37067 = ~pi02717 & w21088;
assign w37068 = ~w37066 & ~w37067;
assign w37069 = pi07695 & ~w20992;
assign w37070 = ~pi02712 & w20992;
assign w37071 = ~w37069 & ~w37070;
assign w37072 = pi07696 & ~w20966;
assign w37073 = ~pi02167 & w20966;
assign w37074 = ~w37072 & ~w37073;
assign w37075 = pi07697 & ~w20966;
assign w37076 = w17620 & w18291;
assign w37077 = ~w37075 & ~w37076;
assign w37078 = pi07698 & ~w20992;
assign w37079 = ~pi02713 & w20992;
assign w37080 = ~w37078 & ~w37079;
assign w37081 = pi07699 & ~w20992;
assign w37082 = ~pi02714 & w20992;
assign w37083 = ~w37081 & ~w37082;
assign w37084 = pi07700 & ~w20992;
assign w37085 = ~pi02715 & w20992;
assign w37086 = ~w37084 & ~w37085;
assign w37087 = pi07701 & ~w20992;
assign w37088 = ~pi02716 & w20992;
assign w37089 = ~w37087 & ~w37088;
assign w37090 = pi07702 & ~w20992;
assign w37091 = ~pi02717 & w20992;
assign w37092 = ~w37090 & ~w37091;
assign w37093 = pi07703 & ~w20939;
assign w37094 = ~pi02711 & w20939;
assign w37095 = ~w37093 & ~w37094;
assign w37096 = pi07704 & ~w20966;
assign w37097 = w17594 & w18291;
assign w37098 = ~w37096 & ~w37097;
assign w37099 = pi07705 & ~w20939;
assign w37100 = ~pi02712 & w20939;
assign w37101 = ~w37099 & ~w37100;
assign w37102 = pi07706 & ~w20939;
assign w37103 = w18617 & w20209;
assign w37104 = ~w37102 & ~w37103;
assign w37105 = pi07707 & ~w20791;
assign w37106 = ~pi02703 & w20791;
assign w37107 = ~w37105 & ~w37106;
assign w37108 = pi07708 & ~w20939;
assign w37109 = w17742 & w18617;
assign w37110 = ~w37108 & ~w37109;
assign w37111 = pi07709 & ~w20791;
assign w37112 = ~pi02721 & w20791;
assign w37113 = ~w37111 & ~w37112;
assign w37114 = pi07710 & ~w20939;
assign w37115 = ~pi02715 & w20939;
assign w37116 = ~w37114 & ~w37115;
assign w37117 = pi07711 & ~w20791;
assign w37118 = w17411 & w19797;
assign w37119 = ~w37117 & ~w37118;
assign w37120 = pi07712 & ~w20791;
assign w37121 = ~pi02718 & w20791;
assign w37122 = ~w37120 & ~w37121;
assign w37123 = pi07713 & ~w20939;
assign w37124 = w16973 & w18617;
assign w37125 = ~w37123 & ~w37124;
assign w37126 = pi07714 & ~w20883;
assign w37127 = ~pi02712 & w20883;
assign w37128 = ~w37126 & ~w37127;
assign w37129 = pi07715 & ~w20791;
assign w37130 = ~pi02167 & w20791;
assign w37131 = ~w37129 & ~w37130;
assign w37132 = pi07716 & ~w20883;
assign w37133 = ~pi02170 & w20883;
assign w37134 = ~w37132 & ~w37133;
assign w37135 = pi07717 & ~w20883;
assign w37136 = ~pi02713 & w20883;
assign w37137 = ~w37135 & ~w37136;
assign w37138 = pi07718 & ~w20791;
assign w37139 = ~pi02164 & w20791;
assign w37140 = ~w37138 & ~w37139;
assign w37141 = pi07719 & ~w20883;
assign w37142 = ~pi02714 & w20883;
assign w37143 = ~w37141 & ~w37142;
assign w37144 = pi07720 & ~w20883;
assign w37145 = ~pi02715 & w20883;
assign w37146 = ~w37144 & ~w37145;
assign w37147 = pi07721 & ~w20883;
assign w37148 = ~pi02716 & w20883;
assign w37149 = ~w37147 & ~w37148;
assign w37150 = pi07722 & ~w20883;
assign w37151 = ~pi02717 & w20883;
assign w37152 = ~w37150 & ~w37151;
assign w37153 = pi07723 & ~w20791;
assign w37154 = ~pi02719 & w20791;
assign w37155 = ~w37153 & ~w37154;
assign w37156 = pi07724 & ~w20553;
assign w37157 = ~pi02721 & w20553;
assign w37158 = ~w37156 & ~w37157;
assign w37159 = pi07725 & ~w20553;
assign w37160 = ~pi02169 & w20553;
assign w37161 = ~w37159 & ~w37160;
assign w37162 = pi07726 & ~w20751;
assign w37163 = ~pi02711 & w20751;
assign w37164 = ~w37162 & ~w37163;
assign w37165 = pi07727 & ~w20553;
assign w37166 = ~pi02718 & w20553;
assign w37167 = ~w37165 & ~w37166;
assign w37168 = pi07728 & ~w20553;
assign w37169 = ~pi02167 & w20553;
assign w37170 = ~w37168 & ~w37169;
assign w37171 = pi07729 & ~w20751;
assign w37172 = w17039 & w20209;
assign w37173 = ~w37171 & ~w37172;
assign w37174 = pi07730 & ~w20751;
assign w37175 = ~pi02713 & w20751;
assign w37176 = ~w37174 & ~w37175;
assign w37177 = pi07731 & ~w20553;
assign w37178 = ~pi02164 & w20553;
assign w37179 = ~w37177 & ~w37178;
assign w37180 = pi07732 & ~w20751;
assign w37181 = ~pi02714 & w20751;
assign w37182 = ~w37180 & ~w37181;
assign w37183 = pi07733 & ~w20751;
assign w37184 = ~pi02715 & w20751;
assign w37185 = ~w37183 & ~w37184;
assign w37186 = pi07734 & ~w20751;
assign w37187 = ~pi02716 & w20751;
assign w37188 = ~w37186 & ~w37187;
assign w37189 = pi07735 & ~w20751;
assign w37190 = ~pi02717 & w20751;
assign w37191 = ~w37189 & ~w37190;
assign w37192 = pi07736 & ~w20553;
assign w37193 = w17305 & w17594;
assign w37194 = ~w37192 & ~w37193;
assign w37195 = pi07737 & ~w20512;
assign w37196 = w17811 & w18022;
assign w37197 = ~w37195 & ~w37196;
assign w37198 = pi07738 & ~w20512;
assign w37199 = w17586 & w18022;
assign w37200 = ~w37198 & ~w37199;
assign w37201 = pi07739 & ~w20512;
assign w37202 = w18022 & w19797;
assign w37203 = ~w37201 & ~w37202;
assign w37204 = pi07740 & ~w20512;
assign w37205 = w18022 & w19273;
assign w37206 = ~w37204 & ~w37205;
assign w37207 = pi07741 & ~w20512;
assign w37208 = w18022 & w19312;
assign w37209 = ~w37207 & ~w37208;
assign w37210 = pi07742 & ~w20394;
assign w37211 = ~pi02711 & w20394;
assign w37212 = ~w37210 & ~w37211;
assign w37213 = pi07743 & ~w20394;
assign w37214 = ~pi02712 & w20394;
assign w37215 = ~w37213 & ~w37214;
assign w37216 = pi07744 & ~w20394;
assign w37217 = ~pi02170 & w20394;
assign w37218 = ~w37216 & ~w37217;
assign w37219 = pi07745 & ~w20394;
assign w37220 = ~pi02713 & w20394;
assign w37221 = ~w37219 & ~w37220;
assign w37222 = pi07746 & ~w20394;
assign w37223 = w17742 & w18454;
assign w37224 = ~w37222 & ~w37223;
assign w37225 = pi07747 & ~w20394;
assign w37226 = ~pi02716 & w20394;
assign w37227 = ~w37225 & ~w37226;
assign w37228 = pi07748 & ~w20512;
assign w37229 = w17594 & w18022;
assign w37230 = ~w37228 & ~w37229;
assign w37231 = pi07749 & ~w20394;
assign w37232 = ~pi02717 & w20394;
assign w37233 = ~w37231 & ~w37232;
assign w37234 = pi07750 & ~w20181;
assign w37235 = ~pi02712 & w20181;
assign w37236 = ~w37234 & ~w37235;
assign w37237 = pi07751 & ~w20181;
assign w37238 = ~pi02170 & w20181;
assign w37239 = ~w37237 & ~w37238;
assign w37240 = pi07752 & ~w20181;
assign w37241 = ~pi02713 & w20181;
assign w37242 = ~w37240 & ~w37241;
assign w37243 = pi07753 & ~w20181;
assign w37244 = w17710 & w18059;
assign w37245 = ~w37243 & ~w37244;
assign w37246 = pi07754 & ~w20181;
assign w37247 = ~pi02716 & w20181;
assign w37248 = ~w37246 & ~w37247;
assign w37249 = pi07755 & ~w20181;
assign w37250 = ~pi02717 & w20181;
assign w37251 = ~w37249 & ~w37250;
assign w37252 = pi07756 & ~w19967;
assign w37253 = ~pi02711 & w19967;
assign w37254 = ~w37252 & ~w37253;
assign w37255 = pi07757 & ~w19967;
assign w37256 = ~pi02712 & w19967;
assign w37257 = ~w37255 & ~w37256;
assign w37258 = pi07758 & ~w19967;
assign w37259 = ~pi02170 & w19967;
assign w37260 = ~w37258 & ~w37259;
assign w37261 = pi07759 & ~w19967;
assign w37262 = ~pi02713 & w19967;
assign w37263 = ~w37261 & ~w37262;
assign w37264 = pi07760 & ~w19967;
assign w37265 = ~pi02715 & w19967;
assign w37266 = ~w37264 & ~w37265;
assign w37267 = pi07761 & ~w19967;
assign w37268 = ~pi02716 & w19967;
assign w37269 = ~w37267 & ~w37268;
assign w37270 = pi07762 & ~w19967;
assign w37271 = ~pi02717 & w19967;
assign w37272 = ~w37270 & ~w37271;
assign w37273 = pi07763 & ~w18761;
assign w37274 = ~pi02712 & w18761;
assign w37275 = ~w37273 & ~w37274;
assign w37276 = pi07764 & ~w18761;
assign w37277 = ~pi02170 & w18761;
assign w37278 = ~w37276 & ~w37277;
assign w37279 = pi07765 & ~w18761;
assign w37280 = ~pi02713 & w18761;
assign w37281 = ~w37279 & ~w37280;
assign w37282 = pi07766 & ~w18761;
assign w37283 = ~pi02715 & w18761;
assign w37284 = ~w37282 & ~w37283;
assign w37285 = pi07767 & ~w18761;
assign w37286 = ~pi02716 & w18761;
assign w37287 = ~w37285 & ~w37286;
assign w37288 = pi07768 & ~w18761;
assign w37289 = ~pi02717 & w18761;
assign w37290 = ~w37288 & ~w37289;
assign w37291 = pi07769 & ~w18382;
assign w37292 = ~pi02711 & w18382;
assign w37293 = ~w37291 & ~w37292;
assign w37294 = pi07770 & ~w18382;
assign w37295 = ~pi02712 & w18382;
assign w37296 = ~w37294 & ~w37295;
assign w37297 = pi07771 & ~w18382;
assign w37298 = ~pi02170 & w18382;
assign w37299 = ~w37297 & ~w37298;
assign w37300 = pi07772 & ~w17950;
assign w37301 = ~pi02703 & w17950;
assign w37302 = ~w37300 & ~w37301;
assign w37303 = pi07773 & ~w18382;
assign w37304 = ~pi02714 & w18382;
assign w37305 = ~w37303 & ~w37304;
assign w37306 = pi07774 & ~w17950;
assign w37307 = ~pi02721 & w17950;
assign w37308 = ~w37306 & ~w37307;
assign w37309 = pi07775 & ~w18382;
assign w37310 = ~pi02716 & w18382;
assign w37311 = ~w37309 & ~w37310;
assign w37312 = pi07776 & ~w18382;
assign w37313 = w16973 & w17631;
assign w37314 = ~w37312 & ~w37313;
assign w37315 = pi07777 & ~w18382;
assign w37316 = ~pi02715 & w18382;
assign w37317 = ~w37315 & ~w37316;
assign w37318 = pi07778 & ~w17950;
assign w37319 = ~pi02718 & w17950;
assign w37320 = ~w37318 & ~w37319;
assign w37321 = pi07779 & ~w17950;
assign w37322 = ~pi02164 & w17950;
assign w37323 = ~w37321 & ~w37322;
assign w37324 = pi07780 & ~w17950;
assign w37325 = ~pi02722 & w17950;
assign w37326 = ~w37324 & ~w37325;
assign w37327 = pi07781 & ~w17674;
assign w37328 = ~pi02711 & w17674;
assign w37329 = ~w37327 & ~w37328;
assign w37330 = pi07782 & ~w17674;
assign w37331 = ~pi02712 & w17674;
assign w37332 = ~w37330 & ~w37331;
assign w37333 = pi07783 & ~w17674;
assign w37334 = ~pi02170 & w17674;
assign w37335 = ~w37333 & ~w37334;
assign w37336 = pi07784 & ~w17950;
assign w37337 = ~pi02719 & w17950;
assign w37338 = ~w37336 & ~w37337;
assign w37339 = pi07785 & ~w17674;
assign w37340 = ~pi02713 & w17674;
assign w37341 = ~w37339 & ~w37340;
assign w37342 = pi07786 & ~w17794;
assign w37343 = ~pi02703 & w17794;
assign w37344 = ~w37342 & ~w37343;
assign w37345 = pi07787 & ~w17674;
assign w37346 = ~pi02715 & w17674;
assign w37347 = ~w37345 & ~w37346;
assign w37348 = pi07788 & ~w17794;
assign w37349 = ~pi02721 & w17794;
assign w37350 = ~w37348 & ~w37349;
assign w37351 = pi07789 & ~w17674;
assign w37352 = ~pi02717 & w17674;
assign w37353 = ~w37351 & ~w37352;
assign w37354 = pi07790 & ~w17794;
assign w37355 = ~pi02169 & w17794;
assign w37356 = ~w37354 & ~w37355;
assign w37357 = pi07791 & ~w17794;
assign w37358 = ~pi02718 & w17794;
assign w37359 = ~w37357 & ~w37358;
assign w37360 = pi07792 & ~w17794;
assign w37361 = ~pi02164 & w17794;
assign w37362 = ~w37360 & ~w37361;
assign w37363 = pi07793 & ~w17794;
assign w37364 = ~pi02722 & w17794;
assign w37365 = ~w37363 & ~w37364;
assign w37366 = pi07794 & ~w17794;
assign w37367 = ~pi02719 & w17794;
assign w37368 = ~w37366 & ~w37367;
assign w37369 = pi07795 & ~w17615;
assign w37370 = ~pi02703 & w17615;
assign w37371 = ~w37369 & ~w37370;
assign w37372 = pi07796 & ~w17615;
assign w37373 = ~pi02721 & w17615;
assign w37374 = ~w37372 & ~w37373;
assign w37375 = pi07797 & ~w17315;
assign w37376 = ~pi02711 & w17315;
assign w37377 = ~w37375 & ~w37376;
assign w37378 = pi07798 & ~w17615;
assign w37379 = ~pi02169 & w17615;
assign w37380 = ~w37378 & ~w37379;
assign w37381 = pi07799 & ~w17615;
assign w37382 = ~pi02718 & w17615;
assign w37383 = ~w37381 & ~w37382;
assign w37384 = pi07800 & ~w17315;
assign w37385 = ~pi02170 & w17315;
assign w37386 = ~w37384 & ~w37385;
assign w37387 = pi07801 & ~w17315;
assign w37388 = w17314 & w17929;
assign w37389 = ~w37387 & ~w37388;
assign w37390 = pi07802 & ~w17315;
assign w37391 = ~pi02714 & w17315;
assign w37392 = ~w37390 & ~w37391;
assign w37393 = pi07803 & ~w17315;
assign w37394 = ~pi02715 & w17315;
assign w37395 = ~w37393 & ~w37394;
assign w37396 = pi07804 & ~w17615;
assign w37397 = ~pi02164 & w17615;
assign w37398 = ~w37396 & ~w37397;
assign w37399 = pi07805 & ~w17315;
assign w37400 = ~pi02717 & w17315;
assign w37401 = ~w37399 & ~w37400;
assign w37402 = ~w16905 & w17125;
assign w37403 = pi07806 & ~w37402;
assign w37404 = ~pi02711 & w37402;
assign w37405 = ~w37403 & ~w37404;
assign w37406 = pi07807 & ~w17615;
assign w37407 = ~pi02722 & w17615;
assign w37408 = ~w37406 & ~w37407;
assign w37409 = pi07808 & ~w37402;
assign w37410 = ~pi02712 & w37402;
assign w37411 = ~w37409 & ~w37410;
assign w37412 = pi07809 & ~w37402;
assign w37413 = w17125 & w20209;
assign w37414 = ~w37412 & ~w37413;
assign w37415 = pi07810 & ~w17615;
assign w37416 = w17594 & w17614;
assign w37417 = ~w37415 & ~w37416;
assign w37418 = pi07811 & ~w37402;
assign w37419 = ~pi02713 & w37402;
assign w37420 = ~w37418 & ~w37419;
assign w37421 = ~w16992 & w17526;
assign w37422 = pi07812 & ~w37421;
assign w37423 = ~pi02703 & w37421;
assign w37424 = ~w37422 & ~w37423;
assign w37425 = pi07813 & ~w37402;
assign w37426 = ~pi02715 & w37402;
assign w37427 = ~w37425 & ~w37426;
assign w37428 = pi07814 & ~w37402;
assign w37429 = ~pi02716 & w37402;
assign w37430 = ~w37428 & ~w37429;
assign w37431 = pi07815 & ~w37402;
assign w37432 = ~pi02717 & w37402;
assign w37433 = ~w37431 & ~w37432;
assign w37434 = pi07816 & ~w37421;
assign w37435 = ~pi02169 & w37421;
assign w37436 = ~w37434 & ~w37435;
assign w37437 = pi07817 & ~w37421;
assign w37438 = ~pi02718 & w37421;
assign w37439 = ~w37437 & ~w37438;
assign w37440 = pi07818 & ~w37421;
assign w37441 = ~pi02164 & w37421;
assign w37442 = ~w37440 & ~w37441;
assign w37443 = pi07819 & ~w37421;
assign w37444 = ~pi02722 & w37421;
assign w37445 = ~w37443 & ~w37444;
assign w37446 = pi07820 & ~w37421;
assign w37447 = ~pi02719 & w37421;
assign w37448 = ~w37446 & ~w37447;
assign w37449 = pi07821 & ~w21559;
assign w37450 = ~pi02703 & w21559;
assign w37451 = ~w37449 & ~w37450;
assign w37452 = pi07822 & ~w21559;
assign w37453 = ~pi02721 & w21559;
assign w37454 = ~w37452 & ~w37453;
assign w37455 = pi07823 & ~w33190;
assign w37456 = ~pi02711 & w33190;
assign w37457 = ~w37455 & ~w37456;
assign w37458 = pi07824 & ~w33190;
assign w37459 = w17020 & w17239;
assign w37460 = ~w37458 & ~w37459;
assign w37461 = pi07825 & ~w33190;
assign w37462 = ~pi02170 & w33190;
assign w37463 = ~w37461 & ~w37462;
assign w37464 = pi07826 & ~w33190;
assign w37465 = ~pi02713 & w33190;
assign w37466 = ~w37464 & ~w37465;
assign w37467 = pi07827 & ~w21559;
assign w37468 = ~pi02718 & w21559;
assign w37469 = ~w37467 & ~w37468;
assign w37470 = pi07828 & ~w21559;
assign w37471 = ~pi02167 & w21559;
assign w37472 = ~w37470 & ~w37471;
assign w37473 = pi07829 & ~w33190;
assign w37474 = ~pi02715 & w33190;
assign w37475 = ~w37473 & ~w37474;
assign w37476 = pi07830 & ~w21559;
assign w37477 = ~pi02164 & w21559;
assign w37478 = ~w37476 & ~w37477;
assign w37479 = pi07831 & ~w33190;
assign w37480 = ~pi02717 & w33190;
assign w37481 = ~w37479 & ~w37480;
assign w37482 = pi07832 & ~w26162;
assign w37483 = ~pi02711 & w26162;
assign w37484 = ~w37482 & ~w37483;
assign w37485 = pi07833 & ~w21559;
assign w37486 = ~pi02722 & w21559;
assign w37487 = ~w37485 & ~w37486;
assign w37488 = pi07834 & ~w26162;
assign w37489 = ~pi02712 & w26162;
assign w37490 = ~w37488 & ~w37489;
assign w37491 = pi07835 & ~w26162;
assign w37492 = ~pi02170 & w26162;
assign w37493 = ~w37491 & ~w37492;
assign w37494 = pi07836 & ~w21559;
assign w37495 = ~pi02719 & w21559;
assign w37496 = ~w37494 & ~w37495;
assign w37497 = pi07837 & ~w26162;
assign w37498 = ~pi02713 & w26162;
assign w37499 = ~w37497 & ~w37498;
assign w37500 = pi07838 & ~w21689;
assign w37501 = ~pi02703 & w21689;
assign w37502 = ~w37500 & ~w37501;
assign w37503 = pi07839 & ~w26162;
assign w37504 = w17167 & w18059;
assign w37505 = ~w37503 & ~w37504;
assign w37506 = pi07840 & ~w26162;
assign w37507 = ~pi02716 & w26162;
assign w37508 = ~w37506 & ~w37507;
assign w37509 = pi07841 & ~w26162;
assign w37510 = ~pi02717 & w26162;
assign w37511 = ~w37509 & ~w37510;
assign w37512 = pi07842 & ~w21689;
assign w37513 = ~pi02169 & w21689;
assign w37514 = ~w37512 & ~w37513;
assign w37515 = pi07843 & ~w21689;
assign w37516 = ~pi02718 & w21689;
assign w37517 = ~w37515 & ~w37516;
assign w37518 = pi07844 & ~w21689;
assign w37519 = ~pi02167 & w21689;
assign w37520 = ~w37518 & ~w37519;
assign w37521 = pi07845 & ~w21689;
assign w37522 = ~pi02164 & w21689;
assign w37523 = ~w37521 & ~w37522;
assign w37524 = pi07846 & ~w17269;
assign w37525 = ~pi02711 & w17269;
assign w37526 = ~w37524 & ~w37525;
assign w37527 = pi07847 & ~w21689;
assign w37528 = ~pi02722 & w21689;
assign w37529 = ~w37527 & ~w37528;
assign w37530 = pi07848 & ~w17269;
assign w37531 = w17020 & w17205;
assign w37532 = ~w37530 & ~w37531;
assign w37533 = pi07849 & ~w17269;
assign w37534 = ~pi02170 & w17269;
assign w37535 = ~w37533 & ~w37534;
assign w37536 = pi07850 & ~w21689;
assign w37537 = ~pi02719 & w21689;
assign w37538 = ~w37536 & ~w37537;
assign w37539 = pi07851 & ~w17269;
assign w37540 = w17205 & w17742;
assign w37541 = ~w37539 & ~w37540;
assign w37542 = ~w16992 & w21154;
assign w37543 = pi07852 & ~w37542;
assign w37544 = ~pi02703 & w37542;
assign w37545 = ~w37543 & ~w37544;
assign w37546 = pi07853 & ~w17269;
assign w37547 = ~pi02715 & w17269;
assign w37548 = ~w37546 & ~w37547;
assign w37549 = pi07854 & ~w37542;
assign w37550 = ~pi02721 & w37542;
assign w37551 = ~w37549 & ~w37550;
assign w37552 = pi07855 & ~w17269;
assign w37553 = ~pi02717 & w17269;
assign w37554 = ~w37552 & ~w37553;
assign w37555 = pi07856 & ~w20501;
assign w37556 = ~pi02711 & w20501;
assign w37557 = ~w37555 & ~w37556;
assign w37558 = pi07857 & ~w37542;
assign w37559 = ~pi02169 & w37542;
assign w37560 = ~w37558 & ~w37559;
assign w37561 = pi07858 & ~w37542;
assign w37562 = ~pi02718 & w37542;
assign w37563 = ~w37561 & ~w37562;
assign w37564 = pi07859 & ~w20501;
assign w37565 = ~pi02170 & w20501;
assign w37566 = ~w37564 & ~w37565;
assign w37567 = pi07860 & ~w20501;
assign w37568 = ~pi02713 & w20501;
assign w37569 = ~w37567 & ~w37568;
assign w37570 = pi07861 & ~w20501;
assign w37571 = ~pi02714 & w20501;
assign w37572 = ~w37570 & ~w37571;
assign w37573 = pi07862 & ~w20501;
assign w37574 = ~pi02715 & w20501;
assign w37575 = ~w37573 & ~w37574;
assign w37576 = pi07863 & ~w37542;
assign w37577 = w19273 & w21154;
assign w37578 = ~w37576 & ~w37577;
assign w37579 = pi07864 & ~w20501;
assign w37580 = ~pi02717 & w20501;
assign w37581 = ~w37579 & ~w37580;
assign w37582 = pi07865 & ~w21022;
assign w37583 = ~pi02711 & w21022;
assign w37584 = ~w37582 & ~w37583;
assign w37585 = pi07866 & ~w37542;
assign w37586 = ~pi02164 & w37542;
assign w37587 = ~w37585 & ~w37586;
assign w37588 = pi07867 & ~w37542;
assign w37589 = ~pi02722 & w37542;
assign w37590 = ~w37588 & ~w37589;
assign w37591 = pi07868 & ~w21022;
assign w37592 = ~pi02170 & w21022;
assign w37593 = ~w37591 & ~w37592;
assign w37594 = pi07869 & ~w37542;
assign w37595 = ~pi02719 & w37542;
assign w37596 = ~w37594 & ~w37595;
assign w37597 = pi07870 & ~w21022;
assign w37598 = ~pi02714 & w21022;
assign w37599 = ~w37597 & ~w37598;
assign w37600 = pi07871 & ~w20721;
assign w37601 = ~pi02703 & w20721;
assign w37602 = ~w37600 & ~w37601;
assign w37603 = pi07872 & ~w21022;
assign w37604 = ~pi02715 & w21022;
assign w37605 = ~w37603 & ~w37604;
assign w37606 = pi07873 & ~w21022;
assign w37607 = ~pi02716 & w21022;
assign w37608 = ~w37606 & ~w37607;
assign w37609 = pi07874 & ~w21022;
assign w37610 = w16973 & w17200;
assign w37611 = ~w37609 & ~w37610;
assign w37612 = pi07875 & ~w20787;
assign w37613 = ~pi02711 & w20787;
assign w37614 = ~w37612 & ~w37613;
assign w37615 = pi07876 & ~w20721;
assign w37616 = ~pi02721 & w20721;
assign w37617 = ~w37615 & ~w37616;
assign w37618 = pi07877 & ~w20721;
assign w37619 = ~pi02169 & w20721;
assign w37620 = ~w37618 & ~w37619;
assign w37621 = pi07878 & ~w20787;
assign w37622 = w17172 & w20209;
assign w37623 = ~w37621 & ~w37622;
assign w37624 = pi07879 & ~w20787;
assign w37625 = ~pi02713 & w20787;
assign w37626 = ~w37624 & ~w37625;
assign w37627 = pi07880 & ~w20787;
assign w37628 = ~pi02714 & w20787;
assign w37629 = ~w37627 & ~w37628;
assign w37630 = pi07881 & ~w20787;
assign w37631 = ~pi02715 & w20787;
assign w37632 = ~w37630 & ~w37631;
assign w37633 = pi07882 & ~w20721;
assign w37634 = ~pi02167 & w20721;
assign w37635 = ~w37633 & ~w37634;
assign w37636 = pi07883 & ~w20787;
assign w37637 = ~pi02717 & w20787;
assign w37638 = ~w37636 & ~w37637;
assign w37639 = pi07884 & ~w20743;
assign w37640 = ~pi02711 & w20743;
assign w37641 = ~w37639 & ~w37640;
assign w37642 = pi07885 & ~w20721;
assign w37643 = ~pi02164 & w20721;
assign w37644 = ~w37642 & ~w37643;
assign w37645 = pi07886 & ~w20743;
assign w37646 = ~pi02712 & w20743;
assign w37647 = ~w37645 & ~w37646;
assign w37648 = pi07887 & ~w20743;
assign w37649 = ~pi02170 & w20743;
assign w37650 = ~w37648 & ~w37649;
assign w37651 = pi07888 & ~w20721;
assign w37652 = ~pi02722 & w20721;
assign w37653 = ~w37651 & ~w37652;
assign w37654 = pi07889 & ~w20743;
assign w37655 = ~pi02713 & w20743;
assign w37656 = ~w37654 & ~w37655;
assign w37657 = pi07890 & ~w20743;
assign w37658 = ~pi02714 & w20743;
assign w37659 = ~w37657 & ~w37658;
assign w37660 = ~w16992 & w18631;
assign w37661 = pi07891 & ~w37660;
assign w37662 = ~pi02703 & w37660;
assign w37663 = ~w37661 & ~w37662;
assign w37664 = pi07892 & ~w37660;
assign w37665 = ~pi02721 & w37660;
assign w37666 = ~w37664 & ~w37665;
assign w37667 = pi07893 & ~w20743;
assign w37668 = ~pi02716 & w20743;
assign w37669 = ~w37667 & ~w37668;
assign w37670 = pi07894 & ~w20743;
assign w37671 = ~pi02717 & w20743;
assign w37672 = ~w37670 & ~w37671;
assign w37673 = pi07895 & ~w18741;
assign w37674 = ~pi02711 & w18741;
assign w37675 = ~w37673 & ~w37674;
assign w37676 = pi07896 & ~w37660;
assign w37677 = ~pi02169 & w37660;
assign w37678 = ~w37676 & ~w37677;
assign w37679 = pi07897 & ~w18741;
assign w37680 = ~pi02170 & w18741;
assign w37681 = ~w37679 & ~w37680;
assign w37682 = pi07898 & ~w18741;
assign w37683 = ~pi02713 & w18741;
assign w37684 = ~w37682 & ~w37683;
assign w37685 = pi07899 & ~w37660;
assign w37686 = ~pi02718 & w37660;
assign w37687 = ~w37685 & ~w37686;
assign w37688 = pi07900 & ~w18741;
assign w37689 = ~pi02714 & w18741;
assign w37690 = ~w37688 & ~w37689;
assign w37691 = pi07901 & ~w18741;
assign w37692 = ~pi02715 & w18741;
assign w37693 = ~w37691 & ~w37692;
assign w37694 = pi07902 & ~w37660;
assign w37695 = ~pi02167 & w37660;
assign w37696 = ~w37694 & ~w37695;
assign w37697 = pi07903 & ~w18741;
assign w37698 = ~pi02717 & w18741;
assign w37699 = ~w37697 & ~w37698;
assign w37700 = pi07904 & ~w20269;
assign w37701 = ~pi02711 & w20269;
assign w37702 = ~w37700 & ~w37701;
assign w37703 = pi07905 & ~w37660;
assign w37704 = ~pi02164 & w37660;
assign w37705 = ~w37703 & ~w37704;
assign w37706 = pi07906 & ~w20269;
assign w37707 = ~pi02170 & w20269;
assign w37708 = ~w37706 & ~w37707;
assign w37709 = pi07907 & ~w37660;
assign w37710 = ~pi02722 & w37660;
assign w37711 = ~w37709 & ~w37710;
assign w37712 = pi07908 & ~w20269;
assign w37713 = ~pi02713 & w20269;
assign w37714 = ~w37712 & ~w37713;
assign w37715 = pi07909 & ~w37660;
assign w37716 = ~pi02719 & w37660;
assign w37717 = ~w37715 & ~w37716;
assign w37718 = pi07910 & ~w20269;
assign w37719 = ~pi02715 & w20269;
assign w37720 = ~w37718 & ~w37719;
assign w37721 = pi07911 & ~w20269;
assign w37722 = w17317 & w17479;
assign w37723 = ~w37721 & ~w37722;
assign w37724 = pi07912 & ~w20204;
assign w37725 = ~pi02703 & w20204;
assign w37726 = ~w37724 & ~w37725;
assign w37727 = pi07913 & ~w20204;
assign w37728 = ~pi02721 & w20204;
assign w37729 = ~w37727 & ~w37728;
assign w37730 = pi07914 & ~w20269;
assign w37731 = ~pi02717 & w20269;
assign w37732 = ~w37730 & ~w37731;
assign w37733 = pi07915 & ~w20193;
assign w37734 = ~pi02711 & w20193;
assign w37735 = ~w37733 & ~w37734;
assign w37736 = pi07916 & ~w20204;
assign w37737 = ~pi02169 & w20204;
assign w37738 = ~w37736 & ~w37737;
assign w37739 = pi07917 & ~w20193;
assign w37740 = ~pi02170 & w20193;
assign w37741 = ~w37739 & ~w37740;
assign w37742 = pi07918 & ~w20193;
assign w37743 = ~pi02713 & w20193;
assign w37744 = ~w37742 & ~w37743;
assign w37745 = pi07919 & ~w20193;
assign w37746 = ~pi02714 & w20193;
assign w37747 = ~w37745 & ~w37746;
assign w37748 = pi07920 & ~w20193;
assign w37749 = ~pi02715 & w20193;
assign w37750 = ~w37748 & ~w37749;
assign w37751 = pi07921 & ~w20204;
assign w37752 = ~pi02167 & w20204;
assign w37753 = ~w37751 & ~w37752;
assign w37754 = pi07922 & ~w20193;
assign w37755 = ~pi02717 & w20193;
assign w37756 = ~w37754 & ~w37755;
assign w37757 = pi07923 & ~w18757;
assign w37758 = ~pi02711 & w18757;
assign w37759 = ~w37757 & ~w37758;
assign w37760 = pi07924 & ~w20204;
assign w37761 = ~pi02164 & w20204;
assign w37762 = ~w37760 & ~w37761;
assign w37763 = pi07925 & ~w18757;
assign w37764 = w17020 & w17114;
assign w37765 = ~w37763 & ~w37764;
assign w37766 = pi07926 & ~w18757;
assign w37767 = ~pi02170 & w18757;
assign w37768 = ~w37766 & ~w37767;
assign w37769 = pi07927 & ~w20204;
assign w37770 = ~pi02722 & w20204;
assign w37771 = ~w37769 & ~w37770;
assign w37772 = pi07928 & ~w18757;
assign w37773 = ~pi02713 & w18757;
assign w37774 = ~w37772 & ~w37773;
assign w37775 = pi07929 & ~w20204;
assign w37776 = ~pi02719 & w20204;
assign w37777 = ~w37775 & ~w37776;
assign w37778 = pi07930 & ~w18757;
assign w37779 = ~pi02715 & w18757;
assign w37780 = ~w37778 & ~w37779;
assign w37781 = pi07931 & ~w18757;
assign w37782 = w17114 & w17317;
assign w37783 = ~w37781 & ~w37782;
assign w37784 = ~w16992 & w20775;
assign w37785 = pi07932 & ~w37784;
assign w37786 = ~pi02703 & w37784;
assign w37787 = ~w37785 & ~w37786;
assign w37788 = pi07933 & ~w18757;
assign w37789 = ~pi02717 & w18757;
assign w37790 = ~w37788 & ~w37789;
assign w37791 = pi07934 & ~w17548;
assign w37792 = ~pi02711 & w17548;
assign w37793 = ~w37791 & ~w37792;
assign w37794 = pi07935 & ~w36472;
assign w37795 = w17532 & w20561;
assign w37796 = ~w37794 & ~w37795;
assign w37797 = pi07936 & ~w37784;
assign w37798 = ~pi02721 & w37784;
assign w37799 = ~w37797 & ~w37798;
assign w37800 = pi07937 & ~w17548;
assign w37801 = w17249 & w20209;
assign w37802 = ~w37800 & ~w37801;
assign w37803 = pi07938 & ~w37784;
assign w37804 = ~pi02169 & w37784;
assign w37805 = ~w37803 & ~w37804;
assign w37806 = pi07939 & ~w17548;
assign w37807 = ~pi02713 & w17548;
assign w37808 = ~w37806 & ~w37807;
assign w37809 = pi07940 & ~w37784;
assign w37810 = ~pi02718 & w37784;
assign w37811 = ~w37809 & ~w37810;
assign w37812 = pi07941 & ~w17548;
assign w37813 = w17249 & w17742;
assign w37814 = ~w37812 & ~w37813;
assign w37815 = pi07942 & ~w17548;
assign w37816 = ~pi02715 & w17548;
assign w37817 = ~w37815 & ~w37816;
assign w37818 = pi07943 & ~w37784;
assign w37819 = ~pi02167 & w37784;
assign w37820 = ~w37818 & ~w37819;
assign w37821 = pi07944 & ~w17548;
assign w37822 = ~pi02717 & w17548;
assign w37823 = ~w37821 & ~w37822;
assign w37824 = pi07945 & ~w17561;
assign w37825 = ~pi02711 & w17561;
assign w37826 = ~w37824 & ~w37825;
assign w37827 = pi07946 & ~w37784;
assign w37828 = w17620 & w20775;
assign w37829 = ~w37827 & ~w37828;
assign w37830 = pi07947 & ~w17561;
assign w37831 = w17047 & w20209;
assign w37832 = ~w37830 & ~w37831;
assign w37833 = pi07948 & ~w37784;
assign w37834 = w17594 & w20775;
assign w37835 = ~w37833 & ~w37834;
assign w37836 = pi07949 & ~w17561;
assign w37837 = ~pi02714 & w17561;
assign w37838 = ~w37836 & ~w37837;
assign w37839 = pi07950 & ~w17561;
assign w37840 = w17047 & w18059;
assign w37841 = ~w37839 & ~w37840;
assign w37842 = pi07951 & ~w17561;
assign w37843 = w17047 & w17317;
assign w37844 = ~w37842 & ~w37843;
assign w37845 = pi07952 & ~w37784;
assign w37846 = ~pi02722 & w37784;
assign w37847 = ~w37845 & ~w37846;
assign w37848 = pi07953 & ~w17561;
assign w37849 = ~pi02717 & w17561;
assign w37850 = ~w37848 & ~w37849;
assign w37851 = pi07954 & ~w17584;
assign w37852 = w17532 & w17583;
assign w37853 = ~w37851 & ~w37852;
assign w37854 = pi07955 & ~w17584;
assign w37855 = w17583 & w17811;
assign w37856 = ~w37854 & ~w37855;
assign w37857 = pi07956 & ~w17584;
assign w37858 = w17583 & w19797;
assign w37859 = ~w37857 & ~w37858;
assign w37860 = pi07957 & ~w17584;
assign w37861 = w17583 & w19273;
assign w37862 = ~w37860 & ~w37861;
assign w37863 = pi07958 & ~w17491;
assign w37864 = ~pi02711 & w17491;
assign w37865 = ~w37863 & ~w37864;
assign w37866 = pi07959 & ~w17491;
assign w37867 = ~pi02712 & w17491;
assign w37868 = ~w37866 & ~w37867;
assign w37869 = pi07960 & ~w17491;
assign w37870 = ~pi02170 & w17491;
assign w37871 = ~w37869 & ~w37870;
assign w37872 = pi07961 & ~w17584;
assign w37873 = w17583 & w19312;
assign w37874 = ~w37872 & ~w37873;
assign w37875 = pi07962 & ~w17491;
assign w37876 = ~pi02714 & w17491;
assign w37877 = ~w37875 & ~w37876;
assign w37878 = pi07963 & ~w17584;
assign w37879 = w17583 & w17594;
assign w37880 = ~w37878 & ~w37879;
assign w37881 = pi07964 & ~w17491;
assign w37882 = ~pi02715 & w17491;
assign w37883 = ~w37881 & ~w37882;
assign w37884 = pi07965 & ~w17491;
assign w37885 = ~pi02716 & w17491;
assign w37886 = ~w37884 & ~w37885;
assign w37887 = pi07966 & ~w21527;
assign w37888 = ~pi02703 & w21527;
assign w37889 = ~w37887 & ~w37888;
assign w37890 = pi07967 & ~w17491;
assign w37891 = ~pi02717 & w17491;
assign w37892 = ~w37890 & ~w37891;
assign w37893 = pi07968 & ~w21527;
assign w37894 = w17811 & w20566;
assign w37895 = ~w37893 & ~w37894;
assign w37896 = pi07969 & ~w21527;
assign w37897 = w17586 & w20566;
assign w37898 = ~w37896 & ~w37897;
assign w37899 = pi07970 & ~w21527;
assign w37900 = ~pi02167 & w21527;
assign w37901 = ~w37899 & ~w37900;
assign w37902 = ~w16905 & w18645;
assign w37903 = pi07971 & ~w37902;
assign w37904 = ~pi02711 & w37902;
assign w37905 = ~w37903 & ~w37904;
assign w37906 = pi07972 & ~w37902;
assign w37907 = ~pi02712 & w37902;
assign w37908 = ~w37906 & ~w37907;
assign w37909 = pi07973 & ~w37902;
assign w37910 = ~pi02170 & w37902;
assign w37911 = ~w37909 & ~w37910;
assign w37912 = pi07974 & ~w21527;
assign w37913 = ~pi02722 & w21527;
assign w37914 = ~w37912 & ~w37913;
assign w37915 = pi07975 & ~w37902;
assign w37916 = ~pi02714 & w37902;
assign w37917 = ~w37915 & ~w37916;
assign w37918 = pi07976 & ~w21527;
assign w37919 = ~pi02719 & w21527;
assign w37920 = ~w37918 & ~w37919;
assign w37921 = pi07977 & ~w37902;
assign w37922 = ~pi02715 & w37902;
assign w37923 = ~w37921 & ~w37922;
assign w37924 = pi07978 & ~w37902;
assign w37925 = ~pi02716 & w37902;
assign w37926 = ~w37924 & ~w37925;
assign w37927 = pi07979 & ~w21220;
assign w37928 = ~pi02703 & w21220;
assign w37929 = ~w37927 & ~w37928;
assign w37930 = pi07980 & ~w37902;
assign w37931 = ~pi02717 & w37902;
assign w37932 = ~w37930 & ~w37931;
assign w37933 = pi07981 & ~w21220;
assign w37934 = ~pi02721 & w21220;
assign w37935 = ~w37933 & ~w37934;
assign w37936 = pi07982 & ~w21220;
assign w37937 = ~pi02718 & w21220;
assign w37938 = ~w37936 & ~w37937;
assign w37939 = pi07983 & ~w27432;
assign w37940 = ~pi02711 & w27432;
assign w37941 = ~w37939 & ~w37940;
assign w37942 = pi07984 & ~w21220;
assign w37943 = ~pi02167 & w21220;
assign w37944 = ~w37942 & ~w37943;
assign w37945 = pi07985 & ~w27432;
assign w37946 = ~pi02712 & w27432;
assign w37947 = ~w37945 & ~w37946;
assign w37948 = pi07986 & ~w27432;
assign w37949 = ~pi02170 & w27432;
assign w37950 = ~w37948 & ~w37949;
assign w37951 = pi07987 & ~w21220;
assign w37952 = ~pi02722 & w21220;
assign w37953 = ~w37951 & ~w37952;
assign w37954 = pi07988 & ~w27432;
assign w37955 = ~pi02714 & w27432;
assign w37956 = ~w37954 & ~w37955;
assign w37957 = pi07989 & ~w27432;
assign w37958 = ~pi02715 & w27432;
assign w37959 = ~w37957 & ~w37958;
assign w37960 = pi07990 & ~w27432;
assign w37961 = ~pi02716 & w27432;
assign w37962 = ~w37960 & ~w37961;
assign w37963 = pi07991 & ~w22146;
assign w37964 = ~pi02703 & w22146;
assign w37965 = ~w37963 & ~w37964;
assign w37966 = pi07992 & ~w27432;
assign w37967 = ~pi02717 & w27432;
assign w37968 = ~w37966 & ~w37967;
assign w37969 = pi07993 & ~w21220;
assign w37970 = ~pi02719 & w21220;
assign w37971 = ~w37969 & ~w37970;
assign w37972 = pi07994 & ~w18727;
assign w37973 = ~pi09962 & w18727;
assign w37974 = ~w37972 & ~w37973;
assign w37975 = pi07995 & ~w22146;
assign w37976 = ~pi02169 & w22146;
assign w37977 = ~w37975 & ~w37976;
assign w37978 = pi07996 & ~w22146;
assign w37979 = ~pi02718 & w22146;
assign w37980 = ~w37978 & ~w37979;
assign w37981 = pi07997 & ~w22146;
assign w37982 = ~pi02167 & w22146;
assign w37983 = ~w37981 & ~w37982;
assign w37984 = pi07998 & ~w22146;
assign w37985 = ~pi02164 & w22146;
assign w37986 = ~w37984 & ~w37985;
assign w37987 = pi07999 & ~w22146;
assign w37988 = ~pi02719 & w22146;
assign w37989 = ~w37987 & ~w37988;
assign w37990 = pi08000 & ~w21496;
assign w37991 = ~pi02703 & w21496;
assign w37992 = ~w37990 & ~w37991;
assign w37993 = pi08001 & ~w21289;
assign w37994 = ~pi02712 & w21289;
assign w37995 = ~w37993 & ~w37994;
assign w37996 = pi08002 & ~w21496;
assign w37997 = ~pi02721 & w21496;
assign w37998 = ~w37996 & ~w37997;
assign w37999 = pi08003 & ~w21289;
assign w38000 = ~pi02170 & w21289;
assign w38001 = ~w37999 & ~w38000;
assign w38002 = pi08004 & ~w21289;
assign w38003 = ~pi02713 & w21289;
assign w38004 = ~w38002 & ~w38003;
assign w38005 = pi08005 & ~w21496;
assign w38006 = ~pi02169 & w21496;
assign w38007 = ~w38005 & ~w38006;
assign w38008 = pi08006 & ~w21289;
assign w38009 = ~pi02714 & w21289;
assign w38010 = ~w38008 & ~w38009;
assign w38011 = pi08007 & ~w21289;
assign w38012 = ~pi02715 & w21289;
assign w38013 = ~w38011 & ~w38012;
assign w38014 = pi08008 & ~w21289;
assign w38015 = ~pi02716 & w21289;
assign w38016 = ~w38014 & ~w38015;
assign w38017 = pi08009 & ~w21289;
assign w38018 = ~pi02717 & w21289;
assign w38019 = ~w38017 & ~w38018;
assign w38020 = pi08010 & ~w21510;
assign w38021 = ~pi02711 & w21510;
assign w38022 = ~w38020 & ~w38021;
assign w38023 = pi08011 & ~w21510;
assign w38024 = ~pi02712 & w21510;
assign w38025 = ~w38023 & ~w38024;
assign w38026 = pi08012 & ~w21510;
assign w38027 = ~pi02170 & w21510;
assign w38028 = ~w38026 & ~w38027;
assign w38029 = pi08013 & ~w21496;
assign w38030 = ~pi02164 & w21496;
assign w38031 = ~w38029 & ~w38030;
assign w38032 = pi08014 & ~w21510;
assign w38033 = ~pi02714 & w21510;
assign w38034 = ~w38032 & ~w38033;
assign w38035 = pi08015 & ~w21496;
assign w38036 = ~pi02719 & w21496;
assign w38037 = ~w38035 & ~w38036;
assign w38038 = pi08016 & ~w21510;
assign w38039 = ~pi02715 & w21510;
assign w38040 = ~w38038 & ~w38039;
assign w38041 = pi08017 & ~w21510;
assign w38042 = ~pi02716 & w21510;
assign w38043 = ~w38041 & ~w38042;
assign w38044 = pi08018 & ~w21496;
assign w38045 = ~pi02722 & w21496;
assign w38046 = ~w38044 & ~w38045;
assign w38047 = pi08019 & ~w21510;
assign w38048 = ~pi02717 & w21510;
assign w38049 = ~w38047 & ~w38048;
assign w38050 = pi08020 & ~w21052;
assign w38051 = ~pi02711 & w21052;
assign w38052 = ~w38050 & ~w38051;
assign w38053 = pi08021 & ~w21052;
assign w38054 = ~pi02170 & w21052;
assign w38055 = ~w38053 & ~w38054;
assign w38056 = pi08022 & ~w21052;
assign w38057 = ~pi02713 & w21052;
assign w38058 = ~w38056 & ~w38057;
assign w38059 = pi08023 & ~w21052;
assign w38060 = ~pi02714 & w21052;
assign w38061 = ~w38059 & ~w38060;
assign w38062 = pi08024 & ~w21052;
assign w38063 = ~pi02716 & w21052;
assign w38064 = ~w38062 & ~w38063;
assign w38065 = pi08025 & ~w21052;
assign w38066 = ~pi02717 & w21052;
assign w38067 = ~w38065 & ~w38066;
assign w38068 = pi08026 & ~w20817;
assign w38069 = ~pi02711 & w20817;
assign w38070 = ~w38068 & ~w38069;
assign w38071 = pi08027 & ~w20795;
assign w38072 = ~pi02703 & w20795;
assign w38073 = ~w38071 & ~w38072;
assign w38074 = pi08028 & ~w20817;
assign w38075 = ~pi02170 & w20817;
assign w38076 = ~w38074 & ~w38075;
assign w38077 = pi08029 & ~w20795;
assign w38078 = ~pi02721 & w20795;
assign w38079 = ~w38077 & ~w38078;
assign w38080 = pi08030 & ~w20817;
assign w38081 = ~pi02713 & w20817;
assign w38082 = ~w38080 & ~w38081;
assign w38083 = pi08031 & ~w20817;
assign w38084 = ~pi02714 & w20817;
assign w38085 = ~w38083 & ~w38084;
assign w38086 = pi08032 & ~w20817;
assign w38087 = w17556 & w18059;
assign w38088 = ~w38086 & ~w38087;
assign w38089 = pi08033 & ~w20795;
assign w38090 = ~pi02169 & w20795;
assign w38091 = ~w38089 & ~w38090;
assign w38092 = pi08034 & ~w20817;
assign w38093 = ~pi02717 & w20817;
assign w38094 = ~w38092 & ~w38093;
assign w38095 = pi08035 & ~w20795;
assign w38096 = ~pi02718 & w20795;
assign w38097 = ~w38095 & ~w38096;
assign w38098 = pi08036 & ~w20795;
assign w38099 = ~pi02167 & w20795;
assign w38100 = ~w38098 & ~w38099;
assign w38101 = pi08037 & ~w20795;
assign w38102 = ~pi02722 & w20795;
assign w38103 = ~w38101 & ~w38102;
assign w38104 = pi08038 & ~w20795;
assign w38105 = ~pi02719 & w20795;
assign w38106 = ~w38104 & ~w38105;
assign w38107 = pi08039 & ~w20680;
assign w38108 = ~pi02711 & w20680;
assign w38109 = ~w38107 & ~w38108;
assign w38110 = pi08040 & ~w20680;
assign w38111 = ~pi02170 & w20680;
assign w38112 = ~w38110 & ~w38111;
assign w38113 = pi08041 & ~w20680;
assign w38114 = ~pi02713 & w20680;
assign w38115 = ~w38113 & ~w38114;
assign w38116 = pi08042 & ~w20680;
assign w38117 = ~pi02714 & w20680;
assign w38118 = ~w38116 & ~w38117;
assign w38119 = pi08043 & ~w20680;
assign w38120 = ~pi02715 & w20680;
assign w38121 = ~w38119 & ~w38120;
assign w38122 = pi08044 & ~w20680;
assign w38123 = ~pi02716 & w20680;
assign w38124 = ~w38122 & ~w38123;
assign w38125 = pi08045 & ~w20680;
assign w38126 = ~pi02717 & w20680;
assign w38127 = ~w38125 & ~w38126;
assign w38128 = pi08046 & ~w20226;
assign w38129 = ~pi02703 & w20226;
assign w38130 = ~w38128 & ~w38129;
assign w38131 = pi08047 & ~w20226;
assign w38132 = w17907 & w19797;
assign w38133 = ~w38131 & ~w38132;
assign w38134 = pi08048 & ~w20226;
assign w38135 = w17586 & w17907;
assign w38136 = ~w38134 & ~w38135;
assign w38137 = pi08049 & ~w20155;
assign w38138 = ~pi02711 & w20155;
assign w38139 = ~w38137 & ~w38138;
assign w38140 = pi08050 & ~w20155;
assign w38141 = ~pi02712 & w20155;
assign w38142 = ~w38140 & ~w38141;
assign w38143 = pi08051 & ~w20155;
assign w38144 = ~pi02170 & w20155;
assign w38145 = ~w38143 & ~w38144;
assign w38146 = pi08052 & ~w20226;
assign w38147 = ~pi02164 & w20226;
assign w38148 = ~w38146 & ~w38147;
assign w38149 = pi08053 & ~w20155;
assign w38150 = ~pi02714 & w20155;
assign w38151 = ~w38149 & ~w38150;
assign w38152 = pi08054 & ~w20226;
assign w38153 = ~pi02722 & w20226;
assign w38154 = ~w38152 & ~w38153;
assign w38155 = pi08055 & ~w20155;
assign w38156 = ~pi02715 & w20155;
assign w38157 = ~w38155 & ~w38156;
assign w38158 = pi08056 & ~w20155;
assign w38159 = ~pi02716 & w20155;
assign w38160 = ~w38158 & ~w38159;
assign w38161 = pi08057 & ~w20226;
assign w38162 = w17594 & w17907;
assign w38163 = ~w38161 & ~w38162;
assign w38164 = pi08058 & ~w20155;
assign w38165 = ~pi02717 & w20155;
assign w38166 = ~w38164 & ~w38165;
assign w38167 = pi08059 & ~w20189;
assign w38168 = w17119 & w17603;
assign w38169 = ~w38167 & ~w38168;
assign w38170 = pi08060 & ~w20000;
assign w38171 = w17532 & w17754;
assign w38172 = ~w38170 & ~w38171;
assign w38173 = pi08061 & ~w20189;
assign w38174 = ~pi02170 & w20189;
assign w38175 = ~w38173 & ~w38174;
assign w38176 = pi08062 & ~w20189;
assign w38177 = ~pi02713 & w20189;
assign w38178 = ~w38176 & ~w38177;
assign w38179 = pi08063 & ~w20189;
assign w38180 = ~pi02714 & w20189;
assign w38181 = ~w38179 & ~w38180;
assign w38182 = pi08064 & ~w20189;
assign w38183 = ~pi02715 & w20189;
assign w38184 = ~w38182 & ~w38183;
assign w38185 = pi08065 & ~w20189;
assign w38186 = ~pi02716 & w20189;
assign w38187 = ~w38185 & ~w38186;
assign w38188 = pi08066 & ~w20189;
assign w38189 = ~pi02717 & w20189;
assign w38190 = ~w38188 & ~w38189;
assign w38191 = pi08067 & ~w20000;
assign w38192 = w17586 & w17754;
assign w38193 = ~w38191 & ~w38192;
assign w38194 = pi08068 & ~w20000;
assign w38195 = w17754 & w19273;
assign w38196 = ~w38194 & ~w38195;
assign w38197 = pi08069 & ~w20000;
assign w38198 = w17620 & w17754;
assign w38199 = ~w38197 & ~w38198;
assign w38200 = pi08070 & ~w20000;
assign w38201 = w17754 & w19312;
assign w38202 = ~w38200 & ~w38201;
assign w38203 = pi08071 & ~w20000;
assign w38204 = w17594 & w17754;
assign w38205 = ~w38203 & ~w38204;
assign w38206 = pi08072 & ~w19545;
assign w38207 = ~pi02703 & w19545;
assign w38208 = ~w38206 & ~w38207;
assign w38209 = pi08073 & ~w19545;
assign w38210 = ~pi02169 & w19545;
assign w38211 = ~w38209 & ~w38210;
assign w38212 = pi08074 & ~w19406;
assign w38213 = ~pi02711 & w19406;
assign w38214 = ~w38212 & ~w38213;
assign w38215 = pi08075 & ~w19545;
assign w38216 = ~pi02718 & w19545;
assign w38217 = ~w38215 & ~w38216;
assign w38218 = pi08076 & ~w19406;
assign w38219 = ~pi02170 & w19406;
assign w38220 = ~w38218 & ~w38219;
assign w38221 = pi08077 & ~w19545;
assign w38222 = ~pi02167 & w19545;
assign w38223 = ~w38221 & ~w38222;
assign w38224 = pi08078 & ~w19406;
assign w38225 = ~pi02713 & w19406;
assign w38226 = ~w38224 & ~w38225;
assign w38227 = pi08079 & ~w19545;
assign w38228 = ~pi02164 & w19545;
assign w38229 = ~w38227 & ~w38228;
assign w38230 = pi08080 & ~w19406;
assign w38231 = ~pi02715 & w19406;
assign w38232 = ~w38230 & ~w38231;
assign w38233 = pi08081 & ~w19406;
assign w38234 = ~pi02716 & w19406;
assign w38235 = ~w38233 & ~w38234;
assign w38236 = pi08082 & ~w19545;
assign w38237 = ~pi02722 & w19545;
assign w38238 = ~w38236 & ~w38237;
assign w38239 = pi08083 & ~w19406;
assign w38240 = ~pi02717 & w19406;
assign w38241 = ~w38239 & ~w38240;
assign w38242 = pi08084 & ~w18804;
assign w38243 = ~pi02711 & w18804;
assign w38244 = ~w38242 & ~w38243;
assign w38245 = pi08085 & ~w19545;
assign w38246 = ~pi02719 & w19545;
assign w38247 = ~w38245 & ~w38246;
assign w38248 = pi08086 & ~w17552;
assign w38249 = ~pi02703 & w17552;
assign w38250 = ~w38248 & ~w38249;
assign w38251 = pi08087 & ~w18804;
assign w38252 = ~pi02170 & w18804;
assign w38253 = ~w38251 & ~w38252;
assign w38254 = pi08088 & ~w18804;
assign w38255 = ~pi02713 & w18804;
assign w38256 = ~w38254 & ~w38255;
assign w38257 = pi08089 & ~w18804;
assign w38258 = ~pi02714 & w18804;
assign w38259 = ~w38257 & ~w38258;
assign w38260 = pi08090 & ~w18804;
assign w38261 = ~pi02715 & w18804;
assign w38262 = ~w38260 & ~w38261;
assign w38263 = pi08091 & ~w17552;
assign w38264 = ~pi02169 & w17552;
assign w38265 = ~w38263 & ~w38264;
assign w38266 = pi08092 & ~w18804;
assign w38267 = ~pi02716 & w18804;
assign w38268 = ~w38266 & ~w38267;
assign w38269 = pi08093 & ~w18804;
assign w38270 = ~pi02717 & w18804;
assign w38271 = ~w38269 & ~w38270;
assign w38272 = pi08094 & ~w17946;
assign w38273 = ~pi02711 & w17946;
assign w38274 = ~w38272 & ~w38273;
assign w38275 = pi08095 & ~w17946;
assign w38276 = w17020 & w17259;
assign w38277 = ~w38275 & ~w38276;
assign w38278 = pi08096 & ~w17946;
assign w38279 = ~pi02170 & w17946;
assign w38280 = ~w38278 & ~w38279;
assign w38281 = pi08097 & ~w17552;
assign w38282 = ~pi02167 & w17552;
assign w38283 = ~w38281 & ~w38282;
assign w38284 = pi08098 & ~w17946;
assign w38285 = ~pi02713 & w17946;
assign w38286 = ~w38284 & ~w38285;
assign w38287 = pi08099 & ~w17552;
assign w38288 = ~pi02164 & w17552;
assign w38289 = ~w38287 & ~w38288;
assign w38290 = pi08100 & ~w17946;
assign w38291 = ~pi02715 & w17946;
assign w38292 = ~w38290 & ~w38291;
assign w38293 = pi08101 & ~w17946;
assign w38294 = w17259 & w17317;
assign w38295 = ~w38293 & ~w38294;
assign w38296 = pi08102 & ~w17552;
assign w38297 = ~pi02719 & w17552;
assign w38298 = ~w38296 & ~w38297;
assign w38299 = pi08103 & ~w17946;
assign w38300 = ~pi02717 & w17946;
assign w38301 = ~w38299 & ~w38300;
assign w38302 = pi08104 & ~w17763;
assign w38303 = ~pi02711 & w17763;
assign w38304 = ~w38302 & ~w38303;
assign w38305 = pi08105 & ~w17763;
assign w38306 = ~pi02170 & w17763;
assign w38307 = ~w38305 & ~w38306;
assign w38308 = pi08106 & ~w17763;
assign w38309 = ~pi02713 & w17763;
assign w38310 = ~w38308 & ~w38309;
assign w38311 = ~w16992 & w17938;
assign w38312 = pi08107 & ~w38311;
assign w38313 = ~pi02703 & w38311;
assign w38314 = ~w38312 & ~w38313;
assign w38315 = pi08108 & ~w38311;
assign w38316 = ~pi02721 & w38311;
assign w38317 = ~w38315 & ~w38316;
assign w38318 = pi08109 & ~w17763;
assign w38319 = ~pi02714 & w17763;
assign w38320 = ~w38318 & ~w38319;
assign w38321 = pi08110 & ~w17763;
assign w38322 = ~pi02715 & w17763;
assign w38323 = ~w38321 & ~w38322;
assign w38324 = pi08111 & ~w38311;
assign w38325 = w17938 & w19797;
assign w38326 = ~w38324 & ~w38325;
assign w38327 = pi08112 & ~w17763;
assign w38328 = ~pi02717 & w17763;
assign w38329 = ~w38327 & ~w38328;
assign w38330 = pi08113 & ~w17536;
assign w38331 = w17535 & w17603;
assign w38332 = ~w38330 & ~w38331;
assign w38333 = pi08114 & ~w38311;
assign w38334 = ~pi02718 & w38311;
assign w38335 = ~w38333 & ~w38334;
assign w38336 = pi08115 & ~w17536;
assign w38337 = w17535 & w20209;
assign w38338 = ~w38336 & ~w38337;
assign w38339 = pi08116 & ~w38311;
assign w38340 = ~pi02167 & w38311;
assign w38341 = ~w38339 & ~w38340;
assign w38342 = pi08117 & ~w17536;
assign w38343 = ~pi02713 & w17536;
assign w38344 = ~w38342 & ~w38343;
assign w38345 = pi08118 & ~w17536;
assign w38346 = ~pi02715 & w17536;
assign w38347 = ~w38345 & ~w38346;
assign w38348 = pi08119 & ~w17536;
assign w38349 = ~pi02716 & w17536;
assign w38350 = ~w38348 & ~w38349;
assign w38351 = pi08120 & ~w38311;
assign w38352 = w17938 & w19312;
assign w38353 = ~w38351 & ~w38352;
assign w38354 = pi08121 & ~w17536;
assign w38355 = ~pi02717 & w17536;
assign w38356 = ~w38354 & ~w38355;
assign w38357 = pi08122 & ~w38311;
assign w38358 = ~pi02164 & w38311;
assign w38359 = ~w38357 & ~w38358;
assign w38360 = pi08123 & ~w17012;
assign w38361 = ~pi02703 & w17012;
assign w38362 = ~w38360 & ~w38361;
assign w38363 = pi08124 & ~w38311;
assign w38364 = w17594 & w17938;
assign w38365 = ~w38363 & ~w38364;
assign w38366 = pi08125 & ~w17012;
assign w38367 = ~pi02721 & w17012;
assign w38368 = ~w38366 & ~w38367;
assign w38369 = pi08126 & ~w17362;
assign w38370 = ~pi02711 & w17362;
assign w38371 = ~w38369 & ~w38370;
assign w38372 = pi08127 & ~w17012;
assign w38373 = ~pi02718 & w17012;
assign w38374 = ~w38372 & ~w38373;
assign w38375 = pi08128 & ~w17362;
assign w38376 = ~pi02170 & w17362;
assign w38377 = ~w38375 & ~w38376;
assign w38378 = pi08129 & ~w17012;
assign w38379 = ~pi02164 & w17012;
assign w38380 = ~w38378 & ~w38379;
assign w38381 = pi08130 & ~w17362;
assign w38382 = ~pi02713 & w17362;
assign w38383 = ~w38381 & ~w38382;
assign w38384 = pi08131 & ~w17362;
assign w38385 = ~pi02715 & w17362;
assign w38386 = ~w38384 & ~w38385;
assign w38387 = pi08132 & ~w17362;
assign w38388 = ~pi02716 & w17362;
assign w38389 = ~w38387 & ~w38388;
assign w38390 = pi08133 & ~w17012;
assign w38391 = ~pi02167 & w17012;
assign w38392 = ~w38390 & ~w38391;
assign w38393 = pi08134 & ~w17012;
assign w38394 = ~pi02722 & w17012;
assign w38395 = ~w38393 & ~w38394;
assign w38396 = pi08135 & ~w17362;
assign w38397 = ~pi02717 & w17362;
assign w38398 = ~w38396 & ~w38397;
assign w38399 = pi08136 & ~w17012;
assign w38400 = w17011 & w17594;
assign w38401 = ~w38399 & ~w38400;
assign w38402 = pi08137 & ~w17109;
assign w38403 = ~pi02703 & w17109;
assign w38404 = ~w38402 & ~w38403;
assign w38405 = pi08138 & ~w17109;
assign w38406 = ~pi02169 & w17109;
assign w38407 = ~w38405 & ~w38406;
assign w38408 = pi08139 & ~w17109;
assign w38409 = ~pi02718 & w17109;
assign w38410 = ~w38408 & ~w38409;
assign w38411 = pi08140 & ~w17109;
assign w38412 = ~pi02167 & w17109;
assign w38413 = ~w38411 & ~w38412;
assign w38414 = pi08141 & ~w17109;
assign w38415 = ~pi02722 & w17109;
assign w38416 = ~w38414 & ~w38415;
assign w38417 = pi08142 & ~w17109;
assign w38418 = ~pi02719 & w17109;
assign w38419 = ~w38417 & ~w38418;
assign w38420 = ~w16992 & w17098;
assign w38421 = pi08143 & ~w38420;
assign w38422 = ~pi02703 & w38420;
assign w38423 = ~w38421 & ~w38422;
assign w38424 = pi08144 & ~w36450;
assign w38425 = ~pi02711 & w36450;
assign w38426 = ~w38424 & ~w38425;
assign w38427 = pi08145 & ~w38420;
assign w38428 = w17098 & w17811;
assign w38429 = ~w38427 & ~w38428;
assign w38430 = pi08146 & ~w38420;
assign w38431 = ~pi02169 & w38420;
assign w38432 = ~w38430 & ~w38431;
assign w38433 = pi08147 & ~w38420;
assign w38434 = w17098 & w17586;
assign w38435 = ~w38433 & ~w38434;
assign w38436 = pi08148 & ~w38420;
assign w38437 = ~pi02167 & w38420;
assign w38438 = ~w38436 & ~w38437;
assign w38439 = pi08149 & ~w38420;
assign w38440 = ~pi02164 & w38420;
assign w38441 = ~w38439 & ~w38440;
assign w38442 = pi08150 & ~w38420;
assign w38443 = ~pi02722 & w38420;
assign w38444 = ~w38442 & ~w38443;
assign w38445 = pi08151 & ~w38420;
assign w38446 = w17098 & w17594;
assign w38447 = ~w38445 & ~w38446;
assign w38448 = ~w16992 & w20244;
assign w38449 = pi08152 & ~w38448;
assign w38450 = w17811 & w20244;
assign w38451 = ~w38449 & ~w38450;
assign w38452 = pi08153 & ~w38448;
assign w38453 = ~pi02169 & w38448;
assign w38454 = ~w38452 & ~w38453;
assign w38455 = pi08154 & ~w38448;
assign w38456 = ~pi02718 & w38448;
assign w38457 = ~w38455 & ~w38456;
assign w38458 = pi08155 & ~w38448;
assign w38459 = ~pi02164 & w38448;
assign w38460 = ~w38458 & ~w38459;
assign w38461 = pi08156 & ~w38448;
assign w38462 = ~pi02722 & w38448;
assign w38463 = ~w38461 & ~w38462;
assign w38464 = pi08157 & ~w38448;
assign w38465 = ~pi02719 & w38448;
assign w38466 = ~w38464 & ~w38465;
assign w38467 = ~w16992 & w18542;
assign w38468 = pi08158 & ~w38467;
assign w38469 = ~pi02721 & w38467;
assign w38470 = ~w38468 & ~w38469;
assign w38471 = pi08159 & ~w38467;
assign w38472 = ~pi02169 & w38467;
assign w38473 = ~w38471 & ~w38472;
assign w38474 = pi08160 & ~w38467;
assign w38475 = ~pi02718 & w38467;
assign w38476 = ~w38474 & ~w38475;
assign w38477 = pi08161 & ~w38467;
assign w38478 = w18542 & w19273;
assign w38479 = ~w38477 & ~w38478;
assign w38480 = pi08162 & ~w38467;
assign w38481 = ~pi02164 & w38467;
assign w38482 = ~w38480 & ~w38481;
assign w38483 = pi08163 & ~w38467;
assign w38484 = ~pi02722 & w38467;
assign w38485 = ~w38483 & ~w38484;
assign w38486 = pi08164 & ~w38467;
assign w38487 = ~pi02719 & w38467;
assign w38488 = ~w38486 & ~w38487;
assign w38489 = pi08165 & ~w26635;
assign w38490 = w17811 & w18662;
assign w38491 = ~w38489 & ~w38490;
assign w38492 = pi08166 & ~w26635;
assign w38493 = w18662 & w19797;
assign w38494 = ~w38492 & ~w38493;
assign w38495 = pi08167 & ~w26635;
assign w38496 = w17586 & w18662;
assign w38497 = ~w38495 & ~w38496;
assign w38498 = pi08168 & ~w26635;
assign w38499 = w17620 & w18662;
assign w38500 = ~w38498 & ~w38499;
assign w38501 = pi08169 & ~w26635;
assign w38502 = w18662 & w19312;
assign w38503 = ~w38501 & ~w38502;
assign w38504 = pi08170 & ~w26635;
assign w38505 = w17594 & w18662;
assign w38506 = ~w38504 & ~w38505;
assign w38507 = pi08171 & ~w23447;
assign w38508 = ~pi02721 & w23447;
assign w38509 = ~w38507 & ~w38508;
assign w38510 = pi08172 & ~w23447;
assign w38511 = ~pi02169 & w23447;
assign w38512 = ~w38510 & ~w38511;
assign w38513 = pi08173 & ~w23447;
assign w38514 = ~pi02718 & w23447;
assign w38515 = ~w38513 & ~w38514;
assign w38516 = pi08174 & ~w23447;
assign w38517 = ~pi02167 & w23447;
assign w38518 = ~w38516 & ~w38517;
assign w38519 = pi08175 & ~w23447;
assign w38520 = ~pi02164 & w23447;
assign w38521 = ~w38519 & ~w38520;
assign w38522 = pi08176 & ~w23447;
assign w38523 = ~pi02722 & w23447;
assign w38524 = ~w38522 & ~w38523;
assign w38525 = pi08177 & ~w23447;
assign w38526 = ~pi02719 & w23447;
assign w38527 = ~w38525 & ~w38526;
assign w38528 = pi08178 & ~w21517;
assign w38529 = ~pi02721 & w21517;
assign w38530 = ~w38528 & ~w38529;
assign w38531 = pi08179 & ~w21517;
assign w38532 = ~pi02169 & w21517;
assign w38533 = ~w38531 & ~w38532;
assign w38534 = pi08180 & ~w21517;
assign w38535 = ~pi02718 & w21517;
assign w38536 = ~w38534 & ~w38535;
assign w38537 = pi08181 & ~w21517;
assign w38538 = w17620 & w18554;
assign w38539 = ~w38537 & ~w38538;
assign w38540 = pi08182 & ~w21517;
assign w38541 = w18554 & w19312;
assign w38542 = ~w38540 & ~w38541;
assign w38543 = pi08183 & ~w21517;
assign w38544 = ~pi02719 & w21517;
assign w38545 = ~w38543 & ~w38544;
assign w38546 = pi08184 & ~w21484;
assign w38547 = ~pi02721 & w21484;
assign w38548 = ~w38546 & ~w38547;
assign w38549 = pi08185 & ~w21484;
assign w38550 = ~pi02169 & w21484;
assign w38551 = ~w38549 & ~w38550;
assign w38552 = pi08186 & ~w21484;
assign w38553 = ~pi02718 & w21484;
assign w38554 = ~w38552 & ~w38553;
assign w38555 = pi08187 & ~w21484;
assign w38556 = ~pi02167 & w21484;
assign w38557 = ~w38555 & ~w38556;
assign w38558 = pi08188 & ~w21484;
assign w38559 = ~pi02164 & w21484;
assign w38560 = ~w38558 & ~w38559;
assign w38561 = pi08189 & ~w21484;
assign w38562 = ~pi02722 & w21484;
assign w38563 = ~w38561 & ~w38562;
assign w38564 = pi08190 & ~w21484;
assign w38565 = ~pi02719 & w21484;
assign w38566 = ~w38564 & ~w38565;
assign w38567 = pi08191 & ~w20906;
assign w38568 = ~pi02721 & w20906;
assign w38569 = ~w38567 & ~w38568;
assign w38570 = pi08192 & ~w20906;
assign w38571 = ~pi02169 & w20906;
assign w38572 = ~w38570 & ~w38571;
assign w38573 = pi08193 & ~w20906;
assign w38574 = w17586 & w18454;
assign w38575 = ~w38573 & ~w38574;
assign w38576 = pi08194 & ~w20906;
assign w38577 = ~pi02164 & w20906;
assign w38578 = ~w38576 & ~w38577;
assign w38579 = pi08195 & ~w20906;
assign w38580 = ~pi02722 & w20906;
assign w38581 = ~w38579 & ~w38580;
assign w38582 = pi08196 & ~w20906;
assign w38583 = w17594 & w18454;
assign w38584 = ~w38582 & ~w38583;
assign w38585 = pi08197 & ~w20856;
assign w38586 = ~pi02721 & w20856;
assign w38587 = ~w38585 & ~w38586;
assign w38588 = pi08198 & ~w20856;
assign w38589 = w17710 & w19797;
assign w38590 = ~w38588 & ~w38589;
assign w38591 = pi08199 & ~w20856;
assign w38592 = ~pi02718 & w20856;
assign w38593 = ~w38591 & ~w38592;
assign w38594 = pi08200 & ~w20856;
assign w38595 = ~pi02167 & w20856;
assign w38596 = ~w38594 & ~w38595;
assign w38597 = pi08201 & ~w20856;
assign w38598 = ~pi02164 & w20856;
assign w38599 = ~w38597 & ~w38598;
assign w38600 = pi08202 & ~w20856;
assign w38601 = ~pi02722 & w20856;
assign w38602 = ~w38600 & ~w38601;
assign w38603 = pi08203 & ~w20856;
assign w38604 = ~pi02719 & w20856;
assign w38605 = ~w38603 & ~w38604;
assign w38606 = pi08204 & ~w20839;
assign w38607 = ~pi02721 & w20839;
assign w38608 = ~w38606 & ~w38607;
assign w38609 = pi08205 & ~w20839;
assign w38610 = ~pi02169 & w20839;
assign w38611 = ~w38609 & ~w38610;
assign w38612 = pi08206 & ~w20839;
assign w38613 = ~pi02718 & w20839;
assign w38614 = ~w38612 & ~w38613;
assign w38615 = pi08207 & ~w20839;
assign w38616 = w17620 & w18468;
assign w38617 = ~w38615 & ~w38616;
assign w38618 = pi08208 & ~w20839;
assign w38619 = ~pi02722 & w20839;
assign w38620 = ~w38618 & ~w38619;
assign w38621 = pi08209 & ~w20839;
assign w38622 = ~pi02719 & w20839;
assign w38623 = ~w38621 & ~w38622;
assign w38624 = pi08210 & ~w20780;
assign w38625 = ~pi02721 & w20780;
assign w38626 = ~w38624 & ~w38625;
assign w38627 = pi08211 & ~w20780;
assign w38628 = ~pi02169 & w20780;
assign w38629 = ~w38627 & ~w38628;
assign w38630 = pi08212 & ~w20780;
assign w38631 = ~pi02718 & w20780;
assign w38632 = ~w38630 & ~w38631;
assign w38633 = pi08213 & ~w20780;
assign w38634 = ~pi02167 & w20780;
assign w38635 = ~w38633 & ~w38634;
assign w38636 = pi08214 & ~w20780;
assign w38637 = ~pi02164 & w20780;
assign w38638 = ~w38636 & ~w38637;
assign w38639 = pi08215 & ~w20780;
assign w38640 = ~pi02722 & w20780;
assign w38641 = ~w38639 & ~w38640;
assign w38642 = pi08216 & ~w20780;
assign w38643 = ~pi02719 & w20780;
assign w38644 = ~w38642 & ~w38643;
assign w38645 = pi08217 & ~w20461;
assign w38646 = ~pi02169 & w20461;
assign w38647 = ~w38645 & ~w38646;
assign w38648 = pi08218 & ~w20461;
assign w38649 = ~pi02721 & w20461;
assign w38650 = ~w38648 & ~w38649;
assign w38651 = pi08219 & ~w20461;
assign w38652 = ~pi02718 & w20461;
assign w38653 = ~w38651 & ~w38652;
assign w38654 = pi08220 & ~w20461;
assign w38655 = ~pi02164 & w20461;
assign w38656 = ~w38654 & ~w38655;
assign w38657 = pi08221 & ~w20461;
assign w38658 = ~pi02722 & w20461;
assign w38659 = ~w38657 & ~w38658;
assign w38660 = pi08222 & ~w20461;
assign w38661 = ~pi02719 & w20461;
assign w38662 = ~w38660 & ~w38661;
assign w38663 = pi08223 & ~w19665;
assign w38664 = w17416 & w17811;
assign w38665 = ~w38663 & ~w38664;
assign w38666 = pi08224 & ~w19665;
assign w38667 = ~pi02169 & w19665;
assign w38668 = ~w38666 & ~w38667;
assign w38669 = pi08225 & ~w19665;
assign w38670 = ~pi02718 & w19665;
assign w38671 = ~w38669 & ~w38670;
assign w38672 = pi08226 & ~w19665;
assign w38673 = w17416 & w19273;
assign w38674 = ~w38672 & ~w38673;
assign w38675 = pi08227 & ~w19665;
assign w38676 = ~pi02164 & w19665;
assign w38677 = ~w38675 & ~w38676;
assign w38678 = pi08228 & ~w19665;
assign w38679 = w17416 & w19312;
assign w38680 = ~w38678 & ~w38679;
assign w38681 = pi08229 & ~w19665;
assign w38682 = ~pi02719 & w19665;
assign w38683 = ~w38681 & ~w38682;
assign w38684 = pi08230 & ~w20162;
assign w38685 = ~pi02703 & w20162;
assign w38686 = ~w38684 & ~w38685;
assign w38687 = pi08231 & ~w20162;
assign w38688 = ~pi02721 & w20162;
assign w38689 = ~w38687 & ~w38688;
assign w38690 = pi08232 & ~w20162;
assign w38691 = w17314 & w19797;
assign w38692 = ~w38690 & ~w38691;
assign w38693 = pi08233 & ~w20162;
assign w38694 = ~pi02167 & w20162;
assign w38695 = ~w38693 & ~w38694;
assign w38696 = pi08234 & ~w20162;
assign w38697 = ~pi02164 & w20162;
assign w38698 = ~w38696 & ~w38697;
assign w38699 = pi08235 & ~w20162;
assign w38700 = ~pi02722 & w20162;
assign w38701 = ~w38699 & ~w38700;
assign w38702 = pi08236 & ~w19791;
assign w38703 = ~pi02703 & w19791;
assign w38704 = ~w38702 & ~w38703;
assign w38705 = pi08237 & ~w19791;
assign w38706 = ~pi02721 & w19791;
assign w38707 = ~w38705 & ~w38706;
assign w38708 = pi08238 & ~w19791;
assign w38709 = ~pi02169 & w19791;
assign w38710 = ~w38708 & ~w38709;
assign w38711 = pi08239 & ~w19791;
assign w38712 = ~pi02167 & w19791;
assign w38713 = ~w38711 & ~w38712;
assign w38714 = pi08240 & ~w19791;
assign w38715 = ~pi02718 & w19791;
assign w38716 = ~w38714 & ~w38715;
assign w38717 = pi08241 & ~w19791;
assign w38718 = ~pi02164 & w19791;
assign w38719 = ~w38717 & ~w38718;
assign w38720 = pi08242 & ~w19791;
assign w38721 = ~pi02722 & w19791;
assign w38722 = ~w38720 & ~w38721;
assign w38723 = pi08243 & ~w19476;
assign w38724 = ~pi02703 & w19476;
assign w38725 = ~w38723 & ~w38724;
assign w38726 = pi08244 & ~w19476;
assign w38727 = ~pi02721 & w19476;
assign w38728 = ~w38726 & ~w38727;
assign w38729 = pi08245 & ~w19476;
assign w38730 = ~pi02169 & w19476;
assign w38731 = ~w38729 & ~w38730;
assign w38732 = pi08246 & ~w19476;
assign w38733 = w17239 & w19273;
assign w38734 = ~w38732 & ~w38733;
assign w38735 = pi08247 & ~w19476;
assign w38736 = ~pi02164 & w19476;
assign w38737 = ~w38735 & ~w38736;
assign w38738 = pi08248 & ~w19476;
assign w38739 = ~pi02722 & w19476;
assign w38740 = ~w38738 & ~w38739;
assign w38741 = pi08249 & ~w19202;
assign w38742 = w17167 & w17532;
assign w38743 = ~w38741 & ~w38742;
assign w38744 = pi08250 & ~w19202;
assign w38745 = ~pi02721 & w19202;
assign w38746 = ~w38744 & ~w38745;
assign w38747 = pi08251 & ~w19202;
assign w38748 = ~pi02169 & w19202;
assign w38749 = ~w38747 & ~w38748;
assign w38750 = pi08252 & ~w19202;
assign w38751 = ~pi02718 & w19202;
assign w38752 = ~w38750 & ~w38751;
assign w38753 = pi08253 & ~w19202;
assign w38754 = ~pi02167 & w19202;
assign w38755 = ~w38753 & ~w38754;
assign w38756 = pi08254 & ~w19202;
assign w38757 = ~pi02164 & w19202;
assign w38758 = ~w38756 & ~w38757;
assign w38759 = pi08255 & ~w19202;
assign w38760 = ~pi02722 & w19202;
assign w38761 = ~w38759 & ~w38760;
assign w38762 = pi08256 & ~w17206;
assign w38763 = ~pi02703 & w17206;
assign w38764 = ~w38762 & ~w38763;
assign w38765 = pi08257 & ~w17206;
assign w38766 = ~pi02721 & w17206;
assign w38767 = ~w38765 & ~w38766;
assign w38768 = pi08258 & ~w17206;
assign w38769 = ~pi02169 & w17206;
assign w38770 = ~w38768 & ~w38769;
assign w38771 = pi08259 & ~w17206;
assign w38772 = ~pi02167 & w17206;
assign w38773 = ~w38771 & ~w38772;
assign w38774 = pi08260 & ~w17206;
assign w38775 = ~pi02164 & w17206;
assign w38776 = ~w38774 & ~w38775;
assign w38777 = pi08261 & ~w17206;
assign w38778 = ~pi02722 & w17206;
assign w38779 = ~w38777 & ~w38778;
assign w38780 = pi08262 & ~w17992;
assign w38781 = ~pi02703 & w17992;
assign w38782 = ~w38780 & ~w38781;
assign w38783 = pi08263 & ~w17992;
assign w38784 = ~pi02721 & w17992;
assign w38785 = ~w38783 & ~w38784;
assign w38786 = pi08264 & ~w17992;
assign w38787 = ~pi02169 & w17992;
assign w38788 = ~w38786 & ~w38787;
assign w38789 = pi08265 & ~w17992;
assign w38790 = ~pi02718 & w17992;
assign w38791 = ~w38789 & ~w38790;
assign w38792 = pi08266 & ~w17992;
assign w38793 = ~pi02167 & w17992;
assign w38794 = ~w38792 & ~w38793;
assign w38795 = pi08267 & ~w17992;
assign w38796 = ~pi02164 & w17992;
assign w38797 = ~w38795 & ~w38796;
assign w38798 = pi08268 & ~w17992;
assign w38799 = ~pi02722 & w17992;
assign w38800 = ~w38798 & ~w38799;
assign w38801 = pi08269 & ~w17790;
assign w38802 = ~pi02703 & w17790;
assign w38803 = ~w38801 & ~w38802;
assign w38804 = pi08270 & ~w17790;
assign w38805 = w17200 & w17811;
assign w38806 = ~w38804 & ~w38805;
assign w38807 = pi08271 & ~w17790;
assign w38808 = ~pi02169 & w17790;
assign w38809 = ~w38807 & ~w38808;
assign w38810 = pi08272 & ~w17790;
assign w38811 = ~pi02167 & w17790;
assign w38812 = ~w38810 & ~w38811;
assign w38813 = pi08273 & ~w17790;
assign w38814 = w17200 & w17620;
assign w38815 = ~w38813 & ~w38814;
assign w38816 = pi08274 & ~w17790;
assign w38817 = ~pi02722 & w17790;
assign w38818 = ~w38816 & ~w38817;
assign w38819 = pi08275 & ~w17873;
assign w38820 = ~pi02703 & w17873;
assign w38821 = ~w38819 & ~w38820;
assign w38822 = pi08276 & ~w17873;
assign w38823 = ~pi02721 & w17873;
assign w38824 = ~w38822 & ~w38823;
assign w38825 = pi08277 & ~w17873;
assign w38826 = ~pi02169 & w17873;
assign w38827 = ~w38825 & ~w38826;
assign w38828 = pi08278 & ~w17873;
assign w38829 = ~pi02718 & w17873;
assign w38830 = ~w38828 & ~w38829;
assign w38831 = pi08279 & ~w17873;
assign w38832 = ~pi02167 & w17873;
assign w38833 = ~w38831 & ~w38832;
assign w38834 = pi08280 & ~w17873;
assign w38835 = w17172 & w17620;
assign w38836 = ~w38834 & ~w38835;
assign w38837 = pi08281 & ~w17873;
assign w38838 = w17172 & w19312;
assign w38839 = ~w38837 & ~w38838;
assign w38840 = pi08282 & ~w17592;
assign w38841 = w17023 & w17532;
assign w38842 = ~w38840 & ~w38841;
assign w38843 = pi08283 & ~w17592;
assign w38844 = w17023 & w17811;
assign w38845 = ~w38843 & ~w38844;
assign w38846 = pi08284 & ~w17592;
assign w38847 = w17023 & w19797;
assign w38848 = ~w38846 & ~w38847;
assign w38849 = pi08285 & ~w17592;
assign w38850 = w17023 & w19273;
assign w38851 = ~w38849 & ~w38850;
assign w38852 = pi08286 & ~w17592;
assign w38853 = w17023 & w17620;
assign w38854 = ~w38852 & ~w38853;
assign w38855 = pi08287 & ~w17592;
assign w38856 = w17023 & w19312;
assign w38857 = ~w38855 & ~w38856;
assign w38858 = ~w16992 & w18740;
assign w38859 = pi08288 & ~w38858;
assign w38860 = w17532 & w18740;
assign w38861 = ~w38859 & ~w38860;
assign w38862 = pi08289 & ~w38858;
assign w38863 = w17811 & w18740;
assign w38864 = ~w38862 & ~w38863;
assign w38865 = pi08290 & ~w38858;
assign w38866 = w18740 & w19797;
assign w38867 = ~w38865 & ~w38866;
assign w38868 = pi08291 & ~w38858;
assign w38869 = w17586 & w18740;
assign w38870 = ~w38868 & ~w38869;
assign w38871 = pi08292 & ~w38858;
assign w38872 = w18740 & w19273;
assign w38873 = ~w38871 & ~w38872;
assign w38874 = pi08293 & ~w38858;
assign w38875 = w17620 & w18740;
assign w38876 = ~w38874 & ~w38875;
assign w38877 = pi08294 & ~w38858;
assign w38878 = w18740 & w19312;
assign w38879 = ~w38877 & ~w38878;
assign w38880 = pi08295 & ~w38858;
assign w38881 = w17594 & w18740;
assign w38882 = ~w38880 & ~w38881;
assign w38883 = pi08296 & ~w17480;
assign w38884 = w17479 & w17811;
assign w38885 = ~w38883 & ~w38884;
assign w38886 = pi08297 & ~w17480;
assign w38887 = ~pi02169 & w17480;
assign w38888 = ~w38886 & ~w38887;
assign w38889 = pi08298 & ~w17480;
assign w38890 = ~pi02167 & w17480;
assign w38891 = ~w38889 & ~w38890;
assign w38892 = pi08299 & ~w17480;
assign w38893 = ~pi02164 & w17480;
assign w38894 = ~w38892 & ~w38893;
assign w38895 = pi08300 & ~w17480;
assign w38896 = ~pi02722 & w17480;
assign w38897 = ~w38895 & ~w38896;
assign w38898 = pi08301 & ~w17399;
assign w38899 = ~pi02703 & w17399;
assign w38900 = ~w38898 & ~w38899;
assign w38901 = pi08302 & ~w17399;
assign w38902 = w17398 & w17811;
assign w38903 = ~w38901 & ~w38902;
assign w38904 = pi08303 & ~w17399;
assign w38905 = ~pi02169 & w17399;
assign w38906 = ~w38904 & ~w38905;
assign w38907 = pi08304 & ~w17399;
assign w38908 = ~pi02718 & w17399;
assign w38909 = ~w38907 & ~w38908;
assign w38910 = pi08305 & ~w17399;
assign w38911 = ~pi02167 & w17399;
assign w38912 = ~w38910 & ~w38911;
assign w38913 = pi08306 & ~w17399;
assign w38914 = ~pi02164 & w17399;
assign w38915 = ~w38913 & ~w38914;
assign w38916 = pi08307 & ~w17399;
assign w38917 = ~pi02719 & w17399;
assign w38918 = ~w38916 & ~w38917;
assign w38919 = pi08308 & ~w17115;
assign w38920 = ~pi02703 & w17115;
assign w38921 = ~w38919 & ~w38920;
assign w38922 = pi08309 & ~w17115;
assign w38923 = w17114 & w17811;
assign w38924 = ~w38922 & ~w38923;
assign w38925 = pi08310 & ~w17115;
assign w38926 = ~pi02169 & w17115;
assign w38927 = ~w38925 & ~w38926;
assign w38928 = pi08311 & ~w17115;
assign w38929 = ~pi02167 & w17115;
assign w38930 = ~w38928 & ~w38929;
assign w38931 = pi08312 & ~w17115;
assign w38932 = ~pi02164 & w17115;
assign w38933 = ~w38931 & ~w38932;
assign w38934 = pi08313 & ~w17115;
assign w38935 = ~pi02722 & w17115;
assign w38936 = ~w38934 & ~w38935;
assign w38937 = pi08314 & ~w17250;
assign w38938 = w17249 & w17532;
assign w38939 = ~w38937 & ~w38938;
assign w38940 = pi08315 & ~w17250;
assign w38941 = ~pi02721 & w17250;
assign w38942 = ~w38940 & ~w38941;
assign w38943 = pi08316 & ~w17250;
assign w38944 = w17249 & w19797;
assign w38945 = ~w38943 & ~w38944;
assign w38946 = pi08317 & ~w17250;
assign w38947 = ~pi02718 & w17250;
assign w38948 = ~w38946 & ~w38947;
assign w38949 = pi08318 & ~w17250;
assign w38950 = ~pi02167 & w17250;
assign w38951 = ~w38949 & ~w38950;
assign w38952 = pi08319 & ~w17250;
assign w38953 = ~pi02164 & w17250;
assign w38954 = ~w38952 & ~w38953;
assign w38955 = pi08320 & ~w17250;
assign w38956 = ~pi02722 & w17250;
assign w38957 = ~w38955 & ~w38956;
assign w38958 = pi08321 & ~w17196;
assign w38959 = ~pi02703 & w17196;
assign w38960 = ~w38958 & ~w38959;
assign w38961 = pi08322 & ~w17196;
assign w38962 = ~pi02721 & w17196;
assign w38963 = ~w38961 & ~w38962;
assign w38964 = pi08323 & ~w17196;
assign w38965 = ~pi02169 & w17196;
assign w38966 = ~w38964 & ~w38965;
assign w38967 = pi08324 & ~w17196;
assign w38968 = ~pi02167 & w17196;
assign w38969 = ~w38967 & ~w38968;
assign w38970 = pi08325 & ~w17196;
assign w38971 = w17047 & w17620;
assign w38972 = ~w38970 & ~w38971;
assign w38973 = pi08326 & ~w17196;
assign w38974 = ~pi02722 & w17196;
assign w38975 = ~w38973 & ~w38974;
assign w38976 = ~w16992 & w17490;
assign w38977 = pi08327 & ~w38976;
assign w38978 = ~pi02721 & w38976;
assign w38979 = ~w38977 & ~w38978;
assign w38980 = pi08328 & ~w38976;
assign w38981 = ~pi02703 & w38976;
assign w38982 = ~w38980 & ~w38981;
assign w38983 = pi08329 & ~w38976;
assign w38984 = ~pi02169 & w38976;
assign w38985 = ~w38983 & ~w38984;
assign w38986 = pi08330 & ~w38976;
assign w38987 = ~pi02718 & w38976;
assign w38988 = ~w38986 & ~w38987;
assign w38989 = pi08331 & ~w38976;
assign w38990 = ~pi02167 & w38976;
assign w38991 = ~w38989 & ~w38990;
assign w38992 = pi08332 & ~w38976;
assign w38993 = ~pi02164 & w38976;
assign w38994 = ~w38992 & ~w38993;
assign w38995 = pi08333 & ~w38976;
assign w38996 = ~pi02722 & w38976;
assign w38997 = ~w38995 & ~w38996;
assign w38998 = pi08334 & ~w25912;
assign w38999 = ~pi02703 & w25912;
assign w39000 = ~w38998 & ~w38999;
assign w39001 = pi08335 & ~w25912;
assign w39002 = w17811 & w18645;
assign w39003 = ~w39001 & ~w39002;
assign w39004 = pi08336 & ~w25912;
assign w39005 = ~pi02718 & w25912;
assign w39006 = ~w39004 & ~w39005;
assign w39007 = pi08337 & ~w25912;
assign w39008 = ~pi02167 & w25912;
assign w39009 = ~w39007 & ~w39008;
assign w39010 = pi08338 & ~w25912;
assign w39011 = ~pi02164 & w25912;
assign w39012 = ~w39010 & ~w39011;
assign w39013 = pi08339 & ~w25912;
assign w39014 = ~pi02722 & w25912;
assign w39015 = ~w39013 & ~w39014;
assign w39016 = pi08340 & ~w21330;
assign w39017 = w17500 & w17532;
assign w39018 = ~w39016 & ~w39017;
assign w39019 = pi08341 & ~w21330;
assign w39020 = ~pi02721 & w21330;
assign w39021 = ~w39019 & ~w39020;
assign w39022 = pi08342 & ~w21330;
assign w39023 = ~pi02169 & w21330;
assign w39024 = ~w39022 & ~w39023;
assign w39025 = pi08343 & ~w21330;
assign w39026 = ~pi02718 & w21330;
assign w39027 = ~w39025 & ~w39026;
assign w39028 = pi08344 & ~w21330;
assign w39029 = ~pi02167 & w21330;
assign w39030 = ~w39028 & ~w39029;
assign w39031 = pi08345 & ~w21330;
assign w39032 = ~pi02164 & w21330;
assign w39033 = ~w39031 & ~w39032;
assign w39034 = pi08346 & ~w21330;
assign w39035 = w17500 & w19312;
assign w39036 = ~w39034 & ~w39035;
assign w39037 = pi08347 & ~w21443;
assign w39038 = ~pi02703 & w21443;
assign w39039 = ~w39037 & ~w39038;
assign w39040 = pi08348 & ~w21443;
assign w39041 = ~pi02721 & w21443;
assign w39042 = ~w39040 & ~w39041;
assign w39043 = pi08349 & ~w21443;
assign w39044 = ~pi02718 & w21443;
assign w39045 = ~w39043 & ~w39044;
assign w39046 = pi08350 & ~w21443;
assign w39047 = ~pi02167 & w21443;
assign w39048 = ~w39046 & ~w39047;
assign w39049 = pi08351 & ~w21443;
assign w39050 = ~pi02164 & w21443;
assign w39051 = ~w39049 & ~w39050;
assign w39052 = pi08352 & ~w21443;
assign w39053 = ~pi02722 & w21443;
assign w39054 = ~w39052 & ~w39053;
assign w39055 = pi08353 & ~w21070;
assign w39056 = ~pi02721 & w21070;
assign w39057 = ~w39055 & ~w39056;
assign w39058 = pi08354 & ~w21360;
assign w39059 = ~pi02703 & w21360;
assign w39060 = ~w39058 & ~w39059;
assign w39061 = pi08355 & ~w21360;
assign w39062 = ~pi02721 & w21360;
assign w39063 = ~w39061 & ~w39062;
assign w39064 = pi08356 & ~w21360;
assign w39065 = ~pi02169 & w21360;
assign w39066 = ~w39064 & ~w39065;
assign w39067 = pi08357 & ~w21360;
assign w39068 = ~pi02718 & w21360;
assign w39069 = ~w39067 & ~w39068;
assign w39070 = pi08358 & ~w21360;
assign w39071 = w18370 & w19273;
assign w39072 = ~w39070 & ~w39071;
assign w39073 = pi08359 & ~w21360;
assign w39074 = ~pi02164 & w21360;
assign w39075 = ~w39073 & ~w39074;
assign w39076 = pi08360 & ~w21360;
assign w39077 = ~pi02722 & w21360;
assign w39078 = ~w39076 & ~w39077;
assign w39079 = pi08361 & ~w21345;
assign w39080 = ~pi02721 & w21345;
assign w39081 = ~w39079 & ~w39080;
assign w39082 = pi08362 & ~w21345;
assign w39083 = ~pi02703 & w21345;
assign w39084 = ~w39082 & ~w39083;
assign w39085 = pi08363 & ~w21345;
assign w39086 = w16999 & w19797;
assign w39087 = ~w39085 & ~w39086;
assign w39088 = pi08364 & ~w21345;
assign w39089 = ~pi02164 & w21345;
assign w39090 = ~w39088 & ~w39089;
assign w39091 = pi08365 & ~w21345;
assign w39092 = ~pi02722 & w21345;
assign w39093 = ~w39091 & ~w39092;
assign w39094 = pi08366 & ~w21345;
assign w39095 = ~pi02167 & w21345;
assign w39096 = ~w39094 & ~w39095;
assign w39097 = pi08367 & ~w21122;
assign w39098 = ~pi02703 & w21122;
assign w39099 = ~w39097 & ~w39098;
assign w39100 = pi08368 & ~w21122;
assign w39101 = ~pi02721 & w21122;
assign w39102 = ~w39100 & ~w39101;
assign w39103 = pi08369 & ~w21122;
assign w39104 = w17556 & w17586;
assign w39105 = ~w39103 & ~w39104;
assign w39106 = pi08370 & ~w21122;
assign w39107 = ~pi02169 & w21122;
assign w39108 = ~w39106 & ~w39107;
assign w39109 = pi08371 & ~w21122;
assign w39110 = w17556 & w19273;
assign w39111 = ~w39109 & ~w39110;
assign w39112 = pi08372 & ~w21122;
assign w39113 = ~pi02164 & w21122;
assign w39114 = ~w39112 & ~w39113;
assign w39115 = pi08373 & ~w21122;
assign w39116 = ~pi02722 & w21122;
assign w39117 = ~w39115 & ~w39116;
assign w39118 = pi08374 & ~w20867;
assign w39119 = w17811 & w17855;
assign w39120 = ~w39118 & ~w39119;
assign w39121 = pi08375 & ~w20867;
assign w39122 = w17532 & w17855;
assign w39123 = ~w39121 & ~w39122;
assign w39124 = pi08376 & ~w20867;
assign w39125 = ~pi02169 & w20867;
assign w39126 = ~w39124 & ~w39125;
assign w39127 = pi08377 & ~w20867;
assign w39128 = ~pi02164 & w20867;
assign w39129 = ~w39127 & ~w39128;
assign w39130 = pi08378 & ~w20867;
assign w39131 = ~pi02167 & w20867;
assign w39132 = ~w39130 & ~w39131;
assign w39133 = pi08379 & ~w20867;
assign w39134 = ~pi02722 & w20867;
assign w39135 = ~w39133 & ~w39134;
assign w39136 = pi08380 & ~w20825;
assign w39137 = ~pi02703 & w20825;
assign w39138 = ~w39136 & ~w39137;
assign w39139 = pi08381 & ~w20825;
assign w39140 = ~pi02721 & w20825;
assign w39141 = ~w39139 & ~w39140;
assign w39142 = pi08382 & ~w20825;
assign w39143 = ~pi02169 & w20825;
assign w39144 = ~w39142 & ~w39143;
assign w39145 = pi08383 & ~w20825;
assign w39146 = ~pi02718 & w20825;
assign w39147 = ~w39145 & ~w39146;
assign w39148 = pi08384 & ~w20825;
assign w39149 = w17461 & w19273;
assign w39150 = ~w39148 & ~w39149;
assign w39151 = pi08385 & ~w20825;
assign w39152 = ~pi02164 & w20825;
assign w39153 = ~w39151 & ~w39152;
assign w39154 = pi08386 & ~w20825;
assign w39155 = ~pi02722 & w20825;
assign w39156 = ~w39154 & ~w39155;
assign w39157 = pi08387 & ~w20835;
assign w39158 = ~pi02703 & w20835;
assign w39159 = ~w39157 & ~w39158;
assign w39160 = pi08388 & ~w20835;
assign w39161 = ~pi02721 & w20835;
assign w39162 = ~w39160 & ~w39161;
assign w39163 = pi08389 & ~w20835;
assign w39164 = ~pi02169 & w20835;
assign w39165 = ~w39163 & ~w39164;
assign w39166 = pi08390 & ~w20835;
assign w39167 = ~pi02167 & w20835;
assign w39168 = ~w39166 & ~w39167;
assign w39169 = pi08391 & ~w20835;
assign w39170 = ~pi02164 & w20835;
assign w39171 = ~w39169 & ~w39170;
assign w39172 = pi08392 & ~w20835;
assign w39173 = ~pi02722 & w20835;
assign w39174 = ~w39172 & ~w39173;
assign w39175 = pi08393 & ~w20843;
assign w39176 = ~pi02703 & w20843;
assign w39177 = ~w39175 & ~w39176;
assign w39178 = pi08394 & ~w20843;
assign w39179 = ~pi02721 & w20843;
assign w39180 = ~w39178 & ~w39179;
assign w39181 = pi08395 & ~w20843;
assign w39182 = ~pi02169 & w20843;
assign w39183 = ~w39181 & ~w39182;
assign w39184 = pi08396 & ~w20843;
assign w39185 = ~pi02167 & w20843;
assign w39186 = ~w39184 & ~w39185;
assign w39187 = pi08397 & ~w20843;
assign w39188 = ~pi02718 & w20843;
assign w39189 = ~w39187 & ~w39188;
assign w39190 = pi08398 & ~w20843;
assign w39191 = ~pi02164 & w20843;
assign w39192 = ~w39190 & ~w39191;
assign w39193 = pi08399 & ~w20843;
assign w39194 = ~pi02722 & w20843;
assign w39195 = ~w39193 & ~w39194;
assign w39196 = pi08400 & ~w20771;
assign w39197 = ~pi02703 & w20771;
assign w39198 = ~w39196 & ~w39197;
assign w39199 = pi08401 & ~w20771;
assign w39200 = ~pi02721 & w20771;
assign w39201 = ~w39199 & ~w39200;
assign w39202 = pi08402 & ~w20771;
assign w39203 = ~pi02169 & w20771;
assign w39204 = ~w39202 & ~w39203;
assign w39205 = pi08403 & ~w20771;
assign w39206 = ~pi02167 & w20771;
assign w39207 = ~w39205 & ~w39206;
assign w39208 = pi08404 & ~w20771;
assign w39209 = ~pi02164 & w20771;
assign w39210 = ~w39208 & ~w39209;
assign w39211 = pi08405 & ~w20771;
assign w39212 = ~pi02722 & w20771;
assign w39213 = ~w39211 & ~w39212;
assign w39214 = pi08406 & ~w19634;
assign w39215 = ~pi02703 & w19634;
assign w39216 = ~w39214 & ~w39215;
assign w39217 = pi08407 & ~w19634;
assign w39218 = ~pi02721 & w19634;
assign w39219 = ~w39217 & ~w39218;
assign w39220 = pi08408 & ~w19634;
assign w39221 = ~pi02169 & w19634;
assign w39222 = ~w39220 & ~w39221;
assign w39223 = pi08409 & ~w19634;
assign w39224 = ~pi02167 & w19634;
assign w39225 = ~w39223 & ~w39224;
assign w39226 = pi08410 & ~w19634;
assign w39227 = ~pi02722 & w19634;
assign w39228 = ~w39226 & ~w39227;
assign w39229 = pi08411 & ~w19634;
assign w39230 = ~pi02718 & w19634;
assign w39231 = ~w39229 & ~w39230;
assign w39232 = pi08412 & ~w19634;
assign w39233 = ~pi02164 & w19634;
assign w39234 = ~w39232 & ~w39233;
assign w39235 = pi08413 & ~w19694;
assign w39236 = ~pi02703 & w19694;
assign w39237 = ~w39235 & ~w39236;
assign w39238 = pi08414 & ~w19694;
assign w39239 = ~pi02721 & w19694;
assign w39240 = ~w39238 & ~w39239;
assign w39241 = pi08415 & ~w19694;
assign w39242 = ~pi02169 & w19694;
assign w39243 = ~w39241 & ~w39242;
assign w39244 = pi08416 & ~w19694;
assign w39245 = ~pi02167 & w19694;
assign w39246 = ~w39244 & ~w39245;
assign w39247 = pi08417 & ~w19694;
assign w39248 = ~pi02164 & w19694;
assign w39249 = ~w39247 & ~w39248;
assign w39250 = pi08418 & ~w19694;
assign w39251 = w17762 & w19312;
assign w39252 = ~w39250 & ~w39251;
assign w39253 = pi08419 & ~w20166;
assign w39254 = ~pi02703 & w20166;
assign w39255 = ~w39253 & ~w39254;
assign w39256 = pi08420 & ~w20166;
assign w39257 = ~pi02721 & w20166;
assign w39258 = ~w39256 & ~w39257;
assign w39259 = pi08421 & ~w20166;
assign w39260 = ~pi02169 & w20166;
assign w39261 = ~w39259 & ~w39260;
assign w39262 = pi08422 & ~w20166;
assign w39263 = ~pi02718 & w20166;
assign w39264 = ~w39262 & ~w39263;
assign w39265 = pi08423 & ~w20166;
assign w39266 = ~pi02167 & w20166;
assign w39267 = ~w39265 & ~w39266;
assign w39268 = pi08424 & ~w20166;
assign w39269 = ~pi02164 & w20166;
assign w39270 = ~w39268 & ~w39269;
assign w39271 = pi08425 & ~w20166;
assign w39272 = ~pi02722 & w20166;
assign w39273 = ~w39271 & ~w39272;
assign w39274 = pi08426 & ~w19145;
assign w39275 = ~pi02721 & w19145;
assign w39276 = ~w39274 & ~w39275;
assign w39277 = pi08427 & ~w19145;
assign w39278 = w17361 & w17532;
assign w39279 = ~w39277 & ~w39278;
assign w39280 = pi08428 & ~w19145;
assign w39281 = ~pi02169 & w19145;
assign w39282 = ~w39280 & ~w39281;
assign w39283 = pi08429 & ~w19145;
assign w39284 = w17361 & w19273;
assign w39285 = ~w39283 & ~w39284;
assign w39286 = pi08430 & ~w19145;
assign w39287 = w17361 & w17620;
assign w39288 = ~w39286 & ~w39287;
assign w39289 = pi08431 & ~w19145;
assign w39290 = w17361 & w19312;
assign w39291 = ~w39289 & ~w39290;
assign w39292 = pi08432 & ~w19380;
assign w39293 = ~pi09961 & w19380;
assign w39294 = ~w39292 & ~w39293;
assign w39295 = pi08433 & ~w19380;
assign w39296 = ~pi09848 & w19380;
assign w39297 = ~w39295 & ~w39296;
assign w39298 = pi08434 & ~w19380;
assign w39299 = ~pi09812 & w19380;
assign w39300 = ~w39298 & ~w39299;
assign w39301 = pi08435 & ~w19380;
assign w39302 = ~pi02704 & w19380;
assign w39303 = ~w39301 & ~w39302;
assign w39304 = pi08436 & ~w19380;
assign w39305 = ~pi02178 & w19380;
assign w39306 = ~w39304 & ~w39305;
assign w39307 = pi08437 & ~w19380;
assign w39308 = w17128 & w19379;
assign w39309 = ~w39307 & ~w39308;
assign w39310 = pi08438 & ~w19380;
assign w39311 = ~pi09954 & w19380;
assign w39312 = ~w39310 & ~w39311;
assign w39313 = pi08439 & ~w18746;
assign w39314 = w18745 & w19365;
assign w39315 = ~w39313 & ~w39314;
assign w39316 = pi08440 & ~w18746;
assign w39317 = ~pi09848 & w18746;
assign w39318 = ~w39316 & ~w39317;
assign w39319 = pi08441 & ~w18746;
assign w39320 = ~pi09812 & w18746;
assign w39321 = ~w39319 & ~w39320;
assign w39322 = pi08442 & ~w18746;
assign w39323 = ~pi02704 & w18746;
assign w39324 = ~w39322 & ~w39323;
assign w39325 = pi08443 & ~w18746;
assign w39326 = ~pi09954 & w18746;
assign w39327 = ~w39325 & ~w39326;
assign w39328 = pi08444 & ~w18746;
assign w39329 = ~pi02720 & w18746;
assign w39330 = ~w39328 & ~w39329;
assign w39331 = pi08445 & ~w17978;
assign w39332 = ~pi09961 & w17978;
assign w39333 = ~w39331 & ~w39332;
assign w39334 = pi08446 & ~w17978;
assign w39335 = ~pi09848 & w17978;
assign w39336 = ~w39334 & ~w39335;
assign w39337 = pi08447 & ~w17978;
assign w39338 = ~pi09812 & w17978;
assign w39339 = ~w39337 & ~w39338;
assign w39340 = pi08448 & ~w17978;
assign w39341 = ~pi02704 & w17978;
assign w39342 = ~w39340 & ~w39341;
assign w39343 = pi08449 & ~w17978;
assign w39344 = ~pi02178 & w17978;
assign w39345 = ~w39343 & ~w39344;
assign w39346 = pi08450 & ~w17978;
assign w39347 = ~pi09954 & w17978;
assign w39348 = ~w39346 & ~w39347;
assign w39349 = pi08451 & ~w17978;
assign w39350 = ~pi02720 & w17978;
assign w39351 = ~w39349 & ~w39350;
assign w39352 = pi08452 & ~w18028;
assign w39353 = ~pi09961 & w18028;
assign w39354 = ~w39352 & ~w39353;
assign w39355 = pi08453 & ~w18028;
assign w39356 = w17186 & w18027;
assign w39357 = ~w39355 & ~w39356;
assign w39358 = pi08454 & ~w18028;
assign w39359 = ~pi09812 & w18028;
assign w39360 = ~w39358 & ~w39359;
assign w39361 = pi08455 & ~w18028;
assign w39362 = w17513 & w18027;
assign w39363 = ~w39361 & ~w39362;
assign w39364 = pi08456 & ~w18028;
assign w39365 = ~pi02720 & w18028;
assign w39366 = ~w39364 & ~w39365;
assign w39367 = pi08457 & ~w18028;
assign w39368 = ~pi02704 & w18028;
assign w39369 = ~w39367 & ~w39368;
assign w39370 = pi08458 & ~w31348;
assign w39371 = ~pi09961 & w31348;
assign w39372 = ~w39370 & ~w39371;
assign w39373 = pi08459 & ~w31348;
assign w39374 = ~pi09848 & w31348;
assign w39375 = ~w39373 & ~w39374;
assign w39376 = pi08460 & ~w31348;
assign w39377 = ~pi02704 & w31348;
assign w39378 = ~w39376 & ~w39377;
assign w39379 = pi08461 & ~w31348;
assign w39380 = ~pi02178 & w31348;
assign w39381 = ~w39379 & ~w39380;
assign w39382 = pi08462 & ~w31348;
assign w39383 = ~pi09954 & w31348;
assign w39384 = ~w39382 & ~w39383;
assign w39385 = pi08463 & ~w31348;
assign w39386 = ~pi02720 & w31348;
assign w39387 = ~w39385 & ~w39386;
assign w39388 = pi08464 & ~w31348;
assign w39389 = ~pi09962 & w31348;
assign w39390 = ~w39388 & ~w39389;
assign w39391 = pi08465 & ~w17232;
assign w39392 = ~pi09848 & w17232;
assign w39393 = ~w39391 & ~w39392;
assign w39394 = pi08466 & ~w17232;
assign w39395 = ~pi09812 & w17232;
assign w39396 = ~w39394 & ~w39395;
assign w39397 = pi08467 & ~w17232;
assign w39398 = ~pi02704 & w17232;
assign w39399 = ~w39397 & ~w39398;
assign w39400 = pi08468 & ~w17232;
assign w39401 = ~pi02720 & w17232;
assign w39402 = ~w39400 & ~w39401;
assign w39403 = pi08469 & ~w17232;
assign w39404 = ~pi09962 & w17232;
assign w39405 = ~w39403 & ~w39404;
assign w39406 = pi08470 & ~w17184;
assign w39407 = w17183 & w19365;
assign w39408 = ~w39406 & ~w39407;
assign w39409 = pi08471 & ~w17184;
assign w39410 = ~pi09812 & w17184;
assign w39411 = ~w39409 & ~w39410;
assign w39412 = pi08472 & ~w17184;
assign w39413 = ~pi02704 & w17184;
assign w39414 = ~w39412 & ~w39413;
assign w39415 = pi08473 & ~w17184;
assign w39416 = ~pi02178 & w17184;
assign w39417 = ~w39415 & ~w39416;
assign w39418 = pi08474 & ~w17184;
assign w39419 = ~pi09954 & w17184;
assign w39420 = ~w39418 & ~w39419;
assign w39421 = pi08475 & ~w17184;
assign w39422 = ~pi02720 & w17184;
assign w39423 = ~w39421 & ~w39422;
assign w39424 = pi08476 & ~w17184;
assign w39425 = w17183 & w17439;
assign w39426 = ~w39424 & ~w39425;
assign w39427 = pi08477 & ~w17386;
assign w39428 = ~pi09961 & w17386;
assign w39429 = ~w39427 & ~w39428;
assign w39430 = pi08478 & ~w17386;
assign w39431 = ~pi02704 & w17386;
assign w39432 = ~w39430 & ~w39431;
assign w39433 = pi08479 & ~w17386;
assign w39434 = ~pi09812 & w17386;
assign w39435 = ~w39433 & ~w39434;
assign w39436 = pi08480 & ~w17386;
assign w39437 = ~pi02178 & w17386;
assign w39438 = ~w39436 & ~w39437;
assign w39439 = pi08481 & ~w17386;
assign w39440 = ~pi02720 & w17386;
assign w39441 = ~w39439 & ~w39440;
assign w39442 = pi08482 & ~w17386;
assign w39443 = ~pi09962 & w17386;
assign w39444 = ~w39442 & ~w39443;
assign w39445 = pi08483 & ~w17350;
assign w39446 = ~pi09961 & w17350;
assign w39447 = ~w39445 & ~w39446;
assign w39448 = pi08484 & ~w17350;
assign w39449 = ~pi09812 & w17350;
assign w39450 = ~w39448 & ~w39449;
assign w39451 = pi08485 & ~w17350;
assign w39452 = ~pi02704 & w17350;
assign w39453 = ~w39451 & ~w39452;
assign w39454 = pi08486 & ~w17350;
assign w39455 = ~pi02178 & w17350;
assign w39456 = ~w39454 & ~w39455;
assign w39457 = pi08487 & ~w17350;
assign w39458 = ~pi09954 & w17350;
assign w39459 = ~w39457 & ~w39458;
assign w39460 = pi08488 & ~w17350;
assign w39461 = ~pi02720 & w17350;
assign w39462 = ~w39460 & ~w39461;
assign w39463 = pi08489 & ~w17350;
assign w39464 = ~pi09962 & w17350;
assign w39465 = ~w39463 & ~w39464;
assign w39466 = pi08490 & ~w17211;
assign w39467 = ~pi09961 & w17211;
assign w39468 = ~w39466 & ~w39467;
assign w39469 = pi08491 & ~w31676;
assign w39470 = ~pi09848 & w31676;
assign w39471 = ~w39469 & ~w39470;
assign w39472 = pi08492 & ~w17211;
assign w39473 = ~pi09848 & w17211;
assign w39474 = ~w39472 & ~w39473;
assign w39475 = pi08493 & ~w17211;
assign w39476 = ~pi09812 & w17211;
assign w39477 = ~w39475 & ~w39476;
assign w39478 = pi08494 & ~w17211;
assign w39479 = ~pi02178 & w17211;
assign w39480 = ~w39478 & ~w39479;
assign w39481 = pi08495 & ~w17211;
assign w39482 = ~pi09954 & w17211;
assign w39483 = ~w39481 & ~w39482;
assign w39484 = pi08496 & ~w17211;
assign w39485 = ~pi02720 & w17211;
assign w39486 = ~w39484 & ~w39485;
assign w39487 = pi08497 & ~w20090;
assign w39488 = w16941 & w19365;
assign w39489 = ~w39487 & ~w39488;
assign w39490 = pi08498 & ~w20090;
assign w39491 = w16941 & w17186;
assign w39492 = ~w39490 & ~w39491;
assign w39493 = pi08499 & ~w20090;
assign w39494 = w16941 & w17193;
assign w39495 = ~w39493 & ~w39494;
assign w39496 = pi08500 & ~w20090;
assign w39497 = ~pi02704 & w20090;
assign w39498 = ~w39496 & ~w39497;
assign w39499 = pi08501 & ~w20090;
assign w39500 = w16941 & w18861;
assign w39501 = ~w39499 & ~w39500;
assign w39502 = pi08502 & ~w20090;
assign w39503 = ~pi09954 & w20090;
assign w39504 = ~w39502 & ~w39503;
assign w39505 = pi08503 & ~w22053;
assign w39506 = ~pi02720 & w22053;
assign w39507 = ~w39505 & ~w39506;
assign w39508 = pi08504 & ~w31676;
assign w39509 = ~pi09961 & w31676;
assign w39510 = ~w39508 & ~w39509;
assign w39511 = pi08505 & ~w31676;
assign w39512 = ~pi09812 & w31676;
assign w39513 = ~w39511 & ~w39512;
assign w39514 = pi08506 & ~w31676;
assign w39515 = ~pi02704 & w31676;
assign w39516 = ~w39514 & ~w39515;
assign w39517 = pi08507 & ~w31676;
assign w39518 = ~pi09954 & w31676;
assign w39519 = ~w39517 & ~w39518;
assign w39520 = pi08508 & ~w31676;
assign w39521 = ~pi02720 & w31676;
assign w39522 = ~w39520 & ~w39521;
assign w39523 = pi08509 & ~w31676;
assign w39524 = ~pi09962 & w31676;
assign w39525 = ~w39523 & ~w39524;
assign w39526 = pi08510 & ~w24403;
assign w39527 = ~pi09848 & w24403;
assign w39528 = ~w39526 & ~w39527;
assign w39529 = pi08511 & ~w24403;
assign w39530 = ~pi09812 & w24403;
assign w39531 = ~w39529 & ~w39530;
assign w39532 = pi08512 & ~w24403;
assign w39533 = ~pi02704 & w24403;
assign w39534 = ~w39532 & ~w39533;
assign w39535 = pi08513 & ~w24403;
assign w39536 = ~pi02178 & w24403;
assign w39537 = ~w39535 & ~w39536;
assign w39538 = pi08514 & ~w24403;
assign w39539 = ~pi02720 & w24403;
assign w39540 = ~w39538 & ~w39539;
assign w39541 = pi08515 & ~w24403;
assign w39542 = ~pi09962 & w24403;
assign w39543 = ~w39541 & ~w39542;
assign w39544 = pi08516 & ~w24004;
assign w39545 = ~pi09961 & w24004;
assign w39546 = ~w39544 & ~w39545;
assign w39547 = pi08517 & ~w24004;
assign w39548 = ~pi09812 & w24004;
assign w39549 = ~w39547 & ~w39548;
assign w39550 = pi08518 & ~w24004;
assign w39551 = ~pi02704 & w24004;
assign w39552 = ~w39550 & ~w39551;
assign w39553 = pi08519 & ~w24004;
assign w39554 = w17837 & w18861;
assign w39555 = ~w39553 & ~w39554;
assign w39556 = pi08520 & ~w24004;
assign w39557 = ~pi02720 & w24004;
assign w39558 = ~w39556 & ~w39557;
assign w39559 = pi08521 & ~w24004;
assign w39560 = ~pi09962 & w24004;
assign w39561 = ~w39559 & ~w39560;
assign w39562 = pi08522 & ~w22053;
assign w39563 = ~pi09961 & w22053;
assign w39564 = ~w39562 & ~w39563;
assign w39565 = pi08523 & ~w22053;
assign w39566 = ~pi02704 & w22053;
assign w39567 = ~w39565 & ~w39566;
assign w39568 = pi08524 & ~w22053;
assign w39569 = w18861 & w20465;
assign w39570 = ~w39568 & ~w39569;
assign w39571 = pi08525 & ~w22053;
assign w39572 = ~pi09954 & w22053;
assign w39573 = ~w39571 & ~w39572;
assign w39574 = pi08526 & ~w22053;
assign w39575 = ~pi09962 & w22053;
assign w39576 = ~w39574 & ~w39575;
assign w39577 = pi08527 & ~w21488;
assign w39578 = ~pi09961 & w21488;
assign w39579 = ~w39577 & ~w39578;
assign w39580 = pi08528 & ~w21488;
assign w39581 = ~pi09848 & w21488;
assign w39582 = ~w39580 & ~w39581;
assign w39583 = pi08529 & ~w21488;
assign w39584 = w17814 & w18861;
assign w39585 = ~w39583 & ~w39584;
assign w39586 = pi08530 & ~w21488;
assign w39587 = w17128 & w17814;
assign w39588 = ~w39586 & ~w39587;
assign w39589 = pi08531 & ~w21488;
assign w39590 = ~pi09962 & w21488;
assign w39591 = ~w39589 & ~w39590;
assign w39592 = pi08532 & ~w21385;
assign w39593 = ~pi09848 & w21385;
assign w39594 = ~w39592 & ~w39593;
assign w39595 = pi08533 & ~w21385;
assign w39596 = ~pi09812 & w21385;
assign w39597 = ~w39595 & ~w39596;
assign w39598 = pi08534 & ~w21385;
assign w39599 = ~pi02704 & w21385;
assign w39600 = ~w39598 & ~w39599;
assign w39601 = pi08535 & ~w21385;
assign w39602 = w17513 & w17822;
assign w39603 = ~w39601 & ~w39602;
assign w39604 = pi08536 & ~w21385;
assign w39605 = w17439 & w17822;
assign w39606 = ~w39604 & ~w39605;
assign w39607 = pi08537 & ~w21367;
assign w39608 = ~pi09961 & w21367;
assign w39609 = ~w39607 & ~w39608;
assign w39610 = pi08538 & ~w21367;
assign w39611 = ~pi09848 & w21367;
assign w39612 = ~w39610 & ~w39611;
assign w39613 = pi08539 & ~w21367;
assign w39614 = ~pi02704 & w21367;
assign w39615 = ~w39613 & ~w39614;
assign w39616 = pi08540 & ~w21367;
assign w39617 = w17513 & w17775;
assign w39618 = ~w39616 & ~w39617;
assign w39619 = pi08541 & ~w22053;
assign w39620 = ~pi09848 & w22053;
assign w39621 = ~w39619 & ~w39620;
assign w39622 = pi08542 & ~w21367;
assign w39623 = ~pi02720 & w21367;
assign w39624 = ~w39622 & ~w39623;
assign w39625 = pi08543 & ~w21356;
assign w39626 = ~pi09961 & w21356;
assign w39627 = ~w39625 & ~w39626;
assign w39628 = pi08544 & ~w21356;
assign w39629 = ~pi09848 & w21356;
assign w39630 = ~w39628 & ~w39629;
assign w39631 = pi08545 & ~w21356;
assign w39632 = ~pi09812 & w21356;
assign w39633 = ~w39631 & ~w39632;
assign w39634 = pi08546 & ~w21356;
assign w39635 = ~pi09954 & w21356;
assign w39636 = ~w39634 & ~w39635;
assign w39637 = pi08547 & ~w21356;
assign w39638 = ~pi02720 & w21356;
assign w39639 = ~w39637 & ~w39638;
assign w39640 = pi08548 & ~w21356;
assign w39641 = ~pi09962 & w21356;
assign w39642 = ~w39640 & ~w39641;
assign w39643 = pi08549 & ~w18210;
assign w39644 = ~pi09812 & w18210;
assign w39645 = ~w39643 & ~w39644;
assign w39646 = pi08550 & ~w18210;
assign w39647 = w17028 & w17311;
assign w39648 = ~w39646 & ~w39647;
assign w39649 = pi08551 & ~w18210;
assign w39650 = ~pi09954 & w18210;
assign w39651 = ~w39649 & ~w39650;
assign w39652 = pi08552 & ~w18210;
assign w39653 = ~pi02720 & w18210;
assign w39654 = ~w39652 & ~w39653;
assign w39655 = pi08553 & ~w18210;
assign w39656 = w17028 & w17439;
assign w39657 = ~w39655 & ~w39656;
assign w39658 = pi08554 & ~w21270;
assign w39659 = ~pi09961 & w21270;
assign w39660 = ~w39658 & ~w39659;
assign w39661 = pi08555 & ~w21270;
assign w39662 = ~pi09848 & w21270;
assign w39663 = ~w39661 & ~w39662;
assign w39664 = pi08556 & ~w21270;
assign w39665 = ~pi02178 & w21270;
assign w39666 = ~w39664 & ~w39665;
assign w39667 = pi08557 & ~w21270;
assign w39668 = w17053 & w17513;
assign w39669 = ~w39667 & ~w39668;
assign w39670 = pi08558 & ~w21270;
assign w39671 = ~pi02720 & w21270;
assign w39672 = ~w39670 & ~w39671;
assign w39673 = pi08559 & ~w21266;
assign w39674 = ~pi09848 & w21266;
assign w39675 = ~w39673 & ~w39674;
assign w39676 = pi08560 & ~w21266;
assign w39677 = w17006 & w17193;
assign w39678 = ~w39676 & ~w39677;
assign w39679 = pi08561 & ~w21266;
assign w39680 = ~pi02704 & w21266;
assign w39681 = ~w39679 & ~w39680;
assign w39682 = pi08562 & ~w27595;
assign w39683 = ~pi02170 & w27595;
assign w39684 = ~w39682 & ~w39683;
assign w39685 = pi08563 & ~w36416;
assign w39686 = ~pi02713 & w36416;
assign w39687 = ~w39685 & ~w39686;
assign w39688 = pi08564 & ~w21266;
assign w39689 = ~pi09954 & w21266;
assign w39690 = ~w39688 & ~w39689;
assign w39691 = pi08565 & ~w21266;
assign w39692 = w17006 & w17128;
assign w39693 = ~w39691 & ~w39692;
assign w39694 = pi08566 & ~w21266;
assign w39695 = ~pi09962 & w21266;
assign w39696 = ~w39694 & ~w39695;
assign w39697 = pi08567 & ~w21202;
assign w39698 = ~pi09961 & w21202;
assign w39699 = ~w39697 & ~w39698;
assign w39700 = pi08568 & ~w21202;
assign w39701 = ~pi09848 & w21202;
assign w39702 = ~w39700 & ~w39701;
assign w39703 = pi08569 & ~w21202;
assign w39704 = ~pi02704 & w21202;
assign w39705 = ~w39703 & ~w39704;
assign w39706 = pi08570 & ~w21202;
assign w39707 = ~pi02178 & w21202;
assign w39708 = ~w39706 & ~w39707;
assign w39709 = pi08571 & ~w21177;
assign w39710 = ~pi09961 & w21177;
assign w39711 = ~w39709 & ~w39710;
assign w39712 = pi08572 & ~w21202;
assign w39713 = ~pi09962 & w21202;
assign w39714 = ~w39712 & ~w39713;
assign w39715 = pi08573 & ~w21177;
assign w39716 = ~pi09848 & w21177;
assign w39717 = ~w39715 & ~w39716;
assign w39718 = pi08574 & ~w21177;
assign w39719 = w17311 & w17406;
assign w39720 = ~w39718 & ~w39719;
assign w39721 = pi08575 & ~w21177;
assign w39722 = ~pi02178 & w21177;
assign w39723 = ~w39721 & ~w39722;
assign w39724 = pi08576 & ~w21177;
assign w39725 = ~pi02720 & w21177;
assign w39726 = ~w39724 & ~w39725;
assign w39727 = pi08577 & ~w21162;
assign w39728 = ~pi09848 & w21162;
assign w39729 = ~w39727 & ~w39728;
assign w39730 = pi08578 & ~w21162;
assign w39731 = ~pi09812 & w21162;
assign w39732 = ~w39730 & ~w39731;
assign w39733 = pi08579 & ~w21162;
assign w39734 = ~pi02704 & w21162;
assign w39735 = ~w39733 & ~w39734;
assign w39736 = pi08580 & ~w21162;
assign w39737 = ~pi02178 & w21162;
assign w39738 = ~w39736 & ~w39737;
assign w39739 = pi08581 & ~w21162;
assign w39740 = ~pi09954 & w21162;
assign w39741 = ~w39739 & ~w39740;
assign w39742 = pi08582 & ~w21162;
assign w39743 = ~pi09962 & w21162;
assign w39744 = ~w39742 & ~w39743;
assign w39745 = pi08583 & ~w21000;
assign w39746 = ~pi09961 & w21000;
assign w39747 = ~w39745 & ~w39746;
assign w39748 = pi08584 & ~w21000;
assign w39749 = ~pi09848 & w21000;
assign w39750 = ~w39748 & ~w39749;
assign w39751 = pi08585 & ~w21000;
assign w39752 = ~pi02178 & w21000;
assign w39753 = ~w39751 & ~w39752;
assign w39754 = pi08586 & ~w21000;
assign w39755 = ~pi09954 & w21000;
assign w39756 = ~w39754 & ~w39755;
assign w39757 = pi08587 & ~w21000;
assign w39758 = ~pi09962 & w21000;
assign w39759 = ~w39757 & ~w39758;
assign w39760 = pi08588 & ~w20974;
assign w39761 = ~pi09961 & w20974;
assign w39762 = ~w39760 & ~w39761;
assign w39763 = pi08589 & ~w20974;
assign w39764 = w17186 & w19596;
assign w39765 = ~w39763 & ~w39764;
assign w39766 = pi08590 & ~w20974;
assign w39767 = ~pi02704 & w20974;
assign w39768 = ~w39766 & ~w39767;
assign w39769 = pi08591 & ~w20974;
assign w39770 = w17513 & w19596;
assign w39771 = ~w39769 & ~w39770;
assign w39772 = pi08592 & ~w20974;
assign w39773 = w17128 & w19596;
assign w39774 = ~w39772 & ~w39773;
assign w39775 = pi08593 & ~w20974;
assign w39776 = w17439 & w19596;
assign w39777 = ~w39775 & ~w39776;
assign w39778 = pi08594 & ~w17280;
assign w39779 = ~pi09961 & w17280;
assign w39780 = ~w39778 & ~w39779;
assign w39781 = pi08595 & ~w17280;
assign w39782 = ~pi09848 & w17280;
assign w39783 = ~w39781 & ~w39782;
assign w39784 = pi08596 & ~w17280;
assign w39785 = ~pi09812 & w17280;
assign w39786 = ~w39784 & ~w39785;
assign w39787 = pi08597 & ~w17280;
assign w39788 = w17279 & w17513;
assign w39789 = ~w39787 & ~w39788;
assign w39790 = pi08598 & ~w17280;
assign w39791 = ~pi02720 & w17280;
assign w39792 = ~w39790 & ~w39791;
assign w39793 = pi08599 & ~w20739;
assign w39794 = ~pi09961 & w20739;
assign w39795 = ~w39793 & ~w39794;
assign w39796 = pi08600 & ~w20739;
assign w39797 = w17193 & w19282;
assign w39798 = ~w39796 & ~w39797;
assign w39799 = pi08601 & ~w20739;
assign w39800 = ~pi02704 & w20739;
assign w39801 = ~w39799 & ~w39800;
assign w39802 = pi08602 & ~w20739;
assign w39803 = ~pi02178 & w20739;
assign w39804 = ~w39802 & ~w39803;
assign w39805 = pi08603 & ~w20739;
assign w39806 = ~pi02720 & w20739;
assign w39807 = ~w39805 & ~w39806;
assign w39808 = pi08604 & ~w20739;
assign w39809 = ~pi09962 & w20739;
assign w39810 = ~w39808 & ~w39809;
assign w39811 = pi08605 & ~w18727;
assign w39812 = ~pi09961 & w18727;
assign w39813 = ~w39811 & ~w39812;
assign w39814 = pi08606 & ~w18727;
assign w39815 = ~pi09848 & w18727;
assign w39816 = ~w39814 & ~w39815;
assign w39817 = pi08607 & ~w18727;
assign w39818 = ~pi09812 & w18727;
assign w39819 = ~w39817 & ~w39818;
assign w39820 = pi08608 & ~w18727;
assign w39821 = w18726 & w18861;
assign w39822 = ~w39820 & ~w39821;
assign w39823 = pi08609 & ~w18727;
assign w39824 = ~pi09954 & w18727;
assign w39825 = ~w39823 & ~w39824;
assign w39826 = pi08610 & ~w18848;
assign w39827 = ~pi09961 & w18848;
assign w39828 = ~w39826 & ~w39827;
assign w39829 = pi08611 & ~w18848;
assign w39830 = ~pi09812 & w18848;
assign w39831 = ~w39829 & ~w39830;
assign w39832 = pi08612 & ~w18848;
assign w39833 = ~pi02704 & w18848;
assign w39834 = ~w39832 & ~w39833;
assign w39835 = pi08613 & ~w18848;
assign w39836 = ~pi09962 & w18848;
assign w39837 = ~w39835 & ~w39836;
assign w39838 = pi08614 & ~w18627;
assign w39839 = ~pi09961 & w18627;
assign w39840 = ~w39838 & ~w39839;
assign w39841 = pi08615 & ~w18627;
assign w39842 = ~pi09812 & w18627;
assign w39843 = ~w39841 & ~w39842;
assign w39844 = pi08616 & ~w18627;
assign w39845 = ~pi02178 & w18627;
assign w39846 = ~w39844 & ~w39845;
assign w39847 = pi08617 & ~w18627;
assign w39848 = ~pi09954 & w18627;
assign w39849 = ~w39847 & ~w39848;
assign w39850 = pi08618 & ~w18627;
assign w39851 = ~pi02720 & w18627;
assign w39852 = ~w39850 & ~w39851;
assign w39853 = pi08619 & ~w18627;
assign w39854 = ~pi09962 & w18627;
assign w39855 = ~w39853 & ~w39854;
assign w39856 = pi08620 & ~w18809;
assign w39857 = ~pi09961 & w18809;
assign w39858 = ~w39856 & ~w39857;
assign w39859 = pi08621 & ~w18809;
assign w39860 = w17186 & w18808;
assign w39861 = ~w39859 & ~w39860;
assign w39862 = pi08622 & ~w18809;
assign w39863 = w17193 & w18808;
assign w39864 = ~w39862 & ~w39863;
assign w39865 = pi08623 & ~w18809;
assign w39866 = ~pi02704 & w18809;
assign w39867 = ~w39865 & ~w39866;
assign w39868 = pi08624 & ~w18809;
assign w39869 = w17513 & w18808;
assign w39870 = ~w39868 & ~w39869;
assign w39871 = pi08625 & ~w18809;
assign w39872 = ~pi02720 & w18809;
assign w39873 = ~w39871 & ~w39872;
assign w39874 = pi08626 & ~w18718;
assign w39875 = ~pi09961 & w18718;
assign w39876 = ~w39874 & ~w39875;
assign w39877 = pi08627 & ~w18718;
assign w39878 = w17186 & w18186;
assign w39879 = ~w39877 & ~w39878;
assign w39880 = pi08628 & ~w18718;
assign w39881 = ~pi09812 & w18718;
assign w39882 = ~w39880 & ~w39881;
assign w39883 = pi08629 & ~w18718;
assign w39884 = ~pi02178 & w18718;
assign w39885 = ~w39883 & ~w39884;
assign w39886 = pi08630 & ~w18718;
assign w39887 = w17513 & w18186;
assign w39888 = ~w39886 & ~w39887;
assign w39889 = pi08631 & ~w18718;
assign w39890 = ~pi02720 & w18718;
assign w39891 = ~w39889 & ~w39890;
assign w39892 = pi08632 & ~w18718;
assign w39893 = ~pi09962 & w18718;
assign w39894 = ~w39892 & ~w39893;
assign w39895 = pi08633 & ~w17085;
assign w39896 = w17084 & w19365;
assign w39897 = ~w39895 & ~w39896;
assign w39898 = pi08634 & ~w17085;
assign w39899 = ~pi09848 & w17085;
assign w39900 = ~w39898 & ~w39899;
assign w39901 = pi08635 & ~w17085;
assign w39902 = w17084 & w17193;
assign w39903 = ~w39901 & ~w39902;
assign w39904 = pi08636 & ~w17085;
assign w39905 = w17084 & w18861;
assign w39906 = ~w39904 & ~w39905;
assign w39907 = pi08637 & ~w17085;
assign w39908 = ~pi09954 & w17085;
assign w39909 = ~w39907 & ~w39908;
assign w39910 = pi08638 & ~w17085;
assign w39911 = ~pi02720 & w17085;
assign w39912 = ~w39910 & ~w39911;
assign w39913 = pi08639 & ~w18427;
assign w39914 = ~pi09961 & w18427;
assign w39915 = ~w39913 & ~w39914;
assign w39916 = pi08640 & ~w18427;
assign w39917 = ~pi09848 & w18427;
assign w39918 = ~w39916 & ~w39917;
assign w39919 = pi08641 & ~w18427;
assign w39920 = ~pi09812 & w18427;
assign w39921 = ~w39919 & ~w39920;
assign w39922 = pi08642 & ~w18427;
assign w39923 = ~pi02178 & w18427;
assign w39924 = ~w39922 & ~w39923;
assign w39925 = pi08643 & ~w18427;
assign w39926 = ~pi09954 & w18427;
assign w39927 = ~w39925 & ~w39926;
assign w39928 = pi08644 & ~w18427;
assign w39929 = ~pi02720 & w18427;
assign w39930 = ~w39928 & ~w39929;
assign w39931 = pi08645 & ~w18427;
assign w39932 = ~pi09962 & w18427;
assign w39933 = ~w39931 & ~w39932;
assign w39934 = pi08646 & ~w17988;
assign w39935 = w17808 & w19365;
assign w39936 = ~w39934 & ~w39935;
assign w39937 = pi08647 & ~w17988;
assign w39938 = ~pi09848 & w17988;
assign w39939 = ~w39937 & ~w39938;
assign w39940 = pi08648 & ~w17988;
assign w39941 = w17193 & w17808;
assign w39942 = ~w39940 & ~w39941;
assign w39943 = pi08649 & ~w17988;
assign w39944 = ~pi02178 & w17988;
assign w39945 = ~w39943 & ~w39944;
assign w39946 = pi08650 & ~w17988;
assign w39947 = w17513 & w17808;
assign w39948 = ~w39946 & ~w39947;
assign w39949 = pi08651 & ~w17988;
assign w39950 = ~pi02720 & w17988;
assign w39951 = ~w39949 & ~w39950;
assign w39952 = pi08652 & ~w17896;
assign w39953 = w17390 & w19365;
assign w39954 = ~w39952 & ~w39953;
assign w39955 = pi08653 & ~w17896;
assign w39956 = ~pi09848 & w17896;
assign w39957 = ~w39955 & ~w39956;
assign w39958 = pi08654 & ~w17896;
assign w39959 = w17193 & w17390;
assign w39960 = ~w39958 & ~w39959;
assign w39961 = pi08655 & ~w17896;
assign w39962 = ~pi02178 & w17896;
assign w39963 = ~w39961 & ~w39962;
assign w39964 = pi08656 & ~w17896;
assign w39965 = w17390 & w17513;
assign w39966 = ~w39964 & ~w39965;
assign w39967 = pi08657 & ~w17896;
assign w39968 = w17128 & w17390;
assign w39969 = ~w39967 & ~w39968;
assign w39970 = pi08658 & ~w17896;
assign w39971 = ~pi09962 & w17896;
assign w39972 = ~w39970 & ~w39971;
assign w39973 = pi08659 & ~w17496;
assign w39974 = ~pi09961 & w17496;
assign w39975 = ~w39973 & ~w39974;
assign w39976 = pi08660 & ~w17496;
assign w39977 = ~pi09848 & w17496;
assign w39978 = ~w39976 & ~w39977;
assign w39979 = pi08661 & ~w17496;
assign w39980 = ~pi09812 & w17496;
assign w39981 = ~w39979 & ~w39980;
assign w39982 = pi08662 & ~w17496;
assign w39983 = ~pi02178 & w17496;
assign w39984 = ~w39982 & ~w39983;
assign w39985 = pi08663 & ~w17496;
assign w39986 = ~pi09954 & w17496;
assign w39987 = ~w39985 & ~w39986;
assign w39988 = pi08664 & ~w17496;
assign w39989 = ~pi09962 & w17496;
assign w39990 = ~w39988 & ~w39989;
assign w39991 = pi08665 & ~w17451;
assign w39992 = w17450 & w19365;
assign w39993 = ~w39991 & ~w39992;
assign w39994 = pi08666 & ~w17451;
assign w39995 = ~pi09848 & w17451;
assign w39996 = ~w39994 & ~w39995;
assign w39997 = pi08667 & ~w17451;
assign w39998 = ~pi09812 & w17451;
assign w39999 = ~w39997 & ~w39998;
assign w40000 = pi08668 & ~w17451;
assign w40001 = ~pi02178 & w17451;
assign w40002 = ~w40000 & ~w40001;
assign w40003 = pi08669 & ~w17451;
assign w40004 = ~pi09954 & w17451;
assign w40005 = ~w40003 & ~w40004;
assign w40006 = pi08670 & ~w17451;
assign w40007 = ~pi02720 & w17451;
assign w40008 = ~w40006 & ~w40007;
assign w40009 = pi08671 & ~w17451;
assign w40010 = ~pi09962 & w17451;
assign w40011 = ~w40009 & ~w40010;
assign w40012 = pi08672 & ~w17437;
assign w40013 = w17436 & w19365;
assign w40014 = ~w40012 & ~w40013;
assign w40015 = pi08673 & ~w17437;
assign w40016 = ~pi09848 & w17437;
assign w40017 = ~w40015 & ~w40016;
assign w40018 = pi08674 & ~w17437;
assign w40019 = ~pi09812 & w17437;
assign w40020 = ~w40018 & ~w40019;
assign w40021 = pi08675 & ~w17437;
assign w40022 = w17436 & w18861;
assign w40023 = ~w40021 & ~w40022;
assign w40024 = pi08676 & ~w17437;
assign w40025 = ~pi09954 & w17437;
assign w40026 = ~w40024 & ~w40025;
assign w40027 = pi08677 & ~w17437;
assign w40028 = ~pi02720 & w17437;
assign w40029 = ~w40027 & ~w40028;
assign w40030 = pi08678 & ~w17354;
assign w40031 = ~pi09961 & w17354;
assign w40032 = ~w40030 & ~w40031;
assign w40033 = pi08679 & ~w17354;
assign w40034 = ~pi09848 & w17354;
assign w40035 = ~w40033 & ~w40034;
assign w40036 = pi08680 & ~w17354;
assign w40037 = w16978 & w17193;
assign w40038 = ~w40036 & ~w40037;
assign w40039 = pi08681 & ~w17354;
assign w40040 = ~pi02178 & w17354;
assign w40041 = ~w40039 & ~w40040;
assign w40042 = pi08682 & ~w17354;
assign w40043 = w16978 & w17513;
assign w40044 = ~w40042 & ~w40043;
assign w40045 = pi08683 & ~w17354;
assign w40046 = ~pi02720 & w17354;
assign w40047 = ~w40045 & ~w40046;
assign w40048 = pi08684 & ~w17354;
assign w40049 = ~pi09962 & w17354;
assign w40050 = ~w40048 & ~w40049;
assign w40051 = pi08685 & ~w17158;
assign w40052 = w16912 & w19365;
assign w40053 = ~w40051 & ~w40052;
assign w40054 = pi08686 & ~w17158;
assign w40055 = ~pi09848 & w17158;
assign w40056 = ~w40054 & ~w40055;
assign w40057 = pi08687 & ~w17158;
assign w40058 = ~pi09812 & w17158;
assign w40059 = ~w40057 & ~w40058;
assign w40060 = pi08688 & ~w17158;
assign w40061 = ~pi02178 & w17158;
assign w40062 = ~w40060 & ~w40061;
assign w40063 = pi08689 & ~w17158;
assign w40064 = ~pi09954 & w17158;
assign w40065 = ~w40063 & ~w40064;
assign w40066 = pi08690 & ~w17158;
assign w40067 = w16912 & w17128;
assign w40068 = ~w40066 & ~w40067;
assign w40069 = pi08691 & ~w17285;
assign w40070 = ~pi09961 & w17285;
assign w40071 = ~w40069 & ~w40070;
assign w40072 = pi08692 & ~w17285;
assign w40073 = ~pi09848 & w17285;
assign w40074 = ~w40072 & ~w40073;
assign w40075 = pi08693 & ~w17285;
assign w40076 = ~pi09812 & w17285;
assign w40077 = ~w40075 & ~w40076;
assign w40078 = pi08694 & ~w17285;
assign w40079 = ~pi02178 & w17285;
assign w40080 = ~w40078 & ~w40079;
assign w40081 = pi08695 & ~w17285;
assign w40082 = ~pi09954 & w17285;
assign w40083 = ~w40081 & ~w40082;
assign w40084 = pi08696 & ~w17285;
assign w40085 = ~pi02720 & w17285;
assign w40086 = ~w40084 & ~w40085;
assign w40087 = pi08697 & ~w17285;
assign w40088 = ~pi09962 & w17285;
assign w40089 = ~w40087 & ~w40088;
assign w40090 = pi08698 & ~w17178;
assign w40091 = ~pi09961 & w17178;
assign w40092 = ~w40090 & ~w40091;
assign w40093 = pi08699 & ~w17178;
assign w40094 = ~pi09848 & w17178;
assign w40095 = ~w40093 & ~w40094;
assign w40096 = pi08700 & ~w17178;
assign w40097 = ~pi09812 & w17178;
assign w40098 = ~w40096 & ~w40097;
assign w40099 = pi08701 & ~w17178;
assign w40100 = ~pi02178 & w17178;
assign w40101 = ~w40099 & ~w40100;
assign w40102 = pi08702 & ~w17178;
assign w40103 = ~pi09954 & w17178;
assign w40104 = ~w40102 & ~w40103;
assign w40105 = pi08703 & ~w17178;
assign w40106 = ~pi02720 & w17178;
assign w40107 = ~w40105 & ~w40106;
assign w40108 = ~w16928 & w18177;
assign w40109 = pi08704 & ~w40108;
assign w40110 = ~pi09961 & w40108;
assign w40111 = ~w40109 & ~w40110;
assign w40112 = pi08705 & ~w40108;
assign w40113 = ~pi09848 & w40108;
assign w40114 = ~w40112 & ~w40113;
assign w40115 = pi08706 & ~w40108;
assign w40116 = ~pi09812 & w40108;
assign w40117 = ~w40115 & ~w40116;
assign w40118 = pi08707 & ~w40108;
assign w40119 = ~pi02178 & w40108;
assign w40120 = ~w40118 & ~w40119;
assign w40121 = pi08708 & ~w40108;
assign w40122 = ~pi09954 & w40108;
assign w40123 = ~w40121 & ~w40122;
assign w40124 = pi08709 & ~w40108;
assign w40125 = ~pi02720 & w40108;
assign w40126 = ~w40124 & ~w40125;
assign w40127 = pi08710 & ~w40108;
assign w40128 = ~pi09962 & w40108;
assign w40129 = ~w40127 & ~w40128;
assign w40130 = pi08711 & ~w23529;
assign w40131 = ~pi09961 & w23529;
assign w40132 = ~w40130 & ~w40131;
assign w40133 = pi08712 & ~w23529;
assign w40134 = w17186 & w17565;
assign w40135 = ~w40133 & ~w40134;
assign w40136 = pi08713 & ~w23529;
assign w40137 = w17193 & w17565;
assign w40138 = ~w40136 & ~w40137;
assign w40139 = pi08714 & ~w23529;
assign w40140 = ~pi02178 & w23529;
assign w40141 = ~w40139 & ~w40140;
assign w40142 = pi08715 & ~w23529;
assign w40143 = ~pi09954 & w23529;
assign w40144 = ~w40142 & ~w40143;
assign w40145 = pi08716 & ~w23529;
assign w40146 = w17128 & w17565;
assign w40147 = ~w40145 & ~w40146;
assign w40148 = pi08717 & ~w21488;
assign w40149 = ~pi09812 & w21488;
assign w40150 = ~w40148 & ~w40149;
assign w40151 = pi08718 & ~w21262;
assign w40152 = w18040 & w19365;
assign w40153 = ~w40151 & ~w40152;
assign w40154 = pi08719 & ~w21262;
assign w40155 = ~pi09848 & w21262;
assign w40156 = ~w40154 & ~w40155;
assign w40157 = pi08720 & ~w21262;
assign w40158 = w17311 & w18040;
assign w40159 = ~w40157 & ~w40158;
assign w40160 = pi08721 & ~w21262;
assign w40161 = ~pi02178 & w21262;
assign w40162 = ~w40160 & ~w40161;
assign w40163 = pi08722 & ~w21262;
assign w40164 = ~pi09954 & w21262;
assign w40165 = ~w40163 & ~w40164;
assign w40166 = pi08723 & ~w21262;
assign w40167 = w17128 & w18040;
assign w40168 = ~w40166 & ~w40167;
assign w40169 = pi08724 & ~w21262;
assign w40170 = ~pi09962 & w21262;
assign w40171 = ~w40169 & ~w40170;
assign w40172 = pi08725 & ~w21341;
assign w40173 = w17917 & w19365;
assign w40174 = ~w40172 & ~w40173;
assign w40175 = pi08726 & ~w21341;
assign w40176 = ~pi09848 & w21341;
assign w40177 = ~w40175 & ~w40176;
assign w40178 = pi08727 & ~w21341;
assign w40179 = w17311 & w17917;
assign w40180 = ~w40178 & ~w40179;
assign w40181 = pi08728 & ~w21341;
assign w40182 = ~pi02178 & w21341;
assign w40183 = ~w40181 & ~w40182;
assign w40184 = pi08729 & ~w21341;
assign w40185 = ~pi09954 & w21341;
assign w40186 = ~w40184 & ~w40185;
assign w40187 = pi08730 & ~w21341;
assign w40188 = ~pi09962 & w21341;
assign w40189 = ~w40187 & ~w40188;
assign w40190 = pi08731 & ~w21378;
assign w40191 = ~pi09961 & w21378;
assign w40192 = ~w40190 & ~w40191;
assign w40193 = pi08732 & ~w21378;
assign w40194 = w17186 & w17668;
assign w40195 = ~w40193 & ~w40194;
assign w40196 = pi08733 & ~w21378;
assign w40197 = w17311 & w17668;
assign w40198 = ~w40196 & ~w40197;
assign w40199 = pi08734 & ~w21378;
assign w40200 = ~pi02178 & w21378;
assign w40201 = ~w40199 & ~w40200;
assign w40202 = pi08735 & ~w21378;
assign w40203 = ~pi09954 & w21378;
assign w40204 = ~w40202 & ~w40203;
assign w40205 = pi08736 & ~w21378;
assign w40206 = ~pi02720 & w21378;
assign w40207 = ~w40205 & ~w40206;
assign w40208 = pi08737 & ~w21378;
assign w40209 = ~pi09962 & w21378;
assign w40210 = ~w40208 & ~w40209;
assign w40211 = pi08738 & ~w20902;
assign w40212 = ~pi09961 & w20902;
assign w40213 = ~w40211 & ~w40212;
assign w40214 = pi08739 & ~w20902;
assign w40215 = w17186 & w17636;
assign w40216 = ~w40214 & ~w40215;
assign w40217 = pi08740 & ~w20902;
assign w40218 = ~pi02704 & w20902;
assign w40219 = ~w40217 & ~w40218;
assign w40220 = pi08741 & ~w20902;
assign w40221 = ~pi02178 & w20902;
assign w40222 = ~w40220 & ~w40221;
assign w40223 = pi08742 & ~w20902;
assign w40224 = w17513 & w17636;
assign w40225 = ~w40223 & ~w40224;
assign w40226 = pi08743 & ~w20902;
assign w40227 = ~pi09962 & w20902;
assign w40228 = ~w40226 & ~w40227;
assign w40229 = pi08744 & ~w21192;
assign w40230 = ~pi09961 & w21192;
assign w40231 = ~w40229 & ~w40230;
assign w40232 = pi08745 & ~w21192;
assign w40233 = w16961 & w17186;
assign w40234 = ~w40232 & ~w40233;
assign w40235 = pi08746 & ~w21192;
assign w40236 = ~pi02704 & w21192;
assign w40237 = ~w40235 & ~w40236;
assign w40238 = pi08747 & ~w21192;
assign w40239 = w16961 & w18861;
assign w40240 = ~w40238 & ~w40239;
assign w40241 = pi08748 & ~w21192;
assign w40242 = w16961 & w17513;
assign w40243 = ~w40241 & ~w40242;
assign w40244 = pi08749 & ~w21192;
assign w40245 = ~pi02720 & w21192;
assign w40246 = ~w40244 & ~w40245;
assign w40247 = pi08750 & ~w21192;
assign w40248 = w16961 & w17439;
assign w40249 = ~w40247 & ~w40248;
assign w40250 = pi08751 & ~w20887;
assign w40251 = ~pi09961 & w20887;
assign w40252 = ~w40250 & ~w40251;
assign w40253 = pi08752 & ~w20887;
assign w40254 = ~pi09848 & w20887;
assign w40255 = ~w40253 & ~w40254;
assign w40256 = pi08753 & ~w20887;
assign w40257 = ~pi02704 & w20887;
assign w40258 = ~w40256 & ~w40257;
assign w40259 = pi08754 & ~w20887;
assign w40260 = ~pi02178 & w20887;
assign w40261 = ~w40259 & ~w40260;
assign w40262 = pi08755 & ~w20887;
assign w40263 = ~pi09954 & w20887;
assign w40264 = ~w40262 & ~w40263;
assign w40265 = pi08756 & ~w20887;
assign w40266 = ~pi09962 & w20887;
assign w40267 = ~w40265 & ~w40266;
assign w40268 = pi08757 & ~w21004;
assign w40269 = w17650 & w19365;
assign w40270 = ~w40268 & ~w40269;
assign w40271 = pi08758 & ~w21004;
assign w40272 = ~pi09848 & w21004;
assign w40273 = ~w40271 & ~w40272;
assign w40274 = pi08759 & ~w21004;
assign w40275 = w17311 & w17650;
assign w40276 = ~w40274 & ~w40275;
assign w40277 = pi08760 & ~w21004;
assign w40278 = ~pi02178 & w21004;
assign w40279 = ~w40277 & ~w40278;
assign w40280 = pi08761 & ~w21004;
assign w40281 = ~pi09954 & w21004;
assign w40282 = ~w40280 & ~w40281;
assign w40283 = pi08762 & ~w21004;
assign w40284 = w17128 & w17650;
assign w40285 = ~w40283 & ~w40284;
assign w40286 = pi08763 & ~w21004;
assign w40287 = ~pi09962 & w21004;
assign w40288 = ~w40286 & ~w40287;
assign w40289 = pi08764 & ~w20799;
assign w40290 = w18622 & w19365;
assign w40291 = ~w40289 & ~w40290;
assign w40292 = pi08765 & ~w20799;
assign w40293 = ~pi09848 & w20799;
assign w40294 = ~w40292 & ~w40293;
assign w40295 = pi08766 & ~w20799;
assign w40296 = w17311 & w18622;
assign w40297 = ~w40295 & ~w40296;
assign w40298 = pi08767 & ~w20799;
assign w40299 = w18622 & w18861;
assign w40300 = ~w40298 & ~w40299;
assign w40301 = pi08768 & ~w20799;
assign w40302 = ~pi09954 & w20799;
assign w40303 = ~w40301 & ~w40302;
assign w40304 = pi08769 & ~w20799;
assign w40305 = ~pi09962 & w20799;
assign w40306 = ~w40304 & ~w40305;
assign w40307 = pi08770 & ~w17191;
assign w40308 = w17190 & w19365;
assign w40309 = ~w40307 & ~w40308;
assign w40310 = pi08771 & ~w17191;
assign w40311 = ~pi09848 & w17191;
assign w40312 = ~w40310 & ~w40311;
assign w40313 = pi08772 & ~w36892;
assign w40314 = ~pi02167 & w36892;
assign w40315 = ~w40313 & ~w40314;
assign w40316 = pi08773 & ~w17191;
assign w40317 = ~pi02704 & w17191;
assign w40318 = ~w40316 & ~w40317;
assign w40319 = pi08774 & ~w17191;
assign w40320 = w17190 & w18861;
assign w40321 = ~w40319 & ~w40320;
assign w40322 = pi08775 & ~w17191;
assign w40323 = ~pi02720 & w17191;
assign w40324 = ~w40322 & ~w40323;
assign w40325 = pi08776 & ~w17191;
assign w40326 = ~pi09954 & w17191;
assign w40327 = ~w40325 & ~w40326;
assign w40328 = pi08777 & ~w17191;
assign w40329 = ~pi09962 & w17191;
assign w40330 = ~w40328 & ~w40329;
assign w40331 = pi08778 & ~w18777;
assign w40332 = ~pi09961 & w18777;
assign w40333 = ~w40331 & ~w40332;
assign w40334 = pi08779 & ~w18777;
assign w40335 = ~pi09848 & w18777;
assign w40336 = ~w40334 & ~w40335;
assign w40337 = pi08780 & ~w18777;
assign w40338 = ~pi02178 & w18777;
assign w40339 = ~w40337 & ~w40338;
assign w40340 = pi08781 & ~w18777;
assign w40341 = ~pi09954 & w18777;
assign w40342 = ~w40340 & ~w40341;
assign w40343 = pi08782 & ~w18777;
assign w40344 = ~pi02720 & w18777;
assign w40345 = ~w40343 & ~w40344;
assign w40346 = pi08783 & ~w18777;
assign w40347 = ~pi09812 & w18777;
assign w40348 = ~w40346 & ~w40347;
assign w40349 = pi08784 & ~w18765;
assign w40350 = ~pi09961 & w18765;
assign w40351 = ~w40349 & ~w40350;
assign w40352 = pi08785 & ~w18765;
assign w40353 = ~pi09848 & w18765;
assign w40354 = ~w40352 & ~w40353;
assign w40355 = pi08786 & ~w18765;
assign w40356 = ~pi02704 & w18765;
assign w40357 = ~w40355 & ~w40356;
assign w40358 = pi08787 & ~w18765;
assign w40359 = ~pi02178 & w18765;
assign w40360 = ~w40358 & ~w40359;
assign w40361 = pi08788 & ~w18765;
assign w40362 = ~pi09954 & w18765;
assign w40363 = ~w40361 & ~w40362;
assign w40364 = pi08789 & ~w18765;
assign w40365 = ~pi02720 & w18765;
assign w40366 = ~w40364 & ~w40365;
assign w40367 = pi08790 & ~w18765;
assign w40368 = ~pi09962 & w18765;
assign w40369 = ~w40367 & ~w40368;
assign w40370 = pi08791 & ~w18732;
assign w40371 = ~pi09961 & w18732;
assign w40372 = ~w40370 & ~w40371;
assign w40373 = pi08792 & ~w18732;
assign w40374 = ~pi09848 & w18732;
assign w40375 = ~w40373 & ~w40374;
assign w40376 = pi08793 & ~w18732;
assign w40377 = w17311 & w18731;
assign w40378 = ~w40376 & ~w40377;
assign w40379 = pi08794 & ~w18732;
assign w40380 = ~pi02178 & w18732;
assign w40381 = ~w40379 & ~w40380;
assign w40382 = pi08795 & ~w18732;
assign w40383 = ~pi09954 & w18732;
assign w40384 = ~w40382 & ~w40383;
assign w40385 = pi08796 & ~w18732;
assign w40386 = ~pi09962 & w18732;
assign w40387 = ~w40385 & ~w40386;
assign w40388 = pi08797 & ~w18684;
assign w40389 = ~pi09961 & w18684;
assign w40390 = ~w40388 & ~w40389;
assign w40391 = pi08798 & ~w18684;
assign w40392 = w17186 & w18683;
assign w40393 = ~w40391 & ~w40392;
assign w40394 = pi08799 & ~w18684;
assign w40395 = ~pi02704 & w18684;
assign w40396 = ~w40394 & ~w40395;
assign w40397 = pi08800 & ~w18684;
assign w40398 = ~pi02178 & w18684;
assign w40399 = ~w40397 & ~w40398;
assign w40400 = pi08801 & ~w18684;
assign w40401 = ~pi09954 & w18684;
assign w40402 = ~w40400 & ~w40401;
assign w40403 = pi08802 & ~w18684;
assign w40404 = w17128 & w18683;
assign w40405 = ~w40403 & ~w40404;
assign w40406 = pi08803 & ~w18684;
assign w40407 = w17439 & w18683;
assign w40408 = ~w40406 & ~w40407;
assign w40409 = pi08804 & ~w18349;
assign w40410 = ~pi09961 & w18349;
assign w40411 = ~w40409 & ~w40410;
assign w40412 = pi08805 & ~w18349;
assign w40413 = ~pi09848 & w18349;
assign w40414 = ~w40412 & ~w40413;
assign w40415 = pi08806 & ~w18349;
assign w40416 = ~pi02704 & w18349;
assign w40417 = ~w40415 & ~w40416;
assign w40418 = pi08807 & ~w18349;
assign w40419 = ~pi02178 & w18349;
assign w40420 = ~w40418 & ~w40419;
assign w40421 = pi08808 & ~w18349;
assign w40422 = ~pi09954 & w18349;
assign w40423 = ~w40421 & ~w40422;
assign w40424 = pi08809 & ~w18349;
assign w40425 = ~pi09962 & w18349;
assign w40426 = ~w40424 & ~w40425;
assign w40427 = pi08810 & ~w17522;
assign w40428 = ~pi09961 & w17522;
assign w40429 = ~w40427 & ~w40428;
assign w40430 = pi08811 & ~w17522;
assign w40431 = ~pi09848 & w17522;
assign w40432 = ~w40430 & ~w40431;
assign w40433 = pi08812 & ~w17522;
assign w40434 = ~pi02704 & w17522;
assign w40435 = ~w40433 & ~w40434;
assign w40436 = pi08813 & ~w17522;
assign w40437 = ~pi02178 & w17522;
assign w40438 = ~w40436 & ~w40437;
assign w40439 = pi08814 & ~w17522;
assign w40440 = ~pi09954 & w17522;
assign w40441 = ~w40439 & ~w40440;
assign w40442 = pi08815 & ~w17522;
assign w40443 = ~pi02720 & w17522;
assign w40444 = ~w40442 & ~w40443;
assign w40445 = pi08816 & ~w17522;
assign w40446 = ~pi09962 & w17522;
assign w40447 = ~w40445 & ~w40446;
assign w40448 = pi08817 & ~w17326;
assign w40449 = ~pi09961 & w17326;
assign w40450 = ~w40448 & ~w40449;
assign w40451 = pi08818 & ~w17326;
assign w40452 = w17186 & w17325;
assign w40453 = ~w40451 & ~w40452;
assign w40454 = pi08819 & ~w17326;
assign w40455 = ~pi02704 & w17326;
assign w40456 = ~w40454 & ~w40455;
assign w40457 = pi08820 & ~w17326;
assign w40458 = ~pi02178 & w17326;
assign w40459 = ~w40457 & ~w40458;
assign w40460 = pi08821 & ~w17326;
assign w40461 = ~pi09954 & w17326;
assign w40462 = ~w40460 & ~w40461;
assign w40463 = pi08822 & ~w17326;
assign w40464 = w17325 & w17439;
assign w40465 = ~w40463 & ~w40464;
assign w40466 = pi08823 & ~w17475;
assign w40467 = ~pi09961 & w17475;
assign w40468 = ~w40466 & ~w40467;
assign w40469 = pi08824 & ~w17475;
assign w40470 = ~pi09848 & w17475;
assign w40471 = ~w40469 & ~w40470;
assign w40472 = pi08825 & ~w17475;
assign w40473 = ~pi02704 & w17475;
assign w40474 = ~w40472 & ~w40473;
assign w40475 = pi08826 & ~w17475;
assign w40476 = ~pi02178 & w17475;
assign w40477 = ~w40475 & ~w40476;
assign w40478 = pi08827 & ~w17475;
assign w40479 = ~pi09954 & w17475;
assign w40480 = ~w40478 & ~w40479;
assign w40481 = pi08828 & ~w17475;
assign w40482 = ~pi02720 & w17475;
assign w40483 = ~w40481 & ~w40482;
assign w40484 = pi08829 & ~w17475;
assign w40485 = ~pi09962 & w17475;
assign w40486 = ~w40484 & ~w40485;
assign w40487 = pi08830 & ~w17321;
assign w40488 = ~pi09961 & w17321;
assign w40489 = ~w40487 & ~w40488;
assign w40490 = pi08831 & ~w17321;
assign w40491 = ~pi09848 & w17321;
assign w40492 = ~w40490 & ~w40491;
assign w40493 = pi08832 & ~w17321;
assign w40494 = ~pi02704 & w17321;
assign w40495 = ~w40493 & ~w40494;
assign w40496 = pi08833 & ~w17321;
assign w40497 = ~pi02178 & w17321;
assign w40498 = ~w40496 & ~w40497;
assign w40499 = pi08834 & ~w17321;
assign w40500 = w17320 & w17513;
assign w40501 = ~w40499 & ~w40500;
assign w40502 = pi08835 & ~w17321;
assign w40503 = w17320 & w17439;
assign w40504 = ~w40502 & ~w40503;
assign w40505 = pi08836 & ~w17345;
assign w40506 = ~pi09961 & w17345;
assign w40507 = ~w40505 & ~w40506;
assign w40508 = pi08837 & ~w17345;
assign w40509 = ~pi09848 & w17345;
assign w40510 = ~w40508 & ~w40509;
assign w40511 = pi08838 & ~w17345;
assign w40512 = ~pi02704 & w17345;
assign w40513 = ~w40511 & ~w40512;
assign w40514 = pi08839 & ~w17345;
assign w40515 = w17344 & w18861;
assign w40516 = ~w40514 & ~w40515;
assign w40517 = pi08840 & ~w17345;
assign w40518 = ~pi09954 & w17345;
assign w40519 = ~w40517 & ~w40518;
assign w40520 = pi08841 & ~w17345;
assign w40521 = ~pi02720 & w17345;
assign w40522 = ~w40520 & ~w40521;
assign w40523 = pi08842 & ~w17345;
assign w40524 = ~pi09962 & w17345;
assign w40525 = ~w40523 & ~w40524;
assign w40526 = pi08843 & ~w17163;
assign w40527 = ~pi09961 & w17163;
assign w40528 = ~w40526 & ~w40527;
assign w40529 = pi08844 & ~w17163;
assign w40530 = ~pi09848 & w17163;
assign w40531 = ~w40529 & ~w40530;
assign w40532 = pi08845 & ~w17163;
assign w40533 = ~pi02704 & w17163;
assign w40534 = ~w40532 & ~w40533;
assign w40535 = pi08846 & ~w17163;
assign w40536 = ~pi02178 & w17163;
assign w40537 = ~w40535 & ~w40536;
assign w40538 = pi08847 & ~w17163;
assign w40539 = ~pi09954 & w17163;
assign w40540 = ~w40538 & ~w40539;
assign w40541 = pi08848 & ~w17163;
assign w40542 = ~pi09962 & w17163;
assign w40543 = ~w40541 & ~w40542;
assign w40544 = pi08849 & ~w17245;
assign w40545 = ~pi09961 & w17245;
assign w40546 = ~w40544 & ~w40545;
assign w40547 = pi08850 & ~w17245;
assign w40548 = ~pi09848 & w17245;
assign w40549 = ~w40547 & ~w40548;
assign w40550 = pi08851 & ~w17245;
assign w40551 = ~pi02704 & w17245;
assign w40552 = ~w40550 & ~w40551;
assign w40553 = pi08852 & ~w17245;
assign w40554 = ~pi02178 & w17245;
assign w40555 = ~w40553 & ~w40554;
assign w40556 = pi08853 & ~w17245;
assign w40557 = ~pi09954 & w17245;
assign w40558 = ~w40556 & ~w40557;
assign w40559 = pi08854 & ~w17245;
assign w40560 = ~pi02720 & w17245;
assign w40561 = ~w40559 & ~w40560;
assign w40562 = pi08855 & ~w17245;
assign w40563 = ~pi09962 & w17245;
assign w40564 = ~w40562 & ~w40563;
assign w40565 = pi08856 & ~w31269;
assign w40566 = ~pi09961 & w31269;
assign w40567 = ~w40565 & ~w40566;
assign w40568 = pi08857 & ~w31269;
assign w40569 = ~pi09848 & w31269;
assign w40570 = ~w40568 & ~w40569;
assign w40571 = pi08858 & ~w31269;
assign w40572 = ~pi02704 & w31269;
assign w40573 = ~w40571 & ~w40572;
assign w40574 = pi08859 & ~w31269;
assign w40575 = ~pi02178 & w31269;
assign w40576 = ~w40574 & ~w40575;
assign w40577 = pi08860 & ~w31269;
assign w40578 = ~pi09954 & w31269;
assign w40579 = ~w40577 & ~w40578;
assign w40580 = pi08861 & ~w31269;
assign w40581 = ~pi09962 & w31269;
assign w40582 = ~w40580 & ~w40581;
assign w40583 = pi08862 & ~w27038;
assign w40584 = ~pi09961 & w27038;
assign w40585 = ~w40583 & ~w40584;
assign w40586 = pi08863 & ~w27038;
assign w40587 = ~pi09848 & w27038;
assign w40588 = ~w40586 & ~w40587;
assign w40589 = pi08864 & ~w27038;
assign w40590 = ~pi02704 & w27038;
assign w40591 = ~w40589 & ~w40590;
assign w40592 = pi08865 & ~w27038;
assign w40593 = ~pi02178 & w27038;
assign w40594 = ~w40592 & ~w40593;
assign w40595 = pi08866 & ~w27038;
assign w40596 = ~pi09954 & w27038;
assign w40597 = ~w40595 & ~w40596;
assign w40598 = pi08867 & ~w27038;
assign w40599 = w17128 & w18217;
assign w40600 = ~w40598 & ~w40599;
assign w40601 = pi08868 & ~w27038;
assign w40602 = ~pi09962 & w27038;
assign w40603 = ~w40601 & ~w40602;
assign w40604 = pi08869 & ~w21224;
assign w40605 = ~pi09961 & w21224;
assign w40606 = ~w40604 & ~w40605;
assign w40607 = pi08870 & ~w21224;
assign w40608 = ~pi09848 & w21224;
assign w40609 = ~w40607 & ~w40608;
assign w40610 = pi08871 & ~w21224;
assign w40611 = ~pi02704 & w21224;
assign w40612 = ~w40610 & ~w40611;
assign w40613 = pi08872 & ~w21224;
assign w40614 = ~pi02178 & w21224;
assign w40615 = ~w40613 & ~w40614;
assign w40616 = pi08873 & ~w21224;
assign w40617 = ~pi09954 & w21224;
assign w40618 = ~w40616 & ~w40617;
assign w40619 = pi08874 & ~w21224;
assign w40620 = ~pi09962 & w21224;
assign w40621 = ~w40619 & ~w40620;
assign w40622 = pi08875 & ~w21432;
assign w40623 = ~pi09961 & w21432;
assign w40624 = ~w40622 & ~w40623;
assign w40625 = pi08876 & ~w21432;
assign w40626 = ~pi09848 & w21432;
assign w40627 = ~w40625 & ~w40626;
assign w40628 = pi08877 & ~w21432;
assign w40629 = w16986 & w17311;
assign w40630 = ~w40628 & ~w40629;
assign w40631 = pi08878 & ~w21432;
assign w40632 = ~pi02178 & w21432;
assign w40633 = ~w40631 & ~w40632;
assign w40634 = pi08879 & ~w21432;
assign w40635 = ~pi09954 & w21432;
assign w40636 = ~w40634 & ~w40635;
assign w40637 = pi08880 & ~w21432;
assign w40638 = ~pi02720 & w21432;
assign w40639 = ~w40637 & ~w40638;
assign w40640 = pi08881 & ~w21432;
assign w40641 = ~pi09962 & w21432;
assign w40642 = ~w40640 & ~w40641;
assign w40643 = pi08882 & ~w21146;
assign w40644 = w17694 & w19365;
assign w40645 = ~w40643 & ~w40644;
assign w40646 = pi08883 & ~w21146;
assign w40647 = w17186 & w17694;
assign w40648 = ~w40646 & ~w40647;
assign w40649 = pi08884 & ~w21146;
assign w40650 = ~pi02704 & w21146;
assign w40651 = ~w40649 & ~w40650;
assign w40652 = pi08885 & ~w21146;
assign w40653 = w17694 & w18861;
assign w40654 = ~w40652 & ~w40653;
assign w40655 = pi08886 & ~w21146;
assign w40656 = ~pi09954 & w21146;
assign w40657 = ~w40655 & ~w40656;
assign w40658 = pi08887 & ~w21146;
assign w40659 = ~pi09962 & w21146;
assign w40660 = ~w40658 & ~w40659;
assign w40661 = pi08888 & ~w20924;
assign w40662 = ~pi09961 & w20924;
assign w40663 = ~w40661 & ~w40662;
assign w40664 = pi08889 & ~w20924;
assign w40665 = ~pi09848 & w20924;
assign w40666 = ~w40664 & ~w40665;
assign w40667 = pi08890 & ~w20924;
assign w40668 = ~pi02704 & w20924;
assign w40669 = ~w40667 & ~w40668;
assign w40670 = pi08891 & ~w20924;
assign w40671 = ~pi02178 & w20924;
assign w40672 = ~w40670 & ~w40671;
assign w40673 = pi08892 & ~w20924;
assign w40674 = ~pi09954 & w20924;
assign w40675 = ~w40673 & ~w40674;
assign w40676 = pi08893 & ~w20924;
assign w40677 = ~pi02720 & w20924;
assign w40678 = ~w40676 & ~w40677;
assign w40679 = pi08894 & ~w20924;
assign w40680 = ~pi09962 & w20924;
assign w40681 = ~w40679 & ~w40680;
assign w40682 = pi08895 & ~w17149;
assign w40683 = ~pi09961 & w17149;
assign w40684 = ~w40682 & ~w40683;
assign w40685 = pi08896 & ~w17149;
assign w40686 = ~pi09848 & w17149;
assign w40687 = ~w40685 & ~w40686;
assign w40688 = pi08897 & ~w17149;
assign w40689 = ~pi02704 & w17149;
assign w40690 = ~w40688 & ~w40689;
assign w40691 = pi08898 & ~w17149;
assign w40692 = ~pi02178 & w17149;
assign w40693 = ~w40691 & ~w40692;
assign w40694 = pi08899 & ~w17149;
assign w40695 = ~pi09954 & w17149;
assign w40696 = ~w40694 & ~w40695;
assign w40697 = pi08900 & ~w17149;
assign w40698 = ~pi09962 & w17149;
assign w40699 = ~w40697 & ~w40698;
assign w40700 = pi08901 & ~w18564;
assign w40701 = ~pi09961 & w18564;
assign w40702 = ~w40700 & ~w40701;
assign w40703 = pi08902 & ~w18564;
assign w40704 = ~pi09848 & w18564;
assign w40705 = ~w40703 & ~w40704;
assign w40706 = pi08903 & ~w18564;
assign w40707 = ~pi02704 & w18564;
assign w40708 = ~w40706 & ~w40707;
assign w40709 = pi08904 & ~w18564;
assign w40710 = ~pi02178 & w18564;
assign w40711 = ~w40709 & ~w40710;
assign w40712 = pi08905 & ~w18564;
assign w40713 = ~pi09954 & w18564;
assign w40714 = ~w40712 & ~w40713;
assign w40715 = pi08906 & ~w18564;
assign w40716 = ~pi02720 & w18564;
assign w40717 = ~w40715 & ~w40716;
assign w40718 = pi08907 & ~w18564;
assign w40719 = ~pi09962 & w18564;
assign w40720 = ~w40718 & ~w40719;
assign w40721 = pi08908 & ~w18814;
assign w40722 = w18813 & w19365;
assign w40723 = ~w40721 & ~w40722;
assign w40724 = pi08909 & ~w18814;
assign w40725 = w17186 & w18813;
assign w40726 = ~w40724 & ~w40725;
assign w40727 = pi08910 & ~w18814;
assign w40728 = w17311 & w18813;
assign w40729 = ~w40727 & ~w40728;
assign w40730 = pi08911 & ~w18814;
assign w40731 = ~pi02178 & w18814;
assign w40732 = ~w40730 & ~w40731;
assign w40733 = pi08912 & ~w18814;
assign w40734 = ~pi09954 & w18814;
assign w40735 = ~w40733 & ~w40734;
assign w40736 = pi08913 & ~w18814;
assign w40737 = ~pi09962 & w18814;
assign w40738 = ~w40736 & ~w40737;
assign w40739 = pi08914 & ~w18782;
assign w40740 = w18781 & w19365;
assign w40741 = ~w40739 & ~w40740;
assign w40742 = pi08915 & ~w18782;
assign w40743 = ~pi09848 & w18782;
assign w40744 = ~w40742 & ~w40743;
assign w40745 = pi08916 & ~w18782;
assign w40746 = ~pi02704 & w18782;
assign w40747 = ~w40745 & ~w40746;
assign w40748 = pi08917 & ~w18782;
assign w40749 = ~pi02178 & w18782;
assign w40750 = ~w40748 & ~w40749;
assign w40751 = pi08918 & ~w18782;
assign w40752 = ~pi09954 & w18782;
assign w40753 = ~w40751 & ~w40752;
assign w40754 = pi08919 & ~w18782;
assign w40755 = ~pi02720 & w18782;
assign w40756 = ~w40754 & ~w40755;
assign w40757 = pi08920 & ~w18782;
assign w40758 = ~pi09962 & w18782;
assign w40759 = ~w40757 & ~w40758;
assign w40760 = pi08921 & ~w17506;
assign w40761 = ~pi09961 & w17506;
assign w40762 = ~w40760 & ~w40761;
assign w40763 = pi08922 & ~w17506;
assign w40764 = w17186 & w17505;
assign w40765 = ~w40763 & ~w40764;
assign w40766 = pi08923 & ~w17506;
assign w40767 = w17311 & w17505;
assign w40768 = ~w40766 & ~w40767;
assign w40769 = pi08924 & ~w17506;
assign w40770 = ~pi02178 & w17506;
assign w40771 = ~w40769 & ~w40770;
assign w40772 = pi08925 & ~w17506;
assign w40773 = w17128 & w17505;
assign w40774 = ~w40772 & ~w40773;
assign w40775 = pi08926 & ~w17506;
assign w40776 = ~pi09962 & w17506;
assign w40777 = ~w40775 & ~w40776;
assign w40778 = pi08927 & ~w18450;
assign w40779 = w18449 & w19365;
assign w40780 = ~w40778 & ~w40779;
assign w40781 = pi08928 & ~w18450;
assign w40782 = ~pi09848 & w18450;
assign w40783 = ~w40781 & ~w40782;
assign w40784 = pi08929 & ~w18450;
assign w40785 = ~pi02704 & w18450;
assign w40786 = ~w40784 & ~w40785;
assign w40787 = pi08930 & ~w18450;
assign w40788 = ~pi02178 & w18450;
assign w40789 = ~w40787 & ~w40788;
assign w40790 = pi08931 & ~w18450;
assign w40791 = ~pi09954 & w18450;
assign w40792 = ~w40790 & ~w40791;
assign w40793 = pi08932 & ~w18450;
assign w40794 = ~pi02720 & w18450;
assign w40795 = ~w40793 & ~w40794;
assign w40796 = pi08933 & ~w18450;
assign w40797 = ~pi09962 & w18450;
assign w40798 = ~w40796 & ~w40797;
assign w40799 = pi08934 & ~w17154;
assign w40800 = ~pi09961 & w17154;
assign w40801 = ~w40799 & ~w40800;
assign w40802 = pi08935 & ~w17154;
assign w40803 = w17153 & w17186;
assign w40804 = ~w40802 & ~w40803;
assign w40805 = pi08936 & ~w17154;
assign w40806 = ~pi02704 & w17154;
assign w40807 = ~w40805 & ~w40806;
assign w40808 = pi08937 & ~w17154;
assign w40809 = ~pi02178 & w17154;
assign w40810 = ~w40808 & ~w40809;
assign w40811 = pi08938 & ~w17154;
assign w40812 = w17153 & w17513;
assign w40813 = ~w40811 & ~w40812;
assign w40814 = pi08939 & ~w17154;
assign w40815 = ~pi09962 & w17154;
assign w40816 = ~w40814 & ~w40815;
assign w40817 = pi08940 & ~w17467;
assign w40818 = ~pi09961 & w17467;
assign w40819 = ~w40817 & ~w40818;
assign w40820 = pi08941 & ~w17467;
assign w40821 = ~pi09848 & w17467;
assign w40822 = ~w40820 & ~w40821;
assign w40823 = pi08942 & ~w17467;
assign w40824 = ~pi02704 & w17467;
assign w40825 = ~w40823 & ~w40824;
assign w40826 = pi08943 & ~w17467;
assign w40827 = ~pi02178 & w17467;
assign w40828 = ~w40826 & ~w40827;
assign w40829 = pi08944 & ~w17467;
assign w40830 = ~pi09954 & w17467;
assign w40831 = ~w40829 & ~w40830;
assign w40832 = pi08945 & ~w17467;
assign w40833 = ~pi02720 & w17467;
assign w40834 = ~w40832 & ~w40833;
assign w40835 = pi08946 & ~w17467;
assign w40836 = ~pi09962 & w17467;
assign w40837 = ~w40835 & ~w40836;
assign w40838 = pi08947 & ~w17421;
assign w40839 = w17339 & w19365;
assign w40840 = ~w40838 & ~w40839;
assign w40841 = pi08948 & ~w17421;
assign w40842 = ~pi09848 & w17421;
assign w40843 = ~w40841 & ~w40842;
assign w40844 = pi08949 & ~w17421;
assign w40845 = ~pi02704 & w17421;
assign w40846 = ~w40844 & ~w40845;
assign w40847 = pi08950 & ~w17421;
assign w40848 = ~pi02178 & w17421;
assign w40849 = ~w40847 & ~w40848;
assign w40850 = pi08951 & ~w17421;
assign w40851 = w17339 & w17513;
assign w40852 = ~w40850 & ~w40851;
assign w40853 = pi08952 & ~w17421;
assign w40854 = ~pi09962 & w17421;
assign w40855 = ~w40853 & ~w40854;
assign w40856 = pi08953 & ~w17301;
assign w40857 = ~pi09961 & w17301;
assign w40858 = ~w40856 & ~w40857;
assign w40859 = pi08954 & ~w17301;
assign w40860 = ~pi09848 & w17301;
assign w40861 = ~w40859 & ~w40860;
assign w40862 = pi08955 & ~w17301;
assign w40863 = ~pi02704 & w17301;
assign w40864 = ~w40862 & ~w40863;
assign w40865 = pi08956 & ~w17301;
assign w40866 = ~pi02178 & w17301;
assign w40867 = ~w40865 & ~w40866;
assign w40868 = pi08957 & ~w17301;
assign w40869 = ~pi09954 & w17301;
assign w40870 = ~w40868 & ~w40869;
assign w40871 = pi08958 & ~w17301;
assign w40872 = w17128 & w17300;
assign w40873 = ~w40871 & ~w40872;
assign w40874 = pi08959 & ~w17301;
assign w40875 = ~pi09962 & w17301;
assign w40876 = ~w40874 & ~w40875;
assign w40877 = pi08960 & ~w17255;
assign w40878 = ~pi09961 & w17255;
assign w40879 = ~w40877 & ~w40878;
assign w40880 = pi08961 & ~w17255;
assign w40881 = ~pi09848 & w17255;
assign w40882 = ~w40880 & ~w40881;
assign w40883 = pi08962 & ~w17255;
assign w40884 = ~pi02704 & w17255;
assign w40885 = ~w40883 & ~w40884;
assign w40886 = pi08963 & ~w17255;
assign w40887 = ~pi02178 & w17255;
assign w40888 = ~w40886 & ~w40887;
assign w40889 = pi08964 & ~w17255;
assign w40890 = ~pi09954 & w17255;
assign w40891 = ~w40889 & ~w40890;
assign w40892 = pi08965 & ~w17255;
assign w40893 = ~pi09962 & w17255;
assign w40894 = ~w40892 & ~w40893;
assign w40895 = pi08966 & ~w17265;
assign w40896 = w17264 & w19365;
assign w40897 = ~w40895 & ~w40896;
assign w40898 = pi08967 & ~w17265;
assign w40899 = w17186 & w17264;
assign w40900 = ~w40898 & ~w40899;
assign w40901 = pi08968 & ~w17265;
assign w40902 = w17264 & w17311;
assign w40903 = ~w40901 & ~w40902;
assign w40904 = pi08969 & ~w17265;
assign w40905 = w17264 & w18861;
assign w40906 = ~w40904 & ~w40905;
assign w40907 = pi08970 & ~w17265;
assign w40908 = w17264 & w17513;
assign w40909 = ~w40907 & ~w40908;
assign w40910 = pi08971 & ~w17265;
assign w40911 = w17128 & w17264;
assign w40912 = ~w40910 & ~w40911;
assign w40913 = pi08972 & ~w17265;
assign w40914 = w17264 & w17439;
assign w40915 = ~w40913 & ~w40914;
assign w40916 = pi08973 & ~w21216;
assign w40917 = w17663 & w19365;
assign w40918 = ~w40916 & ~w40917;
assign w40919 = pi08974 & ~w21216;
assign w40920 = w17186 & w17663;
assign w40921 = ~w40919 & ~w40920;
assign w40922 = pi08975 & ~w21216;
assign w40923 = ~pi02704 & w21216;
assign w40924 = ~w40922 & ~w40923;
assign w40925 = pi08976 & ~w21216;
assign w40926 = ~pi02178 & w21216;
assign w40927 = ~w40925 & ~w40926;
assign w40928 = pi08977 & ~w21216;
assign w40929 = ~pi09954 & w21216;
assign w40930 = ~w40928 & ~w40929;
assign w40931 = pi08978 & ~w21216;
assign w40932 = ~pi09962 & w21216;
assign w40933 = ~w40931 & ~w40932;
assign w40934 = pi08979 & ~w21326;
assign w40935 = ~pi09961 & w21326;
assign w40936 = ~w40934 & ~w40935;
assign w40937 = pi08980 & ~w21326;
assign w40938 = ~pi09848 & w21326;
assign w40939 = ~w40937 & ~w40938;
assign w40940 = pi08981 & ~w21326;
assign w40941 = ~pi02704 & w21326;
assign w40942 = ~w40940 & ~w40941;
assign w40943 = pi08982 & ~w21326;
assign w40944 = ~pi02178 & w21326;
assign w40945 = ~w40943 & ~w40944;
assign w40946 = pi08983 & ~w21326;
assign w40947 = w17513 & w17681;
assign w40948 = ~w40946 & ~w40947;
assign w40949 = pi08984 & ~w21326;
assign w40950 = ~pi02720 & w21326;
assign w40951 = ~w40949 & ~w40950;
assign w40952 = pi08985 & ~w21326;
assign w40953 = ~pi09962 & w21326;
assign w40954 = ~w40952 & ~w40953;
assign w40955 = pi08986 & ~w21352;
assign w40956 = ~pi09961 & w21352;
assign w40957 = ~w40955 & ~w40956;
assign w40958 = pi08987 & ~w21352;
assign w40959 = ~pi09848 & w21352;
assign w40960 = ~w40958 & ~w40959;
assign w40961 = pi08988 & ~w21352;
assign w40962 = w17311 & w17749;
assign w40963 = ~w40961 & ~w40962;
assign w40964 = pi08989 & ~w21352;
assign w40965 = ~pi02178 & w21352;
assign w40966 = ~w40964 & ~w40965;
assign w40967 = pi08990 & ~w21352;
assign w40968 = ~pi09954 & w21352;
assign w40969 = ~w40967 & ~w40968;
assign w40970 = pi08991 & ~w21352;
assign w40971 = ~pi09962 & w21352;
assign w40972 = ~w40970 & ~w40971;
assign w40973 = pi08992 & ~w21307;
assign w40974 = ~pi09961 & w21307;
assign w40975 = ~w40973 & ~w40974;
assign w40976 = pi08993 & ~w21307;
assign w40977 = ~pi09848 & w21307;
assign w40978 = ~w40976 & ~w40977;
assign w40979 = pi08994 & ~w21307;
assign w40980 = ~pi02704 & w21307;
assign w40981 = ~w40979 & ~w40980;
assign w40982 = pi08995 & ~w21307;
assign w40983 = ~pi02178 & w21307;
assign w40984 = ~w40982 & ~w40983;
assign w40985 = pi08996 & ~w21307;
assign w40986 = ~pi09954 & w21307;
assign w40987 = ~w40985 & ~w40986;
assign w40988 = pi08997 & ~w21307;
assign w40989 = w17128 & w17658;
assign w40990 = ~w40988 & ~w40989;
assign w40991 = pi08998 & ~w21307;
assign w40992 = w17439 & w17658;
assign w40993 = ~w40991 & ~w40992;
assign w40994 = pi08999 & ~w21258;
assign w40995 = ~pi09961 & w21258;
assign w40996 = ~w40994 & ~w40995;
assign w40997 = pi09000 & ~w21258;
assign w40998 = ~pi09848 & w21258;
assign w40999 = ~w40997 & ~w40998;
assign w41000 = pi09001 & ~w21258;
assign w41001 = ~pi02704 & w21258;
assign w41002 = ~w41000 & ~w41001;
assign w41003 = pi09002 & ~w21258;
assign w41004 = w18861 & w20561;
assign w41005 = ~w41003 & ~w41004;
assign w41006 = pi09003 & ~w21258;
assign w41007 = ~pi02720 & w21258;
assign w41008 = ~w41006 & ~w41007;
assign w41009 = pi09004 & ~w21258;
assign w41010 = ~pi09962 & w21258;
assign w41011 = ~w41009 & ~w41010;
assign w41012 = pi09005 & ~w21239;
assign w41013 = w19365 & w20470;
assign w41014 = ~w41012 & ~w41013;
assign w41015 = pi09006 & ~w21239;
assign w41016 = ~pi09848 & w21239;
assign w41017 = ~w41015 & ~w41016;
assign w41018 = pi09007 & ~w21239;
assign w41019 = ~pi02178 & w21239;
assign w41020 = ~w41018 & ~w41019;
assign w41021 = pi09008 & ~w21239;
assign w41022 = ~pi09954 & w21239;
assign w41023 = ~w41021 & ~w41022;
assign w41024 = pi09009 & ~w21239;
assign w41025 = ~pi02720 & w21239;
assign w41026 = ~w41024 & ~w41025;
assign w41027 = pi09010 & ~w21239;
assign w41028 = ~pi09962 & w21239;
assign w41029 = ~w41027 & ~w41028;
assign w41030 = pi09011 & ~w21239;
assign w41031 = ~pi02704 & w21239;
assign w41032 = ~w41030 & ~w41031;
assign w41033 = pi09012 & ~w21142;
assign w41034 = ~pi09961 & w21142;
assign w41035 = ~w41033 & ~w41034;
assign w41036 = pi09013 & ~w21142;
assign w41037 = ~pi09848 & w21142;
assign w41038 = ~w41036 & ~w41037;
assign w41039 = pi09014 & ~w21142;
assign w41040 = ~pi02704 & w21142;
assign w41041 = ~w41039 & ~w41040;
assign w41042 = pi09015 & ~w21142;
assign w41043 = w18032 & w18861;
assign w41044 = ~w41042 & ~w41043;
assign w41045 = pi09016 & ~w21142;
assign w41046 = ~pi09954 & w21142;
assign w41047 = ~w41045 & ~w41046;
assign w41048 = pi09017 & ~w21142;
assign w41049 = ~pi09962 & w21142;
assign w41050 = ~w41048 & ~w41049;
assign w41051 = pi09018 & ~w20996;
assign w41052 = ~pi09961 & w20996;
assign w41053 = ~w41051 & ~w41052;
assign w41054 = pi09019 & ~w20996;
assign w41055 = ~pi09848 & w20996;
assign w41056 = ~w41054 & ~w41055;
assign w41057 = pi09020 & ~w20996;
assign w41058 = ~pi02704 & w20996;
assign w41059 = ~w41057 & ~w41058;
assign w41060 = pi09021 & ~w20996;
assign w41061 = ~pi02178 & w20996;
assign w41062 = ~w41060 & ~w41061;
assign w41063 = pi09022 & ~w20996;
assign w41064 = ~pi09954 & w20996;
assign w41065 = ~w41063 & ~w41064;
assign w41066 = pi09023 & ~w20996;
assign w41067 = ~pi02720 & w20996;
assign w41068 = ~w41066 & ~w41067;
assign w41069 = pi09024 & ~w20996;
assign w41070 = ~pi09962 & w20996;
assign w41071 = ~w41069 & ~w41070;
assign w41072 = pi09025 & ~w18514;
assign w41073 = ~pi09961 & w18514;
assign w41074 = ~w41072 & ~w41073;
assign w41075 = pi09026 & ~w18514;
assign w41076 = ~pi09848 & w18514;
assign w41077 = ~w41075 & ~w41076;
assign w41078 = pi09027 & ~w18514;
assign w41079 = ~pi02704 & w18514;
assign w41080 = ~w41078 & ~w41079;
assign w41081 = pi09028 & ~w18514;
assign w41082 = w17540 & w18861;
assign w41083 = ~w41081 & ~w41082;
assign w41084 = pi09029 & ~w18514;
assign w41085 = ~pi09954 & w18514;
assign w41086 = ~w41084 & ~w41085;
assign w41087 = pi09030 & ~w18514;
assign w41088 = ~pi09962 & w18514;
assign w41089 = ~w41087 & ~w41088;
assign w41090 = pi09031 & ~w18950;
assign w41091 = ~pi09961 & w18950;
assign w41092 = ~w41090 & ~w41091;
assign w41093 = pi09032 & ~w18950;
assign w41094 = ~pi09848 & w18950;
assign w41095 = ~w41093 & ~w41094;
assign w41096 = pi09033 & ~w36416;
assign w41097 = w17922 & w18059;
assign w41098 = ~w41096 & ~w41097;
assign w41099 = pi09034 & ~w18950;
assign w41100 = w17311 & w18949;
assign w41101 = ~w41099 & ~w41100;
assign w41102 = pi09035 & ~w18950;
assign w41103 = ~pi02178 & w18950;
assign w41104 = ~w41102 & ~w41103;
assign w41105 = pi09036 & ~w18950;
assign w41106 = ~pi09954 & w18950;
assign w41107 = ~w41105 & ~w41106;
assign w41108 = pi09037 & ~w18950;
assign w41109 = ~pi02720 & w18950;
assign w41110 = ~w41108 & ~w41109;
assign w41111 = pi09038 & ~w18950;
assign w41112 = ~pi09962 & w18950;
assign w41113 = ~w41111 & ~w41112;
assign w41114 = pi09039 & ~w18722;
assign w41115 = ~pi09961 & w18722;
assign w41116 = ~w41114 & ~w41115;
assign w41117 = pi09040 & ~w18722;
assign w41118 = ~pi09848 & w18722;
assign w41119 = ~w41117 & ~w41118;
assign w41120 = pi09041 & ~w18722;
assign w41121 = ~pi02704 & w18722;
assign w41122 = ~w41120 & ~w41121;
assign w41123 = pi09042 & ~w18722;
assign w41124 = ~pi02178 & w18722;
assign w41125 = ~w41123 & ~w41124;
assign w41126 = pi09043 & ~w18722;
assign w41127 = ~pi09954 & w18722;
assign w41128 = ~w41126 & ~w41127;
assign w41129 = pi09044 & ~w18722;
assign w41130 = ~pi09962 & w18722;
assign w41131 = ~w41129 & ~w41130;
assign w41132 = pi09045 & ~w18736;
assign w41133 = ~pi09961 & w18736;
assign w41134 = ~w41132 & ~w41133;
assign w41135 = pi09046 & ~w18736;
assign w41136 = ~pi09848 & w18736;
assign w41137 = ~w41135 & ~w41136;
assign w41138 = pi09047 & ~w18736;
assign w41139 = ~pi02704 & w18736;
assign w41140 = ~w41138 & ~w41139;
assign w41141 = pi09048 & ~w18736;
assign w41142 = w18526 & w18861;
assign w41143 = ~w41141 & ~w41142;
assign w41144 = pi09049 & ~w18736;
assign w41145 = ~pi09954 & w18736;
assign w41146 = ~w41144 & ~w41145;
assign w41147 = pi09050 & ~w18736;
assign w41148 = w17128 & w18526;
assign w41149 = ~w41147 & ~w41148;
assign w41150 = pi09051 & ~w18736;
assign w41151 = ~pi09962 & w18736;
assign w41152 = ~w41150 & ~w41151;
assign w41153 = pi09052 & ~w18292;
assign w41154 = ~pi09961 & w18292;
assign w41155 = ~w41153 & ~w41154;
assign w41156 = pi09053 & ~w18292;
assign w41157 = ~pi09848 & w18292;
assign w41158 = ~w41156 & ~w41157;
assign w41159 = pi09054 & ~w18292;
assign w41160 = w17311 & w18291;
assign w41161 = ~w41159 & ~w41160;
assign w41162 = pi09055 & ~w18292;
assign w41163 = ~pi02178 & w18292;
assign w41164 = ~w41162 & ~w41163;
assign w41165 = pi09056 & ~w18292;
assign w41166 = ~pi09954 & w18292;
assign w41167 = ~w41165 & ~w41166;
assign w41168 = pi09057 & ~w18292;
assign w41169 = ~pi09962 & w18292;
assign w41170 = ~w41168 & ~w41169;
assign w41171 = pi09058 & ~w17412;
assign w41172 = w17411 & w19365;
assign w41173 = ~w41171 & ~w41172;
assign w41174 = pi09059 & ~w17412;
assign w41175 = ~pi09848 & w17412;
assign w41176 = ~w41174 & ~w41175;
assign w41177 = pi09060 & ~w17412;
assign w41178 = ~pi02704 & w17412;
assign w41179 = ~w41177 & ~w41178;
assign w41180 = pi09061 & ~w17412;
assign w41181 = ~pi02178 & w17412;
assign w41182 = ~w41180 & ~w41181;
assign w41183 = pi09062 & ~w17412;
assign w41184 = w17411 & w17513;
assign w41185 = ~w41183 & ~w41184;
assign w41186 = pi09063 & ~w17412;
assign w41187 = ~pi02720 & w17412;
assign w41188 = ~w41186 & ~w41187;
assign w41189 = pi09064 & ~w17412;
assign w41190 = ~pi09962 & w17412;
assign w41191 = ~w41189 & ~w41190;
assign w41192 = pi09065 & ~w17306;
assign w41193 = ~pi09961 & w17306;
assign w41194 = ~w41192 & ~w41193;
assign w41195 = pi09066 & ~w17306;
assign w41196 = ~pi09848 & w17306;
assign w41197 = ~w41195 & ~w41196;
assign w41198 = pi09067 & ~w17306;
assign w41199 = ~pi02704 & w17306;
assign w41200 = ~w41198 & ~w41199;
assign w41201 = pi09068 & ~w17306;
assign w41202 = ~pi02178 & w17306;
assign w41203 = ~w41201 & ~w41202;
assign w41204 = pi09069 & ~w17306;
assign w41205 = w17305 & w17513;
assign w41206 = ~w41204 & ~w41205;
assign w41207 = pi09070 & ~w17306;
assign w41208 = w17305 & w17439;
assign w41209 = ~w41207 & ~w41208;
assign w41210 = pi09071 & ~w21254;
assign w41211 = ~pi09961 & w21254;
assign w41212 = ~w41210 & ~w41211;
assign w41213 = pi09072 & ~w21254;
assign w41214 = ~pi09848 & w21254;
assign w41215 = ~w41213 & ~w41214;
assign w41216 = pi09073 & ~w21254;
assign w41217 = ~pi02704 & w21254;
assign w41218 = ~w41216 & ~w41217;
assign w41219 = pi09074 & ~w21254;
assign w41220 = ~pi02178 & w21254;
assign w41221 = ~w41219 & ~w41220;
assign w41222 = pi09075 & ~w21254;
assign w41223 = ~pi02720 & w21254;
assign w41224 = ~w41222 & ~w41223;
assign w41225 = pi09076 & ~w21254;
assign w41226 = ~pi09954 & w21254;
assign w41227 = ~w41225 & ~w41226;
assign w41228 = pi09077 & ~w21254;
assign w41229 = ~pi09962 & w21254;
assign w41230 = ~w41228 & ~w41229;
assign w41231 = pi09078 & ~w31030;
assign w41232 = ~pi09961 & w31030;
assign w41233 = ~w41231 & ~w41232;
assign w41234 = pi09079 & ~w31030;
assign w41235 = ~pi09848 & w31030;
assign w41236 = ~w41234 & ~w41235;
assign w41237 = pi09080 & ~w31030;
assign w41238 = ~pi02704 & w31030;
assign w41239 = ~w41237 & ~w41238;
assign w41240 = pi09081 & ~w31030;
assign w41241 = ~pi02178 & w31030;
assign w41242 = ~w41240 & ~w41241;
assign w41243 = pi09082 & ~w31030;
assign w41244 = ~pi09954 & w31030;
assign w41245 = ~w41243 & ~w41244;
assign w41246 = pi09083 & ~w31030;
assign w41247 = ~pi09962 & w31030;
assign w41248 = ~w41246 & ~w41247;
assign w41249 = pi09084 & ~w21250;
assign w41250 = ~pi09961 & w21250;
assign w41251 = ~w41249 & ~w41250;
assign w41252 = pi09085 & ~w21250;
assign w41253 = w17186 & w17686;
assign w41254 = ~w41252 & ~w41253;
assign w41255 = pi09086 & ~w21250;
assign w41256 = ~pi02704 & w21250;
assign w41257 = ~w41255 & ~w41256;
assign w41258 = pi09087 & ~w21250;
assign w41259 = ~pi02178 & w21250;
assign w41260 = ~w41258 & ~w41259;
assign w41261 = pi09088 & ~w21250;
assign w41262 = ~pi09954 & w21250;
assign w41263 = ~w41261 & ~w41262;
assign w41264 = pi09089 & ~w21250;
assign w41265 = ~pi02720 & w21250;
assign w41266 = ~w41264 & ~w41265;
assign w41267 = pi09090 & ~w21250;
assign w41268 = ~pi09962 & w21250;
assign w41269 = ~w41267 & ~w41268;
assign w41270 = pi09091 & ~w21399;
assign w41271 = ~pi09961 & w21399;
assign w41272 = ~w41270 & ~w41271;
assign w41273 = pi09092 & ~w21399;
assign w41274 = ~pi09848 & w21399;
assign w41275 = ~w41273 & ~w41274;
assign w41276 = pi09093 & ~w21399;
assign w41277 = ~pi02704 & w21399;
assign w41278 = ~w41276 & ~w41277;
assign w41279 = pi09094 & ~w21399;
assign w41280 = w17614 & w18861;
assign w41281 = ~w41279 & ~w41280;
assign w41282 = pi09095 & ~w21399;
assign w41283 = w17513 & w17614;
assign w41284 = ~w41282 & ~w41283;
assign w41285 = pi09096 & ~w21399;
assign w41286 = w17439 & w17614;
assign w41287 = ~w41285 & ~w41286;
assign w41288 = pi09097 & ~w21403;
assign w41289 = ~pi09961 & w21403;
assign w41290 = ~w41288 & ~w41289;
assign w41291 = pi09098 & ~w21403;
assign w41292 = ~pi09848 & w21403;
assign w41293 = ~w41291 & ~w41292;
assign w41294 = pi09099 & ~w21403;
assign w41295 = ~pi02704 & w21403;
assign w41296 = ~w41294 & ~w41295;
assign w41297 = pi09100 & ~w21403;
assign w41298 = ~pi02178 & w21403;
assign w41299 = ~w41297 & ~w41298;
assign w41300 = pi09101 & ~w21403;
assign w41301 = w17513 & w17526;
assign w41302 = ~w41300 & ~w41301;
assign w41303 = pi09102 & ~w21403;
assign w41304 = ~pi02720 & w21403;
assign w41305 = ~w41303 & ~w41304;
assign w41306 = pi09103 & ~w21403;
assign w41307 = ~pi09962 & w21403;
assign w41308 = ~w41306 & ~w41307;
assign w41309 = pi09104 & ~w21392;
assign w41310 = w17922 & w19365;
assign w41311 = ~w41309 & ~w41310;
assign w41312 = pi09105 & ~w21392;
assign w41313 = w17186 & w17922;
assign w41314 = ~w41312 & ~w41313;
assign w41315 = pi09106 & ~w21392;
assign w41316 = ~pi02704 & w21392;
assign w41317 = ~w41315 & ~w41316;
assign w41318 = pi09107 & ~w21392;
assign w41319 = w17922 & w18861;
assign w41320 = ~w41318 & ~w41319;
assign w41321 = pi09108 & ~w21392;
assign w41322 = w17513 & w17922;
assign w41323 = ~w41321 & ~w41322;
assign w41324 = pi09109 & ~w21392;
assign w41325 = w17439 & w17922;
assign w41326 = ~w41324 & ~w41325;
assign w41327 = pi09110 & ~w21374;
assign w41328 = ~pi09961 & w21374;
assign w41329 = ~w41327 & ~w41328;
assign w41330 = pi09111 & ~w21374;
assign w41331 = ~pi09848 & w21374;
assign w41332 = ~w41330 & ~w41331;
assign w41333 = pi09112 & ~w21374;
assign w41334 = ~pi02704 & w21374;
assign w41335 = ~w41333 & ~w41334;
assign w41336 = pi09113 & ~w21374;
assign w41337 = ~pi02178 & w21374;
assign w41338 = ~w41336 & ~w41337;
assign w41339 = pi09114 & ~w21374;
assign w41340 = ~pi09954 & w21374;
assign w41341 = ~w41339 & ~w41340;
assign w41342 = pi09115 & ~w21374;
assign w41343 = ~pi02720 & w21374;
assign w41344 = ~w41342 & ~w41343;
assign w41345 = pi09116 & ~w21374;
assign w41346 = ~pi09962 & w21374;
assign w41347 = ~w41345 & ~w41346;
assign w41348 = pi09117 & ~w21155;
assign w41349 = ~pi09961 & w21155;
assign w41350 = ~w41348 & ~w41349;
assign w41351 = pi09118 & ~w21155;
assign w41352 = ~pi09848 & w21155;
assign w41353 = ~w41351 & ~w41352;
assign w41354 = pi09119 & ~w21155;
assign w41355 = ~pi02704 & w21155;
assign w41356 = ~w41354 & ~w41355;
assign w41357 = pi09120 & ~w21155;
assign w41358 = ~pi02178 & w21155;
assign w41359 = ~w41357 & ~w41358;
assign w41360 = pi09121 & ~w21155;
assign w41361 = ~pi09954 & w21155;
assign w41362 = ~w41360 & ~w41361;
assign w41363 = pi09122 & ~w21155;
assign w41364 = ~pi09962 & w21155;
assign w41365 = ~w41363 & ~w41364;
assign w41366 = pi09123 & ~w20970;
assign w41367 = ~pi09961 & w20970;
assign w41368 = ~w41366 & ~w41367;
assign w41369 = pi09124 & ~w20970;
assign w41370 = ~pi09848 & w20970;
assign w41371 = ~w41369 & ~w41370;
assign w41372 = pi09125 & ~w20970;
assign w41373 = ~pi02704 & w20970;
assign w41374 = ~w41372 & ~w41373;
assign w41375 = pi09126 & ~w20970;
assign w41376 = ~pi02178 & w20970;
assign w41377 = ~w41375 & ~w41376;
assign w41378 = pi09127 & ~w20970;
assign w41379 = w17513 & w20720;
assign w41380 = ~w41378 & ~w41379;
assign w41381 = pi09128 & ~w20970;
assign w41382 = ~pi02720 & w20970;
assign w41383 = ~w41381 & ~w41382;
assign w41384 = pi09129 & ~w20970;
assign w41385 = w17439 & w20720;
assign w41386 = ~w41384 & ~w41385;
assign w41387 = pi09130 & ~w18632;
assign w41388 = ~pi09961 & w18632;
assign w41389 = ~w41387 & ~w41388;
assign w41390 = pi09131 & ~w18632;
assign w41391 = ~pi09848 & w18632;
assign w41392 = ~w41390 & ~w41391;
assign w41393 = pi09132 & ~w18632;
assign w41394 = ~pi02704 & w18632;
assign w41395 = ~w41393 & ~w41394;
assign w41396 = pi09133 & ~w18632;
assign w41397 = ~pi02178 & w18632;
assign w41398 = ~w41396 & ~w41397;
assign w41399 = pi09134 & ~w18632;
assign w41400 = ~pi09954 & w18632;
assign w41401 = ~w41399 & ~w41400;
assign w41402 = pi09135 & ~w18632;
assign w41403 = ~pi09962 & w18632;
assign w41404 = ~w41402 & ~w41403;
assign w41405 = pi09136 & ~w17335;
assign w41406 = w17334 & w19365;
assign w41407 = ~w41405 & ~w41406;
assign w41408 = pi09137 & ~w17335;
assign w41409 = w17186 & w17334;
assign w41410 = ~w41408 & ~w41409;
assign w41411 = pi09138 & ~w17335;
assign w41412 = ~pi02704 & w17335;
assign w41413 = ~w41411 & ~w41412;
assign w41414 = pi09139 & ~w17335;
assign w41415 = w17334 & w18861;
assign w41416 = ~w41414 & ~w41415;
assign w41417 = pi09140 & ~w17335;
assign w41418 = w17334 & w17513;
assign w41419 = ~w41417 & ~w41418;
assign w41420 = pi09141 & ~w17335;
assign w41421 = w17128 & w17334;
assign w41422 = ~w41420 & ~w41421;
assign w41423 = pi09142 & ~w17335;
assign w41424 = w17334 & w17439;
assign w41425 = ~w41423 & ~w41424;
assign w41426 = ~w16928 & w20775;
assign w41427 = pi09143 & ~w41426;
assign w41428 = ~pi09961 & w41426;
assign w41429 = ~w41427 & ~w41428;
assign w41430 = pi09144 & ~w41426;
assign w41431 = ~pi09848 & w41426;
assign w41432 = ~w41430 & ~w41431;
assign w41433 = pi09145 & ~w41426;
assign w41434 = ~pi02704 & w41426;
assign w41435 = ~w41433 & ~w41434;
assign w41436 = pi09146 & ~w41426;
assign w41437 = ~pi02178 & w41426;
assign w41438 = ~w41436 & ~w41437;
assign w41439 = pi09147 & ~w41426;
assign w41440 = ~pi09954 & w41426;
assign w41441 = ~w41439 & ~w41440;
assign w41442 = pi09148 & ~w41426;
assign w41443 = ~pi09962 & w41426;
assign w41444 = ~w41442 & ~w41443;
assign w41445 = pi09149 & ~w21337;
assign w41446 = ~pi09961 & w21337;
assign w41447 = ~w41445 & ~w41446;
assign w41448 = pi09150 & ~w21337;
assign w41449 = ~pi09848 & w21337;
assign w41450 = ~w41448 & ~w41449;
assign w41451 = pi09151 & ~w21337;
assign w41452 = ~pi02704 & w21337;
assign w41453 = ~w41451 & ~w41452;
assign w41454 = pi09152 & ~w21337;
assign w41455 = ~pi02178 & w21337;
assign w41456 = ~w41454 & ~w41455;
assign w41457 = pi09153 & ~w21337;
assign w41458 = ~pi09954 & w21337;
assign w41459 = ~w41457 & ~w41458;
assign w41460 = pi09154 & ~w21337;
assign w41461 = ~pi02720 & w21337;
assign w41462 = ~w41460 & ~w41461;
assign w41463 = pi09155 & ~w21337;
assign w41464 = ~pi09962 & w21337;
assign w41465 = ~w41463 & ~w41464;
assign w41466 = pi09156 & ~w21150;
assign w41467 = ~pi09961 & w21150;
assign w41468 = ~w41466 & ~w41467;
assign w41469 = pi09157 & ~w21150;
assign w41470 = w17186 & w20566;
assign w41471 = ~w41469 & ~w41470;
assign w41472 = pi09158 & ~w21150;
assign w41473 = w17311 & w20566;
assign w41474 = ~w41472 & ~w41473;
assign w41475 = pi09159 & ~w21150;
assign w41476 = ~pi02178 & w21150;
assign w41477 = ~w41475 & ~w41476;
assign w41478 = pi09160 & ~w21150;
assign w41479 = w17513 & w20566;
assign w41480 = ~w41478 & ~w41479;
assign w41481 = pi09161 & ~w21150;
assign w41482 = w17439 & w20566;
assign w41483 = ~w41481 & ~w41482;
assign w41484 = pi09162 & ~w21181;
assign w41485 = ~pi09961 & w21181;
assign w41486 = ~w41484 & ~w41485;
assign w41487 = pi09163 & ~w21181;
assign w41488 = ~pi09848 & w21181;
assign w41489 = ~w41487 & ~w41488;
assign w41490 = pi09164 & ~w21181;
assign w41491 = ~pi02704 & w21181;
assign w41492 = ~w41490 & ~w41491;
assign w41493 = pi09165 & ~w21181;
assign w41494 = ~pi02178 & w21181;
assign w41495 = ~w41493 & ~w41494;
assign w41496 = pi09166 & ~w21181;
assign w41497 = ~pi09954 & w21181;
assign w41498 = ~w41496 & ~w41497;
assign w41499 = pi09167 & ~w21181;
assign w41500 = ~pi02720 & w21181;
assign w41501 = ~w41499 & ~w41500;
assign w41502 = pi09168 & ~w21181;
assign w41503 = ~pi09962 & w21181;
assign w41504 = ~w41502 & ~w41503;
assign w41505 = pi09169 & ~w16932;
assign w41506 = ~pi09961 & w16932;
assign w41507 = ~w41505 & ~w41506;
assign w41508 = pi09170 & ~w16932;
assign w41509 = ~pi09848 & w16932;
assign w41510 = ~w41508 & ~w41509;
assign w41511 = pi09171 & ~w16932;
assign w41512 = ~pi02704 & w16932;
assign w41513 = ~w41511 & ~w41512;
assign w41514 = pi09172 & ~w16932;
assign w41515 = ~pi02178 & w16932;
assign w41516 = ~w41514 & ~w41515;
assign w41517 = pi09173 & ~w16932;
assign w41518 = ~pi09954 & w16932;
assign w41519 = ~w41517 & ~w41518;
assign w41520 = pi09174 & ~w16932;
assign w41521 = ~pi09962 & w16932;
assign w41522 = ~w41520 & ~w41521;
assign w41523 = ~w16928 & w18772;
assign w41524 = pi09175 & ~w41523;
assign w41525 = ~pi09961 & w41523;
assign w41526 = ~w41524 & ~w41525;
assign w41527 = pi09176 & ~w41523;
assign w41528 = ~pi09848 & w41523;
assign w41529 = ~w41527 & ~w41528;
assign w41530 = pi09177 & ~w41523;
assign w41531 = ~pi02178 & w41523;
assign w41532 = ~w41530 & ~w41531;
assign w41533 = pi09178 & ~w41523;
assign w41534 = w17513 & w18772;
assign w41535 = ~w41533 & ~w41534;
assign w41536 = pi09179 & ~w41523;
assign w41537 = ~pi02720 & w41523;
assign w41538 = ~w41536 & ~w41537;
assign w41539 = pi09180 & ~w41523;
assign w41540 = ~pi09962 & w41523;
assign w41541 = ~w41539 & ~w41540;
assign w41542 = pi09181 & ~w41523;
assign w41543 = ~pi09812 & w41523;
assign w41544 = ~w41542 & ~w41543;
assign w41545 = pi09182 & ~w21303;
assign w41546 = ~pi09961 & w21303;
assign w41547 = ~w41545 & ~w41546;
assign w41548 = pi09183 & ~w21303;
assign w41549 = ~pi09848 & w21303;
assign w41550 = ~w41548 & ~w41549;
assign w41551 = pi09184 & ~w21303;
assign w41552 = w17311 & w18300;
assign w41553 = ~w41551 & ~w41552;
assign w41554 = pi09185 & ~w21303;
assign w41555 = ~pi02178 & w21303;
assign w41556 = ~w41554 & ~w41555;
assign w41557 = pi09186 & ~w21303;
assign w41558 = ~pi09954 & w21303;
assign w41559 = ~w41557 & ~w41558;
assign w41560 = pi09187 & ~w21303;
assign w41561 = ~pi09962 & w21303;
assign w41562 = ~w41560 & ~w41561;
assign w41563 = pi09188 & ~w21322;
assign w41564 = ~pi09961 & w21322;
assign w41565 = ~w41563 & ~w41564;
assign w41566 = pi09189 & ~w21322;
assign w41567 = w17186 & w17907;
assign w41568 = ~w41566 & ~w41567;
assign w41569 = pi09190 & ~w21322;
assign w41570 = ~pi02704 & w21322;
assign w41571 = ~w41569 & ~w41570;
assign w41572 = pi09191 & ~w21322;
assign w41573 = w17907 & w18861;
assign w41574 = ~w41572 & ~w41573;
assign w41575 = pi09192 & ~w21322;
assign w41576 = w17513 & w17907;
assign w41577 = ~w41575 & ~w41576;
assign w41578 = pi09193 & ~w21322;
assign w41579 = ~pi02720 & w21322;
assign w41580 = ~w41578 & ~w41579;
assign w41581 = pi09194 & ~w21322;
assign w41582 = w17439 & w17907;
assign w41583 = ~w41581 & ~w41582;
assign w41584 = pi09195 & ~w20932;
assign w41585 = ~pi09848 & w20932;
assign w41586 = ~w41584 & ~w41585;
assign w41587 = pi09196 & ~w20932;
assign w41588 = w17193 & w17754;
assign w41589 = ~w41587 & ~w41588;
assign w41590 = pi09197 & ~w20932;
assign w41591 = ~pi02178 & w20932;
assign w41592 = ~w41590 & ~w41591;
assign w41593 = pi09198 & ~w20932;
assign w41594 = ~pi09961 & w20932;
assign w41595 = ~w41593 & ~w41594;
assign w41596 = pi09199 & ~w20932;
assign w41597 = ~pi02720 & w20932;
assign w41598 = ~w41596 & ~w41597;
assign w41599 = pi09200 & ~w20932;
assign w41600 = ~pi09962 & w20932;
assign w41601 = ~w41599 & ~w41600;
assign w41602 = pi09201 & ~w29987;
assign w41603 = w17428 & w19365;
assign w41604 = ~w41602 & ~w41603;
assign w41605 = pi09202 & ~w29987;
assign w41606 = ~pi09848 & w29987;
assign w41607 = ~w41605 & ~w41606;
assign w41608 = pi09203 & ~w29987;
assign w41609 = ~pi02704 & w29987;
assign w41610 = ~w41608 & ~w41609;
assign w41611 = pi09204 & ~w29987;
assign w41612 = w17428 & w18861;
assign w41613 = ~w41611 & ~w41612;
assign w41614 = pi09205 & ~w29987;
assign w41615 = ~pi09954 & w29987;
assign w41616 = ~w41614 & ~w41615;
assign w41617 = pi09206 & ~w29987;
assign w41618 = ~pi02720 & w29987;
assign w41619 = ~w41617 & ~w41618;
assign w41620 = pi09207 & ~w29987;
assign w41621 = ~pi09962 & w29987;
assign w41622 = ~w41620 & ~w41621;
assign w41623 = pi09208 & ~w36686;
assign w41624 = ~pi09961 & w36686;
assign w41625 = ~w41623 & ~w41624;
assign w41626 = pi09209 & ~w36686;
assign w41627 = ~pi09848 & w36686;
assign w41628 = ~w41626 & ~w41627;
assign w41629 = pi09210 & ~w36686;
assign w41630 = ~pi02704 & w36686;
assign w41631 = ~w41629 & ~w41630;
assign w41632 = pi09211 & ~w36686;
assign w41633 = ~pi02178 & w36686;
assign w41634 = ~w41632 & ~w41633;
assign w41635 = pi09212 & ~w36686;
assign w41636 = ~pi09954 & w36686;
assign w41637 = ~w41635 & ~w41636;
assign w41638 = pi09213 & ~w36686;
assign w41639 = ~pi09962 & w36686;
assign w41640 = ~w41638 & ~w41639;
assign w41641 = pi09214 & ~w17939;
assign w41642 = ~pi09961 & w17939;
assign w41643 = ~w41641 & ~w41642;
assign w41644 = pi09215 & ~w17939;
assign w41645 = ~pi09848 & w17939;
assign w41646 = ~w41644 & ~w41645;
assign w41647 = pi09216 & ~w17939;
assign w41648 = ~pi02704 & w17939;
assign w41649 = ~w41647 & ~w41648;
assign w41650 = pi09217 & ~w17939;
assign w41651 = ~pi02178 & w17939;
assign w41652 = ~w41650 & ~w41651;
assign w41653 = pi09218 & ~w17939;
assign w41654 = ~pi09954 & w17939;
assign w41655 = ~w41653 & ~w41654;
assign w41656 = pi09219 & ~w17939;
assign w41657 = ~pi02720 & w17939;
assign w41658 = ~w41656 & ~w41657;
assign w41659 = pi09220 & ~w17939;
assign w41660 = ~pi09962 & w17939;
assign w41661 = ~w41659 & ~w41660;
assign w41662 = pi09221 & ~w20215;
assign w41663 = ~pi09961 & w20215;
assign w41664 = ~w41662 & ~w41663;
assign w41665 = pi09222 & ~w20215;
assign w41666 = ~pi09848 & w20215;
assign w41667 = ~w41665 & ~w41666;
assign w41668 = pi09223 & ~w20215;
assign w41669 = ~pi02704 & w20215;
assign w41670 = ~w41668 & ~w41669;
assign w41671 = pi09224 & ~w20215;
assign w41672 = ~pi02178 & w20215;
assign w41673 = ~w41671 & ~w41672;
assign w41674 = pi09225 & ~w20215;
assign w41675 = ~pi09954 & w20215;
assign w41676 = ~w41674 & ~w41675;
assign w41677 = pi09226 & ~w20215;
assign w41678 = ~pi09962 & w20215;
assign w41679 = ~w41677 & ~w41678;
assign w41680 = pi09227 & ~w22185;
assign w41681 = ~pi09961 & w22185;
assign w41682 = ~w41680 & ~w41681;
assign w41683 = pi09228 & ~w22185;
assign w41684 = ~pi09848 & w22185;
assign w41685 = ~w41683 & ~w41684;
assign w41686 = pi09229 & ~w22185;
assign w41687 = ~pi02704 & w22185;
assign w41688 = ~w41686 & ~w41687;
assign w41689 = pi09230 & ~w22185;
assign w41690 = ~pi02178 & w22185;
assign w41691 = ~w41689 & ~w41690;
assign w41692 = pi09231 & ~w22185;
assign w41693 = ~pi09954 & w22185;
assign w41694 = ~w41692 & ~w41693;
assign w41695 = pi09232 & ~w22185;
assign w41696 = ~pi02720 & w22185;
assign w41697 = ~w41695 & ~w41696;
assign w41698 = pi09233 & ~w22185;
assign w41699 = ~pi09962 & w22185;
assign w41700 = ~w41698 & ~w41699;
assign w41701 = pi09234 & ~w18062;
assign w41702 = w17098 & w19365;
assign w41703 = ~w41701 & ~w41702;
assign w41704 = pi09235 & ~w18062;
assign w41705 = ~pi09848 & w18062;
assign w41706 = ~w41704 & ~w41705;
assign w41707 = pi09236 & ~w18062;
assign w41708 = ~pi02704 & w18062;
assign w41709 = ~w41707 & ~w41708;
assign w41710 = pi09237 & ~w18062;
assign w41711 = ~pi02178 & w18062;
assign w41712 = ~w41710 & ~w41711;
assign w41713 = pi09238 & ~w18062;
assign w41714 = ~pi09954 & w18062;
assign w41715 = ~w41713 & ~w41714;
assign w41716 = pi09239 & ~w18062;
assign w41717 = ~pi09962 & w18062;
assign w41718 = ~w41716 & ~w41717;
assign w41719 = pi09240 & ~w20706;
assign w41720 = ~pi09961 & w20706;
assign w41721 = ~w41719 & ~w41720;
assign w41722 = pi09241 & ~w20706;
assign w41723 = ~pi09848 & w20706;
assign w41724 = ~w41722 & ~w41723;
assign w41725 = pi09242 & ~w17173;
assign w41726 = w17172 & w17193;
assign w41727 = ~w41725 & ~w41726;
assign w41728 = pi09243 & ~w20706;
assign w41729 = ~pi02704 & w20706;
assign w41730 = ~w41728 & ~w41729;
assign w41731 = pi09244 & ~w20706;
assign w41732 = ~pi02178 & w20706;
assign w41733 = ~w41731 & ~w41732;
assign w41734 = pi09245 & ~w20706;
assign w41735 = ~pi09954 & w20706;
assign w41736 = ~w41734 & ~w41735;
assign w41737 = pi09246 & ~w20706;
assign w41738 = ~pi02720 & w20706;
assign w41739 = ~w41737 & ~w41738;
assign w41740 = pi09247 & ~w20706;
assign w41741 = w17439 & w20244;
assign w41742 = ~w41740 & ~w41741;
assign w41743 = pi09248 & ~w20366;
assign w41744 = ~pi09961 & w20366;
assign w41745 = ~w41743 & ~w41744;
assign w41746 = pi09249 & ~w20366;
assign w41747 = ~pi09848 & w20366;
assign w41748 = ~w41746 & ~w41747;
assign w41749 = pi09250 & ~w20366;
assign w41750 = ~pi02704 & w20366;
assign w41751 = ~w41749 & ~w41750;
assign w41752 = pi09251 & ~w20366;
assign w41753 = ~pi02178 & w20366;
assign w41754 = ~w41752 & ~w41753;
assign w41755 = pi09252 & ~w20366;
assign w41756 = ~pi09954 & w20366;
assign w41757 = ~w41755 & ~w41756;
assign w41758 = pi09253 & ~w20366;
assign w41759 = ~pi09962 & w20366;
assign w41760 = ~w41758 & ~w41759;
assign w41761 = pi09254 & ~w18753;
assign w41762 = ~pi09961 & w18753;
assign w41763 = ~w41761 & ~w41762;
assign w41764 = pi09255 & ~w18753;
assign w41765 = ~pi09848 & w18753;
assign w41766 = ~w41764 & ~w41765;
assign w41767 = pi09256 & ~w18753;
assign w41768 = ~pi02704 & w18753;
assign w41769 = ~w41767 & ~w41768;
assign w41770 = pi09257 & ~w18753;
assign w41771 = ~pi02178 & w18753;
assign w41772 = ~w41770 & ~w41771;
assign w41773 = pi09258 & ~w18753;
assign w41774 = ~pi09954 & w18753;
assign w41775 = ~w41773 & ~w41774;
assign w41776 = pi09259 & ~w18753;
assign w41777 = w17128 & w18662;
assign w41778 = ~w41776 & ~w41777;
assign w41779 = pi09260 & ~w18753;
assign w41780 = ~pi09962 & w18753;
assign w41781 = ~w41779 & ~w41780;
assign w41782 = pi09261 & ~w20370;
assign w41783 = w18617 & w19365;
assign w41784 = ~w41782 & ~w41783;
assign w41785 = pi09262 & ~w20370;
assign w41786 = ~pi09848 & w20370;
assign w41787 = ~w41785 & ~w41786;
assign w41788 = pi09263 & ~w20370;
assign w41789 = ~pi02704 & w20370;
assign w41790 = ~w41788 & ~w41789;
assign w41791 = pi09264 & ~w20370;
assign w41792 = ~pi02178 & w20370;
assign w41793 = ~w41791 & ~w41792;
assign w41794 = pi09265 & ~w20370;
assign w41795 = ~pi09954 & w20370;
assign w41796 = ~w41794 & ~w41795;
assign w41797 = pi09266 & ~w20370;
assign w41798 = ~pi09962 & w20370;
assign w41799 = ~w41797 & ~w41798;
assign w41800 = pi09267 & ~w18555;
assign w41801 = ~pi09961 & w18555;
assign w41802 = ~w41800 & ~w41801;
assign w41803 = pi09268 & ~w18555;
assign w41804 = ~pi09848 & w18555;
assign w41805 = ~w41803 & ~w41804;
assign w41806 = pi09269 & ~w18555;
assign w41807 = ~pi02704 & w18555;
assign w41808 = ~w41806 & ~w41807;
assign w41809 = pi09270 & ~w18555;
assign w41810 = ~pi02178 & w18555;
assign w41811 = ~w41809 & ~w41810;
assign w41812 = pi09271 & ~w18555;
assign w41813 = ~pi09954 & w18555;
assign w41814 = ~w41812 & ~w41813;
assign w41815 = pi09272 & ~w18555;
assign w41816 = ~pi02720 & w18555;
assign w41817 = ~w41815 & ~w41816;
assign w41818 = pi09273 & ~w18555;
assign w41819 = ~pi09962 & w18555;
assign w41820 = ~w41818 & ~w41819;
assign w41821 = pi09274 & ~w18105;
assign w41822 = ~pi09961 & w18105;
assign w41823 = ~w41821 & ~w41822;
assign w41824 = pi09275 & ~w18105;
assign w41825 = ~pi09848 & w18105;
assign w41826 = ~w41824 & ~w41825;
assign w41827 = pi09276 & ~w18105;
assign w41828 = ~pi02704 & w18105;
assign w41829 = ~w41827 & ~w41828;
assign w41830 = pi09277 & ~w18105;
assign w41831 = ~pi02178 & w18105;
assign w41832 = ~w41830 & ~w41831;
assign w41833 = pi09278 & ~w18105;
assign w41834 = ~pi02720 & w18105;
assign w41835 = ~w41833 & ~w41834;
assign w41836 = pi09279 & ~w18105;
assign w41837 = ~pi09962 & w18105;
assign w41838 = ~w41836 & ~w41837;
assign w41839 = pi09280 & ~w20281;
assign w41840 = ~pi09961 & w20281;
assign w41841 = ~w41839 & ~w41840;
assign w41842 = pi09281 & ~w20281;
assign w41843 = ~pi09848 & w20281;
assign w41844 = ~w41842 & ~w41843;
assign w41845 = pi09282 & ~w20281;
assign w41846 = w17311 & w18454;
assign w41847 = ~w41845 & ~w41846;
assign w41848 = pi09283 & ~w20281;
assign w41849 = ~pi02178 & w20281;
assign w41850 = ~w41848 & ~w41849;
assign w41851 = pi09284 & ~w20281;
assign w41852 = ~pi09954 & w20281;
assign w41853 = ~w41851 & ~w41852;
assign w41854 = pi09285 & ~w20281;
assign w41855 = ~pi02720 & w20281;
assign w41856 = ~w41854 & ~w41855;
assign w41857 = pi09286 & ~w20281;
assign w41858 = ~pi09962 & w20281;
assign w41859 = ~w41857 & ~w41858;
assign w41860 = pi09287 & ~w17711;
assign w41861 = w17710 & w19365;
assign w41862 = ~w41860 & ~w41861;
assign w41863 = pi09288 & ~w17711;
assign w41864 = ~pi09848 & w17711;
assign w41865 = ~w41863 & ~w41864;
assign w41866 = pi09289 & ~w17711;
assign w41867 = ~pi02704 & w17711;
assign w41868 = ~w41866 & ~w41867;
assign w41869 = pi09290 & ~w17711;
assign w41870 = ~pi02178 & w17711;
assign w41871 = ~w41869 & ~w41870;
assign w41872 = pi09291 & ~w17711;
assign w41873 = ~pi09954 & w17711;
assign w41874 = ~w41872 & ~w41873;
assign w41875 = pi09292 & ~w17711;
assign w41876 = ~pi09962 & w17711;
assign w41877 = ~w41875 & ~w41876;
assign w41878 = pi09293 & ~w18469;
assign w41879 = ~pi09961 & w18469;
assign w41880 = ~w41878 & ~w41879;
assign w41881 = pi09294 & ~w18469;
assign w41882 = ~pi09848 & w18469;
assign w41883 = ~w41881 & ~w41882;
assign w41884 = pi09295 & ~w18469;
assign w41885 = ~pi02704 & w18469;
assign w41886 = ~w41884 & ~w41885;
assign w41887 = pi09296 & ~w18469;
assign w41888 = w18468 & w18861;
assign w41889 = ~w41887 & ~w41888;
assign w41890 = pi09297 & ~w18469;
assign w41891 = ~pi09954 & w18469;
assign w41892 = ~w41890 & ~w41891;
assign w41893 = pi09298 & ~w18469;
assign w41894 = ~pi02720 & w18469;
assign w41895 = ~w41893 & ~w41894;
assign w41896 = pi09299 & ~w18469;
assign w41897 = ~pi09962 & w18469;
assign w41898 = ~w41896 & ~w41897;
assign w41899 = pi09300 & ~w17719;
assign w41900 = ~pi09961 & w17719;
assign w41901 = ~w41899 & ~w41900;
assign w41902 = pi09301 & ~w17719;
assign w41903 = ~pi09848 & w17719;
assign w41904 = ~w41902 & ~w41903;
assign w41905 = pi09302 & ~w17719;
assign w41906 = ~pi02704 & w17719;
assign w41907 = ~w41905 & ~w41906;
assign w41908 = pi09303 & ~w17719;
assign w41909 = ~pi02178 & w17719;
assign w41910 = ~w41908 & ~w41909;
assign w41911 = pi09304 & ~w17719;
assign w41912 = ~pi09954 & w17719;
assign w41913 = ~w41911 & ~w41912;
assign w41914 = pi09305 & ~w17719;
assign w41915 = ~pi09962 & w17719;
assign w41916 = ~w41914 & ~w41915;
assign w41917 = pi09306 & ~w17632;
assign w41918 = ~pi09961 & w17632;
assign w41919 = ~w41917 & ~w41918;
assign w41920 = pi09307 & ~w17632;
assign w41921 = ~pi09848 & w17632;
assign w41922 = ~w41920 & ~w41921;
assign w41923 = pi09308 & ~w17632;
assign w41924 = ~pi02704 & w17632;
assign w41925 = ~w41923 & ~w41924;
assign w41926 = pi09309 & ~w17632;
assign w41927 = ~pi02178 & w17632;
assign w41928 = ~w41926 & ~w41927;
assign w41929 = pi09310 & ~w17632;
assign w41930 = ~pi09954 & w17632;
assign w41931 = ~w41929 & ~w41930;
assign w41932 = pi09311 & ~w17632;
assign w41933 = ~pi02720 & w17632;
assign w41934 = ~w41932 & ~w41933;
assign w41935 = pi09312 & ~w17632;
assign w41936 = ~pi09962 & w17632;
assign w41937 = ~w41935 & ~w41936;
assign w41938 = pi09313 & ~w17417;
assign w41939 = ~pi09961 & w17417;
assign w41940 = ~w41938 & ~w41939;
assign w41941 = pi09314 & ~w17417;
assign w41942 = ~pi09848 & w17417;
assign w41943 = ~w41941 & ~w41942;
assign w41944 = pi09315 & ~w17417;
assign w41945 = ~pi02704 & w17417;
assign w41946 = ~w41944 & ~w41945;
assign w41947 = pi09316 & ~w17417;
assign w41948 = ~pi02178 & w17417;
assign w41949 = ~w41947 & ~w41948;
assign w41950 = pi09317 & ~w17417;
assign w41951 = ~pi09954 & w17417;
assign w41952 = ~w41950 & ~w41951;
assign w41953 = pi09318 & ~w17417;
assign w41954 = w17416 & w17439;
assign w41955 = ~w41953 & ~w41954;
assign w41956 = pi09319 & ~w17330;
assign w41957 = ~pi09961 & w17330;
assign w41958 = ~w41956 & ~w41957;
assign w41959 = pi09320 & ~w17330;
assign w41960 = ~pi09848 & w17330;
assign w41961 = ~w41959 & ~w41960;
assign w41962 = pi09321 & ~w17330;
assign w41963 = ~pi02704 & w17330;
assign w41964 = ~w41962 & ~w41963;
assign w41965 = pi09322 & ~w17330;
assign w41966 = ~pi02178 & w17330;
assign w41967 = ~w41965 & ~w41966;
assign w41968 = pi09323 & ~w17330;
assign w41969 = ~pi09954 & w17330;
assign w41970 = ~w41968 & ~w41969;
assign w41971 = pi09324 & ~w17330;
assign w41972 = w17128 & w17314;
assign w41973 = ~w41971 & ~w41972;
assign w41974 = pi09325 & ~w17330;
assign w41975 = ~pi09962 & w17330;
assign w41976 = ~w41974 & ~w41975;
assign w41977 = pi09326 & ~w17126;
assign w41978 = ~pi09961 & w17126;
assign w41979 = ~w41977 & ~w41978;
assign w41980 = pi09327 & ~w17126;
assign w41981 = ~pi09848 & w17126;
assign w41982 = ~w41980 & ~w41981;
assign w41983 = pi09328 & ~w17126;
assign w41984 = w17125 & w17311;
assign w41985 = ~w41983 & ~w41984;
assign w41986 = pi09329 & ~w17126;
assign w41987 = ~pi02178 & w17126;
assign w41988 = ~w41986 & ~w41987;
assign w41989 = pi09330 & ~w17126;
assign w41990 = ~pi09954 & w17126;
assign w41991 = ~w41989 & ~w41990;
assign w41992 = pi09331 & ~w17126;
assign w41993 = ~pi09962 & w17126;
assign w41994 = ~w41992 & ~w41993;
assign w41995 = pi09332 & ~w17240;
assign w41996 = ~pi09961 & w17240;
assign w41997 = ~w41995 & ~w41996;
assign w41998 = pi09333 & ~w17240;
assign w41999 = w17186 & w17239;
assign w42000 = ~w41998 & ~w41999;
assign w42001 = pi09334 & ~w17240;
assign w42002 = ~pi02704 & w17240;
assign w42003 = ~w42001 & ~w42002;
assign w42004 = pi09335 & ~w17240;
assign w42005 = ~pi02178 & w17240;
assign w42006 = ~w42004 & ~w42005;
assign w42007 = pi09336 & ~w17240;
assign w42008 = ~pi09954 & w17240;
assign w42009 = ~w42007 & ~w42008;
assign w42010 = pi09337 & ~w17240;
assign w42011 = ~pi02720 & w17240;
assign w42012 = ~w42010 & ~w42011;
assign w42013 = pi09338 & ~w17240;
assign w42014 = ~pi09962 & w17240;
assign w42015 = ~w42013 & ~w42014;
assign w42016 = pi09339 & ~w17168;
assign w42017 = ~pi09961 & w17168;
assign w42018 = ~w42016 & ~w42017;
assign w42019 = pi09340 & ~w17168;
assign w42020 = ~pi09848 & w17168;
assign w42021 = ~w42019 & ~w42020;
assign w42022 = pi09341 & ~w17168;
assign w42023 = ~pi02704 & w17168;
assign w42024 = ~w42022 & ~w42023;
assign w42025 = pi09342 & ~w17168;
assign w42026 = w17167 & w18861;
assign w42027 = ~w42025 & ~w42026;
assign w42028 = pi09343 & ~w17168;
assign w42029 = ~pi09954 & w17168;
assign w42030 = ~w42028 & ~w42029;
assign w42031 = pi09344 & ~w17168;
assign w42032 = ~pi09962 & w17168;
assign w42033 = ~w42031 & ~w42032;
assign w42034 = ~w16928 & w17205;
assign w42035 = pi09345 & ~w42034;
assign w42036 = ~pi09961 & w42034;
assign w42037 = ~w42035 & ~w42036;
assign w42038 = pi09346 & ~w42034;
assign w42039 = w17186 & w17205;
assign w42040 = ~w42038 & ~w42039;
assign w42041 = pi09347 & ~w36920;
assign w42042 = ~pi02716 & w36920;
assign w42043 = ~w42041 & ~w42042;
assign w42044 = pi09348 & ~w42034;
assign w42045 = w17205 & w17311;
assign w42046 = ~w42044 & ~w42045;
assign w42047 = pi09349 & ~w42034;
assign w42048 = ~pi02178 & w42034;
assign w42049 = ~w42047 & ~w42048;
assign w42050 = pi09350 & ~w42034;
assign w42051 = ~pi09954 & w42034;
assign w42052 = ~w42050 & ~w42051;
assign w42053 = pi09351 & ~w42034;
assign w42054 = ~pi02720 & w42034;
assign w42055 = ~w42053 & ~w42054;
assign w42056 = pi09352 & ~w42034;
assign w42057 = ~pi09962 & w42034;
assign w42058 = ~w42056 & ~w42057;
assign w42059 = pi09353 & ~w17367;
assign w42060 = w17366 & w19365;
assign w42061 = ~w42059 & ~w42060;
assign w42062 = pi09354 & ~w17367;
assign w42063 = w17186 & w17366;
assign w42064 = ~w42062 & ~w42063;
assign w42065 = pi09355 & ~w17367;
assign w42066 = ~pi02704 & w17367;
assign w42067 = ~w42065 & ~w42066;
assign w42068 = pi09356 & ~w17367;
assign w42069 = ~pi02178 & w17367;
assign w42070 = ~w42068 & ~w42069;
assign w42071 = pi09357 & ~w17367;
assign w42072 = ~pi09954 & w17367;
assign w42073 = ~w42071 & ~w42072;
assign w42074 = pi09358 & ~w17367;
assign w42075 = ~pi09962 & w17367;
assign w42076 = ~w42074 & ~w42075;
assign w42077 = pi09359 & ~w17201;
assign w42078 = ~pi09961 & w17201;
assign w42079 = ~w42077 & ~w42078;
assign w42080 = pi09360 & ~w17201;
assign w42081 = w17186 & w17200;
assign w42082 = ~w42080 & ~w42081;
assign w42083 = pi09361 & ~w17201;
assign w42084 = ~pi02704 & w17201;
assign w42085 = ~w42083 & ~w42084;
assign w42086 = pi09362 & ~w17201;
assign w42087 = ~pi02178 & w17201;
assign w42088 = ~w42086 & ~w42087;
assign w42089 = pi09363 & ~w17201;
assign w42090 = ~pi09954 & w17201;
assign w42091 = ~w42089 & ~w42090;
assign w42092 = pi09364 & ~w17201;
assign w42093 = ~pi02720 & w17201;
assign w42094 = ~w42092 & ~w42093;
assign w42095 = pi09365 & ~w17201;
assign w42096 = ~pi09962 & w17201;
assign w42097 = ~w42095 & ~w42096;
assign w42098 = pi09366 & ~w17173;
assign w42099 = ~pi09961 & w17173;
assign w42100 = ~w42098 & ~w42099;
assign w42101 = pi09367 & ~w17173;
assign w42102 = ~pi09848 & w17173;
assign w42103 = ~w42101 & ~w42102;
assign w42104 = pi09368 & ~w17173;
assign w42105 = ~pi02704 & w17173;
assign w42106 = ~w42104 & ~w42105;
assign w42107 = pi09369 & ~w17173;
assign w42108 = ~pi02178 & w17173;
assign w42109 = ~w42107 & ~w42108;
assign w42110 = pi09370 & ~w17173;
assign w42111 = w17172 & w17513;
assign w42112 = ~w42110 & ~w42111;
assign w42113 = pi09371 & ~w17173;
assign w42114 = ~pi09962 & w17173;
assign w42115 = ~w42113 & ~w42114;
assign w42116 = pi09372 & ~w17024;
assign w42117 = ~pi09961 & w17024;
assign w42118 = ~w42116 & ~w42117;
assign w42119 = pi09373 & ~w17024;
assign w42120 = ~pi09848 & w17024;
assign w42121 = ~w42119 & ~w42120;
assign w42122 = pi09374 & ~w17024;
assign w42123 = ~pi02704 & w17024;
assign w42124 = ~w42122 & ~w42123;
assign w42125 = pi09375 & ~w17024;
assign w42126 = ~pi02178 & w17024;
assign w42127 = ~w42125 & ~w42126;
assign w42128 = pi09376 & ~w17024;
assign w42129 = ~pi09954 & w17024;
assign w42130 = ~w42128 & ~w42129;
assign w42131 = pi09377 & ~w17024;
assign w42132 = ~pi02720 & w17024;
assign w42133 = ~w42131 & ~w42132;
assign w42134 = pi09378 & ~w17024;
assign w42135 = ~pi09962 & w17024;
assign w42136 = ~w42134 & ~w42135;
assign w42137 = pi09379 & ~w20919;
assign w42138 = ~pi09961 & w20919;
assign w42139 = ~w42137 & ~w42138;
assign w42140 = pi09380 & ~w20919;
assign w42141 = ~pi09848 & w20919;
assign w42142 = ~w42140 & ~w42141;
assign w42143 = pi09381 & ~w20919;
assign w42144 = ~pi02704 & w20919;
assign w42145 = ~w42143 & ~w42144;
assign w42146 = pi09382 & ~w20919;
assign w42147 = ~pi02178 & w20919;
assign w42148 = ~w42146 & ~w42147;
assign w42149 = pi09383 & ~w20919;
assign w42150 = ~pi09954 & w20919;
assign w42151 = ~w42149 & ~w42150;
assign w42152 = pi09384 & ~w20919;
assign w42153 = ~pi09962 & w20919;
assign w42154 = ~w42152 & ~w42153;
assign w42155 = pi09385 & ~w20821;
assign w42156 = w17479 & w19365;
assign w42157 = ~w42155 & ~w42156;
assign w42158 = pi09386 & ~w20821;
assign w42159 = w17186 & w17479;
assign w42160 = ~w42158 & ~w42159;
assign w42161 = pi09387 & ~w20821;
assign w42162 = w17311 & w17479;
assign w42163 = ~w42161 & ~w42162;
assign w42164 = pi09388 & ~w20821;
assign w42165 = w17479 & w18861;
assign w42166 = ~w42164 & ~w42165;
assign w42167 = pi09389 & ~w20821;
assign w42168 = w17479 & w17513;
assign w42169 = ~w42167 & ~w42168;
assign w42170 = pi09390 & ~w20821;
assign w42171 = w17128 & w17479;
assign w42172 = ~w42170 & ~w42171;
assign w42173 = pi09391 & ~w20821;
assign w42174 = w17439 & w17479;
assign w42175 = ~w42173 & ~w42174;
assign w42176 = pi09392 & ~w21311;
assign w42177 = w17398 & w19365;
assign w42178 = ~w42176 & ~w42177;
assign w42179 = pi09393 & ~w21311;
assign w42180 = ~pi09848 & w21311;
assign w42181 = ~w42179 & ~w42180;
assign w42182 = pi09394 & ~w21311;
assign w42183 = ~pi02704 & w21311;
assign w42184 = ~w42182 & ~w42183;
assign w42185 = pi09395 & ~w21311;
assign w42186 = ~pi02178 & w21311;
assign w42187 = ~w42185 & ~w42186;
assign w42188 = pi09396 & ~w21311;
assign w42189 = ~pi09954 & w21311;
assign w42190 = ~w42188 & ~w42189;
assign w42191 = pi09397 & ~w21311;
assign w42192 = ~pi09962 & w21311;
assign w42193 = ~w42191 & ~w42192;
assign w42194 = pi09398 & ~w24243;
assign w42195 = ~pi09961 & w24243;
assign w42196 = ~w42194 & ~w42195;
assign w42197 = pi09399 & ~w24243;
assign w42198 = ~pi09848 & w24243;
assign w42199 = ~w42197 & ~w42198;
assign w42200 = pi09400 & ~w38467;
assign w42201 = ~pi02703 & w38467;
assign w42202 = ~w42200 & ~w42201;
assign w42203 = pi09401 & ~w24243;
assign w42204 = w17114 & w17311;
assign w42205 = ~w42203 & ~w42204;
assign w42206 = pi09402 & ~w24243;
assign w42207 = ~pi02178 & w24243;
assign w42208 = ~w42206 & ~w42207;
assign w42209 = pi09403 & ~w24243;
assign w42210 = ~pi09954 & w24243;
assign w42211 = ~w42209 & ~w42210;
assign w42212 = pi09404 & ~w24243;
assign w42213 = ~pi02720 & w24243;
assign w42214 = ~w42212 & ~w42213;
assign w42215 = pi09405 & ~w24243;
assign w42216 = ~pi09962 & w24243;
assign w42217 = ~w42215 & ~w42216;
assign w42218 = pi09406 & ~w20875;
assign w42219 = ~pi09961 & w20875;
assign w42220 = ~w42218 & ~w42219;
assign w42221 = pi09407 & ~w20875;
assign w42222 = ~pi09848 & w20875;
assign w42223 = ~w42221 & ~w42222;
assign w42224 = pi09408 & ~w20875;
assign w42225 = ~pi02704 & w20875;
assign w42226 = ~w42224 & ~w42225;
assign w42227 = pi09409 & ~w20875;
assign w42228 = w17249 & w18861;
assign w42229 = ~w42227 & ~w42228;
assign w42230 = pi09410 & ~w20875;
assign w42231 = ~pi09954 & w20875;
assign w42232 = ~w42230 & ~w42231;
assign w42233 = pi09411 & ~w20875;
assign w42234 = ~pi09962 & w20875;
assign w42235 = ~w42233 & ~w42234;
assign w42236 = pi09412 & ~w17048;
assign w42237 = ~pi09961 & w17048;
assign w42238 = ~w42236 & ~w42237;
assign w42239 = pi09413 & ~w17048;
assign w42240 = ~pi09848 & w17048;
assign w42241 = ~w42239 & ~w42240;
assign w42242 = pi09414 & ~w17048;
assign w42243 = ~pi02704 & w17048;
assign w42244 = ~w42242 & ~w42243;
assign w42245 = pi09415 & ~w17048;
assign w42246 = ~pi02178 & w17048;
assign w42247 = ~w42245 & ~w42246;
assign w42248 = pi09416 & ~w17048;
assign w42249 = ~pi09954 & w17048;
assign w42250 = ~w42248 & ~w42249;
assign w42251 = pi09417 & ~w17048;
assign w42252 = ~pi02720 & w17048;
assign w42253 = ~w42251 & ~w42252;
assign w42254 = pi09418 & ~w17048;
assign w42255 = ~pi09962 & w17048;
assign w42256 = ~w42254 & ~w42255;
assign w42257 = pi09419 & ~w20621;
assign w42258 = ~pi09961 & w20621;
assign w42259 = ~w42257 & ~w42258;
assign w42260 = pi09420 & ~w18210;
assign w42261 = ~pi09961 & w18210;
assign w42262 = ~w42260 & ~w42261;
assign w42263 = pi09421 & ~w20621;
assign w42264 = ~pi09812 & w20621;
assign w42265 = ~w42263 & ~w42264;
assign w42266 = pi09422 & ~w20621;
assign w42267 = ~pi02704 & w20621;
assign w42268 = ~w42266 & ~w42267;
assign w42269 = pi09423 & ~w20621;
assign w42270 = ~pi02178 & w20621;
assign w42271 = ~w42269 & ~w42270;
assign w42272 = pi09424 & ~w20621;
assign w42273 = ~pi02720 & w20621;
assign w42274 = ~w42272 & ~w42273;
assign w42275 = pi09425 & ~w20621;
assign w42276 = ~pi09962 & w20621;
assign w42277 = ~w42275 & ~w42276;
assign w42278 = pi09426 & ~w20694;
assign w42279 = ~pi09961 & w20694;
assign w42280 = ~w42278 & ~w42279;
assign w42281 = pi09427 & ~w20694;
assign w42282 = ~pi09812 & w20694;
assign w42283 = ~w42281 & ~w42282;
assign w42284 = pi09428 & ~w20694;
assign w42285 = ~pi02704 & w20694;
assign w42286 = ~w42284 & ~w42285;
assign w42287 = pi09429 & ~w20694;
assign w42288 = ~pi02178 & w20694;
assign w42289 = ~w42287 & ~w42288;
assign w42290 = pi09430 & ~w20694;
assign w42291 = ~pi09954 & w20694;
assign w42292 = ~w42290 & ~w42291;
assign w42293 = pi09431 & ~w20694;
assign w42294 = ~pi02720 & w20694;
assign w42295 = ~w42293 & ~w42294;
assign w42296 = pi09432 & ~w20694;
assign w42297 = ~pi09962 & w20694;
assign w42298 = ~w42296 & ~w42297;
assign w42299 = pi09433 & ~w17501;
assign w42300 = ~pi09961 & w17501;
assign w42301 = ~w42299 & ~w42300;
assign w42302 = pi09434 & ~w17501;
assign w42303 = w17193 & w17500;
assign w42304 = ~w42302 & ~w42303;
assign w42305 = pi09435 & ~w17501;
assign w42306 = ~pi02704 & w17501;
assign w42307 = ~w42305 & ~w42306;
assign w42308 = pi09436 & ~w17501;
assign w42309 = ~pi02178 & w17501;
assign w42310 = ~w42308 & ~w42309;
assign w42311 = pi09437 & ~w17501;
assign w42312 = w17128 & w17500;
assign w42313 = ~w42311 & ~w42312;
assign w42314 = pi09438 & ~w17501;
assign w42315 = w17439 & w17500;
assign w42316 = ~w42314 & ~w42315;
assign w42317 = pi09439 & ~w21185;
assign w42318 = ~pi09961 & w21185;
assign w42319 = ~w42317 & ~w42318;
assign w42320 = pi09440 & ~w21185;
assign w42321 = ~pi09812 & w21185;
assign w42322 = ~w42320 & ~w42321;
assign w42323 = pi09441 & ~w21185;
assign w42324 = ~pi02704 & w21185;
assign w42325 = ~w42323 & ~w42324;
assign w42326 = pi09442 & ~w21185;
assign w42327 = ~pi02178 & w21185;
assign w42328 = ~w42326 & ~w42327;
assign w42329 = pi09443 & ~w21185;
assign w42330 = ~pi09954 & w21185;
assign w42331 = ~w42329 & ~w42330;
assign w42332 = pi09444 & ~w21185;
assign w42333 = ~pi02720 & w21185;
assign w42334 = ~w42332 & ~w42333;
assign w42335 = pi09445 & ~w21185;
assign w42336 = ~pi09962 & w21185;
assign w42337 = ~w42335 & ~w42336;
assign w42338 = pi09446 & ~w19497;
assign w42339 = ~pi09961 & w19497;
assign w42340 = ~w42338 & ~w42339;
assign w42341 = pi09447 & ~w19497;
assign w42342 = ~pi09812 & w19497;
assign w42343 = ~w42341 & ~w42342;
assign w42344 = pi09448 & ~w19497;
assign w42345 = ~pi02704 & w19497;
assign w42346 = ~w42344 & ~w42345;
assign w42347 = pi09449 & ~w19497;
assign w42348 = ~pi02178 & w19497;
assign w42349 = ~w42347 & ~w42348;
assign w42350 = pi09450 & ~w19497;
assign w42351 = ~pi02720 & w19497;
assign w42352 = ~w42350 & ~w42351;
assign w42353 = pi09451 & ~w19497;
assign w42354 = w17439 & w18370;
assign w42355 = ~w42353 & ~w42354;
assign w42356 = pi09452 & ~w17000;
assign w42357 = ~pi09961 & w17000;
assign w42358 = ~w42356 & ~w42357;
assign w42359 = pi09453 & ~w17000;
assign w42360 = ~pi09812 & w17000;
assign w42361 = ~w42359 & ~w42360;
assign w42362 = pi09454 & ~w17000;
assign w42363 = ~pi02704 & w17000;
assign w42364 = ~w42362 & ~w42363;
assign w42365 = pi09455 & ~w17000;
assign w42366 = ~pi02178 & w17000;
assign w42367 = ~w42365 & ~w42366;
assign w42368 = pi09456 & ~w17000;
assign w42369 = ~pi09954 & w17000;
assign w42370 = ~w42368 & ~w42369;
assign w42371 = pi09457 & ~w17000;
assign w42372 = ~pi02720 & w17000;
assign w42373 = ~w42371 & ~w42372;
assign w42374 = pi09458 & ~w17000;
assign w42375 = ~pi09962 & w17000;
assign w42376 = ~w42374 & ~w42375;
assign w42377 = pi09459 & ~w21228;
assign w42378 = ~pi09961 & w21228;
assign w42379 = ~w42377 & ~w42378;
assign w42380 = pi09460 & ~w21228;
assign w42381 = ~pi09812 & w21228;
assign w42382 = ~w42380 & ~w42381;
assign w42383 = pi09461 & ~w21228;
assign w42384 = ~pi02704 & w21228;
assign w42385 = ~w42383 & ~w42384;
assign w42386 = pi09462 & ~w21228;
assign w42387 = ~pi02178 & w21228;
assign w42388 = ~w42386 & ~w42387;
assign w42389 = pi09463 & ~w21228;
assign w42390 = ~pi02720 & w21228;
assign w42391 = ~w42389 & ~w42390;
assign w42392 = pi09464 & ~w21228;
assign w42393 = ~pi09962 & w21228;
assign w42394 = ~w42392 & ~w42393;
assign w42395 = pi09465 & ~w20988;
assign w42396 = ~pi09961 & w20988;
assign w42397 = ~w42395 & ~w42396;
assign w42398 = pi09466 & ~w20988;
assign w42399 = ~pi09812 & w20988;
assign w42400 = ~w42398 & ~w42399;
assign w42401 = pi09467 & ~w20988;
assign w42402 = ~pi02704 & w20988;
assign w42403 = ~w42401 & ~w42402;
assign w42404 = pi09468 & ~w20988;
assign w42405 = ~pi02178 & w20988;
assign w42406 = ~w42404 & ~w42405;
assign w42407 = pi09469 & ~w20988;
assign w42408 = w17513 & w17855;
assign w42409 = ~w42407 & ~w42408;
assign w42410 = pi09470 & ~w20988;
assign w42411 = ~pi02720 & w20988;
assign w42412 = ~w42410 & ~w42411;
assign w42413 = pi09471 & ~w20988;
assign w42414 = w17439 & w17855;
assign w42415 = ~w42413 & ~w42414;
assign w42416 = pi09472 & ~w21177;
assign w42417 = w17406 & w17439;
assign w42418 = ~w42416 & ~w42417;
assign w42419 = pi09473 & ~w17462;
assign w42420 = ~pi09848 & w17462;
assign w42421 = ~w42419 & ~w42420;
assign w42422 = pi09474 & ~w17462;
assign w42423 = w17193 & w17461;
assign w42424 = ~w42422 & ~w42423;
assign w42425 = pi09475 & ~w17462;
assign w42426 = ~pi02704 & w17462;
assign w42427 = ~w42425 & ~w42426;
assign w42428 = pi09476 & ~w17462;
assign w42429 = ~pi09954 & w17462;
assign w42430 = ~w42428 & ~w42429;
assign w42431 = pi09477 & ~w17462;
assign w42432 = ~pi02720 & w17462;
assign w42433 = ~w42431 & ~w42432;
assign w42434 = pi09478 & ~w17462;
assign w42435 = ~pi09962 & w17462;
assign w42436 = ~w42434 & ~w42435;
assign w42437 = pi09479 & ~w17120;
assign w42438 = ~pi09848 & w17120;
assign w42439 = ~w42437 & ~w42438;
assign w42440 = pi09480 & ~w17120;
assign w42441 = ~pi09812 & w17120;
assign w42442 = ~w42440 & ~w42441;
assign w42443 = pi09481 & ~w17120;
assign w42444 = ~pi02704 & w17120;
assign w42445 = ~w42443 & ~w42444;
assign w42446 = pi09482 & ~w17120;
assign w42447 = ~pi02178 & w17120;
assign w42448 = ~w42446 & ~w42447;
assign w42449 = pi09483 & ~w17120;
assign w42450 = w17119 & w17513;
assign w42451 = ~w42449 & ~w42450;
assign w42452 = pi09484 & ~w17120;
assign w42453 = ~pi02720 & w17120;
assign w42454 = ~w42452 & ~w42453;
assign w42455 = pi09485 & ~w17120;
assign w42456 = ~pi09962 & w17120;
assign w42457 = ~w42455 & ~w42456;
assign w42458 = pi09486 & ~w21246;
assign w42459 = ~pi09848 & w21246;
assign w42460 = ~w42458 & ~w42459;
assign w42461 = pi09487 & ~w21246;
assign w42462 = w16922 & w17193;
assign w42463 = ~w42461 & ~w42462;
assign w42464 = pi09488 & ~w21246;
assign w42465 = ~pi02704 & w21246;
assign w42466 = ~w42464 & ~w42465;
assign w42467 = pi09489 & ~w21246;
assign w42468 = ~pi09954 & w21246;
assign w42469 = ~w42467 & ~w42468;
assign w42470 = pi09490 & ~w21246;
assign w42471 = ~pi02720 & w21246;
assign w42472 = ~w42470 & ~w42471;
assign w42473 = pi09491 & ~w21246;
assign w42474 = ~pi09962 & w21246;
assign w42475 = ~w42473 & ~w42474;
assign w42476 = pi09492 & ~w17227;
assign w42477 = ~pi09848 & w17227;
assign w42478 = ~w42476 & ~w42477;
assign w42479 = pi09493 & ~w17227;
assign w42480 = ~pi09812 & w17227;
assign w42481 = ~w42479 & ~w42480;
assign w42482 = pi09494 & ~w17227;
assign w42483 = ~pi02704 & w17227;
assign w42484 = ~w42482 & ~w42483;
assign w42485 = pi09495 & ~w18627;
assign w42486 = ~pi09848 & w18627;
assign w42487 = ~w42485 & ~w42486;
assign w42488 = pi09496 & ~w17227;
assign w42489 = ~pi02178 & w17227;
assign w42490 = ~w42488 & ~w42489;
assign w42491 = pi09497 & ~w17227;
assign w42492 = w17226 & w17513;
assign w42493 = ~w42491 & ~w42492;
assign w42494 = pi09498 & ~w17227;
assign w42495 = ~pi02720 & w17227;
assign w42496 = ~w42494 & ~w42495;
assign w42497 = pi09499 & ~w17260;
assign w42498 = ~pi09961 & w17260;
assign w42499 = ~w42497 & ~w42498;
assign w42500 = pi09500 & ~w17260;
assign w42501 = ~pi09848 & w17260;
assign w42502 = ~w42500 & ~w42501;
assign w42503 = pi09501 & ~w17260;
assign w42504 = ~pi09812 & w17260;
assign w42505 = ~w42503 & ~w42504;
assign w42506 = pi09502 & ~w17260;
assign w42507 = ~pi02178 & w17260;
assign w42508 = ~w42506 & ~w42507;
assign w42509 = pi09503 & ~w17260;
assign w42510 = ~pi09954 & w17260;
assign w42511 = ~w42509 & ~w42510;
assign w42512 = pi09504 & ~w17260;
assign w42513 = ~pi02720 & w17260;
assign w42514 = ~w42512 & ~w42513;
assign w42515 = pi09505 & ~w21500;
assign w42516 = ~pi02707 & w21500;
assign w42517 = ~w42515 & ~w42516;
assign w42518 = ~w16928 & w17762;
assign w42519 = pi09506 & ~w42518;
assign w42520 = w17186 & w17762;
assign w42521 = ~w42519 & ~w42520;
assign w42522 = pi09507 & ~w42518;
assign w42523 = w17193 & w17762;
assign w42524 = ~w42522 & ~w42523;
assign w42525 = pi09508 & ~w42518;
assign w42526 = ~pi02704 & w42518;
assign w42527 = ~w42525 & ~w42526;
assign w42528 = pi09509 & ~w42518;
assign w42529 = w17762 & w18861;
assign w42530 = ~w42528 & ~w42529;
assign w42531 = pi09510 & ~w42518;
assign w42532 = ~pi09954 & w42518;
assign w42533 = ~w42531 & ~w42532;
assign w42534 = pi09511 & ~w42518;
assign w42535 = w17128 & w17762;
assign w42536 = ~w42534 & ~w42535;
assign w42537 = pi09512 & ~w20735;
assign w42538 = ~pi09961 & w20735;
assign w42539 = ~w42537 & ~w42538;
assign w42540 = pi09513 & ~w20735;
assign w42541 = w17186 & w17535;
assign w42542 = ~w42540 & ~w42541;
assign w42543 = pi09514 & ~w20735;
assign w42544 = ~pi09812 & w20735;
assign w42545 = ~w42543 & ~w42544;
assign w42546 = pi09515 & ~w20735;
assign w42547 = ~pi02178 & w20735;
assign w42548 = ~w42546 & ~w42547;
assign w42549 = pi09516 & ~w20735;
assign w42550 = ~pi09954 & w20735;
assign w42551 = ~w42549 & ~w42550;
assign w42552 = pi09517 & ~w20735;
assign w42553 = ~pi02720 & w20735;
assign w42554 = ~w42552 & ~w42553;
assign w42555 = pi09518 & ~w42518;
assign w42556 = w17762 & w19365;
assign w42557 = ~w42555 & ~w42556;
assign w42558 = pi09519 & ~w1193;
assign w42559 = ~pi09519 & ~pi10388;
assign w42560 = pi01216 & ~pi01454;
assign w42561 = w1192 & w42560;
assign w42562 = w11467 & w42559;
assign w42563 = w42561 & w42562;
assign w42564 = w16764 & w42563;
assign w42565 = ~w42558 & ~w42564;
assign w42566 = pi09520 & ~w30616;
assign w42567 = ~pi02708 & w30616;
assign w42568 = ~w42566 & ~w42567;
assign w42569 = pi09521 & ~w31720;
assign w42570 = ~pi02705 & w31720;
assign w42571 = ~w42569 & ~w42570;
assign w42572 = pi09522 & ~w21228;
assign w42573 = ~pi09848 & w21228;
assign w42574 = ~w42572 & ~w42573;
assign w42575 = pi09523 & ~w26184;
assign w42576 = ~pi02712 & w26184;
assign w42577 = ~w42575 & ~w42576;
assign w42578 = pi09524 & ~w20215;
assign w42579 = ~pi09812 & w20215;
assign w42580 = ~w42578 & ~w42579;
assign w42581 = pi09525 & ~w32538;
assign w42582 = ~pi02707 & w32538;
assign w42583 = ~w42581 & ~w42582;
assign w42584 = pi09526 & ~w28918;
assign w42585 = w18861 & w19459;
assign w42586 = ~w42584 & ~w42585;
assign w42587 = pi09527 & ~w28959;
assign w42588 = ~pi02178 & w28959;
assign w42589 = ~w42587 & ~w42588;
assign w42590 = pi09528 & ~w27595;
assign w42591 = ~pi02711 & w27595;
assign w42592 = ~w42590 & ~w42591;
assign w42593 = pi09529 & ~w38976;
assign w42594 = ~pi02719 & w38976;
assign w42595 = ~w42593 & ~w42594;
assign w42596 = pi09530 & ~w28959;
assign w42597 = ~pi09961 & w28959;
assign w42598 = ~w42596 & ~w42597;
assign w42599 = pi09531 & ~w32538;
assign w42600 = w17205 & w18689;
assign w42601 = ~w42599 & ~w42600;
assign w42602 = pi09532 & ~w30594;
assign w42603 = ~pi02706 & w30594;
assign w42604 = ~w42602 & ~w42603;
assign w42605 = pi09533 & ~w34012;
assign w42606 = ~pi02715 & w34012;
assign w42607 = ~w42605 & ~w42606;
assign w42608 = pi09534 & ~w20919;
assign w42609 = ~pi09812 & w20919;
assign w42610 = ~w42608 & ~w42609;
assign w42611 = pi09535 & ~w22807;
assign w42612 = ~pi02160 & w22807;
assign w42613 = ~w42611 & ~w42612;
assign w42614 = pi09536 & ~w31680;
assign w42615 = ~pi02708 & w31680;
assign w42616 = ~w42614 & ~w42615;
assign w42617 = pi09537 & ~w21929;
assign w42618 = ~pi02703 & w21929;
assign w42619 = ~w42617 & ~w42618;
assign w42620 = pi09538 & ~w28937;
assign w42621 = ~pi02178 & w28937;
assign w42622 = ~w42620 & ~w42621;
assign w42623 = pi09539 & ~w30616;
assign w42624 = w17148 & w17925;
assign w42625 = ~w42623 & ~w42624;
assign w42626 = pi09540 & ~w42518;
assign w42627 = w17439 & w17762;
assign w42628 = ~w42626 & ~w42627;
assign w42629 = pi09541 & ~w33190;
assign w42630 = ~pi02714 & w33190;
assign w42631 = ~w42629 & ~w42630;
assign w42632 = pi09542 & ~w31672;
assign w42633 = ~pi02718 & w31672;
assign w42634 = ~w42632 & ~w42633;
assign w42635 = pi09543 & ~w26158;
assign w42636 = ~pi02721 & w26158;
assign w42637 = ~w42635 & ~w42636;
assign w42638 = pi09544 & ~w26139;
assign w42639 = ~pi02712 & w26139;
assign w42640 = ~w42638 & ~w42639;
assign w42641 = pi09545 & ~w26139;
assign w42642 = ~pi02715 & w26139;
assign w42643 = ~w42641 & ~w42642;
assign w42644 = pi09546 & ~w22748;
assign w42645 = w18234 & w18431;
assign w42646 = ~w42644 & ~w42645;
assign w42647 = pi09547 & ~w28792;
assign w42648 = ~pi09961 & w28792;
assign w42649 = ~w42647 & ~w42648;
assign w42650 = pi09548 & ~w33186;
assign w42651 = ~pi02718 & w33186;
assign w42652 = ~w42650 & ~w42651;
assign w42653 = pi09549 & ~w20932;
assign w42654 = ~pi09954 & w20932;
assign w42655 = ~w42653 & ~w42654;
assign w42656 = pi09550 & ~w30575;
assign w42657 = ~pi02708 & w30575;
assign w42658 = ~w42656 & ~w42657;
assign w42659 = pi09551 & ~w31656;
assign w42660 = ~pi02723 & w31656;
assign w42661 = ~w42659 & ~w42660;
assign w42662 = pi09552 & ~w31448;
assign w42663 = ~pi02706 & w31448;
assign w42664 = ~w42662 & ~w42663;
assign w42665 = pi09553 & ~w25565;
assign w42666 = w17929 & w17965;
assign w42667 = ~w42665 & ~w42666;
assign w42668 = pi09554 & ~w36686;
assign w42669 = ~pi09812 & w36686;
assign w42670 = ~w42668 & ~w42669;
assign w42671 = pi09555 & ~w28918;
assign w42672 = w19365 & w19459;
assign w42673 = ~w42671 & ~w42672;
assign w42674 = pi09556 & ~w35966;
assign w42675 = ~pi02170 & w35966;
assign w42676 = ~w42674 & ~w42675;
assign w42677 = pi09557 & ~w32497;
assign w42678 = ~pi02708 & w32497;
assign w42679 = ~w42677 & ~w42678;
assign w42680 = pi09558 & ~w35919;
assign w42681 = ~pi02170 & w35919;
assign w42682 = ~w42680 & ~w42681;
assign w42683 = pi09559 & ~w21492;
assign w42684 = ~pi02160 & w21492;
assign w42685 = ~w42683 & ~w42684;
assign w42686 = pi09560 & ~w38448;
assign w42687 = ~pi02703 & w38448;
assign w42688 = ~w42686 & ~w42687;
assign w42689 = pi09561 & ~w26102;
assign w42690 = ~pi02713 & w26102;
assign w42691 = ~w42689 & ~w42690;
assign w42692 = pi09562 & ~w26102;
assign w42693 = ~pi02715 & w26102;
assign w42694 = ~w42692 & ~w42693;
assign w42695 = pi09563 & ~w35929;
assign w42696 = ~pi02722 & w35929;
assign w42697 = ~w42695 & ~w42696;
assign w42698 = pi09564 & ~w37402;
assign w42699 = ~pi02714 & w37402;
assign w42700 = ~w42698 & ~w42699;
assign w42701 = pi09565 & ~w21540;
assign w42702 = ~pi02716 & w21540;
assign w42703 = ~w42701 & ~w42702;
assign w42704 = pi09566 & ~w22767;
assign w42705 = w18234 & w18247;
assign w42706 = ~w42704 & ~w42705;
assign w42707 = pi09567 & ~w28874;
assign w42708 = ~pi02178 & w28874;
assign w42709 = ~w42707 & ~w42708;
assign w42710 = pi09568 & ~w22748;
assign w42711 = ~pi02710 & w22748;
assign w42712 = ~w42710 & ~w42711;
assign w42713 = pi09569 & ~w30575;
assign w42714 = ~pi02706 & w30575;
assign w42715 = ~w42713 & ~w42714;
assign w42716 = pi09570 & ~w28874;
assign w42717 = w19365 & w19492;
assign w42718 = ~w42716 & ~w42717;
assign w42719 = pi09571 & ~w30553;
assign w42720 = ~pi02706 & w30553;
assign w42721 = ~w42719 & ~w42720;
assign w42722 = pi09572 & ~w31656;
assign w42723 = ~pi02710 & w31656;
assign w42724 = ~w42722 & ~w42723;
assign w42725 = pi09573 & ~w36888;
assign w42726 = ~pi02714 & w36888;
assign w42727 = ~w42725 & ~w42726;
assign w42728 = pi09574 & ~w26098;
assign w42729 = ~pi02721 & w26098;
assign w42730 = ~w42728 & ~w42729;
assign w42731 = pi09575 & ~w28852;
assign w42732 = w18861 & w19518;
assign w42733 = ~w42731 & ~w42732;
assign w42734 = pi09576 & ~w36892;
assign w42735 = ~pi02718 & w36892;
assign w42736 = ~w42734 & ~w42735;
assign w42737 = pi09577 & ~w26076;
assign w42738 = ~pi02712 & w26076;
assign w42739 = ~w42737 & ~w42738;
assign w42740 = pi09578 & ~w28833;
assign w42741 = ~pi02178 & w28833;
assign w42742 = ~w42740 & ~w42741;
assign w42743 = pi09579 & ~w22726;
assign w42744 = ~pi02160 & w22726;
assign w42745 = ~w42743 & ~w42744;
assign w42746 = pi09580 & ~w22707;
assign w42747 = ~pi02710 & w22707;
assign w42748 = ~w42746 & ~w42747;
assign w42749 = pi09581 & ~w26057;
assign w42750 = w18059 & w19852;
assign w42751 = ~w42749 & ~w42750;
assign w42752 = pi09582 & ~w22707;
assign w42753 = ~pi02160 & w22707;
assign w42754 = ~w42752 & ~w42753;
assign w42755 = pi09583 & ~w28833;
assign w42756 = ~pi09961 & w28833;
assign w42757 = ~w42755 & ~w42756;
assign w42758 = pi09584 & ~w26057;
assign w42759 = ~pi02712 & w26057;
assign w42760 = ~w42758 & ~w42759;
assign w42761 = pi09585 & ~w22663;
assign w42762 = ~pi02160 & w22663;
assign w42763 = ~w42761 & ~w42762;
assign w42764 = pi09586 & ~w22685;
assign w42765 = w18234 & w18822;
assign w42766 = ~w42764 & ~w42765;
assign w42767 = pi09587 & ~w35501;
assign w42768 = ~pi02717 & w35501;
assign w42769 = ~w42767 & ~w42768;
assign w42770 = pi09588 & ~w26035;
assign w42771 = ~pi02721 & w26035;
assign w42772 = ~w42770 & ~w42771;
assign w42773 = pi09589 & ~w22663;
assign w42774 = ~pi02710 & w22663;
assign w42775 = ~w42773 & ~w42774;
assign w42776 = pi09590 & ~w28811;
assign w42777 = ~pi02178 & w28811;
assign w42778 = ~w42776 & ~w42777;
assign w42779 = pi09591 & ~w30534;
assign w42780 = ~pi02708 & w30534;
assign w42781 = ~w42779 & ~w42780;
assign w42782 = pi09592 & ~w26016;
assign w42783 = ~pi02721 & w26016;
assign w42784 = ~w42782 & ~w42783;
assign w42785 = pi09593 & ~w30534;
assign w42786 = ~pi02706 & w30534;
assign w42787 = ~w42785 & ~w42786;
assign w42788 = pi09594 & ~w26016;
assign w42789 = ~pi02164 & w26016;
assign w42790 = ~w42788 & ~w42789;
assign w42791 = pi09595 & ~w22644;
assign w42792 = ~pi02705 & w22644;
assign w42793 = ~w42791 & ~w42792;
assign w42794 = pi09596 & ~w36391;
assign w42795 = ~pi02713 & w36391;
assign w42796 = ~w42794 & ~w42795;
assign w42797 = pi09597 & ~w28792;
assign w42798 = ~pi02178 & w28792;
assign w42799 = ~w42797 & ~w42798;
assign w42800 = pi09598 & ~w22644;
assign w42801 = ~pi02723 & w22644;
assign w42802 = ~w42800 & ~w42801;
assign w42803 = pi09599 & ~w22521;
assign w42804 = ~pi02723 & w22521;
assign w42805 = ~w42803 & ~w42804;
assign w42806 = pi09600 & ~w25994;
assign w42807 = ~pi02721 & w25994;
assign w42808 = ~w42806 & ~w42807;
assign w42809 = pi09601 & ~w22603;
assign w42810 = ~pi02705 & w22603;
assign w42811 = ~w42809 & ~w42810;
assign w42812 = pi09602 & ~w30512;
assign w42813 = ~pi02706 & w30512;
assign w42814 = ~w42812 & ~w42813;
assign w42815 = pi09603 & ~w22622;
assign w42816 = ~pi02723 & w22622;
assign w42817 = ~w42815 & ~w42816;
assign w42818 = pi09604 & ~w25975;
assign w42819 = ~pi02715 & w25975;
assign w42820 = ~w42818 & ~w42819;
assign w42821 = pi09605 & ~w22603;
assign w42822 = ~pi02723 & w22603;
assign w42823 = ~w42821 & ~w42822;
assign w42824 = pi09606 & ~w33829;
assign w42825 = ~pi02169 & w33829;
assign w42826 = ~w42824 & ~w42825;
assign w42827 = pi09607 & ~w22562;
assign w42828 = ~pi02723 & w22562;
assign w42829 = ~w42827 & ~w42828;
assign w42830 = pi09608 & ~w25953;
assign w42831 = ~pi02712 & w25953;
assign w42832 = ~w42830 & ~w42831;
assign w42833 = pi09609 & ~w25975;
assign w42834 = ~pi02712 & w25975;
assign w42835 = ~w42833 & ~w42834;
assign w42836 = pi09610 & ~w22581;
assign w42837 = w17671 & w18944;
assign w42838 = ~w42836 & ~w42837;
assign w42839 = pi09611 & ~w28770;
assign w42840 = ~pi02178 & w28770;
assign w42841 = ~w42839 & ~w42840;
assign w42842 = pi09612 & ~w20425;
assign w42843 = ~pi02703 & w20425;
assign w42844 = ~w42842 & ~w42843;
assign w42845 = pi09613 & ~w35473;
assign w42846 = ~pi02714 & w35473;
assign w42847 = ~w42845 & ~w42846;
assign w42848 = pi09614 & ~w25908;
assign w42849 = ~pi02722 & w25908;
assign w42850 = ~w42848 & ~w42849;
assign w42851 = pi09615 & ~w36391;
assign w42852 = ~pi02711 & w36391;
assign w42853 = ~w42851 & ~w42852;
assign w42854 = pi09616 & ~w28751;
assign w42855 = ~pi02178 & w28751;
assign w42856 = ~w42854 & ~w42855;
assign w42857 = pi09617 & ~w28751;
assign w42858 = ~pi09961 & w28751;
assign w42859 = ~w42857 & ~w42858;
assign w42860 = pi09618 & ~w35473;
assign w42861 = ~pi02717 & w35473;
assign w42862 = ~w42860 & ~w42861;
assign w42863 = pi09619 & ~w30493;
assign w42864 = ~pi02708 & w30493;
assign w42865 = ~w42863 & ~w42864;
assign w42866 = pi09620 & ~w25908;
assign w42867 = ~pi02167 & w25908;
assign w42868 = ~w42866 & ~w42867;
assign w42869 = pi09621 & ~w31656;
assign w42870 = ~pi02705 & w31656;
assign w42871 = ~w42869 & ~w42870;
assign w42872 = pi09622 & ~w30493;
assign w42873 = w17925 & w19306;
assign w42874 = ~w42872 & ~w42873;
assign w42875 = pi09623 & ~w37421;
assign w42876 = ~pi02167 & w37421;
assign w42877 = ~w42875 & ~w42876;
assign w42878 = pi09624 & ~w22562;
assign w42879 = ~pi02705 & w22562;
assign w42880 = ~w42878 & ~w42879;
assign w42881 = pi09625 & ~w22540;
assign w42882 = ~pi02723 & w22540;
assign w42883 = ~w42881 & ~w42882;
assign w42884 = pi09626 & ~w25908;
assign w42885 = ~pi02721 & w25908;
assign w42886 = ~w42884 & ~w42885;
assign w42887 = pi09627 & ~w28729;
assign w42888 = w18861 & w19606;
assign w42889 = ~w42887 & ~w42888;
assign w42890 = pi09628 & ~w31634;
assign w42891 = ~pi02705 & w31634;
assign w42892 = ~w42890 & ~w42891;
assign w42893 = pi09629 & ~w22477;
assign w42894 = ~pi02705 & w22477;
assign w42895 = ~w42893 & ~w42894;
assign w42896 = pi09630 & ~w22436;
assign w42897 = ~pi02723 & w22436;
assign w42898 = ~w42896 & ~w42897;
assign w42899 = pi09631 & ~w22521;
assign w42900 = ~pi02705 & w22521;
assign w42901 = ~w42899 & ~w42900;
assign w42902 = pi09632 & ~w37421;
assign w42903 = ~pi02721 & w37421;
assign w42904 = ~w42902 & ~w42903;
assign w42905 = pi09633 & ~w25871;
assign w42906 = ~pi02716 & w25871;
assign w42907 = ~w42905 & ~w42906;
assign w42908 = pi09634 & ~w22477;
assign w42909 = ~pi02723 & w22477;
assign w42910 = ~w42908 & ~w42909;
assign w42911 = pi09635 & ~w25871;
assign w42912 = ~pi02714 & w25871;
assign w42913 = ~w42911 & ~w42912;
assign w42914 = pi09636 & ~w30471;
assign w42915 = ~pi02706 & w30471;
assign w42916 = ~w42914 & ~w42915;
assign w42917 = pi09637 & ~w28710;
assign w42918 = ~pi02178 & w28710;
assign w42919 = ~w42917 & ~w42918;
assign w42920 = pi09638 & ~w25867;
assign w42921 = ~pi02721 & w25867;
assign w42922 = ~w42920 & ~w42921;
assign w42923 = pi09639 & ~w28710;
assign w42924 = ~pi09961 & w28710;
assign w42925 = ~w42923 & ~w42924;
assign w42926 = pi09640 & ~w28669;
assign w42927 = w18861 & w19645;
assign w42928 = ~w42926 & ~w42927;
assign w42929 = pi09641 & ~w28688;
assign w42930 = ~pi02178 & w28688;
assign w42931 = ~w42929 & ~w42930;
assign w42932 = pi09642 & ~w25848;
assign w42933 = ~pi02715 & w25848;
assign w42934 = ~w42932 & ~w42933;
assign w42935 = pi09643 & ~w31615;
assign w42936 = ~pi02723 & w31615;
assign w42937 = ~w42935 & ~w42936;
assign w42938 = pi09644 & ~w25826;
assign w42939 = ~pi02712 & w25826;
assign w42940 = ~w42938 & ~w42939;
assign w42941 = pi09645 & ~w30411;
assign w42942 = w17320 & w17925;
assign w42943 = ~w42941 & ~w42942;
assign w42944 = pi09646 & ~w30452;
assign w42945 = ~pi02708 & w30452;
assign w42946 = ~w42944 & ~w42945;
assign w42947 = pi09647 & ~w25848;
assign w42948 = ~pi02712 & w25848;
assign w42949 = ~w42947 & ~w42948;
assign w42950 = pi09648 & ~w30452;
assign w42951 = ~pi02706 & w30452;
assign w42952 = ~w42950 & ~w42951;
assign w42953 = pi09649 & ~w25807;
assign w42954 = ~pi02712 & w25807;
assign w42955 = ~w42953 & ~w42954;
assign w42956 = pi09650 & ~w42034;
assign w42957 = ~pi09812 & w42034;
assign w42958 = ~w42956 & ~w42957;
assign w42959 = pi09651 & ~w25807;
assign w42960 = ~pi02715 & w25807;
assign w42961 = ~w42959 & ~w42960;
assign w42962 = pi09652 & ~w22455;
assign w42963 = ~pi02723 & w22455;
assign w42964 = ~w42962 & ~w42963;
assign w42965 = pi09653 & ~w28669;
assign w42966 = ~pi09961 & w28669;
assign w42967 = ~w42965 & ~w42966;
assign w42968 = pi09654 & ~w30430;
assign w42969 = w17344 & w17925;
assign w42970 = ~w42968 & ~w42969;
assign w42971 = pi09655 & ~w31615;
assign w42972 = ~pi02705 & w31615;
assign w42973 = ~w42971 & ~w42972;
assign w42974 = pi09656 & ~w30411;
assign w42975 = ~pi02708 & w30411;
assign w42976 = ~w42974 & ~w42975;
assign w42977 = pi09657 & ~w28647;
assign w42978 = ~pi02178 & w28647;
assign w42979 = ~w42977 & ~w42978;
assign w42980 = pi09658 & ~w32504;
assign w42981 = ~pi02703 & w32504;
assign w42982 = ~w42980 & ~w42981;
assign w42983 = pi09659 & ~w30370;
assign w42984 = ~pi02708 & w30370;
assign w42985 = ~w42983 & ~w42984;
assign w42986 = pi09660 & ~w30200;
assign w42987 = ~pi02160 & w30200;
assign w42988 = ~w42986 & ~w42987;
assign w42989 = pi09661 & ~w28628;
assign w42990 = ~pi02178 & w28628;
assign w42991 = ~w42989 & ~w42990;
assign w42992 = pi09662 & ~w32415;
assign w42993 = w17125 & w18067;
assign w42994 = ~w42992 & ~w42993;
assign w42995 = pi09663 & ~w25785;
assign w42996 = ~pi02721 & w25785;
assign w42997 = ~w42995 & ~w42996;
assign w42998 = pi09664 & ~w30389;
assign w42999 = ~pi02706 & w30389;
assign w43000 = ~w42998 & ~w42999;
assign w43001 = pi09665 & ~w32466;
assign w43002 = ~pi02707 & w32466;
assign w43003 = ~w43001 & ~w43002;
assign w43004 = pi09666 & ~w28628;
assign w43005 = ~pi09961 & w28628;
assign w43006 = ~w43004 & ~w43005;
assign w43007 = pi09667 & ~w28565;
assign w43008 = ~pi02178 & w28565;
assign w43009 = ~w43007 & ~w43008;
assign w43010 = pi09668 & ~w31593;
assign w43011 = ~pi02705 & w31593;
assign w43012 = ~w43010 & ~w43011;
assign w43013 = pi09669 & ~w31568;
assign w43014 = ~pi02723 & w31568;
assign w43015 = ~w43013 & ~w43014;
assign w43016 = pi09670 & ~w28606;
assign w43017 = ~pi02178 & w28606;
assign w43018 = ~w43016 & ~w43017;
assign w43019 = pi09671 & ~w25766;
assign w43020 = ~pi02164 & w25766;
assign w43021 = ~w43019 & ~w43020;
assign w43022 = pi09672 & ~w30370;
assign w43023 = w17325 & w17925;
assign w43024 = ~w43022 & ~w43023;
assign w43025 = pi09673 & ~w30348;
assign w43026 = ~pi02706 & w30348;
assign w43027 = ~w43025 & ~w43026;
assign w43028 = pi09674 & ~w33297;
assign w43029 = ~pi02703 & w33297;
assign w43030 = ~w43028 & ~w43029;
assign w43031 = pi09675 & ~w35473;
assign w43032 = w17148 & w20209;
assign w43033 = ~w43031 & ~w43032;
assign w43034 = pi09676 & ~w22332;
assign w43035 = w17671 & w19106;
assign w43036 = ~w43034 & ~w43035;
assign w43037 = pi09677 & ~w25766;
assign w43038 = ~pi02721 & w25766;
assign w43039 = ~w43037 & ~w43038;
assign w43040 = pi09678 & ~w28587;
assign w43041 = ~pi02178 & w28587;
assign w43042 = ~w43040 & ~w43041;
assign w43043 = pi09679 & ~w28587;
assign w43044 = ~pi09961 & w28587;
assign w43045 = ~w43043 & ~w43044;
assign w43046 = pi09680 & ~w33936;
assign w43047 = ~pi02714 & w33936;
assign w43048 = ~w43046 & ~w43047;
assign w43049 = pi09681 & ~w25710;
assign w43050 = w17103 & w17317;
assign w43051 = ~w43049 & ~w43050;
assign w43052 = pi09682 & ~w25744;
assign w43053 = w17020 & w17078;
assign w43054 = ~w43052 & ~w43053;
assign w43055 = pi09683 & ~w31537;
assign w43056 = w17334 & w17925;
assign w43057 = ~w43055 & ~w43056;
assign w43058 = pi09684 & ~w30329;
assign w43059 = ~pi02708 & w30329;
assign w43060 = ~w43058 & ~w43059;
assign w43061 = pi09685 & ~w25710;
assign w43062 = w17103 & w17929;
assign w43063 = ~w43061 & ~w43062;
assign w43064 = pi09686 & ~w35102;
assign w43065 = w19306 & w19312;
assign w43066 = ~w43064 & ~w43065;
assign w43067 = pi09687 & ~w22436;
assign w43068 = ~pi02705 & w22436;
assign w43069 = ~w43067 & ~w43068;
assign w43070 = pi09688 & ~w31530;
assign w43071 = ~pi02722 & w31530;
assign w43072 = ~w43070 & ~w43071;
assign w43073 = pi09689 & ~w28546;
assign w43074 = ~pi02178 & w28546;
assign w43075 = ~w43073 & ~w43074;
assign w43076 = pi09690 & ~w30329;
assign w43077 = ~pi02706 & w30329;
assign w43078 = ~w43076 & ~w43077;
assign w43079 = pi09691 & ~w28546;
assign w43080 = w19365 & w19740;
assign w43081 = ~w43079 & ~w43080;
assign w43082 = pi09692 & ~w28505;
assign w43083 = w19365 & w19826;
assign w43084 = ~w43082 & ~w43083;
assign w43085 = pi09693 & ~w32497;
assign w43086 = ~pi02707 & w32497;
assign w43087 = ~w43085 & ~w43086;
assign w43088 = pi09694 & ~w30285;
assign w43089 = ~pi02707 & w30285;
assign w43090 = ~w43088 & ~w43089;
assign w43091 = pi09695 & ~w35463;
assign w43092 = ~pi02703 & w35463;
assign w43093 = ~w43091 & ~w43092;
assign w43094 = pi09696 & ~w28524;
assign w43095 = w18861 & w19818;
assign w43096 = ~w43094 & ~w43095;
assign w43097 = pi09697 & ~w30307;
assign w43098 = ~pi02706 & w30307;
assign w43099 = ~w43097 & ~w43098;
assign w43100 = pi09698 & ~w25703;
assign w43101 = ~pi02721 & w25703;
assign w43102 = ~w43100 & ~w43101;
assign w43103 = pi09699 & ~w20713;
assign w43104 = ~pi02718 & w20713;
assign w43105 = ~w43103 & ~w43104;
assign w43106 = pi09700 & ~w25684;
assign w43107 = ~pi02712 & w25684;
assign w43108 = ~w43106 & ~w43107;
assign w43109 = pi09701 & ~w25684;
assign w43110 = ~pi02715 & w25684;
assign w43111 = ~w43109 & ~w43110;
assign w43112 = pi09702 & ~w22414;
assign w43113 = ~pi02723 & w22414;
assign w43114 = ~w43112 & ~w43113;
assign w43115 = pi09703 & ~w30285;
assign w43116 = ~pi02708 & w30285;
assign w43117 = ~w43115 & ~w43116;
assign w43118 = pi09704 & ~w28505;
assign w43119 = ~pi02178 & w28505;
assign w43120 = ~w43118 & ~w43119;
assign w43121 = pi09705 & ~w31537;
assign w43122 = ~pi02160 & w31537;
assign w43123 = ~w43121 & ~w43122;
assign w43124 = pi09706 & ~w25662;
assign w43125 = ~pi02712 & w25662;
assign w43126 = ~w43124 & ~w43125;
assign w43127 = pi09707 & ~w28483;
assign w43128 = ~pi02178 & w28483;
assign w43129 = ~w43127 & ~w43128;
assign w43130 = pi09708 & ~w28379;
assign w43131 = ~pi09954 & w28379;
assign w43132 = ~w43130 & ~w43131;
assign w43133 = pi09709 & ~w28439;
assign w43134 = ~pi09954 & w28439;
assign w43135 = ~w43133 & ~w43134;
assign w43136 = pi09710 & ~w30263;
assign w43137 = ~pi02707 & w30263;
assign w43138 = ~w43136 & ~w43137;
assign w43139 = pi09711 & ~w28464;
assign w43140 = ~pi02178 & w28464;
assign w43141 = ~w43139 & ~w43140;
assign w43142 = pi09712 & ~w22395;
assign w43143 = ~pi02723 & w22395;
assign w43144 = ~w43142 & ~w43143;
assign w43145 = pi09713 & ~w30244;
assign w43146 = ~pi02709 & w30244;
assign w43147 = ~w43145 & ~w43146;
assign w43148 = pi09714 & ~w28464;
assign w43149 = ~pi09961 & w28464;
assign w43150 = ~w43148 & ~w43149;
assign w43151 = pi09715 & ~w25643;
assign w43152 = w17626 & w18059;
assign w43153 = ~w43151 & ~w43152;
assign w43154 = pi09716 & ~w22395;
assign w43155 = w18578 & w19130;
assign w43156 = ~w43154 & ~w43155;
assign w43157 = pi09717 & ~w30244;
assign w43158 = ~pi02707 & w30244;
assign w43159 = ~w43157 & ~w43158;
assign w43160 = pi09718 & ~w25643;
assign w43161 = ~pi02712 & w25643;
assign w43162 = ~w43160 & ~w43161;
assign w43163 = pi09719 & ~w31505;
assign w43164 = w18364 & w18631;
assign w43165 = ~w43163 & ~w43164;
assign w43166 = pi09720 & ~w28420;
assign w43167 = ~pi09954 & w28420;
assign w43168 = ~w43166 & ~w43167;
assign w43169 = pi09721 & ~w28398;
assign w43170 = ~pi09954 & w28398;
assign w43171 = ~w43169 & ~w43170;
assign w43172 = pi09722 & ~w28420;
assign w43173 = ~pi09848 & w28420;
assign w43174 = ~w43172 & ~w43173;
assign w43175 = pi09723 & ~w30222;
assign w43176 = ~pi02707 & w30222;
assign w43177 = ~w43175 & ~w43176;
assign w43178 = pi09724 & ~w25621;
assign w43179 = ~pi02721 & w25621;
assign w43180 = ~w43178 & ~w43179;
assign w43181 = pi09725 & ~w25602;
assign w43182 = w17912 & w18059;
assign w43183 = ~w43181 & ~w43182;
assign w43184 = pi09726 & ~w30200;
assign w43185 = ~pi02710 & w30200;
assign w43186 = ~w43184 & ~w43185;
assign w43187 = pi09727 & ~w31505;
assign w43188 = ~pi02706 & w31505;
assign w43189 = ~w43187 & ~w43188;
assign w43190 = pi09728 & ~w22373;
assign w43191 = ~pi02723 & w22373;
assign w43192 = ~w43190 & ~w43191;
assign w43193 = pi09729 & ~w25602;
assign w43194 = ~pi02712 & w25602;
assign w43195 = ~w43193 & ~w43194;
assign w43196 = pi09730 & ~w33968;
assign w43197 = ~pi02719 & w33968;
assign w43198 = ~w43196 & ~w43197;
assign w43199 = pi09731 & ~w33297;
assign w43200 = ~pi02167 & w33297;
assign w43201 = ~w43199 & ~w43200;
assign w43202 = pi09732 & ~w31473;
assign w43203 = ~pi02710 & w31473;
assign w43204 = ~w43202 & ~w43203;
assign w43205 = pi09733 & ~w33256;
assign w43206 = w17762 & w18578;
assign w43207 = ~w43205 & ~w43206;
assign w43208 = pi09734 & ~w35102;
assign w43209 = ~pi02718 & w35102;
assign w43210 = ~w43208 & ~w43209;
assign w43211 = pi09735 & ~w33968;
assign w43212 = ~pi02169 & w33968;
assign w43213 = ~w43211 & ~w43212;
assign w43214 = pi09736 & ~w35102;
assign w43215 = w17620 & w19306;
assign w43216 = ~w43214 & ~w43215;
assign w43217 = pi09737 & ~w33984;
assign w43218 = ~pi02714 & w33984;
assign w43219 = ~w43217 & ~w43218;
assign w43220 = pi09738 & ~w34592;
assign w43221 = w17532 & w17600;
assign w43222 = ~w43220 & ~w43221;
assign w43223 = pi09739 & ~w30178;
assign w43224 = ~pi02160 & w30178;
assign w43225 = ~w43223 & ~w43224;
assign w43226 = pi09740 & ~w33275;
assign w43227 = ~pi02705 & w33275;
assign w43228 = ~w43226 & ~w43227;
assign w43229 = pi09741 & ~w32456;
assign w43230 = ~pi02167 & w32456;
assign w43231 = ~w43229 & ~w43230;
assign w43232 = pi09742 & ~w31473;
assign w43233 = ~pi02723 & w31473;
assign w43234 = ~w43232 & ~w43233;
assign w43235 = pi09743 & ~w22354;
assign w43236 = ~pi02723 & w22354;
assign w43237 = ~w43235 & ~w43236;
assign w43238 = pi09744 & ~w34573;
assign w43239 = w17565 & w17742;
assign w43240 = ~w43238 & ~w43239;
assign w43241 = pi09745 & ~w33984;
assign w43242 = ~pi02712 & w33984;
assign w43243 = ~w43241 & ~w43242;
assign w43244 = pi09746 & ~w32456;
assign w43245 = ~pi02703 & w32456;
assign w43246 = ~w43244 & ~w43245;
assign w43247 = pi09747 & ~w41523;
assign w43248 = ~pi02704 & w41523;
assign w43249 = ~w43247 & ~w43248;
assign w43250 = pi09748 & ~w28357;
assign w43251 = ~pi09954 & w28357;
assign w43252 = ~w43250 & ~w43251;
assign w43253 = pi09749 & ~w28379;
assign w43254 = w17186 & w19988;
assign w43255 = ~w43253 & ~w43254;
assign w43256 = pi09750 & ~w34573;
assign w43257 = w17565 & w17603;
assign w43258 = ~w43256 & ~w43257;
assign w43259 = pi09751 & ~w25558;
assign w43260 = ~pi02718 & w25558;
assign w43261 = ~w43259 & ~w43260;
assign w43262 = pi09752 & ~w33955;
assign w43263 = ~pi02711 & w33955;
assign w43264 = ~w43262 & ~w43263;
assign w43265 = pi09753 & ~w22354;
assign w43266 = ~pi02705 & w22354;
assign w43267 = ~w43265 & ~w43266;
assign w43268 = pi09754 & ~w33256;
assign w43269 = ~pi02723 & w33256;
assign w43270 = ~w43268 & ~w43269;
assign w43271 = pi09755 & ~w32422;
assign w43272 = ~pi02718 & w32422;
assign w43273 = ~w43271 & ~w43272;
assign w43274 = pi09756 & ~w41426;
assign w43275 = w17128 & w20775;
assign w43276 = ~w43274 & ~w43275;
assign w43277 = pi09757 & ~w21385;
assign w43278 = ~pi02178 & w21385;
assign w43279 = ~w43277 & ~w43278;
assign w43280 = pi09758 & ~w17007;
assign w43281 = w17006 & w17742;
assign w43282 = ~w43280 & ~w43281;
assign w43283 = pi09759 & ~w35042;
assign w43284 = ~pi02713 & w35042;
assign w43285 = ~w43283 & ~w43284;
assign w43286 = pi09760 & ~w35042;
assign w43287 = ~pi02717 & w35042;
assign w43288 = ~w43286 & ~w43287;
assign w43289 = pi09761 & ~w34551;
assign w43290 = w17603 & w18177;
assign w43291 = ~w43289 & ~w43290;
assign w43292 = pi09762 & ~w35086;
assign w43293 = ~pi02716 & w35086;
assign w43294 = ~w43292 & ~w43293;
assign w43295 = pi09763 & ~w34491;
assign w43296 = w17284 & w17603;
assign w43297 = ~w43295 & ~w43296;
assign w43298 = pi09764 & ~w34514;
assign w43299 = w17177 & w17603;
assign w43300 = ~w43298 & ~w43299;
assign w43301 = pi09765 & ~w31477;
assign w43302 = ~pi02703 & w31477;
assign w43303 = ~w43301 & ~w43302;
assign w43304 = pi09766 & ~w35086;
assign w43305 = ~pi02713 & w35086;
assign w43306 = ~w43304 & ~w43305;
assign w43307 = pi09767 & ~w33186;
assign w43308 = ~pi02722 & w33186;
assign w43309 = ~w43307 & ~w43308;
assign w43310 = pi09768 & ~w33936;
assign w43311 = ~pi02711 & w33936;
assign w43312 = ~w43310 & ~w43311;
assign w43313 = pi09769 & ~w34514;
assign w43314 = ~pi02716 & w34514;
assign w43315 = ~w43313 & ~w43314;
assign w43316 = pi09770 & ~w31030;
assign w43317 = ~pi09812 & w31030;
assign w43318 = ~w43316 & ~w43317;
assign w43319 = pi09771 & ~w35441;
assign w43320 = ~pi02713 & w35441;
assign w43321 = ~w43319 & ~w43320;
assign w43322 = pi09772 & ~w20090;
assign w43323 = w16941 & w17439;
assign w43324 = ~w43322 & ~w43323;
assign w43325 = pi09773 & ~w35064;
assign w43326 = w16973 & w18683;
assign w43327 = ~w43325 & ~w43326;
assign w43328 = pi09774 & ~w34510;
assign w43329 = ~pi02167 & w34510;
assign w43330 = ~w43328 & ~w43329;
assign w43331 = pi09775 & ~w31269;
assign w43332 = ~pi09812 & w31269;
assign w43333 = ~w43331 & ~w43332;
assign w43334 = pi09776 & ~w31477;
assign w43335 = ~pi02721 & w31477;
assign w43336 = ~w43334 & ~w43335;
assign w43337 = pi09777 & ~w21216;
assign w43338 = w17193 & w17663;
assign w43339 = ~w43337 & ~w43338;
assign w43340 = pi09778 & ~w32422;
assign w43341 = ~pi02703 & w32422;
assign w43342 = ~w43340 & ~w43341;
assign w43343 = pi09779 & ~w21246;
assign w43344 = w16922 & w19365;
assign w43345 = ~w43343 & ~w43344;
assign w43346 = pi09780 & ~w35419;
assign w43347 = w16973 & w17694;
assign w43348 = ~w43346 & ~w43347;
assign w43349 = pi09781 & ~w17061;
assign w43350 = ~pi02723 & w17061;
assign w43351 = ~w43349 & ~w43350;
assign w43352 = pi09782 & ~w38448;
assign w43353 = w19273 & w20244;
assign w43354 = ~w43352 & ~w43353;
assign w43355 = pi09783 & ~w40108;
assign w43356 = ~pi02704 & w40108;
assign w43357 = ~w43355 & ~w43356;
assign w43358 = pi09784 & ~w37902;
assign w43359 = ~pi02713 & w37902;
assign w43360 = ~w43358 & ~w43359;
assign w43361 = pi09785 & ~w30153;
assign w43362 = w17671 & w18009;
assign w43363 = ~w43361 & ~w43362;
assign w43364 = pi09786 & ~w28338;
assign w43365 = ~pi09954 & w28338;
assign w43366 = ~w43364 & ~w43365;
assign w43367 = pi09787 & ~w17126;
assign w43368 = ~pi09812 & w17126;
assign w43369 = ~w43367 & ~w43368;
assign w43370 = pi09788 & ~w34491;
assign w43371 = ~pi02714 & w34491;
assign w43372 = ~w43370 & ~w43371;
assign w43373 = pi09789 & ~w25565;
assign w43374 = ~pi02711 & w25565;
assign w43375 = ~w43373 & ~w43374;
assign w43376 = pi09790 & ~w21527;
assign w43377 = ~pi02164 & w21527;
assign w43378 = ~w43376 & ~w43377;
assign w43379 = pi09791 & ~w33914;
assign w43380 = w17603 & w17734;
assign w43381 = ~w43379 & ~w43380;
assign w43382 = pi09792 & ~w41426;
assign w43383 = ~pi09812 & w41426;
assign w43384 = ~w43382 & ~w43383;
assign w43385 = pi09793 & ~w33194;
assign w43386 = ~pi02710 & w33194;
assign w43387 = ~w43385 & ~w43386;
assign w43388 = pi09794 & ~w35005;
assign w43389 = ~pi02722 & w35005;
assign w43390 = ~w43388 & ~w43389;
assign w43391 = pi09795 & ~w20713;
assign w43392 = ~pi02721 & w20713;
assign w43393 = ~w43391 & ~w43392;
assign w43394 = pi09796 & ~w28338;
assign w43395 = ~pi09848 & w28338;
assign w43396 = ~w43394 & ~w43395;
assign w43397 = pi09797 & ~w35929;
assign w43398 = ~pi02721 & w35929;
assign w43399 = ~w43397 & ~w43398;
assign w43400 = w1242 & w11485;
assign w43401 = pi09798 & ~w43400;
assign w43402 = pi10595 & w43400;
assign w43403 = ~w43401 & ~w43402;
assign w43404 = w1230 & w11485;
assign w43405 = pi09799 & ~w43404;
assign w43406 = pi10596 & w43404;
assign w43407 = ~w43405 & ~w43406;
assign w43408 = pi09800 & ~w43404;
assign w43409 = pi10592 & w43404;
assign w43410 = ~w43408 & ~w43409;
assign w43411 = w1217 & w19266;
assign w43412 = pi09801 & ~w43411;
assign w43413 = pi10602 & w43411;
assign w43414 = ~w43412 & ~w43413;
assign w43415 = pi09802 & ~w22154;
assign w43416 = ~pi09802 & ~pi09867;
assign w43417 = ~w16788 & ~w43416;
assign w43418 = w16800 & w43417;
assign w43419 = ~w43415 & ~w43418;
assign w43420 = w1235 & w11485;
assign w43421 = pi09803 & ~w43420;
assign w43422 = pi10593 & w43420;
assign w43423 = ~w43421 & ~w43422;
assign w43424 = pi09804 & ~w43420;
assign w43425 = pi10591 & w43420;
assign w43426 = ~w43424 & ~w43425;
assign w43427 = w1275 & w11485;
assign w43428 = pi09805 & ~w43427;
assign w43429 = pi10593 & w43427;
assign w43430 = ~w43428 & ~w43429;
assign w43431 = pi09976 & w12912;
assign w43432 = pi09894 & w12906;
assign w43433 = pi09902 & w12902;
assign w43434 = pi00857 & pi09806;
assign w43435 = pi09985 & w12908;
assign w43436 = pi02803 & w12910;
assign w43437 = pi02050 & w12897;
assign w43438 = pi01473 & w12915;
assign w43439 = pi09892 & w12854;
assign w43440 = ~w14236 & ~w43434;
assign w43441 = ~w43432 & w43440;
assign w43442 = ~w43433 & ~w43435;
assign w43443 = ~w43436 & w43442;
assign w43444 = ~w43437 & w43441;
assign w43445 = ~w43438 & w43444;
assign w43446 = ~w43431 & w43443;
assign w43447 = ~w43439 & w43446;
assign w43448 = w43445 & w43447;
assign w43449 = pi09885 & w12854;
assign w43450 = pi02798 & w12910;
assign w43451 = pi09897 & w12902;
assign w43452 = pi00857 & pi09807;
assign w43453 = pi09942 & w12908;
assign w43454 = pi09876 & w12906;
assign w43455 = pi01469 & w12915;
assign w43456 = pi02788 & w12897;
assign w43457 = pi09946 & w12912;
assign w43458 = ~w14236 & ~w43452;
assign w43459 = ~w43450 & w43458;
assign w43460 = ~w43451 & ~w43453;
assign w43461 = ~w43454 & w43460;
assign w43462 = ~w43455 & w43459;
assign w43463 = ~w43456 & w43462;
assign w43464 = ~w43449 & w43461;
assign w43465 = ~w43457 & w43464;
assign w43466 = w43463 & w43465;
assign w43467 = pi09808 & ~w43427;
assign w43468 = pi10596 & w43427;
assign w43469 = ~w43467 & ~w43468;
assign w43470 = pi09809 & ~w43427;
assign w43471 = pi10591 & w43427;
assign w43472 = ~w43470 & ~w43471;
assign w43473 = w1237 & w19266;
assign w43474 = pi09810 & ~w43473;
assign w43475 = pi10602 & w43473;
assign w43476 = ~w43474 & ~w43475;
assign w43477 = pi09811 & ~w43473;
assign w43478 = pi10599 & w43473;
assign w43479 = ~w43477 & ~w43478;
assign w43480 = pi00138 & w19710;
assign w43481 = pi10602 & w19704;
assign w43482 = ~pi09812 & w19713;
assign w43483 = ~w43480 & ~w43481;
assign w43484 = ~w43482 & w43483;
assign w43485 = w1266 & w16143;
assign w43486 = pi09813 & ~w43485;
assign w43487 = pi10608 & w43485;
assign w43488 = ~w43486 & ~w43487;
assign w43489 = pi09814 & ~w43485;
assign w43490 = pi10606 & w43485;
assign w43491 = ~w43489 & ~w43490;
assign w43492 = w1222 & w19266;
assign w43493 = pi09815 & ~w43492;
assign w43494 = ~pi10602 & w43492;
assign w43495 = ~w43493 & ~w43494;
assign w43496 = w1222 & w11485;
assign w43497 = pi09816 & ~w43496;
assign w43498 = pi10597 & w43496;
assign w43499 = ~w43497 & ~w43498;
assign w43500 = pi09817 & ~w43496;
assign w43501 = pi10594 & w43496;
assign w43502 = ~w43500 & ~w43501;
assign w43503 = pi09818 & w12993;
assign w43504 = ~w12989 & w43503;
assign w43505 = w12989 & ~w43503;
assign w43506 = ~w43504 & ~w43505;
assign w43507 = pi00188 & pi09969;
assign w43508 = pi09819 & pi09963;
assign w43509 = w72 & w43508;
assign w43510 = ~w43507 & ~w43509;
assign w43511 = pi09912 & w17066;
assign w43512 = ~pi09819 & ~w43511;
assign w43513 = pi09819 & w43511;
assign w43514 = w43510 & ~w43512;
assign w43515 = ~w43513 & w43514;
assign w43516 = ~pi01305 & ~w14146;
assign w43517 = pi01309 & ~w43516;
assign w43518 = ~pi01306 & ~w43517;
assign w43519 = ~pi00957 & ~w43518;
assign w43520 = pi00962 & ~w43519;
assign w43521 = w11342 & ~w43520;
assign w43522 = pi09820 & ~w11342;
assign w43523 = ~w43521 & ~w43522;
assign w43524 = w671 & ~w793;
assign w43525 = ~pi09822 & ~w21569;
assign w43526 = ~w21570 & ~w43525;
assign w43527 = w21576 & w43526;
assign w43528 = pi09823 & ~w19704;
assign w43529 = w1209 & w19704;
assign w43530 = ~pi10578 & pi10662;
assign w43531 = w43529 & w43530;
assign w43532 = ~w43528 & ~w43531;
assign w43533 = pi09824 & ~w11342;
assign w43534 = pi00486 & pi01249;
assign w43535 = w11342 & w43534;
assign w43536 = ~w43533 & ~w43535;
assign w43537 = ~pi09825 & ~w16030;
assign w43538 = w12993 & ~w16223;
assign w43539 = ~w43537 & w43538;
assign w43540 = pi09826 & ~w43496;
assign w43541 = pi10590 & w43496;
assign w43542 = ~w43540 & ~w43541;
assign w43543 = pi09827 & ~w43496;
assign w43544 = pi10591 & w43496;
assign w43545 = ~w43543 & ~w43544;
assign w43546 = pi09828 & ~w43496;
assign w43547 = pi10592 & w43496;
assign w43548 = ~w43546 & ~w43547;
assign w43549 = pi09829 & ~w43496;
assign w43550 = pi10593 & w43496;
assign w43551 = ~w43549 & ~w43550;
assign w43552 = pi09830 & ~w43496;
assign w43553 = pi10595 & w43496;
assign w43554 = ~w43552 & ~w43553;
assign w43555 = pi09831 & ~w43496;
assign w43556 = pi10596 & w43496;
assign w43557 = ~w43555 & ~w43556;
assign w43558 = pi09832 & ~w43492;
assign w43559 = pi10598 & w43492;
assign w43560 = ~w43558 & ~w43559;
assign w43561 = pi09833 & ~w43492;
assign w43562 = ~pi10599 & w43492;
assign w43563 = ~w43561 & ~w43562;
assign w43564 = pi09834 & ~w43492;
assign w43565 = ~pi10600 & w43492;
assign w43566 = ~w43564 & ~w43565;
assign w43567 = pi09835 & ~w43492;
assign w43568 = ~pi10601 & w43492;
assign w43569 = ~w43567 & ~w43568;
assign w43570 = pi09836 & ~w43492;
assign w43571 = ~pi10604 & w43492;
assign w43572 = ~w43570 & ~w43571;
assign w43573 = pi09837 & ~w43492;
assign w43574 = ~pi10605 & w43492;
assign w43575 = ~w43573 & ~w43574;
assign w43576 = pi09838 & ~w43492;
assign w43577 = ~pi10603 & w43492;
assign w43578 = ~w43576 & ~w43577;
assign w43579 = pi09839 & w19713;
assign w43580 = ~w19710 & ~w43579;
assign w43581 = w1266 & w11485;
assign w43582 = pi09840 & ~w43581;
assign w43583 = ~pi10591 & w43581;
assign w43584 = ~w43582 & ~w43583;
assign w43585 = pi09841 & ~w43581;
assign w43586 = ~pi10592 & w43581;
assign w43587 = ~w43585 & ~w43586;
assign w43588 = pi09842 & ~w43581;
assign w43589 = pi10593 & w43581;
assign w43590 = ~w43588 & ~w43589;
assign w43591 = pi09843 & ~w43581;
assign w43592 = ~pi10594 & w43581;
assign w43593 = ~w43591 & ~w43592;
assign w43594 = pi09844 & ~w43581;
assign w43595 = ~pi10595 & w43581;
assign w43596 = ~w43594 & ~w43595;
assign w43597 = pi09845 & ~w43581;
assign w43598 = ~pi10590 & w43581;
assign w43599 = ~w43597 & ~w43598;
assign w43600 = pi09846 & ~w43485;
assign w43601 = pi10607 & w43485;
assign w43602 = ~w43600 & ~w43601;
assign w43603 = pi09847 & ~w43485;
assign w43604 = pi10609 & w43485;
assign w43605 = ~w43603 & ~w43604;
assign w43606 = pi00137 & w19710;
assign w43607 = pi10601 & w19704;
assign w43608 = ~pi09848 & w19713;
assign w43609 = ~w43606 & ~w43607;
assign w43610 = ~w43608 & w43609;
assign w43611 = w1237 & w11485;
assign w43612 = pi09849 & ~w43611;
assign w43613 = pi10590 & w43611;
assign w43614 = ~w43612 & ~w43613;
assign w43615 = pi09850 & ~w43611;
assign w43616 = pi10591 & w43611;
assign w43617 = ~w43615 & ~w43616;
assign w43618 = pi09851 & ~w43611;
assign w43619 = pi10592 & w43611;
assign w43620 = ~w43618 & ~w43619;
assign w43621 = pi09852 & ~w43611;
assign w43622 = ~pi10593 & w43611;
assign w43623 = ~w43621 & ~w43622;
assign w43624 = pi09853 & ~w43611;
assign w43625 = ~pi10594 & w43611;
assign w43626 = ~w43624 & ~w43625;
assign w43627 = pi09854 & ~w43473;
assign w43628 = pi10598 & w43473;
assign w43629 = ~w43627 & ~w43628;
assign w43630 = w16004 & ~w16224;
assign w43631 = ~w16225 & ~w43630;
assign w43632 = ~pi09856 & ~w16223;
assign w43633 = w12993 & ~w16224;
assign w43634 = ~w43632 & w43633;
assign w43635 = pi09857 & ~w43473;
assign w43636 = pi10601 & w43473;
assign w43637 = ~w43635 & ~w43636;
assign w43638 = pi09858 & ~w43473;
assign w43639 = pi10600 & w43473;
assign w43640 = ~w43638 & ~w43639;
assign w43641 = pi09859 & ~w43427;
assign w43642 = ~pi10590 & w43427;
assign w43643 = ~w43641 & ~w43642;
assign w43644 = pi09860 & ~w43427;
assign w43645 = pi10592 & w43427;
assign w43646 = ~w43644 & ~w43645;
assign w43647 = pi09861 & ~w43427;
assign w43648 = pi10594 & w43427;
assign w43649 = ~w43647 & ~w43648;
assign w43650 = pi09862 & ~w43427;
assign w43651 = pi10595 & w43427;
assign w43652 = ~w43650 & ~w43651;
assign w43653 = w1275 & w19266;
assign w43654 = pi10598 & w43653;
assign w43655 = pi09863 & ~w43653;
assign w43656 = ~w43654 & ~w43655;
assign w43657 = pi09864 & ~w43427;
assign w43658 = pi10597 & w43427;
assign w43659 = ~w43657 & ~w43658;
assign w43660 = ~pi10379 & pi10418;
assign w43661 = pi00539 & ~pi10418;
assign w43662 = ~pi00845 & ~pi10481;
assign w43663 = ~w43660 & ~w43661;
assign w43664 = w43662 & w43663;
assign w43665 = pi01170 & ~pi09924;
assign w43666 = ~w43664 & w43665;
assign w43667 = pi10000 & ~w43666;
assign w43668 = ~pi09865 & ~w11194;
assign w43669 = pi00439 & w11194;
assign w43670 = ~w43667 & ~w43668;
assign w43671 = ~w43669 & w43670;
assign w43672 = pi01455 & w16808;
assign w43673 = ~pi09866 & ~w43672;
assign w43674 = ~w16797 & ~w43673;
assign w43675 = ~pi09867 & ~w16807;
assign w43676 = pi09867 & w22154;
assign w43677 = ~w43675 & ~w43676;
assign w43678 = pi09868 & ~w43420;
assign w43679 = pi10590 & w43420;
assign w43680 = ~w43678 & ~w43679;
assign w43681 = pi09869 & ~w43420;
assign w43682 = ~pi10592 & w43420;
assign w43683 = ~w43681 & ~w43682;
assign w43684 = pi09870 & ~w43420;
assign w43685 = ~pi10594 & w43420;
assign w43686 = ~w43684 & ~w43685;
assign w43687 = pi09871 & ~w43420;
assign w43688 = pi10595 & w43420;
assign w43689 = ~w43687 & ~w43688;
assign w43690 = pi09872 & ~w43420;
assign w43691 = pi10597 & w43420;
assign w43692 = ~w43690 & ~w43691;
assign w43693 = pi09873 & ~w43420;
assign w43694 = pi10596 & w43420;
assign w43695 = ~w43693 & ~w43694;
assign w43696 = pi09874 & ~w43411;
assign w43697 = pi10598 & w43411;
assign w43698 = ~w43696 & ~w43697;
assign w43699 = w1235 & w16143;
assign w43700 = pi10606 & w43699;
assign w43701 = pi09875 & ~w43699;
assign w43702 = ~w43700 & ~w43701;
assign w43703 = pi09876 & ~w43411;
assign w43704 = pi10599 & w43411;
assign w43705 = ~w43703 & ~w43704;
assign w43706 = pi09877 & ~w43404;
assign w43707 = pi10590 & w43404;
assign w43708 = ~w43706 & ~w43707;
assign w43709 = pi09878 & ~w43411;
assign w43710 = pi10600 & w43411;
assign w43711 = ~w43709 & ~w43710;
assign w43712 = pi09879 & ~w43404;
assign w43713 = pi10591 & w43404;
assign w43714 = ~w43712 & ~w43713;
assign w43715 = pi09880 & ~w43411;
assign w43716 = pi10601 & w43411;
assign w43717 = ~w43715 & ~w43716;
assign w43718 = pi09881 & ~w43404;
assign w43719 = pi10593 & w43404;
assign w43720 = ~w43718 & ~w43719;
assign w43721 = pi09882 & ~w43404;
assign w43722 = pi10594 & w43404;
assign w43723 = ~w43721 & ~w43722;
assign w43724 = pi09883 & ~w43404;
assign w43725 = pi10595 & w43404;
assign w43726 = ~w43724 & ~w43725;
assign w43727 = w1232 & w11485;
assign w43728 = pi09884 & ~w43727;
assign w43729 = pi10590 & w43727;
assign w43730 = ~w43728 & ~w43729;
assign w43731 = pi09885 & ~w43727;
assign w43732 = pi10591 & w43727;
assign w43733 = ~w43731 & ~w43732;
assign w43734 = pi09886 & ~w43727;
assign w43735 = pi10592 & w43727;
assign w43736 = ~w43734 & ~w43735;
assign w43737 = pi09887 & ~w43727;
assign w43738 = pi10593 & w43727;
assign w43739 = ~w43737 & ~w43738;
assign w43740 = pi09888 & ~w43404;
assign w43741 = pi10597 & w43404;
assign w43742 = ~w43740 & ~w43741;
assign w43743 = pi09889 & ~w43727;
assign w43744 = pi10594 & w43727;
assign w43745 = ~w43743 & ~w43744;
assign w43746 = pi09890 & ~w43727;
assign w43747 = pi10595 & w43727;
assign w43748 = ~w43746 & ~w43747;
assign w43749 = pi09891 & ~w43411;
assign w43750 = pi10603 & w43411;
assign w43751 = ~w43749 & ~w43750;
assign w43752 = pi09892 & ~w43727;
assign w43753 = pi10596 & w43727;
assign w43754 = ~w43752 & ~w43753;
assign w43755 = pi09893 & ~w43727;
assign w43756 = pi10597 & w43727;
assign w43757 = ~w43755 & ~w43756;
assign w43758 = pi09894 & ~w43411;
assign w43759 = pi10604 & w43411;
assign w43760 = ~w43758 & ~w43759;
assign w43761 = pi09895 & ~w43411;
assign w43762 = pi10605 & w43411;
assign w43763 = ~w43761 & ~w43762;
assign w43764 = w1217 & w16143;
assign w43765 = pi09896 & ~w43764;
assign w43766 = pi10606 & w43764;
assign w43767 = ~w43765 & ~w43766;
assign w43768 = pi09897 & ~w43764;
assign w43769 = pi10607 & w43764;
assign w43770 = ~w43768 & ~w43769;
assign w43771 = pi09898 & ~w43764;
assign w43772 = pi10608 & w43764;
assign w43773 = ~w43771 & ~w43772;
assign w43774 = pi09899 & ~w43764;
assign w43775 = pi10609 & w43764;
assign w43776 = ~w43774 & ~w43775;
assign w43777 = pi09900 & ~w43764;
assign w43778 = pi10610 & w43764;
assign w43779 = ~w43777 & ~w43778;
assign w43780 = pi09901 & ~w43764;
assign w43781 = pi10611 & w43764;
assign w43782 = ~w43780 & ~w43781;
assign w43783 = pi09902 & ~w43764;
assign w43784 = pi10612 & w43764;
assign w43785 = ~w43783 & ~w43784;
assign w43786 = pi09903 & ~w43764;
assign w43787 = pi10613 & w43764;
assign w43788 = ~w43786 & ~w43787;
assign w43789 = w1244 & w11485;
assign w43790 = pi09904 & ~w43789;
assign w43791 = pi10590 & w43789;
assign w43792 = ~w43790 & ~w43791;
assign w43793 = pi09905 & ~w43789;
assign w43794 = pi10591 & w43789;
assign w43795 = ~w43793 & ~w43794;
assign w43796 = pi09906 & ~w43789;
assign w43797 = pi10592 & w43789;
assign w43798 = ~w43796 & ~w43797;
assign w43799 = pi09907 & ~w43789;
assign w43800 = pi10593 & w43789;
assign w43801 = ~w43799 & ~w43800;
assign w43802 = pi09908 & ~w43789;
assign w43803 = pi10594 & w43789;
assign w43804 = ~w43802 & ~w43803;
assign w43805 = pi09909 & ~w43789;
assign w43806 = pi10595 & w43789;
assign w43807 = ~w43805 & ~w43806;
assign w43808 = pi09910 & ~w43789;
assign w43809 = pi10596 & w43789;
assign w43810 = ~w43808 & ~w43809;
assign w43811 = pi09911 & ~w43789;
assign w43812 = pi10597 & w43789;
assign w43813 = ~w43811 & ~w43812;
assign w43814 = ~pi09912 & ~w17066;
assign w43815 = w43510 & ~w43511;
assign w43816 = ~w43814 & w43815;
assign w43817 = pi09913 & ~w43400;
assign w43818 = pi10590 & w43400;
assign w43819 = ~w43817 & ~w43818;
assign w43820 = pi09914 & ~w43400;
assign w43821 = pi10591 & w43400;
assign w43822 = ~w43820 & ~w43821;
assign w43823 = pi09915 & ~w43400;
assign w43824 = pi10592 & w43400;
assign w43825 = ~w43823 & ~w43824;
assign w43826 = pi09916 & ~w43400;
assign w43827 = pi10593 & w43400;
assign w43828 = ~w43826 & ~w43827;
assign w43829 = pi09917 & ~w43400;
assign w43830 = pi10594 & w43400;
assign w43831 = ~w43829 & ~w43830;
assign w43832 = pi09918 & ~w43400;
assign w43833 = pi10596 & w43400;
assign w43834 = ~w43832 & ~w43833;
assign w43835 = pi09919 & ~w43400;
assign w43836 = pi10597 & w43400;
assign w43837 = ~w43835 & ~w43836;
assign w43838 = pi09889 & w12854;
assign w43839 = pi09900 & w12902;
assign w43840 = pi09939 & w12908;
assign w43841 = pi00857 & pi09920;
assign w43842 = pi02789 & w12897;
assign w43843 = pi01472 & w12915;
assign w43844 = pi09801 & w12906;
assign w43845 = pi02801 & w12910;
assign w43846 = pi09975 & w12912;
assign w43847 = ~w43839 & ~w43841;
assign w43848 = ~w43840 & ~w43844;
assign w43849 = ~w43845 & w43848;
assign w43850 = ~w43842 & w43847;
assign w43851 = ~w43843 & w43850;
assign w43852 = ~w43838 & w43849;
assign w43853 = ~w43846 & w43852;
assign w43854 = w43851 & w43853;
assign w43855 = pi09886 & w12854;
assign w43856 = pi09898 & w12902;
assign w43857 = pi09878 & w12906;
assign w43858 = pi00857 & pi09921;
assign w43859 = pi01470 & w12915;
assign w43860 = pi02053 & w12897;
assign w43861 = pi09982 & w12908;
assign w43862 = pi02799 & w12910;
assign w43863 = pi09943 & w12912;
assign w43864 = ~w43856 & ~w43858;
assign w43865 = ~w43857 & ~w43861;
assign w43866 = ~w43862 & w43865;
assign w43867 = ~w43859 & w43864;
assign w43868 = ~w43860 & w43867;
assign w43869 = ~w43855 & w43866;
assign w43870 = ~w43863 & w43869;
assign w43871 = w43868 & w43870;
assign w43872 = pi09945 & w12912;
assign w43873 = pi09891 & w12906;
assign w43874 = pi02802 & w12910;
assign w43875 = pi00857 & pi09922;
assign w43876 = pi01476 & w12915;
assign w43877 = pi02790 & w12897;
assign w43878 = pi09984 & w12908;
assign w43879 = pi09901 & w12902;
assign w43880 = pi09890 & w12854;
assign w43881 = ~w43873 & ~w43875;
assign w43882 = ~w43874 & ~w43878;
assign w43883 = ~w43879 & w43882;
assign w43884 = ~w43876 & w43881;
assign w43885 = ~w43877 & w43884;
assign w43886 = ~w43872 & w43883;
assign w43887 = ~w43880 & w43886;
assign w43888 = w43885 & w43887;
assign w43889 = pi09923 & ~w2431;
assign w43890 = ~pi00188 & ~w43889;
assign w43891 = pi10518 & ~w43664;
assign w43892 = ~pi00445 & ~pi01271;
assign w43893 = pi00445 & pi01271;
assign w43894 = ~w43892 & ~w43893;
assign w43895 = pi00446 & w43894;
assign w43896 = pi01270 & ~w43894;
assign w43897 = ~pi00446 & ~pi01270;
assign w43898 = pi09865 & ~pi09924;
assign w43899 = ~w43897 & w43898;
assign w43900 = ~w43895 & w43899;
assign w43901 = ~w43896 & w43900;
assign w43902 = pi10000 & ~w43901;
assign w43903 = ~pi09924 & ~pi10000;
assign w43904 = w43891 & ~w43903;
assign w43905 = ~w43902 & w43904;
assign w43906 = pi02665 & ~pi09925;
assign w43907 = pi10418 & w43906;
assign w43908 = pi10002 & w43907;
assign w43909 = pi09930 & w43908;
assign w43910 = ~pi09925 & ~w43909;
assign w43911 = w12845 & ~w43910;
assign w43912 = ~pi09926 & ~w17065;
assign w43913 = ~w17066 & ~w43912;
assign w43914 = w43510 & w43913;
assign w43915 = ~pi10389 & pi10467;
assign w43916 = ~w12722 & w43915;
assign w43917 = pi09927 & ~w43916;
assign w43918 = pi09927 & ~w16775;
assign w43919 = pi09996 & ~w43918;
assign w43920 = pi00062 & w43919;
assign w43921 = ~w43917 & ~w43920;
assign w43922 = pi10450 & pi10494;
assign w43923 = w12878 & ~w43922;
assign w43924 = ~pi10345 & ~w43923;
assign w43925 = pi00090 & pi09928;
assign w43926 = ~w43924 & ~w43925;
assign w43927 = pi09929 & ~w11160;
assign w43928 = pi00033 & w16188;
assign w43929 = pi10399 & w13021;
assign w43930 = ~w43928 & w43929;
assign w43931 = ~w43927 & ~w43930;
assign w43932 = ~pi09930 & ~w43908;
assign w43933 = w12845 & ~w43909;
assign w43934 = ~w43932 & w43933;
assign w43935 = pi00025 & ~pi00963;
assign w43936 = w504 & ~w43935;
assign w43937 = ~pi00028 & w14204;
assign w43938 = ~w43936 & ~w43937;
assign w43939 = w715 & w43938;
assign w43940 = w1242 & w19266;
assign w43941 = pi09934 & ~w43940;
assign w43942 = pi10603 & w43940;
assign w43943 = ~w43941 & ~w43942;
assign w43944 = pi09935 & ~w43940;
assign w43945 = pi10601 & w43940;
assign w43946 = ~w43944 & ~w43945;
assign w43947 = pi09936 & ~w43940;
assign w43948 = pi10599 & w43940;
assign w43949 = ~w43947 & ~w43948;
assign w43950 = w1244 & w19266;
assign w43951 = pi09937 & ~w43950;
assign w43952 = pi10605 & w43950;
assign w43953 = ~w43951 & ~w43952;
assign w43954 = pi09938 & ~w43950;
assign w43955 = pi10602 & w43950;
assign w43956 = ~w43954 & ~w43955;
assign w43957 = pi10667 & w11484;
assign w43958 = w1217 & w43957;
assign w43959 = pi09939 & ~w43958;
assign w43960 = pi10618 & w43958;
assign w43961 = ~w43959 & ~w43960;
assign w43962 = pi09940 & ~w43950;
assign w43963 = pi10599 & w43950;
assign w43964 = ~w43962 & ~w43963;
assign w43965 = pi09941 & ~w43958;
assign w43966 = pi10617 & w43958;
assign w43967 = ~w43965 & ~w43966;
assign w43968 = pi09942 & ~w43958;
assign w43969 = pi10615 & w43958;
assign w43970 = ~w43968 & ~w43969;
assign w43971 = w1232 & w19266;
assign w43972 = pi09943 & ~w43971;
assign w43973 = pi10600 & w43971;
assign w43974 = ~w43972 & ~w43973;
assign w43975 = w1230 & w19266;
assign w43976 = pi09944 & ~w43975;
assign w43977 = pi10603 & w43975;
assign w43978 = ~w43976 & ~w43977;
assign w43979 = pi09945 & ~w43971;
assign w43980 = pi10603 & w43971;
assign w43981 = ~w43979 & ~w43980;
assign w43982 = pi09946 & ~w43971;
assign w43983 = pi10599 & w43971;
assign w43984 = ~w43982 & ~w43983;
assign w43985 = pi09947 & ~w43971;
assign w43986 = pi10598 & w43971;
assign w43987 = ~w43985 & ~w43986;
assign w43988 = pi09948 & ~w43975;
assign w43989 = pi10598 & w43975;
assign w43990 = ~w43988 & ~w43989;
assign w43991 = w1235 & w19266;
assign w43992 = pi09949 & ~w43991;
assign w43993 = pi10604 & w43991;
assign w43994 = ~w43992 & ~w43993;
assign w43995 = pi09950 & ~w43991;
assign w43996 = pi10603 & w43991;
assign w43997 = ~w43995 & ~w43996;
assign w43998 = pi09951 & ~w43991;
assign w43999 = pi10601 & w43991;
assign w44000 = ~w43998 & ~w43999;
assign w44001 = pi09952 & ~w43991;
assign w44002 = pi10598 & w43991;
assign w44003 = ~w44001 & ~w44002;
assign w44004 = ~pi09953 & ~w19704;
assign w44005 = ~w19707 & ~w19710;
assign w44006 = ~w44004 & w44005;
assign w44007 = ~pi09954 & w19713;
assign w44008 = pi10605 & w19704;
assign w44009 = ~w44007 & ~w44008;
assign w44010 = pi09818 & w12989;
assign w44011 = ~pi09955 & ~w44010;
assign w44012 = pi09955 & w44010;
assign w44013 = w12993 & ~w44011;
assign w44014 = ~w44012 & w44013;
assign w44015 = pi09956 & ~w11342;
assign w44016 = ~pi09824 & w11342;
assign w44017 = ~w44015 & ~w44016;
assign w44018 = pi09957 & ~w11342;
assign w44019 = ~pi09959 & w11342;
assign w44020 = ~w44018 & ~w44019;
assign w44021 = ~pi09958 & ~w44012;
assign w44022 = pi09958 & w44012;
assign w44023 = w12993 & ~w44022;
assign w44024 = ~w44021 & w44023;
assign w44025 = pi09959 & ~w11342;
assign w44026 = pi09820 & w11342;
assign w44027 = ~w44025 & ~w44026;
assign w44028 = pi09960 & w44023;
assign w44029 = w12989 & w14879;
assign w44030 = ~w44028 & ~w44029;
assign w44031 = ~pi09961 & w19713;
assign w44032 = pi10600 & w19704;
assign w44033 = ~w44031 & ~w44032;
assign w44034 = ~pi09962 & w19713;
assign w44035 = pi10599 & w19704;
assign w44036 = ~w44034 & ~w44035;
assign w44037 = ~pi09963 & ~w75;
assign w44038 = ~w17065 & ~w44037;
assign w44039 = ~w43507 & ~w44038;
assign w44040 = ~w43509 & ~w44039;
assign w44041 = ~pi09865 & w11194;
assign w44042 = ~pi10424 & pi10463;
assign w44043 = ~pi09965 & ~w44042;
assign w44044 = w12119 & ~w44043;
assign w44045 = ~w44041 & w44044;
assign w44046 = pi09966 & w19711;
assign w44047 = ~w19712 & ~w44046;
assign w44048 = pi09967 & ~w43991;
assign w44049 = pi10600 & w43991;
assign w44050 = ~w44048 & ~w44049;
assign w44051 = pi09968 & ~w43991;
assign w44052 = pi10599 & w43991;
assign w44053 = ~w44051 & ~w44052;
assign w44054 = pi09969 & ~w43991;
assign w44055 = pi10602 & w43991;
assign w44056 = ~w44054 & ~w44055;
assign w44057 = pi09970 & ~w43991;
assign w44058 = pi10605 & w43991;
assign w44059 = ~w44057 & ~w44058;
assign w44060 = pi09971 & ~w43975;
assign w44061 = pi10599 & w43975;
assign w44062 = ~w44060 & ~w44061;
assign w44063 = pi09972 & ~w43975;
assign w44064 = pi10600 & w43975;
assign w44065 = ~w44063 & ~w44064;
assign w44066 = pi09973 & ~w43971;
assign w44067 = pi10601 & w43971;
assign w44068 = ~w44066 & ~w44067;
assign w44069 = pi09974 & ~w43975;
assign w44070 = pi10601 & w43975;
assign w44071 = ~w44069 & ~w44070;
assign w44072 = pi09975 & ~w43971;
assign w44073 = pi10602 & w43971;
assign w44074 = ~w44072 & ~w44073;
assign w44075 = pi09976 & ~w43971;
assign w44076 = pi10604 & w43971;
assign w44077 = ~w44075 & ~w44076;
assign w44078 = pi09977 & ~w43971;
assign w44079 = pi10605 & w43971;
assign w44080 = ~w44078 & ~w44079;
assign w44081 = pi09978 & ~w43975;
assign w44082 = pi10602 & w43975;
assign w44083 = ~w44081 & ~w44082;
assign w44084 = pi09979 & ~w43975;
assign w44085 = pi10604 & w43975;
assign w44086 = ~w44084 & ~w44085;
assign w44087 = pi09980 & ~w43975;
assign w44088 = pi10605 & w43975;
assign w44089 = ~w44087 & ~w44088;
assign w44090 = pi09981 & ~w43958;
assign w44091 = pi10614 & w43958;
assign w44092 = ~w44090 & ~w44091;
assign w44093 = pi09982 & ~w43958;
assign w44094 = pi10616 & w43958;
assign w44095 = ~w44093 & ~w44094;
assign w44096 = pi09983 & ~w43950;
assign w44097 = pi10598 & w43950;
assign w44098 = ~w44096 & ~w44097;
assign w44099 = pi09984 & ~w43958;
assign w44100 = pi10619 & w43958;
assign w44101 = ~w44099 & ~w44100;
assign w44102 = pi09985 & ~w43958;
assign w44103 = pi10620 & w43958;
assign w44104 = ~w44102 & ~w44103;
assign w44105 = pi09986 & ~w43950;
assign w44106 = pi10600 & w43950;
assign w44107 = ~w44105 & ~w44106;
assign w44108 = pi09987 & ~w43950;
assign w44109 = pi10601 & w43950;
assign w44110 = ~w44108 & ~w44109;
assign w44111 = pi09988 & ~w43958;
assign w44112 = pi10621 & w43958;
assign w44113 = ~w44111 & ~w44112;
assign w44114 = pi09989 & ~w43950;
assign w44115 = pi10603 & w43950;
assign w44116 = ~w44114 & ~w44115;
assign w44117 = pi09990 & ~w43950;
assign w44118 = pi10604 & w43950;
assign w44119 = ~w44117 & ~w44118;
assign w44120 = pi09991 & ~w43940;
assign w44121 = pi10598 & w43940;
assign w44122 = ~w44120 & ~w44121;
assign w44123 = pi09992 & ~w43940;
assign w44124 = pi10600 & w43940;
assign w44125 = ~w44123 & ~w44124;
assign w44126 = pi09993 & ~w43940;
assign w44127 = pi10602 & w43940;
assign w44128 = ~w44126 & ~w44127;
assign w44129 = pi09994 & ~w43940;
assign w44130 = pi10604 & w43940;
assign w44131 = ~w44129 & ~w44130;
assign w44132 = pi09995 & ~w43940;
assign w44133 = pi10605 & w43940;
assign w44134 = ~w44132 & ~w44133;
assign w44135 = ~pi00062 & ~pi09996;
assign w44136 = ~w43920 & ~w44135;
assign w44137 = ~pi09997 & ~w43919;
assign w44138 = pi00062 & ~w44137;
assign w44139 = pi09998 & ~w19704;
assign w44140 = pi10578 & pi10662;
assign w44141 = w43529 & w44140;
assign w44142 = pi10667 & w44141;
assign w44143 = ~w44139 & ~w44142;
assign w44144 = pi00869 & ~w1448;
assign w44145 = ~pi00869 & ~pi09999;
assign w44146 = ~w44144 & ~w44145;
assign w44147 = ~pi10000 & ~w11126;
assign w44148 = ~pi10378 & pi10418;
assign w44149 = pi00053 & ~pi10418;
assign w44150 = w43662 & ~w44148;
assign w44151 = ~w44149 & w44150;
assign w44152 = ~w11180 & ~w44147;
assign w44153 = ~w44151 & w44152;
assign w44154 = w43891 & w44153;
assign w44155 = pi10428 & pi10459;
assign w44156 = ~pi10001 & ~w44155;
assign w44157 = ~pi10439 & ~w44156;
assign w44158 = ~pi10002 & ~w43907;
assign w44159 = w12845 & ~w43908;
assign w44160 = ~w44158 & w44159;
assign w44161 = pi10003 & ~w16006;
assign w44162 = ~pi10632 & w16006;
assign w44163 = ~w44161 & ~w44162;
assign w44164 = w12984 & w12988;
assign w44165 = pi10004 & ~w44164;
assign w44166 = ~w828 & ~w44165;
assign w44167 = w11707 & w11708;
assign w44168 = pi10005 & ~w44167;
assign w44169 = ~w12877 & ~w44168;
assign w44170 = ~pi10006 & ~pi10454;
assign w44171 = ~w11127 & ~w14863;
assign w44172 = ~pi00062 & ~pi00438;
assign w44173 = ~w44171 & w44172;
assign w44174 = ~w44170 & ~w44173;
assign w44175 = w1242 & w43957;
assign w44176 = pi10007 & ~w44175;
assign w44177 = pi10619 & w44175;
assign w44178 = ~w44176 & ~w44177;
assign w44179 = pi10008 & ~w44175;
assign w44180 = pi10621 & w44175;
assign w44181 = ~w44179 & ~w44180;
assign w44182 = pi10009 & ~w44175;
assign w44183 = pi10618 & w44175;
assign w44184 = ~w44182 & ~w44183;
assign w44185 = pi10010 & ~w44175;
assign w44186 = pi10616 & w44175;
assign w44187 = ~w44185 & ~w44186;
assign w44188 = pi10011 & ~w44175;
assign w44189 = pi10614 & w44175;
assign w44190 = ~w44188 & ~w44189;
assign w44191 = w1242 & w16143;
assign w44192 = pi10012 & ~w44191;
assign w44193 = pi10612 & w44191;
assign w44194 = ~w44192 & ~w44193;
assign w44195 = w1244 & w43957;
assign w44196 = pi10013 & ~w44195;
assign w44197 = pi10616 & w44195;
assign w44198 = ~w44196 & ~w44197;
assign w44199 = pi10014 & ~w44191;
assign w44200 = pi10607 & w44191;
assign w44201 = ~w44199 & ~w44200;
assign w44202 = pi10015 & ~w44195;
assign w44203 = pi10620 & w44195;
assign w44204 = ~w44202 & ~w44203;
assign w44205 = pi10440 & ~w1210;
assign w44206 = ~pi10016 & ~w44205;
assign w44207 = pi10017 & ~w44195;
assign w44208 = pi10619 & w44195;
assign w44209 = ~w44207 & ~w44208;
assign w44210 = w1244 & w16143;
assign w44211 = pi10018 & ~w44210;
assign w44212 = pi10612 & w44210;
assign w44213 = ~w44211 & ~w44212;
assign w44214 = pi10019 & ~w44210;
assign w44215 = pi10609 & w44210;
assign w44216 = ~w44214 & ~w44215;
assign w44217 = w1230 & w43957;
assign w44218 = pi10021 & ~w44217;
assign w44219 = pi10617 & w44217;
assign w44220 = ~w44218 & ~w44219;
assign w44221 = pi10022 & ~w44217;
assign w44222 = pi10621 & w44217;
assign w44223 = ~w44221 & ~w44222;
assign w44224 = pi10023 & ~w44217;
assign w44225 = pi10614 & w44217;
assign w44226 = ~w44224 & ~w44225;
assign w44227 = w1230 & w16143;
assign w44228 = pi10024 & ~w44227;
assign w44229 = pi10613 & w44227;
assign w44230 = ~w44228 & ~w44229;
assign w44231 = pi10025 & ~w44227;
assign w44232 = pi10612 & w44227;
assign w44233 = ~w44231 & ~w44232;
assign w44234 = pi10026 & ~w44227;
assign w44235 = pi10607 & w44227;
assign w44236 = ~w44234 & ~w44235;
assign w44237 = pi10027 & ~w44227;
assign w44238 = pi10606 & w44227;
assign w44239 = ~w44237 & ~w44238;
assign w44240 = pi10028 & ~w19704;
assign w44241 = pi10665 & w44141;
assign w44242 = ~w44240 & ~w44241;
assign w44243 = pi10029 & ~w19704;
assign w44244 = pi10666 & w44141;
assign w44245 = ~w44243 & ~w44244;
assign w44246 = pi10266 & ~pi10406;
assign w44247 = ~w12722 & w44246;
assign w44248 = ~pi10030 & ~w44247;
assign w44249 = ~w14857 & ~w44248;
assign w44250 = pi10031 & pi10356;
assign w44251 = ~w11335 & ~w44250;
assign w44252 = pi09809 & pi09860;
assign w44253 = ~w14192 & ~w44252;
assign w44254 = w11341 & w44253;
assign w44255 = ~w44251 & ~w44254;
assign w44256 = pi10032 & ~w16271;
assign w44257 = ~pi10638 & w16271;
assign w44258 = ~w44256 & ~w44257;
assign w44259 = pi10033 & ~w16271;
assign w44260 = ~pi10625 & w16271;
assign w44261 = ~w44259 & ~w44260;
assign w44262 = pi10034 & ~w16271;
assign w44263 = ~pi10631 & w16271;
assign w44264 = ~w44262 & ~w44263;
assign w44265 = pi10035 & ~w16271;
assign w44266 = ~pi10628 & w16271;
assign w44267 = ~w44265 & ~w44266;
assign w44268 = pi10036 & ~w16271;
assign w44269 = ~pi10644 & w16271;
assign w44270 = ~w44268 & ~w44269;
assign w44271 = pi10037 & ~w16271;
assign w44272 = ~pi10650 & w16271;
assign w44273 = ~w44271 & ~w44272;
assign w44274 = pi10038 & ~w16271;
assign w44275 = ~pi10640 & w16271;
assign w44276 = ~w44274 & ~w44275;
assign w44277 = pi10039 & ~w16271;
assign w44278 = ~pi10633 & w16271;
assign w44279 = ~w44277 & ~w44278;
assign w44280 = pi10040 & ~w16219;
assign w44281 = ~pi10629 & w16219;
assign w44282 = ~w44280 & ~w44281;
assign w44283 = pi10041 & ~w16271;
assign w44284 = ~pi10622 & w16271;
assign w44285 = ~w44283 & ~w44284;
assign w44286 = pi10042 & ~w16219;
assign w44287 = ~pi10652 & w16219;
assign w44288 = ~w44286 & ~w44287;
assign w44289 = pi10043 & ~w16219;
assign w44290 = ~pi10644 & w16219;
assign w44291 = ~w44289 & ~w44290;
assign w44292 = pi10044 & ~w16219;
assign w44293 = ~pi10647 & w16219;
assign w44294 = ~w44292 & ~w44293;
assign w44295 = pi10045 & ~w16219;
assign w44296 = ~pi10648 & w16219;
assign w44297 = ~w44295 & ~w44296;
assign w44298 = pi10046 & ~w16219;
assign w44299 = ~pi10649 & w16219;
assign w44300 = ~w44298 & ~w44299;
assign w44301 = pi10048 & ~w16006;
assign w44302 = ~pi10634 & w16006;
assign w44303 = ~w44301 & ~w44302;
assign w44304 = pi10049 & ~w16225;
assign w44305 = ~pi10632 & w16225;
assign w44306 = ~w44304 & ~w44305;
assign w44307 = pi10050 & w523;
assign w44308 = ~pi09872 & ~pi09967;
assign w44309 = pi10452 & ~pi10587;
assign w44310 = w44308 & w44309;
assign w44311 = ~w535 & w44310;
assign w44312 = ~w44307 & ~w44311;
assign w44313 = pi10051 & ~w16225;
assign w44314 = ~pi10648 & w16225;
assign w44315 = ~w44313 & ~w44314;
assign w44316 = pi10052 & ~w16225;
assign w44317 = ~pi10629 & w16225;
assign w44318 = ~w44316 & ~w44317;
assign w44319 = pi10053 & ~w16219;
assign w44320 = ~pi10637 & w16219;
assign w44321 = ~w44319 & ~w44320;
assign w44322 = pi10054 & ~w16006;
assign w44323 = ~pi10622 & w16006;
assign w44324 = ~w44322 & ~w44323;
assign w44325 = pi10055 & ~w16006;
assign w44326 = ~pi10633 & w16006;
assign w44327 = ~w44325 & ~w44326;
assign w44328 = pi10056 & ~w16006;
assign w44329 = ~pi10638 & w16006;
assign w44330 = ~w44328 & ~w44329;
assign w44331 = pi10057 & ~w16006;
assign w44332 = ~pi10639 & w16006;
assign w44333 = ~w44331 & ~w44332;
assign w44334 = pi10058 & ~w16006;
assign w44335 = ~pi10641 & w16006;
assign w44336 = ~w44334 & ~w44335;
assign w44337 = pi10059 & ~w16006;
assign w44338 = ~pi10642 & w16006;
assign w44339 = ~w44337 & ~w44338;
assign w44340 = pi10060 & ~w16006;
assign w44341 = ~pi10643 & w16006;
assign w44342 = ~w44340 & ~w44341;
assign w44343 = pi10061 & ~w16006;
assign w44344 = ~pi10644 & w16006;
assign w44345 = ~w44343 & ~w44344;
assign w44346 = pi10062 & ~w16006;
assign w44347 = ~pi10646 & w16006;
assign w44348 = ~w44346 & ~w44347;
assign w44349 = pi10063 & ~w16006;
assign w44350 = ~pi10648 & w16006;
assign w44351 = ~w44349 & ~w44350;
assign w44352 = pi10064 & ~w16006;
assign w44353 = ~pi10624 & w16006;
assign w44354 = ~w44352 & ~w44353;
assign w44355 = pi10065 & ~w16006;
assign w44356 = ~pi10653 & w16006;
assign w44357 = ~w44355 & ~w44356;
assign w44358 = pi10066 & ~w16006;
assign w44359 = ~pi10627 & w16006;
assign w44360 = ~w44358 & ~w44359;
assign w44361 = pi10067 & ~w16006;
assign w44362 = ~pi10628 & w16006;
assign w44363 = ~w44361 & ~w44362;
assign w44364 = pi10068 & ~w16006;
assign w44365 = ~pi10629 & w16006;
assign w44366 = ~w44364 & ~w44365;
assign w44367 = pi10069 & ~w16006;
assign w44368 = ~pi10631 & w16006;
assign w44369 = ~w44367 & ~w44368;
assign w44370 = pi10070 & ~w16214;
assign w44371 = ~pi10632 & w16214;
assign w44372 = ~w44370 & ~w44371;
assign w44373 = pi10071 & ~w16214;
assign w44374 = ~pi10634 & w16214;
assign w44375 = ~w44373 & ~w44374;
assign w44376 = pi10072 & ~w16214;
assign w44377 = ~pi10623 & w16214;
assign w44378 = ~w44376 & ~w44377;
assign w44379 = pi10073 & ~w16214;
assign w44380 = ~pi10643 & w16214;
assign w44381 = ~w44379 & ~w44380;
assign w44382 = pi10074 & ~w16214;
assign w44383 = ~pi10647 & w16214;
assign w44384 = ~w44382 & ~w44383;
assign w44385 = pi10075 & ~w16214;
assign w44386 = ~pi10650 & w16214;
assign w44387 = ~w44385 & ~w44386;
assign w44388 = pi10076 & ~w16214;
assign w44389 = ~pi10652 & w16214;
assign w44390 = ~w44388 & ~w44389;
assign w44391 = pi10077 & ~w16214;
assign w44392 = ~pi10626 & w16214;
assign w44393 = ~w44391 & ~w44392;
assign w44394 = pi10078 & ~w16214;
assign w44395 = ~pi10627 & w16214;
assign w44396 = ~w44394 & ~w44395;
assign w44397 = pi10079 & ~w16214;
assign w44398 = ~pi10630 & w16214;
assign w44399 = ~w44397 & ~w44398;
assign w44400 = pi10080 & ~w16014;
assign w44401 = ~pi10622 & w16014;
assign w44402 = ~w44400 & ~w44401;
assign w44403 = pi10081 & ~w16014;
assign w44404 = ~pi10632 & w16014;
assign w44405 = ~w44403 & ~w44404;
assign w44406 = pi10082 & ~w16014;
assign w44407 = ~pi10635 & w16014;
assign w44408 = ~w44406 & ~w44407;
assign w44409 = pi10083 & ~w16014;
assign w44410 = ~pi10637 & w16014;
assign w44411 = ~w44409 & ~w44410;
assign w44412 = pi10084 & ~w16014;
assign w44413 = ~pi10638 & w16014;
assign w44414 = ~w44412 & ~w44413;
assign w44415 = pi10085 & ~w16014;
assign w44416 = ~pi10641 & w16014;
assign w44417 = ~w44415 & ~w44416;
assign w44418 = pi10086 & ~w16014;
assign w44419 = ~pi10645 & w16014;
assign w44420 = ~w44418 & ~w44419;
assign w44421 = pi10087 & ~w16014;
assign w44422 = ~pi10646 & w16014;
assign w44423 = ~w44421 & ~w44422;
assign w44424 = pi10088 & ~w16014;
assign w44425 = ~pi10648 & w16014;
assign w44426 = ~w44424 & ~w44425;
assign w44427 = pi10089 & ~w16014;
assign w44428 = ~pi10624 & w16014;
assign w44429 = ~w44427 & ~w44428;
assign w44430 = pi10090 & ~w16014;
assign w44431 = ~pi10653 & w16014;
assign w44432 = ~w44430 & ~w44431;
assign w44433 = pi10091 & ~w16014;
assign w44434 = ~pi10626 & w16014;
assign w44435 = ~w44433 & ~w44434;
assign w44436 = pi10092 & ~w16014;
assign w44437 = ~pi10629 & w16014;
assign w44438 = ~w44436 & ~w44437;
assign w44439 = pi10093 & ~w16014;
assign w44440 = ~pi10631 & w16014;
assign w44441 = ~w44439 & ~w44440;
assign w44442 = pi10094 & ~w16261;
assign w44443 = ~pi10634 & w16261;
assign w44444 = ~w44442 & ~w44443;
assign w44445 = pi10095 & ~w16261;
assign w44446 = ~pi10638 & w16261;
assign w44447 = ~w44445 & ~w44446;
assign w44448 = pi10096 & ~w16261;
assign w44449 = ~pi10640 & w16261;
assign w44450 = ~w44448 & ~w44449;
assign w44451 = pi10097 & ~w16261;
assign w44452 = ~pi10641 & w16261;
assign w44453 = ~w44451 & ~w44452;
assign w44454 = pi10098 & ~w16261;
assign w44455 = ~pi10623 & w16261;
assign w44456 = ~w44454 & ~w44455;
assign w44457 = pi10099 & ~w16261;
assign w44458 = ~pi10646 & w16261;
assign w44459 = ~w44457 & ~w44458;
assign w44460 = pi10100 & ~w16261;
assign w44461 = ~pi10647 & w16261;
assign w44462 = ~w44460 & ~w44461;
assign w44463 = pi10101 & ~w16261;
assign w44464 = ~pi10648 & w16261;
assign w44465 = ~w44463 & ~w44464;
assign w44466 = pi10102 & ~w16261;
assign w44467 = ~pi10652 & w16261;
assign w44468 = ~w44466 & ~w44467;
assign w44469 = pi10103 & ~w16261;
assign w44470 = ~pi10653 & w16261;
assign w44471 = ~w44469 & ~w44470;
assign w44472 = pi10104 & ~w16261;
assign w44473 = ~pi10627 & w16261;
assign w44474 = ~w44472 & ~w44473;
assign w44475 = pi10105 & ~w16261;
assign w44476 = ~pi10630 & w16261;
assign w44477 = ~w44475 & ~w44476;
assign w44478 = pi10106 & ~w16251;
assign w44479 = ~pi10639 & w16251;
assign w44480 = ~w44478 & ~w44479;
assign w44481 = pi10107 & ~w16251;
assign w44482 = ~pi10641 & w16251;
assign w44483 = ~w44481 & ~w44482;
assign w44484 = pi10108 & ~w16251;
assign w44485 = ~pi10642 & w16251;
assign w44486 = ~w44484 & ~w44485;
assign w44487 = pi10109 & ~w16251;
assign w44488 = ~pi10644 & w16251;
assign w44489 = ~w44487 & ~w44488;
assign w44490 = pi10110 & ~w16251;
assign w44491 = ~pi10630 & w16251;
assign w44492 = ~w44490 & ~w44491;
assign w44493 = pi10111 & ~w16244;
assign w44494 = ~pi10644 & w16244;
assign w44495 = ~w44493 & ~w44494;
assign w44496 = pi10112 & ~w16244;
assign w44497 = ~pi10646 & w16244;
assign w44498 = ~w44496 & ~w44497;
assign w44499 = pi10113 & ~w16244;
assign w44500 = ~pi10647 & w16244;
assign w44501 = ~w44499 & ~w44500;
assign w44502 = pi10114 & ~w16244;
assign w44503 = ~pi10648 & w16244;
assign w44504 = ~w44502 & ~w44503;
assign w44505 = pi10115 & ~w16244;
assign w44506 = ~pi10652 & w16244;
assign w44507 = ~w44505 & ~w44506;
assign w44508 = pi10116 & ~w16237;
assign w44509 = ~pi10632 & w16237;
assign w44510 = ~w44508 & ~w44509;
assign w44511 = pi10117 & ~w16237;
assign w44512 = ~pi10633 & w16237;
assign w44513 = ~w44511 & ~w44512;
assign w44514 = pi10118 & ~w16237;
assign w44515 = ~pi10634 & w16237;
assign w44516 = ~w44514 & ~w44515;
assign w44517 = pi10119 & ~w16237;
assign w44518 = ~pi10637 & w16237;
assign w44519 = ~w44517 & ~w44518;
assign w44520 = pi10120 & ~w16237;
assign w44521 = ~pi10638 & w16237;
assign w44522 = ~w44520 & ~w44521;
assign w44523 = pi10121 & ~w16237;
assign w44524 = ~pi10640 & w16237;
assign w44525 = ~w44523 & ~w44524;
assign w44526 = pi10122 & ~w16237;
assign w44527 = ~pi10623 & w16237;
assign w44528 = ~w44526 & ~w44527;
assign w44529 = pi10123 & ~w16237;
assign w44530 = ~pi10642 & w16237;
assign w44531 = ~w44529 & ~w44530;
assign w44532 = pi10124 & ~w16237;
assign w44533 = ~pi10643 & w16237;
assign w44534 = ~w44532 & ~w44533;
assign w44535 = pi10125 & ~w16237;
assign w44536 = ~pi10645 & w16237;
assign w44537 = ~w44535 & ~w44536;
assign w44538 = pi10126 & ~w16237;
assign w44539 = ~pi10649 & w16237;
assign w44540 = ~w44538 & ~w44539;
assign w44541 = pi10127 & ~w16237;
assign w44542 = ~pi10624 & w16237;
assign w44543 = ~w44541 & ~w44542;
assign w44544 = pi10128 & ~w16237;
assign w44545 = ~pi10652 & w16237;
assign w44546 = ~w44544 & ~w44545;
assign w44547 = pi10129 & ~w16237;
assign w44548 = ~pi10653 & w16237;
assign w44549 = ~w44547 & ~w44548;
assign w44550 = pi10130 & ~w16237;
assign w44551 = ~pi10631 & w16237;
assign w44552 = ~w44550 & ~w44551;
assign w44553 = pi10131 & ~w16233;
assign w44554 = ~pi10632 & w16233;
assign w44555 = ~w44553 & ~w44554;
assign w44556 = pi10132 & ~w16233;
assign w44557 = ~pi10634 & w16233;
assign w44558 = ~w44556 & ~w44557;
assign w44559 = pi10133 & ~w16233;
assign w44560 = ~pi10635 & w16233;
assign w44561 = ~w44559 & ~w44560;
assign w44562 = pi10134 & ~w16233;
assign w44563 = ~pi10636 & w16233;
assign w44564 = ~w44562 & ~w44563;
assign w44565 = pi10135 & ~w16233;
assign w44566 = ~pi10641 & w16233;
assign w44567 = ~w44565 & ~w44566;
assign w44568 = pi10136 & ~w16233;
assign w44569 = ~pi10642 & w16233;
assign w44570 = ~w44568 & ~w44569;
assign w44571 = pi10137 & ~w16233;
assign w44572 = ~pi10646 & w16233;
assign w44573 = ~w44571 & ~w44572;
assign w44574 = pi10138 & ~w16233;
assign w44575 = ~pi10648 & w16233;
assign w44576 = ~w44574 & ~w44575;
assign w44577 = pi10139 & ~w16233;
assign w44578 = ~pi10649 & w16233;
assign w44579 = ~w44577 & ~w44578;
assign w44580 = pi10140 & ~w16233;
assign w44581 = ~pi10651 & w16233;
assign w44582 = ~w44580 & ~w44581;
assign w44583 = pi10141 & ~w16233;
assign w44584 = ~pi10652 & w16233;
assign w44585 = ~w44583 & ~w44584;
assign w44586 = pi10142 & ~w16233;
assign w44587 = ~pi10653 & w16233;
assign w44588 = ~w44586 & ~w44587;
assign w44589 = pi10143 & ~w16233;
assign w44590 = ~pi10626 & w16233;
assign w44591 = ~w44589 & ~w44590;
assign w44592 = pi10144 & ~w16233;
assign w44593 = ~pi10627 & w16233;
assign w44594 = ~w44592 & ~w44593;
assign w44595 = pi10145 & ~w16233;
assign w44596 = ~pi10628 & w16233;
assign w44597 = ~w44595 & ~w44596;
assign w44598 = pi10146 & ~w16233;
assign w44599 = ~pi10630 & w16233;
assign w44600 = ~w44598 & ~w44599;
assign w44601 = pi10147 & ~w16032;
assign w44602 = ~pi10636 & w16032;
assign w44603 = ~w44601 & ~w44602;
assign w44604 = pi10148 & ~w16032;
assign w44605 = ~pi10637 & w16032;
assign w44606 = ~w44604 & ~w44605;
assign w44607 = pi10149 & ~w16032;
assign w44608 = ~pi10638 & w16032;
assign w44609 = ~w44607 & ~w44608;
assign w44610 = pi10150 & ~w16032;
assign w44611 = ~pi10623 & w16032;
assign w44612 = ~w44610 & ~w44611;
assign w44613 = pi10151 & ~w16032;
assign w44614 = ~pi10642 & w16032;
assign w44615 = ~w44613 & ~w44614;
assign w44616 = pi10152 & ~w16032;
assign w44617 = ~pi10643 & w16032;
assign w44618 = ~w44616 & ~w44617;
assign w44619 = pi10153 & ~w16225;
assign w44620 = ~pi10643 & w16225;
assign w44621 = ~w44619 & ~w44620;
assign w44622 = pi10154 & ~w16032;
assign w44623 = ~pi10645 & w16032;
assign w44624 = ~w44622 & ~w44623;
assign w44625 = pi10155 & ~w16032;
assign w44626 = ~pi10648 & w16032;
assign w44627 = ~w44625 & ~w44626;
assign w44628 = pi10156 & ~w16032;
assign w44629 = ~pi10650 & w16032;
assign w44630 = ~w44628 & ~w44629;
assign w44631 = pi10157 & ~w16032;
assign w44632 = ~pi10652 & w16032;
assign w44633 = ~w44631 & ~w44632;
assign w44634 = pi10158 & ~w16032;
assign w44635 = ~pi10628 & w16032;
assign w44636 = ~w44634 & ~w44635;
assign w44637 = pi10159 & ~w16032;
assign w44638 = ~pi10629 & w16032;
assign w44639 = ~w44637 & ~w44638;
assign w44640 = pi10160 & ~w16032;
assign w44641 = ~pi10631 & w16032;
assign w44642 = ~w44640 & ~w44641;
assign w44643 = pi10161 & ~w16229;
assign w44644 = ~pi10635 & w16229;
assign w44645 = ~w44643 & ~w44644;
assign w44646 = pi10162 & ~w16229;
assign w44647 = ~pi10637 & w16229;
assign w44648 = ~w44646 & ~w44647;
assign w44649 = pi10163 & ~w16229;
assign w44650 = ~pi10645 & w16229;
assign w44651 = ~w44649 & ~w44650;
assign w44652 = pi10164 & ~w16229;
assign w44653 = ~pi10646 & w16229;
assign w44654 = ~w44652 & ~w44653;
assign w44655 = pi10165 & ~w16229;
assign w44656 = ~pi10647 & w16229;
assign w44657 = ~w44655 & ~w44656;
assign w44658 = pi10166 & ~w16229;
assign w44659 = ~pi10650 & w16229;
assign w44660 = ~w44658 & ~w44659;
assign w44661 = pi10167 & ~w16229;
assign w44662 = ~pi10624 & w16229;
assign w44663 = ~w44661 & ~w44662;
assign w44664 = pi10168 & ~w16229;
assign w44665 = ~pi10626 & w16229;
assign w44666 = ~w44664 & ~w44665;
assign w44667 = pi10169 & ~w16229;
assign w44668 = ~pi10627 & w16229;
assign w44669 = ~w44667 & ~w44668;
assign w44670 = pi10170 & ~w16229;
assign w44671 = ~pi10629 & w16229;
assign w44672 = ~w44670 & ~w44671;
assign w44673 = pi10171 & ~w16054;
assign w44674 = ~pi10622 & w16054;
assign w44675 = ~w44673 & ~w44674;
assign w44676 = pi10172 & ~w16054;
assign w44677 = ~pi10634 & w16054;
assign w44678 = ~w44676 & ~w44677;
assign w44679 = pi10173 & ~w16054;
assign w44680 = ~pi10636 & w16054;
assign w44681 = ~w44679 & ~w44680;
assign w44682 = pi10174 & ~w16054;
assign w44683 = ~pi10637 & w16054;
assign w44684 = ~w44682 & ~w44683;
assign w44685 = pi10175 & ~w16054;
assign w44686 = ~pi10638 & w16054;
assign w44687 = ~w44685 & ~w44686;
assign w44688 = pi10176 & ~w16054;
assign w44689 = ~pi10642 & w16054;
assign w44690 = ~w44688 & ~w44689;
assign w44691 = pi10177 & ~w16054;
assign w44692 = ~pi10651 & w16054;
assign w44693 = ~w44691 & ~w44692;
assign w44694 = pi10178 & ~w16054;
assign w44695 = ~pi10624 & w16054;
assign w44696 = ~w44694 & ~w44695;
assign w44697 = pi10179 & ~w16054;
assign w44698 = ~pi10652 & w16054;
assign w44699 = ~w44697 & ~w44698;
assign w44700 = pi10180 & ~w16054;
assign w44701 = ~pi10626 & w16054;
assign w44702 = ~w44700 & ~w44701;
assign w44703 = pi10181 & ~w16054;
assign w44704 = ~pi10627 & w16054;
assign w44705 = ~w44703 & ~w44704;
assign w44706 = pi10182 & ~w16054;
assign w44707 = ~pi10628 & w16054;
assign w44708 = ~w44706 & ~w44707;
assign w44709 = pi10183 & ~w16054;
assign w44710 = ~pi10631 & w16054;
assign w44711 = ~w44709 & ~w44710;
assign w44712 = pi10184 & ~w14866;
assign w44713 = ~pi10632 & w14866;
assign w44714 = ~w44712 & ~w44713;
assign w44715 = pi10185 & ~w14866;
assign w44716 = ~pi10637 & w14866;
assign w44717 = ~w44715 & ~w44716;
assign w44718 = pi10186 & ~w14866;
assign w44719 = ~pi10641 & w14866;
assign w44720 = ~w44718 & ~w44719;
assign w44721 = pi10187 & ~w14866;
assign w44722 = ~pi10644 & w14866;
assign w44723 = ~w44721 & ~w44722;
assign w44724 = pi10188 & ~w14866;
assign w44725 = ~pi10646 & w14866;
assign w44726 = ~w44724 & ~w44725;
assign w44727 = pi10189 & ~w14866;
assign w44728 = ~pi10648 & w14866;
assign w44729 = ~w44727 & ~w44728;
assign w44730 = pi10190 & ~w14866;
assign w44731 = ~pi10651 & w14866;
assign w44732 = ~w44730 & ~w44731;
assign w44733 = pi10191 & ~w14866;
assign w44734 = ~pi10624 & w14866;
assign w44735 = ~w44733 & ~w44734;
assign w44736 = pi10192 & ~w14866;
assign w44737 = ~pi10653 & w14866;
assign w44738 = ~w44736 & ~w44737;
assign w44739 = pi10193 & ~w14866;
assign w44740 = ~pi10631 & w14866;
assign w44741 = ~w44739 & ~w44740;
assign w44742 = pi10194 & ~w16225;
assign w44743 = ~pi10636 & w16225;
assign w44744 = ~w44742 & ~w44743;
assign w44745 = pi10195 & ~w16225;
assign w44746 = ~pi10638 & w16225;
assign w44747 = ~w44745 & ~w44746;
assign w44748 = pi10196 & ~w16225;
assign w44749 = ~pi10642 & w16225;
assign w44750 = ~w44748 & ~w44749;
assign w44751 = pi10197 & ~w16225;
assign w44752 = ~pi10644 & w16225;
assign w44753 = ~w44751 & ~w44752;
assign w44754 = pi10198 & ~w16225;
assign w44755 = ~pi10645 & w16225;
assign w44756 = ~w44754 & ~w44755;
assign w44757 = pi10199 & ~w16225;
assign w44758 = ~pi10646 & w16225;
assign w44759 = ~w44757 & ~w44758;
assign w44760 = pi10200 & ~w16225;
assign w44761 = ~pi10649 & w16225;
assign w44762 = ~w44760 & ~w44761;
assign w44763 = pi10201 & ~w16225;
assign w44764 = ~pi10650 & w16225;
assign w44765 = ~w44763 & ~w44764;
assign w44766 = pi10202 & ~w16225;
assign w44767 = ~pi10651 & w16225;
assign w44768 = ~w44766 & ~w44767;
assign w44769 = pi10203 & ~w16225;
assign w44770 = ~pi10631 & w16225;
assign w44771 = ~w44769 & ~w44770;
assign w44772 = pi10204 & ~w16219;
assign w44773 = ~pi10622 & w16219;
assign w44774 = ~w44772 & ~w44773;
assign w44775 = pi10205 & ~w16219;
assign w44776 = ~pi10635 & w16219;
assign w44777 = ~w44775 & ~w44776;
assign w44778 = pi10206 & ~w16219;
assign w44779 = ~pi10640 & w16219;
assign w44780 = ~w44778 & ~w44779;
assign w44781 = pi10207 & ~w16219;
assign w44782 = ~pi10642 & w16219;
assign w44783 = ~w44781 & ~w44782;
assign w44784 = pi10208 & ~w16219;
assign w44785 = ~pi10643 & w16219;
assign w44786 = ~w44784 & ~w44785;
assign w44787 = pi10209 & ~w16219;
assign w44788 = ~pi10645 & w16219;
assign w44789 = ~w44787 & ~w44788;
assign w44790 = pi10210 & ~w16219;
assign w44791 = ~pi10650 & w16219;
assign w44792 = ~w44790 & ~w44791;
assign w44793 = pi10211 & ~w16219;
assign w44794 = ~pi10651 & w16219;
assign w44795 = ~w44793 & ~w44794;
assign w44796 = pi10212 & ~w16219;
assign w44797 = ~pi10624 & w16219;
assign w44798 = ~w44796 & ~w44797;
assign w44799 = pi10213 & ~w16219;
assign w44800 = ~pi10653 & w16219;
assign w44801 = ~w44799 & ~w44800;
assign w44802 = pi10214 & ~w16219;
assign w44803 = ~pi10625 & w16219;
assign w44804 = ~w44802 & ~w44803;
assign w44805 = pi10215 & ~w16219;
assign w44806 = ~pi10627 & w16219;
assign w44807 = ~w44805 & ~w44806;
assign w44808 = pi10216 & ~w16219;
assign w44809 = ~pi10630 & w16219;
assign w44810 = ~w44808 & ~w44809;
assign w44811 = pi10217 & ~w16271;
assign w44812 = ~pi10632 & w16271;
assign w44813 = ~w44811 & ~w44812;
assign w44814 = pi10218 & ~w16271;
assign w44815 = ~pi10637 & w16271;
assign w44816 = ~w44814 & ~w44815;
assign w44817 = pi10219 & ~w16271;
assign w44818 = ~pi10639 & w16271;
assign w44819 = ~w44817 & ~w44818;
assign w44820 = pi10220 & ~w16271;
assign w44821 = ~pi10641 & w16271;
assign w44822 = ~w44820 & ~w44821;
assign w44823 = pi10221 & ~w16271;
assign w44824 = ~pi10623 & w16271;
assign w44825 = ~w44823 & ~w44824;
assign w44826 = pi10222 & ~w16271;
assign w44827 = ~pi10643 & w16271;
assign w44828 = ~w44826 & ~w44827;
assign w44829 = pi10223 & ~w16271;
assign w44830 = ~pi10645 & w16271;
assign w44831 = ~w44829 & ~w44830;
assign w44832 = pi10224 & ~w16271;
assign w44833 = ~pi10646 & w16271;
assign w44834 = ~w44832 & ~w44833;
assign w44835 = pi10225 & ~w16271;
assign w44836 = ~pi10649 & w16271;
assign w44837 = ~w44835 & ~w44836;
assign w44838 = pi10226 & ~w16271;
assign w44839 = ~pi10651 & w16271;
assign w44840 = ~w44838 & ~w44839;
assign w44841 = pi10227 & ~w16271;
assign w44842 = ~pi10624 & w16271;
assign w44843 = ~w44841 & ~w44842;
assign w44844 = pi10228 & ~w16271;
assign w44845 = ~pi10653 & w16271;
assign w44846 = ~w44844 & ~w44845;
assign w44847 = pi10229 & ~w16271;
assign w44848 = ~pi10626 & w16271;
assign w44849 = ~w44847 & ~w44848;
assign w44850 = pi10230 & ~w16271;
assign w44851 = ~pi10629 & w16271;
assign w44852 = ~w44850 & ~w44851;
assign w44853 = ~pi10231 & ~w11341;
assign w44854 = ~w11342 & ~w44853;
assign w44855 = pi10232 & ~w19704;
assign w44856 = pi10664 & w44141;
assign w44857 = ~w44855 & ~w44856;
assign w44858 = pi10233 & ~w44191;
assign w44859 = pi10611 & w44191;
assign w44860 = ~w44858 & ~w44859;
assign w44861 = pi10234 & ~w44227;
assign w44862 = pi10608 & w44227;
assign w44863 = ~w44861 & ~w44862;
assign w44864 = pi10235 & ~w44227;
assign w44865 = pi10609 & w44227;
assign w44866 = ~w44864 & ~w44865;
assign w44867 = pi10236 & ~w44227;
assign w44868 = pi10611 & w44227;
assign w44869 = ~w44867 & ~w44868;
assign w44870 = pi10237 & ~w44227;
assign w44871 = pi10610 & w44227;
assign w44872 = ~w44870 & ~w44871;
assign w44873 = pi10238 & ~w44217;
assign w44874 = pi10616 & w44217;
assign w44875 = ~w44873 & ~w44874;
assign w44876 = pi10239 & ~w44217;
assign w44877 = pi10615 & w44217;
assign w44878 = ~w44876 & ~w44877;
assign w44879 = pi10240 & ~w44217;
assign w44880 = pi10619 & w44217;
assign w44881 = ~w44879 & ~w44880;
assign w44882 = pi10241 & ~w44217;
assign w44883 = pi10618 & w44217;
assign w44884 = ~w44882 & ~w44883;
assign w44885 = pi10242 & ~w44217;
assign w44886 = pi10620 & w44217;
assign w44887 = ~w44885 & ~w44886;
assign w44888 = pi10243 & ~w44210;
assign w44889 = pi10606 & w44210;
assign w44890 = ~w44888 & ~w44889;
assign w44891 = pi10244 & ~w44210;
assign w44892 = pi10607 & w44210;
assign w44893 = ~w44891 & ~w44892;
assign w44894 = pi10245 & ~w44210;
assign w44895 = pi10608 & w44210;
assign w44896 = ~w44894 & ~w44895;
assign w44897 = pi10246 & ~w44210;
assign w44898 = pi10610 & w44210;
assign w44899 = ~w44897 & ~w44898;
assign w44900 = pi10247 & ~w44210;
assign w44901 = pi10611 & w44210;
assign w44902 = ~w44900 & ~w44901;
assign w44903 = pi10248 & ~w44210;
assign w44904 = pi10613 & w44210;
assign w44905 = ~w44903 & ~w44904;
assign w44906 = pi10249 & ~w44195;
assign w44907 = pi10614 & w44195;
assign w44908 = ~w44906 & ~w44907;
assign w44909 = pi10250 & ~w44195;
assign w44910 = pi10615 & w44195;
assign w44911 = ~w44909 & ~w44910;
assign w44912 = pi10251 & ~w44195;
assign w44913 = pi10617 & w44195;
assign w44914 = ~w44912 & ~w44913;
assign w44915 = pi10252 & ~w44195;
assign w44916 = pi10618 & w44195;
assign w44917 = ~w44915 & ~w44916;
assign w44918 = pi10253 & ~w44195;
assign w44919 = pi10621 & w44195;
assign w44920 = ~w44918 & ~w44919;
assign w44921 = pi10254 & ~w44191;
assign w44922 = pi10606 & w44191;
assign w44923 = ~w44921 & ~w44922;
assign w44924 = pi10255 & ~w44191;
assign w44925 = pi10608 & w44191;
assign w44926 = ~w44924 & ~w44925;
assign w44927 = pi10256 & ~w44191;
assign w44928 = pi10609 & w44191;
assign w44929 = ~w44927 & ~w44928;
assign w44930 = pi10257 & ~w44191;
assign w44931 = pi10610 & w44191;
assign w44932 = ~w44930 & ~w44931;
assign w44933 = pi10258 & ~w44191;
assign w44934 = pi10613 & w44191;
assign w44935 = ~w44933 & ~w44934;
assign w44936 = pi10259 & ~w44175;
assign w44937 = pi10615 & w44175;
assign w44938 = ~w44936 & ~w44937;
assign w44939 = pi10260 & ~w44175;
assign w44940 = pi10617 & w44175;
assign w44941 = ~w44939 & ~w44940;
assign w44942 = pi10261 & ~w44175;
assign w44943 = pi10620 & w44175;
assign w44944 = ~w44942 & ~w44943;
assign w44945 = pi10262 & ~w16054;
assign w44946 = ~pi10653 & w16054;
assign w44947 = ~w44945 & ~w44946;
assign w44948 = ~pi00832 & ~pi09841;
assign w44949 = pi00833 & ~pi09842;
assign w44950 = ~pi00831 & ~pi09840;
assign w44951 = ~pi00833 & pi09842;
assign w44952 = pi00832 & pi09841;
assign w44953 = pi00835 & pi09844;
assign w44954 = ~pi00834 & ~pi09843;
assign w44955 = pi00831 & pi09840;
assign w44956 = ~pi00827 & ~pi09845;
assign w44957 = pi00834 & pi09843;
assign w44958 = ~pi00835 & ~pi09844;
assign w44959 = pi00827 & pi09845;
assign w44960 = ~w288 & ~w44948;
assign w44961 = ~w44949 & ~w44950;
assign w44962 = ~w44951 & ~w44952;
assign w44963 = ~w44953 & ~w44954;
assign w44964 = ~w44955 & ~w44956;
assign w44965 = ~w44957 & ~w44958;
assign w44966 = ~w44959 & w44965;
assign w44967 = w44963 & w44964;
assign w44968 = w44961 & w44962;
assign w44969 = w44960 & w44968;
assign w44970 = w44966 & w44967;
assign w44971 = ~w11884 & w44970;
assign w44972 = w44969 & w44971;
assign w44973 = pi00007 & pi00032;
assign w44974 = ~pi10263 & w44973;
assign w44975 = ~w44972 & ~w44974;
assign w44976 = pi10436 & w13021;
assign w44977 = pi10264 & ~w11160;
assign w44978 = ~w44976 & ~w44977;
assign w44979 = pi10470 & pi10493;
assign w44980 = pi10265 & ~w44979;
assign w44981 = ~w575 & ~w44980;
assign w44982 = pi10267 & ~w14866;
assign w44983 = ~pi10643 & w14866;
assign w44984 = ~w44982 & ~w44983;
assign w44985 = pi10268 & ~w14866;
assign w44986 = ~pi10639 & w14866;
assign w44987 = ~w44985 & ~w44986;
assign w44988 = pi10269 & ~w14866;
assign w44989 = ~pi10635 & w14866;
assign w44990 = ~w44988 & ~w44989;
assign w44991 = pi10270 & ~w16054;
assign w44992 = ~pi10629 & w16054;
assign w44993 = ~w44991 & ~w44992;
assign w44994 = pi10271 & ~w14866;
assign w44995 = ~pi10622 & w14866;
assign w44996 = ~w44994 & ~w44995;
assign w44997 = pi10272 & ~w16006;
assign w44998 = ~pi10635 & w16006;
assign w44999 = ~w44997 & ~w44998;
assign w45000 = pi10273 & ~w16054;
assign w45001 = ~pi10639 & w16054;
assign w45002 = ~w45000 & ~w45001;
assign w45003 = pi10274 & ~w16054;
assign w45004 = ~pi10644 & w16054;
assign w45005 = ~w45003 & ~w45004;
assign w45006 = pi10275 & ~w16054;
assign w45007 = ~pi10649 & w16054;
assign w45008 = ~w45006 & ~w45007;
assign w45009 = pi10276 & ~w16054;
assign w45010 = ~pi10643 & w16054;
assign w45011 = ~w45009 & ~w45010;
assign w45012 = pi10277 & ~w16229;
assign w45013 = ~pi10631 & w16229;
assign w45014 = ~w45012 & ~w45013;
assign w45015 = pi10278 & ~w16054;
assign w45016 = ~pi10635 & w16054;
assign w45017 = ~w45015 & ~w45016;
assign w45018 = pi10279 & ~w16054;
assign w45019 = ~pi10632 & w16054;
assign w45020 = ~w45018 & ~w45019;
assign w45021 = pi10280 & ~w16229;
assign w45022 = ~pi10653 & w16229;
assign w45023 = ~w45021 & ~w45022;
assign w45024 = pi10281 & ~w16229;
assign w45025 = ~pi10651 & w16229;
assign w45026 = ~w45024 & ~w45025;
assign w45027 = pi10282 & ~w16229;
assign w45028 = ~pi10648 & w16229;
assign w45029 = ~w45027 & ~w45028;
assign w45030 = pi10283 & ~w16229;
assign w45031 = ~pi10633 & w16229;
assign w45032 = ~w45030 & ~w45031;
assign w45033 = pi10284 & ~w16229;
assign w45034 = ~pi10643 & w16229;
assign w45035 = ~w45033 & ~w45034;
assign w45036 = pi10285 & ~w16229;
assign w45037 = ~pi10636 & w16229;
assign w45038 = ~w45036 & ~w45037;
assign w45039 = pi10286 & ~w16237;
assign w45040 = ~pi10628 & w16237;
assign w45041 = ~w45039 & ~w45040;
assign w45042 = pi10287 & ~w16032;
assign w45043 = ~pi10625 & w16032;
assign w45044 = ~w45042 & ~w45043;
assign w45045 = pi10288 & ~w16233;
assign w45046 = ~pi10631 & w16233;
assign w45047 = ~w45045 & ~w45046;
assign w45048 = pi10289 & ~w16032;
assign w45049 = ~pi10649 & w16032;
assign w45050 = ~w45048 & ~w45049;
assign w45051 = pi10290 & ~w16032;
assign w45052 = ~pi10624 & w16032;
assign w45053 = ~w45051 & ~w45052;
assign w45054 = pi10291 & ~w16032;
assign w45055 = ~pi10644 & w16032;
assign w45056 = ~w45054 & ~w45055;
assign w45057 = pi10292 & ~w16032;
assign w45058 = ~pi10646 & w16032;
assign w45059 = ~w45057 & ~w45058;
assign w45060 = pi10293 & ~w16032;
assign w45061 = ~pi10622 & w16032;
assign w45062 = ~w45060 & ~w45061;
assign w45063 = pi10294 & ~w16032;
assign w45064 = ~pi10634 & w16032;
assign w45065 = ~w45063 & ~w45064;
assign w45066 = pi10295 & ~w16032;
assign w45067 = ~pi10639 & w16032;
assign w45068 = ~w45066 & ~w45067;
assign w45069 = pi10296 & ~w16233;
assign w45070 = ~pi10629 & w16233;
assign w45071 = ~w45069 & ~w45070;
assign w45072 = pi10297 & ~w16233;
assign w45073 = ~pi10625 & w16233;
assign w45074 = ~w45072 & ~w45073;
assign w45075 = pi10298 & ~w16233;
assign w45076 = ~pi10622 & w16233;
assign w45077 = ~w45075 & ~w45076;
assign w45078 = pi10299 & ~w16233;
assign w45079 = ~pi10650 & w16233;
assign w45080 = ~w45078 & ~w45079;
assign w45081 = pi10300 & ~w16233;
assign w45082 = ~pi10623 & w16233;
assign w45083 = ~w45081 & ~w45082;
assign w45084 = pi10301 & ~w16233;
assign w45085 = ~pi10643 & w16233;
assign w45086 = ~w45084 & ~w45085;
assign w45087 = pi10302 & ~w16233;
assign w45088 = ~pi10633 & w16233;
assign w45089 = ~w45087 & ~w45088;
assign w45090 = pi10303 & ~w16233;
assign w45091 = ~pi10640 & w16233;
assign w45092 = ~w45090 & ~w45091;
assign w45093 = pi10304 & ~w16244;
assign w45094 = ~pi10625 & w16244;
assign w45095 = ~w45093 & ~w45094;
assign w45096 = pi10305 & ~w16237;
assign w45097 = ~pi10644 & w16237;
assign w45098 = ~w45096 & ~w45097;
assign w45099 = pi10306 & ~w16237;
assign w45100 = ~pi10651 & w16237;
assign w45101 = ~w45099 & ~w45100;
assign w45102 = pi10307 & ~w16237;
assign w45103 = ~pi10646 & w16237;
assign w45104 = ~w45102 & ~w45103;
assign w45105 = pi10308 & ~w16237;
assign w45106 = ~pi10641 & w16237;
assign w45107 = ~w45105 & ~w45106;
assign w45108 = pi10309 & ~w16237;
assign w45109 = ~pi10636 & w16237;
assign w45110 = ~w45108 & ~w45109;
assign w45111 = pi10310 & ~w16244;
assign w45112 = ~pi10630 & w16244;
assign w45113 = ~w45111 & ~w45112;
assign w45114 = pi10311 & ~w16244;
assign w45115 = ~pi10629 & w16244;
assign w45116 = ~w45114 & ~w45115;
assign w45117 = pi10312 & ~w16244;
assign w45118 = ~pi10650 & w16244;
assign w45119 = ~w45117 & ~w45118;
assign w45120 = pi10313 & ~w16251;
assign w45121 = ~pi10622 & w16251;
assign w45122 = ~w45120 & ~w45121;
assign w45123 = pi10314 & ~w16251;
assign w45124 = ~pi10646 & w16251;
assign w45125 = ~w45123 & ~w45124;
assign w45126 = pi10315 & ~w16251;
assign w45127 = ~pi10631 & w16251;
assign w45128 = ~w45126 & ~w45127;
assign w45129 = pi10316 & ~w16244;
assign w45130 = ~pi10645 & w16244;
assign w45131 = ~w45129 & ~w45130;
assign w45132 = pi10317 & ~w16251;
assign w45133 = ~pi10640 & w16251;
assign w45134 = ~w45132 & ~w45133;
assign w45135 = pi10318 & ~w16261;
assign w45136 = ~pi10629 & w16261;
assign w45137 = ~w45135 & ~w45136;
assign w45138 = pi10319 & ~w16261;
assign w45139 = ~pi10650 & w16261;
assign w45140 = ~w45138 & ~w45139;
assign w45141 = pi10320 & ~w16261;
assign w45142 = ~pi10644 & w16261;
assign w45143 = ~w45141 & ~w45142;
assign w45144 = pi10321 & ~w16261;
assign w45145 = ~pi10635 & w16261;
assign w45146 = ~w45144 & ~w45145;
assign w45147 = pi10322 & ~w16261;
assign w45148 = ~pi10639 & w16261;
assign w45149 = ~w45147 & ~w45148;
assign w45150 = pi10323 & ~w16261;
assign w45151 = ~pi10632 & w16261;
assign w45152 = ~w45150 & ~w45151;
assign w45153 = pi10324 & ~w16014;
assign w45154 = ~pi10627 & w16014;
assign w45155 = ~w45153 & ~w45154;
assign w45156 = pi10325 & ~w16014;
assign w45157 = ~pi10630 & w16014;
assign w45158 = ~w45156 & ~w45157;
assign w45159 = pi10326 & ~w16014;
assign w45160 = ~pi10633 & w16014;
assign w45161 = ~w45159 & ~w45160;
assign w45162 = pi10327 & ~w16006;
assign w45163 = ~pi10652 & w16006;
assign w45164 = ~w45162 & ~w45163;
assign w45165 = pi10328 & ~w16014;
assign w45166 = ~pi10651 & w16014;
assign w45167 = ~w45165 & ~w45166;
assign w45168 = pi10329 & ~w16014;
assign w45169 = ~pi10623 & w16014;
assign w45170 = ~w45168 & ~w45169;
assign w45171 = pi10330 & ~w16014;
assign w45172 = ~pi10643 & w16014;
assign w45173 = ~w45171 & ~w45172;
assign w45174 = pi10331 & ~w16014;
assign w45175 = ~pi10642 & w16014;
assign w45176 = ~w45174 & ~w45175;
assign w45177 = pi10332 & ~w16014;
assign w45178 = ~pi10639 & w16014;
assign w45179 = ~w45177 & ~w45178;
assign w45180 = pi10333 & ~w16214;
assign w45181 = ~pi10628 & w16214;
assign w45182 = ~w45180 & ~w45181;
assign w45183 = pi10334 & ~w16214;
assign w45184 = ~pi10648 & w16214;
assign w45185 = ~w45183 & ~w45184;
assign w45186 = pi10335 & ~w16214;
assign w45187 = ~pi10651 & w16214;
assign w45188 = ~w45186 & ~w45187;
assign w45189 = pi10336 & ~w16214;
assign w45190 = ~pi10646 & w16214;
assign w45191 = ~w45189 & ~w45190;
assign w45192 = pi10337 & ~w16214;
assign w45193 = ~pi10633 & w16214;
assign w45194 = ~w45192 & ~w45193;
assign w45195 = pi10338 & ~w16214;
assign w45196 = ~pi10622 & w16214;
assign w45197 = ~w45195 & ~w45196;
assign w45198 = pi10339 & ~w16006;
assign w45199 = ~pi10630 & w16006;
assign w45200 = ~w45198 & ~w45199;
assign w45201 = pi10340 & ~w16006;
assign w45202 = ~pi10626 & w16006;
assign w45203 = ~w45201 & ~w45202;
assign w45204 = pi10341 & ~w16006;
assign w45205 = ~pi10637 & w16006;
assign w45206 = ~w45204 & ~w45205;
assign w45207 = pi10342 & ~w16006;
assign w45208 = ~pi10645 & w16006;
assign w45209 = ~w45207 & ~w45208;
assign w45210 = pi10343 & ~w16006;
assign w45211 = ~pi10650 & w16006;
assign w45212 = ~w45210 & ~w45211;
assign w45213 = pi10344 & ~w16006;
assign w45214 = ~pi10647 & w16006;
assign w45215 = ~w45213 & ~w45214;
assign w45216 = pi10527 & ~w12874;
assign w45217 = pi10441 & ~pi10494;
assign w45218 = ~pi10345 & ~w1194;
assign w45219 = ~pi09519 & ~w45217;
assign w45220 = ~w45216 & w45219;
assign w45221 = ~w45218 & w45220;
assign w45222 = pi10346 & ~w16006;
assign w45223 = ~pi10623 & w16006;
assign w45224 = ~w45222 & ~w45223;
assign w45225 = ~pi10347 & ~w1583;
assign w45226 = ~pi10577 & ~w1584;
assign w45227 = ~w45225 & w45226;
assign w45228 = ~pi10398 & ~pi10461;
assign w45229 = ~pi10400 & ~pi10455;
assign w45230 = ~pi10407 & ~pi10456;
assign w45231 = ~pi10352 & ~w1371;
assign w45232 = w830 & ~w45231;
assign w45233 = ~w11127 & w45232;
assign w45234 = ~pi10353 & ~w1581;
assign w45235 = ~pi10577 & ~w1582;
assign w45236 = ~w45234 & w45235;
assign w45237 = ~pi02657 & pi02658;
assign w45238 = ~pi02660 & pi10453;
assign w45239 = ~pi10355 & ~w45238;
assign w45240 = ~w45237 & ~w45239;
assign w45241 = w11341 & ~w14191;
assign w45242 = ~pi10356 & ~w45241;
assign w45243 = ~pi10425 & pi10460;
assign w45244 = ~pi10357 & ~w45243;
assign w45245 = ~pi10439 & ~w45244;
assign w45246 = ~pi00140 & w16775;
assign w45247 = ~pi00045 & ~pi00046;
assign w45248 = ~pi10050 & ~pi10476;
assign w45249 = w45247 & w45248;
assign w45250 = w45246 & ~w45249;
assign w45251 = ~pi10397 & ~pi10448;
assign w45252 = ~pi00062 & w2041;
assign w45253 = ~pi10361 & ~w1582;
assign w45254 = ~pi10577 & ~w1583;
assign w45255 = ~w45253 & w45254;
assign w45256 = pi10363 & ~w11160;
assign w45257 = pi00035 & w13022;
assign w45258 = ~pi10500 & w11160;
assign w45259 = ~w45257 & w45258;
assign w45260 = ~w45256 & ~w45259;
assign w45261 = pi00484 & w12879;
assign w45262 = ~pi10364 & ~w12877;
assign w45263 = ~w12879 & ~w12881;
assign w45264 = ~w45262 & w45263;
assign w45265 = ~w45261 & ~w45264;
assign w45266 = pi00869 & ~w1435;
assign w45267 = ~pi00869 & ~pi10369;
assign w45268 = ~w45266 & ~w45267;
assign w45269 = ~pi00044 & w14204;
assign w45270 = pi00025 & w43936;
assign w45271 = ~w45269 & ~w45270;
assign w45272 = w739 & w45271;
assign w45273 = w45246 & w45249;
assign w45274 = ~pi00029 & w14204;
assign w45275 = w770 & ~w45274;
assign w45276 = pi00477 & w12879;
assign w45277 = pi10374 & w45263;
assign w45278 = ~pi10374 & w12876;
assign w45279 = w12881 & w45278;
assign w45280 = ~w45276 & ~w45279;
assign w45281 = ~w45277 & w45280;
assign w45282 = pi01252 & ~pi10377;
assign w45283 = ~w1576 & w45282;
assign w45284 = ~pi00053 & pi10423;
assign w45285 = pi10519 & w45284;
assign w45286 = ~pi10378 & ~w45285;
assign w45287 = ~pi00845 & ~w45286;
assign w45288 = ~pi00539 & pi10423;
assign w45289 = pi10490 & w45288;
assign w45290 = ~pi10379 & ~w45289;
assign w45291 = ~pi00845 & ~w45290;
assign w45292 = pi10433 & ~w12854;
assign w45293 = ~pi00845 & w16299;
assign w45294 = pi01165 & ~w11126;
assign w45295 = ~w45293 & w45294;
assign w45296 = ~pi10381 & ~w45295;
assign w45297 = pi10418 & pi10488;
assign w45298 = ~w45296 & ~w45297;
assign w45299 = pi10382 & ~w12877;
assign w45300 = ~pi10451 & ~w45299;
assign w45301 = pi10384 & ~w11160;
assign w45302 = pi00035 & w16188;
assign w45303 = pi00476 & w11160;
assign w45304 = ~w45302 & w45303;
assign w45305 = ~w45301 & ~w45304;
assign w45306 = ~pi10385 & ~w1580;
assign w45307 = ~pi10577 & ~w1581;
assign w45308 = ~w45306 & w45307;
assign w45309 = ~pi10386 & ~w1579;
assign w45310 = ~pi10577 & ~w1580;
assign w45311 = ~w45309 & w45310;
assign w45312 = ~pi10387 & ~pi10514;
assign w45313 = ~w537 & ~w45312;
assign w45314 = ~pi10478 & pi10479;
assign w45315 = ~w42559 & ~w45314;
assign w45316 = ~pi10467 & ~pi10515;
assign w45317 = ~pi10362 & ~pi10389;
assign w45318 = ~w45316 & ~w45317;
assign w45319 = ~pi10390 & ~pi10446;
assign w45320 = ~pi10457 & ~w45319;
assign w45321 = ~pi10391 & ~w1578;
assign w45322 = ~pi10577 & ~w1579;
assign w45323 = ~w45321 & w45322;
assign w45324 = pi10393 & ~w1194;
assign w45325 = pi09953 & ~pi10540;
assign w45326 = ~pi10345 & w12874;
assign w45327 = w45325 & w45326;
assign w45328 = ~w45324 & ~w45327;
assign w45329 = pi00865 & ~pi10528;
assign w45330 = ~pi10394 & pi10528;
assign w45331 = ~w45329 & ~w45330;
assign w45332 = pi00863 & ~pi10528;
assign w45333 = ~pi10395 & pi10528;
assign w45334 = ~w45332 & ~w45333;
assign w45335 = pi00864 & ~pi10528;
assign w45336 = ~pi10396 & pi10528;
assign w45337 = ~w45335 & ~w45336;
assign w45338 = pi00862 & ~pi10528;
assign w45339 = ~pi10401 & pi10528;
assign w45340 = ~w45338 & ~w45339;
assign w45341 = pi00968 & ~pi10528;
assign w45342 = ~pi10402 & pi10528;
assign w45343 = ~w45341 & ~w45342;
assign w45344 = pi00969 & ~pi10528;
assign w45345 = ~pi10403 & pi10528;
assign w45346 = ~w45344 & ~w45345;
assign w45347 = pi02726 & ~pi10528;
assign w45348 = ~pi10404 & pi10528;
assign w45349 = ~w45347 & ~w45348;
assign w45350 = pi00860 & ~pi10528;
assign w45351 = ~pi10405 & pi10528;
assign w45352 = ~w45350 & ~w45351;
assign w45353 = ~pi10373 & ~pi10406;
assign w45354 = ~pi10266 & pi10542;
assign w45355 = ~w45353 & ~w45354;
assign w45356 = pi10408 & ~w1371;
assign w45357 = pi00062 & w45325;
assign w45358 = w16783 & w45357;
assign w45359 = ~w45356 & ~w45358;
assign w45360 = pi00869 & ~w1432;
assign w45361 = ~pi00869 & ~pi10409;
assign w45362 = ~w45360 & ~w45361;
assign w45363 = pi00859 & ~pi10528;
assign w45364 = ~pi10410 & pi10528;
assign w45365 = ~w45363 & ~w45364;
assign w45366 = pi00861 & ~pi10528;
assign w45367 = ~pi10411 & pi10528;
assign w45368 = ~w45366 & ~w45367;
assign w45369 = pi00848 & ~pi10528;
assign w45370 = ~pi10412 & pi10528;
assign w45371 = ~w45369 & ~w45370;
assign w45372 = pi02725 & ~pi10528;
assign w45373 = ~pi10413 & pi10528;
assign w45374 = ~w45372 & ~w45373;
assign w45375 = pi02157 & ~pi10528;
assign w45376 = ~pi10414 & pi10528;
assign w45377 = ~w45375 & ~w45376;
assign w45378 = pi02730 & ~pi10528;
assign w45379 = ~pi10415 & pi10528;
assign w45380 = ~w45378 & ~w45379;
assign w45381 = pi02728 & ~pi10528;
assign w45382 = ~pi10416 & pi10528;
assign w45383 = ~w45381 & ~w45382;
assign w45384 = pi02727 & ~pi10528;
assign w45385 = ~pi10417 & pi10528;
assign w45386 = ~w45384 & ~w45385;
assign w45387 = pi00053 & pi10418;
assign w45388 = ~w45294 & ~w45387;
assign w45389 = ~pi00869 & ~pi10419;
assign w45390 = ~pi00240 & pi00869;
assign w45391 = ~w45389 & ~w45390;
assign w45392 = pi01251 & ~pi01252;
assign w45393 = pi00357 & ~w45392;
assign w45394 = ~pi00133 & w12877;
assign w45395 = ~w45393 & w45394;
assign w45396 = ~pi10477 & ~pi10482;
assign w45397 = ~pi10521 & ~pi10522;
assign w45398 = ~pi10536 & ~pi10537;
assign w45399 = w45397 & w45398;
assign w45400 = w45396 & w45399;
assign w45401 = w45395 & ~w45400;
assign w45402 = ~pi00869 & ~pi10422;
assign w45403 = ~pi00233 & pi00869;
assign w45404 = ~w45402 & ~w45403;
assign w45405 = ~pi10423 & ~w11126;
assign w45406 = w12844 & ~w45405;
assign w45407 = pi00435 & ~pi10430;
assign w45408 = w10682 & ~w45407;
assign w45409 = ~pi00000 & w45400;
assign w45410 = w45395 & w45409;
assign w45411 = pi10432 & ~pi10539;
assign w45412 = ~pi00062 & pi09997;
assign w45413 = ~w45411 & ~w45412;
assign w45414 = ~pi00963 & ~pi09967;
assign w45415 = ~pi10434 & w45414;
assign w45416 = pi00007 & pi00038;
assign w45417 = ~w45415 & w45416;
assign w45418 = ~pi00841 & pi10435;
assign w45419 = ~pi10446 & w45418;
assign w45420 = pi01272 & ~w45419;
assign w45421 = ~pi00815 & ~pi09875;
assign w45422 = ~pi09967 & pi10587;
assign w45423 = ~w45421 & w45422;
assign w45424 = ~pi10437 & ~w45423;
assign w45425 = ~pi00869 & ~w45424;
assign w45426 = pi09823 & w45325;
assign w45427 = ~w16891 & ~w16904;
assign w45428 = ~w16927 & ~w16991;
assign w45429 = ~w45426 & w45428;
assign w45430 = w45427 & w45429;
assign w45431 = pi01272 & ~pi10443;
assign w45432 = ~pi10469 & ~w45431;
assign w45433 = ~pi10585 & w12874;
assign w45434 = ~w142 & ~w45433;
assign w45435 = pi10471 & ~w1193;
assign w45436 = ~pi00090 & pi09928;
assign w45437 = ~w45435 & ~w45436;
assign w45438 = ~pi10473 & w1204;
assign w45439 = ~w1208 & w45438;
assign w45440 = pi10439 & ~pi10475;
assign w45441 = ~w2178 & ~w45440;
assign w45442 = ~pi10476 & ~pi10523;
assign w45443 = ~pi10470 & ~w45442;
assign w45444 = ~pi00869 & ~pi10477;
assign w45445 = ~pi00434 & pi00869;
assign w45446 = ~w45444 & ~w45445;
assign w45447 = ~pi00845 & pi10481;
assign w45448 = ~pi10381 & ~w45447;
assign w45449 = ~pi00869 & ~pi10482;
assign w45450 = pi00869 & ~pi10437;
assign w45451 = ~w45449 & ~w45450;
assign w45452 = pi00232 & pi00869;
assign w45453 = ~pi00869 & ~pi10521;
assign w45454 = ~w45452 & ~w45453;
assign w45455 = ~pi00869 & ~pi10522;
assign w45456 = ~pi00000 & pi00869;
assign w45457 = ~w45455 & ~w45456;
assign w45458 = ~pi10470 & pi10523;
assign w45459 = pi10004 & ~w45458;
assign w45460 = pi00204 & pi00869;
assign w45461 = ~pi00869 & ~pi10524;
assign w45462 = ~w45460 & ~w45461;
assign w45463 = pi01253 & pi01261;
assign w45464 = pi00053 & pi10535;
assign w45465 = pi01165 & pi10381;
assign w45466 = ~w45464 & ~w45465;
assign w45467 = pi00869 & pi10005;
assign w45468 = ~pi00869 & ~pi10536;
assign w45469 = ~w45467 & ~w45468;
assign w45470 = pi00869 & pi09923;
assign w45471 = ~pi00869 & ~pi10537;
assign w45472 = ~w45470 & ~w45471;
assign w45473 = ~pi00869 & ~pi10538;
assign w45474 = ~pi00357 & pi00869;
assign w45475 = ~w45473 & ~w45474;
assign w45476 = pi00869 & pi00970;
assign w45477 = ~pi00869 & ~pi10541;
assign w45478 = ~w45476 & ~w45477;
assign w45479 = pi04204 & w3562;
assign w45480 = pi07065 & w3466;
assign w45481 = pi07889 & w3560;
assign w45482 = pi04001 & w3574;
assign w45483 = pi09685 & w3071;
assign w45484 = pi07197 & w3225;
assign w45485 = pi07265 & w3358;
assign w45486 = pi03798 & w3137;
assign w45487 = pi03662 & w3362;
assign w45488 = pi02273 & w3418;
assign w45489 = pi06568 & w3344;
assign w45490 = pi03740 & w3322;
assign w45491 = pi02559 & w3184;
assign w45492 = pi07717 & w3584;
assign w45493 = pi01905 & w3424;
assign w45494 = pi07100 & w3340;
assign w45495 = pi03577 & w3544;
assign w45496 = pi04139 & w3328;
assign w45497 = pi06817 & w3199;
assign w45498 = pi06758 & w3450;
assign w45499 = pi03598 & w3268;
assign w45500 = pi02631 & w3188;
assign w45501 = pi04038 & w3181;
assign w45502 = pi01707 & w3384;
assign w45503 = pi07289 & w3276;
assign w45504 = pi06693 & w3460;
assign w45505 = pi06684 & w3356;
assign w45506 = pi03558 & w3197;
assign w45507 = pi03962 & w3394;
assign w45508 = pi06804 & w3203;
assign w45509 = pi07335 & w3165;
assign w45510 = pi07527 & w3596;
assign w45511 = pi04007 & w3494;
assign w45512 = pi04086 & w3326;
assign w45513 = pi09553 & w3456;
assign w45514 = pi07598 & w3616;
assign w45515 = pi03844 & w3548;
assign w45516 = pi04270 & w3556;
assign w45517 = pi06843 & w3227;
assign w45518 = pi07632 & w3446;
assign w45519 = pi07381 & w3194;
assign w45520 = pi07274 & w3448;
assign w45521 = pi02046 & w3520;
assign w45522 = pi02525 & w3594;
assign w45523 = pi07752 & w3320;
assign w45524 = pi03675 & w3404;
assign w45525 = pi01705 & w3332;
assign w45526 = pi06737 & w3314;
assign w45527 = pi03831 & w3310;
assign w45528 = pi06483 & w3232;
assign w45529 = pi06876 & w3153;
assign w45530 = pi04014 & w3428;
assign w45531 = pi08130 & w3242;
assign w45532 = pi08563 & w3207;
assign w45533 = pi03818 & w3260;
assign w45534 = pi06811 & w3129;
assign w45535 = pi06654 & w3480;
assign w45536 = pi03517 & w3306;
assign w45537 = pi02641 & w3438;
assign w45538 = pi06794 & w3392;
assign w45539 = pi06765 & w3236;
assign w45540 = pi07626 & w3606;
assign w45541 = pi07837 & w3318;
assign w45542 = pi06647 & w3288;
assign w45543 = pi03981 & w3118;
assign w45544 = pi03811 & w3292;
assign w45545 = pi03772 & w3536;
assign w45546 = pi07306 & w3508;
assign w45547 = pi04126 & w3115;
assign w45548 = pi07319 & w3312;
assign w45549 = pi07908 & w3148;
assign w45550 = pi03889 & w3576;
assign w45551 = pi02507 & w3580;
assign w45552 = pi04080 & w3290;
assign w45553 = pi07540 & w3093;
assign w45554 = pi08041 & w3524;
assign w45555 = pi07078 & w3139;
assign w45556 = pi03915 & w3348;
assign w45557 = pi04133 & w3190;
assign w45558 = pi07350 & w3201;
assign w45559 = pi03837 & w3244;
assign w45560 = pi03949 & w3498;
assign w45561 = pi06832 & w3422;
assign w45562 = pi06518 & w3308;
assign w45563 = pi03896 & w3209;
assign w45564 = pi06527 & w3436;
assign w45565 = pi07297 & w3434;
assign w45566 = pi07521 & w3352;
assign w45567 = pi07113 & w3286;
assign w45568 = pi04329 & w3488;
assign w45569 = pi06490 & w3240;
assign w45570 = pi02579 & w3254;
assign w45571 = pi07091 & w3572;
assign w45572 = pi07055 & w3234;
assign w45573 = pi04314 & w3211;
assign w45574 = pi06557 & w3604;
assign w45575 = pi09766 & w3398;
assign w45576 = pi02301 & w3406;
assign w45577 = pi07670 & w3366;
assign w45578 = pi07138 & w3410;
assign w45579 = pi04224 & w3258;
assign w45580 = pi09784 & w3602;
assign w45581 = pi03903 & w3338;
assign w45582 = pi06858 & w3462;
assign w45583 = pi06720 & w3540;
assign w45584 = pi07358 & w3372;
assign w45585 = pi07939 & w3324;
assign w45586 = pi01600 & w3158;
assign w45587 = pi06579 & w3492;
assign w45588 = pi06974 & w3256;
assign w45589 = pi08022 & w3368;
assign w45590 = pi03863 & w3350;
assign w45591 = pi07826 & w3096;
assign w45592 = pi03727 & w3534;
assign w45593 = pi03681 & w3330;
assign w45594 = pi06634 & w3550;
assign w45595 = pi08004 & w3179;
assign w45596 = pi06674 & w3378;
assign w45597 = pi04120 & w3086;
assign w45598 = pi04217 & w3302;
assign w45599 = pi04230 & w3122;
assign w45600 = pi06547 & w3598;
assign w45601 = pi02805 & w3127;
assign w45602 = pi07222 & w3221;
assign w45603 = pi08062 & w3246;
assign w45604 = pi03694 & w3530;
assign w45605 = pi07918 & w3294;
assign w45606 = pi07785 & w3546;
assign w45607 = pi07401 & w3430;
assign w45608 = pi03936 & w3592;
assign w45609 = pi02484 & w3173;
assign w45610 = pi06497 & w3266;
assign w45611 = pi03701 & w3250;
assign w45612 = pi03588 & w3500;
assign w45613 = pi02107 & w3376;
assign w45614 = pi07236 & w3620;
assign w45615 = pi06996 & w3442;
assign w45616 = pi07494 & w3270;
assign w45617 = pi06614 & w3554;
assign w45618 = pi07558 & w3426;
assign w45619 = pi03531 & w3380;
assign w45620 = pi03753 & w3103;
assign w45621 = pi06641 & w3568;
assign w45622 = pi07371 & w3600;
assign w45623 = pi07811 & w3280;
assign w45624 = pi06983 & w3518;
assign w45625 = pi03507 & w3614;
assign w45626 = pi04770 & w3386;
assign w45627 = pi07039 & w3300;
assign w45628 = pi03733 & w3400;
assign w45629 = pi06934 & w3186;
assign w45630 = pi06896 & w3082;
assign w45631 = pi07280 & w3566;
assign w45632 = pi07313 & w3167;
assign w45633 = pi01822 & w3264;
assign w45634 = pi07584 & w3532;
assign w45635 = pi07759 & w3478;
assign w45636 = pi04278 & w3388;
assign w45637 = pi02424 & w3238;
assign w45638 = pi04198 & w3412;
assign w45639 = pi08098 & w3558;
assign w45640 = pi04165 & w3146;
assign w45641 = pi03850 & w3490;
assign w45642 = pi07898 & w3342;
assign w45643 = pi03805 & w3262;
assign w45644 = pi07574 & w3474;
assign w45645 = pi01573 & w3432;
assign w45646 = pi04047 & w3502;
assign w45647 = pi07730 & w3106;
assign w45648 = pi02511 & w3382;
assign w45649 = pi08106 & w3408;
assign w45650 = pi06712 & w3414;
assign w45651 = pi07129 & w3552;
assign w45652 = pi06620 & w3452;
assign w45653 = pi07698 & w3468;
assign w45654 = pi07566 & w3516;
assign w45655 = pi08030 & w3160;
assign w45656 = pi06746 & w3538;
assign w45657 = pi06781 & w3354;
assign w45658 = pi06472 & w3486;
assign w45659 = pi06850 & w3304;
assign w45660 = pi07801 & w3542;
assign w45661 = pi03649 & w3470;
assign w45662 = pi06909 & w3278;
assign w45663 = pi04172 & w3564;
assign w45664 = pi04054 & w3454;
assign w45665 = pi06627 & w3528;
assign w45666 = pi01809 & w3476;
assign w45667 = pi04146 & w3484;
assign w45668 = pi07429 & w3458;
assign w45669 = pi02755 & w3162;
assign w45670 = pi07245 & w3272;
assign w45671 = pi08078 & w3110;
assign w45672 = pi06869 & w3496;
assign w45673 = pi07156 & w3135;
assign w45674 = pi07174 & w3156;
assign w45675 = pi07210 & w3472;
assign w45676 = pi07660 & w3608;
assign w45677 = pi07182 & w3205;
assign w45678 = pi07860 & w3402;
assign w45679 = pi03566 & w3336;
assign w45680 = pi06700 & w3586;
assign w45681 = pi06661 & w3217;
assign w45682 = pi04533 & w3578;
assign w45683 = pi07928 & w3316;
assign w45684 = pi03857 & w3526;
assign w45685 = pi07365 & w3374;
assign w45686 = pi04179 & w3370;
assign w45687 = pi07606 & w3175;
assign w45688 = pi07149 & w3420;
assign w45689 = pi06957 & w3078;
assign w45690 = pi07534 & w3125;
assign w45691 = pi04191 & w3512;
assign w45692 = pi07392 & w3590;
assign w45693 = pi01974 & w3064;
assign w45694 = pi04106 & w3214;
assign w45695 = pi03538 & w3346;
assign w45696 = pi07879 & w3229;
assign w45697 = pi07649 & w3440;
assign w45698 = pi06607 & w3219;
assign w45699 = pi04024 & w3522;
assign w45700 = pi06948 & w3284;
assign w45701 = pi07765 & w3282;
assign w45702 = pi07446 & w3192;
assign w45703 = pi01724 & w3612;
assign w45704 = pi07465 & w3390;
assign w45705 = pi06510 & w3143;
assign w45706 = pi04296 & w3588;
assign w45707 = pi06726 & w3482;
assign w45708 = pi07641 & w3570;
assign w45709 = pi08117 & w3510;
assign w45710 = pi06668 & w3112;
assign w45711 = pi06772 & w3298;
assign w45712 = pi09759 & w3506;
assign w45713 = pi06922 & w3514;
assign w45714 = pi08088 & w3150;
assign w45715 = pi07410 & w3171;
assign w45716 = pi07745 & w3444;
assign w45717 = pi04250 & w3504;
assign w45718 = pi09596 & w3464;
assign w45719 = pi04211 & w3169;
assign w45720 = pi04185 & w3618;
assign w45721 = pi03766 & w3274;
assign w45722 = pi09561 & w3334;
assign w45723 = pi09771 & w3364;
assign w45724 = pi04304 & w3396;
assign w45725 = pi03824 & w3610;
assign w45726 = pi04323 & w3582;
assign w45727 = pi07618 & w3223;
assign w45728 = pi06599 & w3252;
assign w45729 = pi04288 & w3177;
assign w45730 = pi03642 & w3416;
assign w45731 = pi07455 & w3360;
assign w45732 = pi03955 & w3132;
assign w45733 = pi06537 & w3248;
assign w45734 = pi03790 & w3296;
assign w45735 = ~w45479 & ~w45480;
assign w45736 = ~w45481 & ~w45482;
assign w45737 = ~w45483 & ~w45484;
assign w45738 = ~w45485 & ~w45486;
assign w45739 = ~w45487 & ~w45488;
assign w45740 = ~w45489 & ~w45490;
assign w45741 = ~w45491 & ~w45492;
assign w45742 = ~w45493 & ~w45494;
assign w45743 = ~w45495 & ~w45496;
assign w45744 = ~w45497 & ~w45498;
assign w45745 = ~w45499 & ~w45500;
assign w45746 = ~w45501 & ~w45502;
assign w45747 = ~w45503 & ~w45504;
assign w45748 = ~w45505 & ~w45506;
assign w45749 = ~w45507 & ~w45508;
assign w45750 = ~w45509 & ~w45510;
assign w45751 = ~w45511 & ~w45512;
assign w45752 = ~w45513 & ~w45514;
assign w45753 = ~w45515 & ~w45516;
assign w45754 = ~w45517 & ~w45518;
assign w45755 = ~w45519 & ~w45520;
assign w45756 = ~w45521 & ~w45522;
assign w45757 = ~w45523 & ~w45524;
assign w45758 = ~w45525 & ~w45526;
assign w45759 = ~w45527 & ~w45528;
assign w45760 = ~w45529 & ~w45530;
assign w45761 = ~w45531 & ~w45532;
assign w45762 = ~w45533 & ~w45534;
assign w45763 = ~w45535 & ~w45536;
assign w45764 = ~w45537 & ~w45538;
assign w45765 = ~w45539 & ~w45540;
assign w45766 = ~w45541 & ~w45542;
assign w45767 = ~w45543 & ~w45544;
assign w45768 = ~w45545 & ~w45546;
assign w45769 = ~w45547 & ~w45548;
assign w45770 = ~w45549 & ~w45550;
assign w45771 = ~w45551 & ~w45552;
assign w45772 = ~w45553 & ~w45554;
assign w45773 = ~w45555 & ~w45556;
assign w45774 = ~w45557 & ~w45558;
assign w45775 = ~w45559 & ~w45560;
assign w45776 = ~w45561 & ~w45562;
assign w45777 = ~w45563 & ~w45564;
assign w45778 = ~w45565 & ~w45566;
assign w45779 = ~w45567 & ~w45568;
assign w45780 = ~w45569 & ~w45570;
assign w45781 = ~w45571 & ~w45572;
assign w45782 = ~w45573 & ~w45574;
assign w45783 = ~w45575 & ~w45576;
assign w45784 = ~w45577 & ~w45578;
assign w45785 = ~w45579 & ~w45580;
assign w45786 = ~w45581 & ~w45582;
assign w45787 = ~w45583 & ~w45584;
assign w45788 = ~w45585 & ~w45586;
assign w45789 = ~w45587 & ~w45588;
assign w45790 = ~w45589 & ~w45590;
assign w45791 = ~w45591 & ~w45592;
assign w45792 = ~w45593 & ~w45594;
assign w45793 = ~w45595 & ~w45596;
assign w45794 = ~w45597 & ~w45598;
assign w45795 = ~w45599 & ~w45600;
assign w45796 = ~w45601 & ~w45602;
assign w45797 = ~w45603 & ~w45604;
assign w45798 = ~w45605 & ~w45606;
assign w45799 = ~w45607 & ~w45608;
assign w45800 = ~w45609 & ~w45610;
assign w45801 = ~w45611 & ~w45612;
assign w45802 = ~w45613 & ~w45614;
assign w45803 = ~w45615 & ~w45616;
assign w45804 = ~w45617 & ~w45618;
assign w45805 = ~w45619 & ~w45620;
assign w45806 = ~w45621 & ~w45622;
assign w45807 = ~w45623 & ~w45624;
assign w45808 = ~w45625 & ~w45626;
assign w45809 = ~w45627 & ~w45628;
assign w45810 = ~w45629 & ~w45630;
assign w45811 = ~w45631 & ~w45632;
assign w45812 = ~w45633 & ~w45634;
assign w45813 = ~w45635 & ~w45636;
assign w45814 = ~w45637 & ~w45638;
assign w45815 = ~w45639 & ~w45640;
assign w45816 = ~w45641 & ~w45642;
assign w45817 = ~w45643 & ~w45644;
assign w45818 = ~w45645 & ~w45646;
assign w45819 = ~w45647 & ~w45648;
assign w45820 = ~w45649 & ~w45650;
assign w45821 = ~w45651 & ~w45652;
assign w45822 = ~w45653 & ~w45654;
assign w45823 = ~w45655 & ~w45656;
assign w45824 = ~w45657 & ~w45658;
assign w45825 = ~w45659 & ~w45660;
assign w45826 = ~w45661 & ~w45662;
assign w45827 = ~w45663 & ~w45664;
assign w45828 = ~w45665 & ~w45666;
assign w45829 = ~w45667 & ~w45668;
assign w45830 = ~w45669 & ~w45670;
assign w45831 = ~w45671 & ~w45672;
assign w45832 = ~w45673 & ~w45674;
assign w45833 = ~w45675 & ~w45676;
assign w45834 = ~w45677 & ~w45678;
assign w45835 = ~w45679 & ~w45680;
assign w45836 = ~w45681 & ~w45682;
assign w45837 = ~w45683 & ~w45684;
assign w45838 = ~w45685 & ~w45686;
assign w45839 = ~w45687 & ~w45688;
assign w45840 = ~w45689 & ~w45690;
assign w45841 = ~w45691 & ~w45692;
assign w45842 = ~w45693 & ~w45694;
assign w45843 = ~w45695 & ~w45696;
assign w45844 = ~w45697 & ~w45698;
assign w45845 = ~w45699 & ~w45700;
assign w45846 = ~w45701 & ~w45702;
assign w45847 = ~w45703 & ~w45704;
assign w45848 = ~w45705 & ~w45706;
assign w45849 = ~w45707 & ~w45708;
assign w45850 = ~w45709 & ~w45710;
assign w45851 = ~w45711 & ~w45712;
assign w45852 = ~w45713 & ~w45714;
assign w45853 = ~w45715 & ~w45716;
assign w45854 = ~w45717 & ~w45718;
assign w45855 = ~w45719 & ~w45720;
assign w45856 = ~w45721 & ~w45722;
assign w45857 = ~w45723 & ~w45724;
assign w45858 = ~w45725 & ~w45726;
assign w45859 = ~w45727 & ~w45728;
assign w45860 = ~w45729 & ~w45730;
assign w45861 = ~w45731 & ~w45732;
assign w45862 = ~w45733 & ~w45734;
assign w45863 = w45861 & w45862;
assign w45864 = w45859 & w45860;
assign w45865 = w45857 & w45858;
assign w45866 = w45855 & w45856;
assign w45867 = w45853 & w45854;
assign w45868 = w45851 & w45852;
assign w45869 = w45849 & w45850;
assign w45870 = w45847 & w45848;
assign w45871 = w45845 & w45846;
assign w45872 = w45843 & w45844;
assign w45873 = w45841 & w45842;
assign w45874 = w45839 & w45840;
assign w45875 = w45837 & w45838;
assign w45876 = w45835 & w45836;
assign w45877 = w45833 & w45834;
assign w45878 = w45831 & w45832;
assign w45879 = w45829 & w45830;
assign w45880 = w45827 & w45828;
assign w45881 = w45825 & w45826;
assign w45882 = w45823 & w45824;
assign w45883 = w45821 & w45822;
assign w45884 = w45819 & w45820;
assign w45885 = w45817 & w45818;
assign w45886 = w45815 & w45816;
assign w45887 = w45813 & w45814;
assign w45888 = w45811 & w45812;
assign w45889 = w45809 & w45810;
assign w45890 = w45807 & w45808;
assign w45891 = w45805 & w45806;
assign w45892 = w45803 & w45804;
assign w45893 = w45801 & w45802;
assign w45894 = w45799 & w45800;
assign w45895 = w45797 & w45798;
assign w45896 = w45795 & w45796;
assign w45897 = w45793 & w45794;
assign w45898 = w45791 & w45792;
assign w45899 = w45789 & w45790;
assign w45900 = w45787 & w45788;
assign w45901 = w45785 & w45786;
assign w45902 = w45783 & w45784;
assign w45903 = w45781 & w45782;
assign w45904 = w45779 & w45780;
assign w45905 = w45777 & w45778;
assign w45906 = w45775 & w45776;
assign w45907 = w45773 & w45774;
assign w45908 = w45771 & w45772;
assign w45909 = w45769 & w45770;
assign w45910 = w45767 & w45768;
assign w45911 = w45765 & w45766;
assign w45912 = w45763 & w45764;
assign w45913 = w45761 & w45762;
assign w45914 = w45759 & w45760;
assign w45915 = w45757 & w45758;
assign w45916 = w45755 & w45756;
assign w45917 = w45753 & w45754;
assign w45918 = w45751 & w45752;
assign w45919 = w45749 & w45750;
assign w45920 = w45747 & w45748;
assign w45921 = w45745 & w45746;
assign w45922 = w45743 & w45744;
assign w45923 = w45741 & w45742;
assign w45924 = w45739 & w45740;
assign w45925 = w45737 & w45738;
assign w45926 = w45735 & w45736;
assign w45927 = w45925 & w45926;
assign w45928 = w45923 & w45924;
assign w45929 = w45921 & w45922;
assign w45930 = w45919 & w45920;
assign w45931 = w45917 & w45918;
assign w45932 = w45915 & w45916;
assign w45933 = w45913 & w45914;
assign w45934 = w45911 & w45912;
assign w45935 = w45909 & w45910;
assign w45936 = w45907 & w45908;
assign w45937 = w45905 & w45906;
assign w45938 = w45903 & w45904;
assign w45939 = w45901 & w45902;
assign w45940 = w45899 & w45900;
assign w45941 = w45897 & w45898;
assign w45942 = w45895 & w45896;
assign w45943 = w45893 & w45894;
assign w45944 = w45891 & w45892;
assign w45945 = w45889 & w45890;
assign w45946 = w45887 & w45888;
assign w45947 = w45885 & w45886;
assign w45948 = w45883 & w45884;
assign w45949 = w45881 & w45882;
assign w45950 = w45879 & w45880;
assign w45951 = w45877 & w45878;
assign w45952 = w45875 & w45876;
assign w45953 = w45873 & w45874;
assign w45954 = w45871 & w45872;
assign w45955 = w45869 & w45870;
assign w45956 = w45867 & w45868;
assign w45957 = w45865 & w45866;
assign w45958 = w45863 & w45864;
assign w45959 = w45957 & w45958;
assign w45960 = w45955 & w45956;
assign w45961 = w45953 & w45954;
assign w45962 = w45951 & w45952;
assign w45963 = w45949 & w45950;
assign w45964 = w45947 & w45948;
assign w45965 = w45945 & w45946;
assign w45966 = w45943 & w45944;
assign w45967 = w45941 & w45942;
assign w45968 = w45939 & w45940;
assign w45969 = w45937 & w45938;
assign w45970 = w45935 & w45936;
assign w45971 = w45933 & w45934;
assign w45972 = w45931 & w45932;
assign w45973 = w45929 & w45930;
assign w45974 = w45927 & w45928;
assign w45975 = w45973 & w45974;
assign w45976 = w45971 & w45972;
assign w45977 = w45969 & w45970;
assign w45978 = w45967 & w45968;
assign w45979 = w45965 & w45966;
assign w45980 = w45963 & w45964;
assign w45981 = w45961 & w45962;
assign w45982 = w45959 & w45960;
assign w45983 = w45981 & w45982;
assign w45984 = w45979 & w45980;
assign w45985 = w45977 & w45978;
assign w45986 = w45975 & w45976;
assign w45987 = w45985 & w45986;
assign w45988 = w45983 & w45984;
assign w45989 = w45987 & w45988;
assign w45990 = ~pi10577 & ~w45989;
assign w45991 = pi03758 & w3526;
assign w45992 = pi06914 & w3300;
assign w45993 = pi04096 & w3522;
assign w45994 = pi07324 & w3620;
assign w45995 = pi02204 & w3197;
assign w45996 = pi06409 & w3392;
assign w45997 = pi08153 & w3366;
assign w45998 = pi04342 & w3115;
assign w45999 = pi07711 & w3171;
assign w46000 = pi08271 & w3580;
assign w46001 = pi07857 & w3386;
assign w46002 = pi08005 & w3474;
assign w46003 = pi08251 & w3318;
assign w46004 = pi02230 & w3175;
assign w46005 = pi03654 & w3260;
assign w46006 = pi05840 & w3248;
assign w46007 = pi08342 & w3578;
assign w46008 = pi08033 & w3532;
assign w46009 = pi06863 & w3442;
assign w46010 = pi07842 & w3270;
assign w46011 = pi04072 & w3428;
assign w46012 = pi06357 & w3450;
assign w46013 = pi02192 & w3544;
assign w46014 = pi03987 & w3132;
assign w46015 = pi04501 & w3582;
assign w46016 = pi07053 & w3286;
assign w46017 = pi05733 & w3266;
assign w46018 = pi08047 & w3616;
assign w46019 = pi06109 & w3288;
assign w46020 = pi06456 & w3129;
assign w46021 = pi06978 & w3139;
assign w46022 = pi02219 & w3380;
assign w46023 = pi04335 & w3086;
assign w46024 = pi06751 & w3186;
assign w46025 = pi08316 & w3324;
assign w46026 = pi06169 & w3378;
assign w46027 = pi08211 & w3282;
assign w46028 = pi03615 & w3296;
assign w46029 = pi06089 & w3568;
assign w46030 = pi06939 & w3234;
assign w46031 = pi02532 & w3254;
assign w46032 = pi03451 & w3530;
assign w46033 = pi06180 & w3356;
assign w46034 = pi07397 & w3448;
assign w46035 = pi04383 & w3370;
assign w46036 = pi04236 & w3290;
assign w46037 = pi03622 & w3137;
assign w46038 = pi03782 & w3350;
assign w46039 = pi07612 & w3374;
assign w46040 = pi04403 & w3412;
assign w46041 = pi07642 & w3600;
assign w46042 = pi08232 & w3542;
assign w46043 = pi06068 & w3528;
assign w46044 = pi06371 & w3236;
assign w46045 = pi05994 & w3219;
assign w46046 = pi08395 & w3110;
assign w46047 = pi08198 & w3320;
assign w46048 = pi07291 & w3221;
assign w46049 = pi03635 & w3292;
assign w46050 = pi08428 & w3242;
assign w46051 = pi07995 & w3516;
assign w46052 = pi02058 & w3534;
assign w46053 = pi04436 & w3122;
assign w46054 = pi08205 & w3478;
assign w46055 = pi06277 & w3540;
assign w46056 = pi08159 & w3594;
assign w46057 = pi08258 & w3188;
assign w46058 = pi07238 & w3225;
assign w46059 = pi07443 & w3434;
assign w46060 = pi05693 & w3232;
assign w46061 = pi07956 & w3093;
assign w46062 = pi02231 & w3306;
assign w46063 = pi08290 & w3342;
assign w46064 = pi06834 & w3518;
assign w46065 = pi06538 & w3304;
assign w46066 = pi03869 & w3576;
assign w46067 = pi06396 & w3354;
assign w46068 = pi07790 & w3360;
assign w46069 = pi03523 & w3400;
assign w46070 = pi02179 & w3500;
assign w46071 = pi07345 & w3376;
assign w46072 = pi04321 & w3602;
assign w46073 = pi03491 & w3064;
assign w46074 = pi03706 & w3244;
assign w46075 = pi03479 & w3250;
assign w46076 = pi06318 & w3314;
assign w46077 = pi07816 & w3464;
assign w46078 = pi04481 & w3588;
assign w46079 = pi05820 & w3436;
assign w46080 = pi02171 & w3268;
assign w46081 = pi06926 & w3398;
assign w46082 = pi07020 & w3340;
assign w46083 = pi07139 & w3135;
assign w46084 = pi08389 & w3246;
assign w46085 = pi04429 & w3258;
assign w46086 = pi02218 & w3346;
assign w46087 = pi04410 & w3562;
assign w46088 = pi03405 & w3330;
assign w46089 = pi07417 & w3566;
assign w46090 = pi08185 & w3106;
assign w46091 = pi05927 & w3344;
assign w46092 = pi03719 & w3548;
assign w46093 = pi04449 & w3504;
assign w46094 = pi08264 & w3402;
assign w46095 = pi08091 & w3606;
assign w46096 = pi04376 & w3564;
assign w46097 = pi04151 & w3502;
assign w46098 = pi01754 & w3201;
assign w46099 = pi08356 & w3438;
assign w46100 = pi04355 & w3328;
assign w46101 = pi08217 & w3264;
assign w46102 = pi06129 & w3480;
assign w46103 = pi04390 & w3618;
assign w46104 = pi06574 & w3496;
assign w46105 = pi08382 & w3418;
assign w46106 = pi06426 & w3203;
assign w46107 = pi06888 & w3432;
assign w46108 = pi09606 & w3272;
assign w46109 = pi06298 & w3482;
assign w46110 = pi08297 & w3148;
assign w46111 = pi06732 & w3514;
assign w46112 = pi08073 & w3223;
assign w46113 = pi06952 & w3466;
assign w46114 = pi07259 & w3472;
assign w46115 = pi08329 & w3158;
assign w46116 = pi07674 & w3426;
assign w46117 = pi07111 & w3410;
assign w46118 = pi03909 & w3348;
assign w46119 = pi06029 & w3554;
assign w46120 = pi08224 & w3546;
assign w46121 = pi07916 & w3596;
assign w46122 = pi07503 & w3312;
assign w46123 = pi08166 & w3468;
assign w46124 = pi02207 & w3614;
assign w46125 = pi03667 & w3610;
assign w46126 = pi04423 & w3302;
assign w46127 = pi04307 & w3214;
assign w46128 = pi08277 & w3229;
assign w46129 = pi06780 & w3284;
assign w46130 = pi07464 & w3508;
assign w46131 = pi02199 & w3336;
assign w46132 = pi02654 & w3207;
assign w46133 = pi06082 & w3550;
assign w46134 = pi08172 & w3173;
assign w46135 = pi06823 & w3256;
assign w46136 = pi03882 & w3338;
assign w46137 = pi01496 & w3570;
assign w46138 = pi04348 & w3190;
assign w46139 = pi06502 & w3422;
assign w46140 = pi04281 & w3334;
assign w46141 = pi08284 & w3560;
assign w46142 = pi03352 & w3470;
assign w46143 = pi07938 & w3125;
assign w46144 = pi07739 & w3458;
assign w46145 = pi07877 & w3382;
assign w46146 = pi08111 & w3446;
assign w46147 = pi06558 & w3462;
assign w46148 = pi03745 & w3490;
assign w46149 = pi04455 & w3184;
assign w46150 = pi04059 & w3574;
assign w46151 = pi04361 & w3484;
assign w46152 = pi03628 & w3262;
assign w46153 = pi06154 & w3112;
assign w46154 = pi07378 & w3358;
assign w46155 = pi07435 & w3276;
assign w46156 = pi06383 & w3298;
assign w46157 = pi07099 & w3552;
assign w46158 = pi08179 & w3584;
assign w46159 = pi07680 & w3590;
assign w46160 = pi04112 & w3181;
assign w46161 = pi07198 & w3156;
assign w46162 = pi08303 & w3294;
assign w46163 = pi08146 & w3608;
assign w46164 = pi05972 & w3252;
assign w46165 = pi05879 & w3604;
assign w46166 = pi06706 & w3278;
assign w46167 = pi07168 & w3364;
assign w46168 = pi08238 & w3280;
assign w46169 = pi04494 & w3211;
assign w46170 = pi08408 & w3558;
assign w46171 = pi08370 & w3160;
assign w46172 = pi02028 & w3536;
assign w46173 = pi04255 & w3326;
assign w46174 = pi04368 & w3146;
assign w46175 = pi03687 & w3310;
assign w46176 = pi03544 & w3322;
assign w46177 = pi08192 & w3444;
assign w46178 = pi07211 & w3205;
assign w46179 = pi03875 & w3209;
assign w46180 = pi02646 & w3238;
assign w46181 = pi04488 & w3396;
assign w46182 = pi05946 & w3492;
assign w46183 = pi08138 & w3440;
assign w46184 = pi06331 & w3538;
assign w46185 = pi04462 & w3556;
assign w46186 = pi01816 & w3308;
assign w46187 = pi07798 & w3390;
assign w46188 = pi07123 & w3420;
assign w46189 = pi04468 & w3388;
assign w46190 = pi02177 & w3162;
assign w46191 = pi06049 & w3452;
assign w46192 = pi08415 & w3408;
assign w46193 = pi03993 & w3394;
assign w46194 = pi04475 & w3177;
assign w46195 = pi04507 & w3488;
assign w46196 = pi07006 & w3572;
assign w46197 = pi03925 & w3456;
assign w46198 = pi05720 & w3240;
assign w46199 = pi08310 & w3316;
assign w46200 = pi03967 & w3498;
assign w46201 = pi04033 & w3118;
assign w46202 = pi08402 & w3150;
assign w46203 = pi05859 & w3598;
assign w46204 = pi08421 & w3510;
assign w46205 = pi03199 & w3520;
assign w46206 = pi03941 & w3592;
assign w46207 = pi06793 & w3078;
assign w46208 = pi07549 & w3165;
assign w46209 = pi06992 & w3406;
assign w46210 = pi08323 & w3332;
assign w46211 = pi05673 & w3486;
assign w46212 = pi08363 & w3368;
assign w46213 = pi05959 & w3612;
assign w46214 = pi07484 & w3167;
assign w46215 = pi04158 & w3454;
assign w46216 = pi08376 & w3524;
assign w46217 = pi01851 & w3143;
assign w46218 = pi04416 & w3169;
assign w46219 = pi03567 & w3103;
assign w46220 = pi07725 & w3476;
assign w46221 = pi03583 & w3274;
assign w46222 = pi06519 & w3227;
assign w46223 = pi03609 & w3424;
assign w46224 = pi03346 & w3416;
assign w46225 = pi02633 & w3179;
assign w46226 = pi01627 & w3372;
assign w46227 = pi03365 & w3362;
assign w46228 = pi01656 & w3217;
assign w46229 = pi01617 & w3153;
assign w46230 = pi06196 & w3460;
assign w46231 = pi06966 & w3127;
assign w46232 = pi02639 & w3506;
assign w46233 = pi06881 & w3384;
assign w46234 = pi07896 & w3352;
assign w46235 = pi06471 & w3199;
assign w46236 = pi07662 & w3194;
assign w46237 = pi04396 & w3512;
assign w46238 = pi04020 & w3071;
assign w46239 = pi08245 & w3096;
assign w46240 = pi01765 & w3192;
assign w46241 = pi09735 & w3082;
assign w46242 = pi04066 & w3494;
assign w46243 = pi06255 & w3414;
assign w46244 = pi06209 & w3586;
assign w46245 = pi07690 & w3430;
assign w46246 = pi02113 & w3404;
assign w46247 = ~w45991 & ~w45992;
assign w46248 = ~w45993 & ~w45994;
assign w46249 = ~w45995 & ~w45996;
assign w46250 = ~w45997 & ~w45998;
assign w46251 = ~w45999 & ~w46000;
assign w46252 = ~w46001 & ~w46002;
assign w46253 = ~w46003 & ~w46004;
assign w46254 = ~w46005 & ~w46006;
assign w46255 = ~w46007 & ~w46008;
assign w46256 = ~w46009 & ~w46010;
assign w46257 = ~w46011 & ~w46012;
assign w46258 = ~w46013 & ~w46014;
assign w46259 = ~w46015 & ~w46016;
assign w46260 = ~w46017 & ~w46018;
assign w46261 = ~w46019 & ~w46020;
assign w46262 = ~w46021 & ~w46022;
assign w46263 = ~w46023 & ~w46024;
assign w46264 = ~w46025 & ~w46026;
assign w46265 = ~w46027 & ~w46028;
assign w46266 = ~w46029 & ~w46030;
assign w46267 = ~w46031 & ~w46032;
assign w46268 = ~w46033 & ~w46034;
assign w46269 = ~w46035 & ~w46036;
assign w46270 = ~w46037 & ~w46038;
assign w46271 = ~w46039 & ~w46040;
assign w46272 = ~w46041 & ~w46042;
assign w46273 = ~w46043 & ~w46044;
assign w46274 = ~w46045 & ~w46046;
assign w46275 = ~w46047 & ~w46048;
assign w46276 = ~w46049 & ~w46050;
assign w46277 = ~w46051 & ~w46052;
assign w46278 = ~w46053 & ~w46054;
assign w46279 = ~w46055 & ~w46056;
assign w46280 = ~w46057 & ~w46058;
assign w46281 = ~w46059 & ~w46060;
assign w46282 = ~w46061 & ~w46062;
assign w46283 = ~w46063 & ~w46064;
assign w46284 = ~w46065 & ~w46066;
assign w46285 = ~w46067 & ~w46068;
assign w46286 = ~w46069 & ~w46070;
assign w46287 = ~w46071 & ~w46072;
assign w46288 = ~w46073 & ~w46074;
assign w46289 = ~w46075 & ~w46076;
assign w46290 = ~w46077 & ~w46078;
assign w46291 = ~w46079 & ~w46080;
assign w46292 = ~w46081 & ~w46082;
assign w46293 = ~w46083 & ~w46084;
assign w46294 = ~w46085 & ~w46086;
assign w46295 = ~w46087 & ~w46088;
assign w46296 = ~w46089 & ~w46090;
assign w46297 = ~w46091 & ~w46092;
assign w46298 = ~w46093 & ~w46094;
assign w46299 = ~w46095 & ~w46096;
assign w46300 = ~w46097 & ~w46098;
assign w46301 = ~w46099 & ~w46100;
assign w46302 = ~w46101 & ~w46102;
assign w46303 = ~w46103 & ~w46104;
assign w46304 = ~w46105 & ~w46106;
assign w46305 = ~w46107 & ~w46108;
assign w46306 = ~w46109 & ~w46110;
assign w46307 = ~w46111 & ~w46112;
assign w46308 = ~w46113 & ~w46114;
assign w46309 = ~w46115 & ~w46116;
assign w46310 = ~w46117 & ~w46118;
assign w46311 = ~w46119 & ~w46120;
assign w46312 = ~w46121 & ~w46122;
assign w46313 = ~w46123 & ~w46124;
assign w46314 = ~w46125 & ~w46126;
assign w46315 = ~w46127 & ~w46128;
assign w46316 = ~w46129 & ~w46130;
assign w46317 = ~w46131 & ~w46132;
assign w46318 = ~w46133 & ~w46134;
assign w46319 = ~w46135 & ~w46136;
assign w46320 = ~w46137 & ~w46138;
assign w46321 = ~w46139 & ~w46140;
assign w46322 = ~w46141 & ~w46142;
assign w46323 = ~w46143 & ~w46144;
assign w46324 = ~w46145 & ~w46146;
assign w46325 = ~w46147 & ~w46148;
assign w46326 = ~w46149 & ~w46150;
assign w46327 = ~w46151 & ~w46152;
assign w46328 = ~w46153 & ~w46154;
assign w46329 = ~w46155 & ~w46156;
assign w46330 = ~w46157 & ~w46158;
assign w46331 = ~w46159 & ~w46160;
assign w46332 = ~w46161 & ~w46162;
assign w46333 = ~w46163 & ~w46164;
assign w46334 = ~w46165 & ~w46166;
assign w46335 = ~w46167 & ~w46168;
assign w46336 = ~w46169 & ~w46170;
assign w46337 = ~w46171 & ~w46172;
assign w46338 = ~w46173 & ~w46174;
assign w46339 = ~w46175 & ~w46176;
assign w46340 = ~w46177 & ~w46178;
assign w46341 = ~w46179 & ~w46180;
assign w46342 = ~w46181 & ~w46182;
assign w46343 = ~w46183 & ~w46184;
assign w46344 = ~w46185 & ~w46186;
assign w46345 = ~w46187 & ~w46188;
assign w46346 = ~w46189 & ~w46190;
assign w46347 = ~w46191 & ~w46192;
assign w46348 = ~w46193 & ~w46194;
assign w46349 = ~w46195 & ~w46196;
assign w46350 = ~w46197 & ~w46198;
assign w46351 = ~w46199 & ~w46200;
assign w46352 = ~w46201 & ~w46202;
assign w46353 = ~w46203 & ~w46204;
assign w46354 = ~w46205 & ~w46206;
assign w46355 = ~w46207 & ~w46208;
assign w46356 = ~w46209 & ~w46210;
assign w46357 = ~w46211 & ~w46212;
assign w46358 = ~w46213 & ~w46214;
assign w46359 = ~w46215 & ~w46216;
assign w46360 = ~w46217 & ~w46218;
assign w46361 = ~w46219 & ~w46220;
assign w46362 = ~w46221 & ~w46222;
assign w46363 = ~w46223 & ~w46224;
assign w46364 = ~w46225 & ~w46226;
assign w46365 = ~w46227 & ~w46228;
assign w46366 = ~w46229 & ~w46230;
assign w46367 = ~w46231 & ~w46232;
assign w46368 = ~w46233 & ~w46234;
assign w46369 = ~w46235 & ~w46236;
assign w46370 = ~w46237 & ~w46238;
assign w46371 = ~w46239 & ~w46240;
assign w46372 = ~w46241 & ~w46242;
assign w46373 = ~w46243 & ~w46244;
assign w46374 = ~w46245 & ~w46246;
assign w46375 = w46373 & w46374;
assign w46376 = w46371 & w46372;
assign w46377 = w46369 & w46370;
assign w46378 = w46367 & w46368;
assign w46379 = w46365 & w46366;
assign w46380 = w46363 & w46364;
assign w46381 = w46361 & w46362;
assign w46382 = w46359 & w46360;
assign w46383 = w46357 & w46358;
assign w46384 = w46355 & w46356;
assign w46385 = w46353 & w46354;
assign w46386 = w46351 & w46352;
assign w46387 = w46349 & w46350;
assign w46388 = w46347 & w46348;
assign w46389 = w46345 & w46346;
assign w46390 = w46343 & w46344;
assign w46391 = w46341 & w46342;
assign w46392 = w46339 & w46340;
assign w46393 = w46337 & w46338;
assign w46394 = w46335 & w46336;
assign w46395 = w46333 & w46334;
assign w46396 = w46331 & w46332;
assign w46397 = w46329 & w46330;
assign w46398 = w46327 & w46328;
assign w46399 = w46325 & w46326;
assign w46400 = w46323 & w46324;
assign w46401 = w46321 & w46322;
assign w46402 = w46319 & w46320;
assign w46403 = w46317 & w46318;
assign w46404 = w46315 & w46316;
assign w46405 = w46313 & w46314;
assign w46406 = w46311 & w46312;
assign w46407 = w46309 & w46310;
assign w46408 = w46307 & w46308;
assign w46409 = w46305 & w46306;
assign w46410 = w46303 & w46304;
assign w46411 = w46301 & w46302;
assign w46412 = w46299 & w46300;
assign w46413 = w46297 & w46298;
assign w46414 = w46295 & w46296;
assign w46415 = w46293 & w46294;
assign w46416 = w46291 & w46292;
assign w46417 = w46289 & w46290;
assign w46418 = w46287 & w46288;
assign w46419 = w46285 & w46286;
assign w46420 = w46283 & w46284;
assign w46421 = w46281 & w46282;
assign w46422 = w46279 & w46280;
assign w46423 = w46277 & w46278;
assign w46424 = w46275 & w46276;
assign w46425 = w46273 & w46274;
assign w46426 = w46271 & w46272;
assign w46427 = w46269 & w46270;
assign w46428 = w46267 & w46268;
assign w46429 = w46265 & w46266;
assign w46430 = w46263 & w46264;
assign w46431 = w46261 & w46262;
assign w46432 = w46259 & w46260;
assign w46433 = w46257 & w46258;
assign w46434 = w46255 & w46256;
assign w46435 = w46253 & w46254;
assign w46436 = w46251 & w46252;
assign w46437 = w46249 & w46250;
assign w46438 = w46247 & w46248;
assign w46439 = w46437 & w46438;
assign w46440 = w46435 & w46436;
assign w46441 = w46433 & w46434;
assign w46442 = w46431 & w46432;
assign w46443 = w46429 & w46430;
assign w46444 = w46427 & w46428;
assign w46445 = w46425 & w46426;
assign w46446 = w46423 & w46424;
assign w46447 = w46421 & w46422;
assign w46448 = w46419 & w46420;
assign w46449 = w46417 & w46418;
assign w46450 = w46415 & w46416;
assign w46451 = w46413 & w46414;
assign w46452 = w46411 & w46412;
assign w46453 = w46409 & w46410;
assign w46454 = w46407 & w46408;
assign w46455 = w46405 & w46406;
assign w46456 = w46403 & w46404;
assign w46457 = w46401 & w46402;
assign w46458 = w46399 & w46400;
assign w46459 = w46397 & w46398;
assign w46460 = w46395 & w46396;
assign w46461 = w46393 & w46394;
assign w46462 = w46391 & w46392;
assign w46463 = w46389 & w46390;
assign w46464 = w46387 & w46388;
assign w46465 = w46385 & w46386;
assign w46466 = w46383 & w46384;
assign w46467 = w46381 & w46382;
assign w46468 = w46379 & w46380;
assign w46469 = w46377 & w46378;
assign w46470 = w46375 & w46376;
assign w46471 = w46469 & w46470;
assign w46472 = w46467 & w46468;
assign w46473 = w46465 & w46466;
assign w46474 = w46463 & w46464;
assign w46475 = w46461 & w46462;
assign w46476 = w46459 & w46460;
assign w46477 = w46457 & w46458;
assign w46478 = w46455 & w46456;
assign w46479 = w46453 & w46454;
assign w46480 = w46451 & w46452;
assign w46481 = w46449 & w46450;
assign w46482 = w46447 & w46448;
assign w46483 = w46445 & w46446;
assign w46484 = w46443 & w46444;
assign w46485 = w46441 & w46442;
assign w46486 = w46439 & w46440;
assign w46487 = w46485 & w46486;
assign w46488 = w46483 & w46484;
assign w46489 = w46481 & w46482;
assign w46490 = w46479 & w46480;
assign w46491 = w46477 & w46478;
assign w46492 = w46475 & w46476;
assign w46493 = w46473 & w46474;
assign w46494 = w46471 & w46472;
assign w46495 = w46493 & w46494;
assign w46496 = w46491 & w46492;
assign w46497 = w46489 & w46490;
assign w46498 = w46487 & w46488;
assign w46499 = w46497 & w46498;
assign w46500 = w46495 & w46496;
assign w46501 = w46499 & w46500;
assign w46502 = ~pi10577 & ~w46501;
assign w46503 = pi02309 & w3514;
assign w46504 = pi08233 & w3542;
assign w46505 = pi07844 & w3270;
assign w46506 = pi03884 & w3338;
assign w46507 = pi04363 & w3484;
assign w46508 = pi06260 & w3414;
assign w46509 = pi06411 & w3392;
assign w46510 = pi08292 & w3342;
assign w46511 = pi07348 & w3376;
assign w46512 = pi05932 & w3344;
assign w46513 = pi08423 & w3510;
assign w46514 = pi04025 & w3071;
assign w46515 = pi04431 & w3258;
assign w46516 = pi08116 & w3446;
assign w46517 = pi06753 & w3186;
assign w46518 = pi07728 & w3476;
assign w46519 = pi01761 & w3288;
assign w46520 = pi05978 & w3252;
assign w46521 = pi06386 & w3298;
assign w46522 = pi04490 & w3396;
assign w46523 = pi04099 & w3522;
assign w46524 = pi06281 & w3540;
assign w46525 = pi03877 & w3209;
assign w46526 = pi03234 & w3544;
assign w46527 = pi07902 & w3352;
assign w46528 = pi06085 & w3550;
assign w46529 = pi01670 & w3360;
assign w46530 = pi03747 & w3490;
assign w46531 = pi04061 & w3574;
assign w46532 = pi04074 & w3428;
assign w46533 = pi02459 & w3478;
assign w46534 = pi04425 & w3302;
assign w46535 = pi03188 & w3346;
assign w46536 = pi07117 & w3410;
assign w46537 = pi03611 & w3424;
assign w46538 = pi03624 & w3137;
assign w46539 = pi07581 & w3201;
assign w46540 = pi02292 & w3616;
assign w46541 = pi07882 & w3382;
assign w46542 = pi08279 & w3229;
assign w46543 = pi04268 & w3468;
assign w46544 = pi03989 & w3132;
assign w46545 = pi06215 & w3586;
assign w46546 = pi07422 & w3566;
assign w46547 = pi03525 & w3400;
assign w46548 = pi03911 & w3348;
assign w46549 = pi06333 & w3538;
assign w46550 = pi04286 & w3334;
assign w46551 = pi08213 & w3282;
assign w46552 = pi04313 & w3214;
assign w46553 = pi06052 & w3452;
assign w46554 = pi03930 & w3456;
assign w46555 = pi08318 & w3324;
assign w46556 = pi03970 & w3498;
assign w46557 = pi08068 & w3175;
assign w46558 = pi08371 & w3160;
assign w46559 = pi01711 & w3192;
assign w46560 = pi04377 & w3564;
assign w46561 = pi08366 & w3368;
assign w46562 = pi05695 & w3232;
assign w46563 = pi05864 & w3598;
assign w46564 = pi04418 & w3169;
assign w46565 = pi04464 & w3556;
assign w46566 = pi08140 & w3440;
assign w46567 = pi04114 & w3181;
assign w46568 = pi05965 & w3612;
assign w46569 = pi09623 & w3464;
assign w46570 = pi04344 & w3115;
assign w46571 = pi03995 & w3394;
assign w46572 = pi08324 & w3332;
assign w46573 = pi04350 & w3190;
assign w46574 = pi08187 & w3106;
assign w46575 = pi03617 & w3296;
assign w46576 = pi07997 & w3516;
assign w46577 = pi04412 & w3562;
assign w46578 = pi03221 & w3336;
assign w46579 = pi03400 & w3404;
assign w46580 = pi07448 & w3434;
assign w46581 = pi08772 & w3600;
assign w46582 = pi04509 & w3488;
assign w46583 = pi07740 & w3458;
assign w46584 = pi09774 & w3442;
assign w46585 = pi04450 & w3504;
assign w46586 = pi04398 & w3512;
assign w46587 = pi07921 & w3596;
assign w46588 = pi06544 & w3304;
assign w46589 = pi08036 & w3532;
assign w46590 = pi04483 & w3588;
assign w46591 = pi02073 & w3250;
assign w46592 = pi08097 & w3606;
assign w46593 = pi04370 & w3146;
assign w46594 = pi06033 & w3554;
assign w46595 = pi01580 & w3112;
assign w46596 = pi08331 & w3158;
assign w46597 = pi04153 & w3502;
assign w46598 = pi07327 & w3620;
assign w46599 = pi02267 & w3240;
assign w46600 = pi06431 & w3203;
assign w46601 = pi01871 & w3139;
assign w46602 = pi05882 & w3604;
assign w46603 = pi06997 & w3406;
assign w46604 = pi07984 & w3426;
assign w46605 = pi03149 & w3614;
assign w46606 = pi07508 & w3312;
assign w46607 = pi08305 & w3294;
assign w46608 = pi07614 & w3374;
assign w46609 = pi04068 & w3494;
assign w46610 = pi03407 & w3330;
assign w46611 = pi02581 & w3506;
assign w46612 = pi07668 & w3194;
assign w46613 = pi08266 & w3402;
assign w46614 = pi08429 & w3242;
assign w46615 = pi04470 & w3388;
assign w46616 = pi06133 & w3480;
assign w46617 = pi07467 & w3508;
assign w46618 = pi03788 & w3350;
assign w46619 = pi05783 & w3143;
assign w46620 = pi03689 & w3310;
assign w46621 = pi02302 & w3234;
assign w46622 = pi05679 & w3486;
assign w46623 = pi05951 & w3492;
assign w46624 = pi04357 & w3328;
assign w46625 = pi06299 & w3482;
assign w46626 = pi09741 & w3356;
assign w46627 = pi06476 & w3199;
assign w46628 = pi07023 & w3340;
assign w46629 = pi08239 & w3280;
assign w46630 = pi07400 & w3448;
assign w46631 = pi04457 & w3184;
assign w46632 = pi07171 & w3364;
assign w46633 = pi07696 & w3430;
assign w46634 = pi01874 & w3462;
assign w46635 = pi08416 & w3408;
assign w46636 = pi03604 & w3536;
assign w46637 = pi06837 & w3518;
assign w46638 = pi02476 & w3278;
assign w46639 = pi07957 & w3093;
assign w46640 = pi08403 & w3150;
assign w46641 = pi06175 & w3378;
assign w46642 = pi04258 & w3326;
assign w46643 = pi06597 & w3153;
assign w46644 = pi08378 & w3524;
assign w46645 = pi08285 & w3560;
assign w46646 = pi02355 & w3264;
assign w46647 = pi06576 & w3496;
assign w46648 = pi01757 & w3436;
assign w46649 = pi03630 & w3262;
assign w46650 = pi03202 & w3520;
assign w46651 = pi07215 & w3205;
assign w46652 = pi04337 & w3086;
assign w46653 = pi07124 & w3420;
assign w46654 = pi08358 & w3438;
assign w46655 = pi02759 & w3290;
assign w46656 = pi07552 & w3165;
assign w46657 = pi07970 & w3238;
assign w46658 = pi03510 & w3534;
assign w46659 = pi02628 & w3300;
assign w46660 = pi04438 & w3122;
assign w46661 = pi03708 & w3244;
assign w46662 = pi08350 & w3179;
assign w46663 = pi02642 & w3474;
assign w46664 = pi03721 & w3548;
assign w46665 = pi04444 & w3162;
assign w46666 = pi06362 & w3450;
assign w46667 = pi04503 & w3582;
assign w46668 = pi03162 & w3306;
assign w46669 = pi02643 & w3584;
assign w46670 = pi03370 & w3362;
assign w46671 = pi08161 & w3594;
assign w46672 = pi07058 & w3286;
assign w46673 = pi02051 & w3322;
assign w46674 = pi01628 & w3390;
assign w46675 = pi09620 & w3118;
assign w46676 = pi06375 & w3236;
assign w46677 = pi07943 & w3125;
assign w46678 = pi08409 & w3558;
assign w46679 = pi04160 & w3454;
assign w46680 = pi06685 & w3082;
assign w46681 = pi03669 & w3610;
assign w46682 = pi08246 & w3096;
assign w46683 = pi06201 & w3460;
assign w46684 = pi08272 & w3580;
assign w46685 = pi03760 & w3526;
assign w46686 = pi08133 & w3570;
assign w46687 = pi07487 & w3167;
assign w46688 = pi07437 & w3276;
assign w46689 = pi07242 & w3225;
assign w46690 = pi07202 & w3156;
assign w46691 = pi03453 & w3530;
assign w46692 = pi08396 & w3110;
assign w46693 = pi04477 & w3177;
assign w46694 = pi06825 & w3256;
assign w46695 = pi05998 & w3219;
assign w46696 = pi08174 & w3173;
assign w46697 = pi03656 & w3260;
assign w46698 = pi09731 & w3129;
assign w46699 = pi08298 & w3148;
assign w46700 = pi08077 & w3223;
assign w46701 = pi07228 & w3254;
assign w46702 = pi08337 & w3602;
assign w46703 = pi07383 & w3358;
assign w46704 = pi04385 & w3370;
assign w46705 = pi08384 & w3418;
assign w46706 = pi08226 & w3546;
assign w46707 = pi02318 & w3398;
assign w46708 = pi04405 & w3412;
assign w46709 = pi03943 & w3592;
assign w46710 = pi02102 & w3127;
assign w46711 = pi08259 & w3188;
assign w46712 = pi03181 & w3380;
assign w46713 = pi03572 & w3103;
assign w46714 = pi05803 & w3308;
assign w46715 = pi07828 & w3207;
assign w46716 = pi01726 & w3078;
assign w46717 = pi04391 & w3618;
assign w46718 = pi06146 & w3217;
assign w46719 = pi07333 & w3272;
assign w46720 = pi07594 & w3372;
assign w46721 = pi02114 & w3266;
assign w46722 = pi06504 & w3422;
assign w46723 = pi03270 & w3268;
assign w46724 = pi07681 & w3590;
assign w46725 = pi03587 & w3274;
assign w46726 = pi07010 & w3572;
assign w46727 = pi08148 & w3608;
assign w46728 = pi07863 & w3386;
assign w46729 = pi05844 & w3248;
assign w46730 = pi08390 & w3246;
assign w46731 = pi03493 & w3064;
assign w46732 = pi08311 & w3316;
assign w46733 = pi03261 & w3500;
assign w46734 = pi03354 & w3470;
assign w46735 = pi09782 & w3366;
assign w46736 = pi07715 & w3171;
assign w46737 = pi06524 & w3227;
assign w46738 = pi03348 & w3416;
assign w46739 = pi07142 & w3135;
assign w46740 = pi03214 & w3197;
assign w46741 = pi06070 & w3528;
assign w46742 = pi03871 & w3576;
assign w46743 = pi08344 & w3578;
assign w46744 = pi06320 & w3314;
assign w46745 = pi08200 & w3320;
assign w46746 = pi02019 & w3466;
assign w46747 = pi08253 & w3318;
assign w46748 = pi06398 & w3354;
assign w46749 = pi01792 & w3284;
assign w46750 = pi06883 & w3384;
assign w46751 = pi07103 & w3552;
assign w46752 = pi04496 & w3211;
assign w46753 = pi01984 & w3472;
assign w46754 = pi02475 & w3444;
assign w46755 = pi03637 & w3292;
assign w46756 = pi06474 & w3432;
assign w46757 = pi07301 & w3221;
assign w46758 = pi01827 & w3568;
assign w46759 = ~w46503 & ~w46504;
assign w46760 = ~w46505 & ~w46506;
assign w46761 = ~w46507 & ~w46508;
assign w46762 = ~w46509 & ~w46510;
assign w46763 = ~w46511 & ~w46512;
assign w46764 = ~w46513 & ~w46514;
assign w46765 = ~w46515 & ~w46516;
assign w46766 = ~w46517 & ~w46518;
assign w46767 = ~w46519 & ~w46520;
assign w46768 = ~w46521 & ~w46522;
assign w46769 = ~w46523 & ~w46524;
assign w46770 = ~w46525 & ~w46526;
assign w46771 = ~w46527 & ~w46528;
assign w46772 = ~w46529 & ~w46530;
assign w46773 = ~w46531 & ~w46532;
assign w46774 = ~w46533 & ~w46534;
assign w46775 = ~w46535 & ~w46536;
assign w46776 = ~w46537 & ~w46538;
assign w46777 = ~w46539 & ~w46540;
assign w46778 = ~w46541 & ~w46542;
assign w46779 = ~w46543 & ~w46544;
assign w46780 = ~w46545 & ~w46546;
assign w46781 = ~w46547 & ~w46548;
assign w46782 = ~w46549 & ~w46550;
assign w46783 = ~w46551 & ~w46552;
assign w46784 = ~w46553 & ~w46554;
assign w46785 = ~w46555 & ~w46556;
assign w46786 = ~w46557 & ~w46558;
assign w46787 = ~w46559 & ~w46560;
assign w46788 = ~w46561 & ~w46562;
assign w46789 = ~w46563 & ~w46564;
assign w46790 = ~w46565 & ~w46566;
assign w46791 = ~w46567 & ~w46568;
assign w46792 = ~w46569 & ~w46570;
assign w46793 = ~w46571 & ~w46572;
assign w46794 = ~w46573 & ~w46574;
assign w46795 = ~w46575 & ~w46576;
assign w46796 = ~w46577 & ~w46578;
assign w46797 = ~w46579 & ~w46580;
assign w46798 = ~w46581 & ~w46582;
assign w46799 = ~w46583 & ~w46584;
assign w46800 = ~w46585 & ~w46586;
assign w46801 = ~w46587 & ~w46588;
assign w46802 = ~w46589 & ~w46590;
assign w46803 = ~w46591 & ~w46592;
assign w46804 = ~w46593 & ~w46594;
assign w46805 = ~w46595 & ~w46596;
assign w46806 = ~w46597 & ~w46598;
assign w46807 = ~w46599 & ~w46600;
assign w46808 = ~w46601 & ~w46602;
assign w46809 = ~w46603 & ~w46604;
assign w46810 = ~w46605 & ~w46606;
assign w46811 = ~w46607 & ~w46608;
assign w46812 = ~w46609 & ~w46610;
assign w46813 = ~w46611 & ~w46612;
assign w46814 = ~w46613 & ~w46614;
assign w46815 = ~w46615 & ~w46616;
assign w46816 = ~w46617 & ~w46618;
assign w46817 = ~w46619 & ~w46620;
assign w46818 = ~w46621 & ~w46622;
assign w46819 = ~w46623 & ~w46624;
assign w46820 = ~w46625 & ~w46626;
assign w46821 = ~w46627 & ~w46628;
assign w46822 = ~w46629 & ~w46630;
assign w46823 = ~w46631 & ~w46632;
assign w46824 = ~w46633 & ~w46634;
assign w46825 = ~w46635 & ~w46636;
assign w46826 = ~w46637 & ~w46638;
assign w46827 = ~w46639 & ~w46640;
assign w46828 = ~w46641 & ~w46642;
assign w46829 = ~w46643 & ~w46644;
assign w46830 = ~w46645 & ~w46646;
assign w46831 = ~w46647 & ~w46648;
assign w46832 = ~w46649 & ~w46650;
assign w46833 = ~w46651 & ~w46652;
assign w46834 = ~w46653 & ~w46654;
assign w46835 = ~w46655 & ~w46656;
assign w46836 = ~w46657 & ~w46658;
assign w46837 = ~w46659 & ~w46660;
assign w46838 = ~w46661 & ~w46662;
assign w46839 = ~w46663 & ~w46664;
assign w46840 = ~w46665 & ~w46666;
assign w46841 = ~w46667 & ~w46668;
assign w46842 = ~w46669 & ~w46670;
assign w46843 = ~w46671 & ~w46672;
assign w46844 = ~w46673 & ~w46674;
assign w46845 = ~w46675 & ~w46676;
assign w46846 = ~w46677 & ~w46678;
assign w46847 = ~w46679 & ~w46680;
assign w46848 = ~w46681 & ~w46682;
assign w46849 = ~w46683 & ~w46684;
assign w46850 = ~w46685 & ~w46686;
assign w46851 = ~w46687 & ~w46688;
assign w46852 = ~w46689 & ~w46690;
assign w46853 = ~w46691 & ~w46692;
assign w46854 = ~w46693 & ~w46694;
assign w46855 = ~w46695 & ~w46696;
assign w46856 = ~w46697 & ~w46698;
assign w46857 = ~w46699 & ~w46700;
assign w46858 = ~w46701 & ~w46702;
assign w46859 = ~w46703 & ~w46704;
assign w46860 = ~w46705 & ~w46706;
assign w46861 = ~w46707 & ~w46708;
assign w46862 = ~w46709 & ~w46710;
assign w46863 = ~w46711 & ~w46712;
assign w46864 = ~w46713 & ~w46714;
assign w46865 = ~w46715 & ~w46716;
assign w46866 = ~w46717 & ~w46718;
assign w46867 = ~w46719 & ~w46720;
assign w46868 = ~w46721 & ~w46722;
assign w46869 = ~w46723 & ~w46724;
assign w46870 = ~w46725 & ~w46726;
assign w46871 = ~w46727 & ~w46728;
assign w46872 = ~w46729 & ~w46730;
assign w46873 = ~w46731 & ~w46732;
assign w46874 = ~w46733 & ~w46734;
assign w46875 = ~w46735 & ~w46736;
assign w46876 = ~w46737 & ~w46738;
assign w46877 = ~w46739 & ~w46740;
assign w46878 = ~w46741 & ~w46742;
assign w46879 = ~w46743 & ~w46744;
assign w46880 = ~w46745 & ~w46746;
assign w46881 = ~w46747 & ~w46748;
assign w46882 = ~w46749 & ~w46750;
assign w46883 = ~w46751 & ~w46752;
assign w46884 = ~w46753 & ~w46754;
assign w46885 = ~w46755 & ~w46756;
assign w46886 = ~w46757 & ~w46758;
assign w46887 = w46885 & w46886;
assign w46888 = w46883 & w46884;
assign w46889 = w46881 & w46882;
assign w46890 = w46879 & w46880;
assign w46891 = w46877 & w46878;
assign w46892 = w46875 & w46876;
assign w46893 = w46873 & w46874;
assign w46894 = w46871 & w46872;
assign w46895 = w46869 & w46870;
assign w46896 = w46867 & w46868;
assign w46897 = w46865 & w46866;
assign w46898 = w46863 & w46864;
assign w46899 = w46861 & w46862;
assign w46900 = w46859 & w46860;
assign w46901 = w46857 & w46858;
assign w46902 = w46855 & w46856;
assign w46903 = w46853 & w46854;
assign w46904 = w46851 & w46852;
assign w46905 = w46849 & w46850;
assign w46906 = w46847 & w46848;
assign w46907 = w46845 & w46846;
assign w46908 = w46843 & w46844;
assign w46909 = w46841 & w46842;
assign w46910 = w46839 & w46840;
assign w46911 = w46837 & w46838;
assign w46912 = w46835 & w46836;
assign w46913 = w46833 & w46834;
assign w46914 = w46831 & w46832;
assign w46915 = w46829 & w46830;
assign w46916 = w46827 & w46828;
assign w46917 = w46825 & w46826;
assign w46918 = w46823 & w46824;
assign w46919 = w46821 & w46822;
assign w46920 = w46819 & w46820;
assign w46921 = w46817 & w46818;
assign w46922 = w46815 & w46816;
assign w46923 = w46813 & w46814;
assign w46924 = w46811 & w46812;
assign w46925 = w46809 & w46810;
assign w46926 = w46807 & w46808;
assign w46927 = w46805 & w46806;
assign w46928 = w46803 & w46804;
assign w46929 = w46801 & w46802;
assign w46930 = w46799 & w46800;
assign w46931 = w46797 & w46798;
assign w46932 = w46795 & w46796;
assign w46933 = w46793 & w46794;
assign w46934 = w46791 & w46792;
assign w46935 = w46789 & w46790;
assign w46936 = w46787 & w46788;
assign w46937 = w46785 & w46786;
assign w46938 = w46783 & w46784;
assign w46939 = w46781 & w46782;
assign w46940 = w46779 & w46780;
assign w46941 = w46777 & w46778;
assign w46942 = w46775 & w46776;
assign w46943 = w46773 & w46774;
assign w46944 = w46771 & w46772;
assign w46945 = w46769 & w46770;
assign w46946 = w46767 & w46768;
assign w46947 = w46765 & w46766;
assign w46948 = w46763 & w46764;
assign w46949 = w46761 & w46762;
assign w46950 = w46759 & w46760;
assign w46951 = w46949 & w46950;
assign w46952 = w46947 & w46948;
assign w46953 = w46945 & w46946;
assign w46954 = w46943 & w46944;
assign w46955 = w46941 & w46942;
assign w46956 = w46939 & w46940;
assign w46957 = w46937 & w46938;
assign w46958 = w46935 & w46936;
assign w46959 = w46933 & w46934;
assign w46960 = w46931 & w46932;
assign w46961 = w46929 & w46930;
assign w46962 = w46927 & w46928;
assign w46963 = w46925 & w46926;
assign w46964 = w46923 & w46924;
assign w46965 = w46921 & w46922;
assign w46966 = w46919 & w46920;
assign w46967 = w46917 & w46918;
assign w46968 = w46915 & w46916;
assign w46969 = w46913 & w46914;
assign w46970 = w46911 & w46912;
assign w46971 = w46909 & w46910;
assign w46972 = w46907 & w46908;
assign w46973 = w46905 & w46906;
assign w46974 = w46903 & w46904;
assign w46975 = w46901 & w46902;
assign w46976 = w46899 & w46900;
assign w46977 = w46897 & w46898;
assign w46978 = w46895 & w46896;
assign w46979 = w46893 & w46894;
assign w46980 = w46891 & w46892;
assign w46981 = w46889 & w46890;
assign w46982 = w46887 & w46888;
assign w46983 = w46981 & w46982;
assign w46984 = w46979 & w46980;
assign w46985 = w46977 & w46978;
assign w46986 = w46975 & w46976;
assign w46987 = w46973 & w46974;
assign w46988 = w46971 & w46972;
assign w46989 = w46969 & w46970;
assign w46990 = w46967 & w46968;
assign w46991 = w46965 & w46966;
assign w46992 = w46963 & w46964;
assign w46993 = w46961 & w46962;
assign w46994 = w46959 & w46960;
assign w46995 = w46957 & w46958;
assign w46996 = w46955 & w46956;
assign w46997 = w46953 & w46954;
assign w46998 = w46951 & w46952;
assign w46999 = w46997 & w46998;
assign w47000 = w46995 & w46996;
assign w47001 = w46993 & w46994;
assign w47002 = w46991 & w46992;
assign w47003 = w46989 & w46990;
assign w47004 = w46987 & w46988;
assign w47005 = w46985 & w46986;
assign w47006 = w46983 & w46984;
assign w47007 = w47005 & w47006;
assign w47008 = w47003 & w47004;
assign w47009 = w47001 & w47002;
assign w47010 = w46999 & w47000;
assign w47011 = w47009 & w47010;
assign w47012 = w47007 & w47008;
assign w47013 = w47011 & w47012;
assign w47014 = ~pi10577 & ~w47013;
assign w47015 = pi04049 & w3502;
assign w47016 = pi09604 & w3454;
assign w47017 = pi02006 & w3470;
assign w47018 = pi07041 & w3300;
assign w47019 = pi07720 & w3584;
assign w47020 = pi06728 & w3482;
assign w47021 = pi07628 & w3606;
assign w47022 = pi06925 & w3514;
assign w47023 = pi07025 & w3432;
assign w47024 = pi06860 & w3462;
assign w47025 = pi06806 & w3203;
assign w47026 = pi06686 & w3356;
assign w47027 = pi07299 & w3434;
assign w47028 = pi01878 & w3604;
assign w47029 = pi06669 & w3112;
assign w47030 = pi06951 & w3284;
assign w47031 = pi01681 & w3252;
assign w47032 = pi02772 & w3370;
assign w47033 = pi06622 & w3452;
assign w47034 = pi07608 & w3175;
assign w47035 = pi01976 & w3250;
assign w47036 = pi06812 & w3129;
assign w47037 = pi03644 & w3416;
assign w47038 = pi06740 & w3314;
assign w47039 = pi07561 & w3426;
assign w47040 = pi04232 & w3122;
assign w47041 = pi07080 & w3139;
assign w47042 = pi03800 & w3137;
assign w47043 = pi01947 & w3103;
assign w47044 = pi03540 & w3346;
assign w47045 = pi01958 & w3248;
assign w47046 = pi01787 & w3262;
assign w47047 = pi06747 & w3538;
assign w47048 = pi08064 & w3246;
assign w47049 = pi06998 & w3442;
assign w47050 = pi06977 & w3256;
assign w47051 = pi07150 & w3420;
assign w47052 = pi06871 & w3496;
assign w47053 = pi07308 & w3508;
assign w47054 = pi03735 & w3400;
assign w47055 = pi07872 & w3580;
assign w47056 = pi04298 & w3588;
assign w47057 = pi06498 & w3266;
assign w47058 = pi07276 & w3448;
assign w47059 = pi03569 & w3336;
assign w47060 = pi03976 & w3071;
assign w47061 = pi07663 & w3608;
assign w47062 = pi06851 & w3304;
assign w47063 = pi02667 & w3412;
assign w47064 = pi08043 & w3524;
assign w47065 = pi06591 & w3612;
assign w47066 = pi09725 & w3592;
assign w47067 = pi01762 & w3310;
assign w47068 = pi07977 & w3602;
assign w47069 = pi09033 & w3207;
assign w47070 = pi08055 & w3418;
assign w47071 = pi02497 & w3232;
assign w47072 = pi06615 & w3554;
assign w47073 = pi07829 & w3096;
assign w47074 = pi09545 & w3214;
assign w47075 = pi07643 & w3570;
assign w47076 = pi07576 & w3474;
assign w47077 = pi07212 & w3472;
assign w47078 = pi04272 & w3556;
assign w47079 = pi03826 & w3610;
assign w47080 = pi09562 & w3334;
assign w47081 = pi07516 & w3382;
assign w47082 = pi02290 & w3590;
assign w47083 = pi03553 & w3520;
assign w47084 = pi07586 & w3532;
assign w47085 = pi07920 & w3294;
assign w47086 = pi04306 & w3396;
assign w47087 = pi07177 & w3156;
assign w47088 = pi07184 & w3205;
assign w47089 = pi07290 & w3276;
assign w47090 = pi01500 & w3422;
assign w47091 = pi04141 & w3328;
assign w47092 = pi03865 & w3350;
assign w47093 = pi03927 & w3456;
assign w47094 = pi01902 & w3450;
assign w47095 = pi06877 & w3153;
assign w47096 = pi06899 & w3082;
assign w47097 = pi02293 & w3308;
assign w47098 = pi03905 & w3338;
assign w47099 = pi06959 & w3078;
assign w47100 = pi03579 & w3544;
assign w47101 = pi09715 & w3498;
assign w47102 = pi02431 & w3560;
assign w47103 = pi07352 & w3201;
assign w47104 = pi02774 & w3564;
assign w47105 = pi07102 & w3340;
assign w47106 = pi09701 & w3394;
assign w47107 = pi07691 & w3594;
assign w47108 = pi07787 & w3546;
assign w47109 = pi06663 & w3217;
assign w47110 = pi06609 & w3219;
assign w47111 = pi07282 & w3566;
assign w47112 = pi03839 & w3244;
assign w47113 = pi07477 & w3464;
assign w47114 = pi01712 & w3171;
assign w47115 = pi06492 & w3240;
assign w47116 = pi07086 & w3406;
assign w47117 = pi04291 & w3177;
assign w47118 = pi03590 & w3500;
assign w47119 = pi03683 & w3330;
assign w47120 = pi08100 & w3558;
assign w47121 = pi01741 & w3476;
assign w47122 = pi01935 & w3274;
assign w47123 = pi07760 & w3478;
assign w47124 = pi06582 & w3492;
assign w47125 = pi07766 & w3282;
assign w47126 = pi06677 & w3378;
assign w47127 = pi07753 & w3320;
assign w47128 = pi04206 & w3562;
assign w47129 = pi02780 & w3484;
assign w47130 = pi06783 & w3354;
assign w47131 = pi01802 & w3260;
assign w47132 = pi04193 & w3512;
assign w47133 = pi07862 & w3402;
assign w47134 = pi04167 & w3146;
assign w47135 = pi02062 & w3306;
assign w47136 = pi03696 & w3530;
assign w47137 = pi07506 & w3386;
assign w47138 = pi07164 & w3364;
assign w47139 = pi01896 & w3598;
assign w47140 = pi04040 & w3181;
assign w47141 = pi02055 & w3380;
assign w47142 = pi07803 & w3542;
assign w47143 = pi01737 & w3526;
assign w47144 = pi07620 & w3223;
assign w47145 = pi08118 & w3510;
assign w47146 = pi07067 & w3466;
assign w47147 = pi07672 & w3366;
assign w47148 = pi01999 & w3362;
assign w47149 = pi06767 & w3236;
assign w47150 = pi06531 & w3436;
assign w47151 = pi04331 & w3488;
assign w47152 = pi08080 & w3110;
assign w47153 = pi09642 & w3428;
assign w47154 = pi07360 & w3372;
assign w47155 = pi06511 & w3143;
assign w47156 = pi06714 & w3414;
assign w47157 = pi07337 & w3165;
assign w47158 = pi03852 & w3490;
assign w47159 = pi01965 & w3534;
assign w47160 = pi06819 & w3199;
assign w47161 = pi07777 & w3264;
assign w47162 = pi06642 & w3568;
assign w47163 = pi06773 & w3298;
assign w47164 = pi02762 & w3258;
assign w47165 = pi02756 & w3504;
assign w47166 = pi07158 & w3135;
assign w47167 = pi01996 & w3404;
assign w47168 = pi04316 & w3211;
assign w47169 = pi03715 & w3064;
assign w47170 = pi07315 & w3167;
assign w47171 = pi07950 & w3332;
assign w47172 = pi08131 & w3242;
assign w47173 = pi06721 & w3540;
assign w47174 = pi07190 & w3254;
assign w47175 = pi04280 & w3388;
assign w47176 = pi08090 & w3150;
assign w47177 = pi06628 & w3528;
assign w47178 = pi07653 & w3440;
assign w47179 = pi07267 & w3358;
assign w47180 = pi06655 & w3480;
assign w47181 = pi07839 & w3318;
assign w47182 = pi03957 & w3132;
assign w47183 = pi07132 & w3552;
assign w47184 = pi03983 & w3118;
assign w47185 = pi07199 & w3225;
assign w47186 = pi09533 & w3460;
assign w47187 = pi07094 & w3572;
assign w47188 = pi07458 & w3360;
assign w47189 = pi02486 & w3600;
assign w47190 = pi06938 & w3186;
assign w47191 = pi06985 & w3518;
assign w47192 = pi07710 & w3173;
assign w47193 = pi08016 & w3438;
assign w47194 = pi08007 & w3179;
assign w47195 = pi03774 & w3536;
assign w47196 = pi07964 & w3158;
assign w47197 = pi03813 & w3292;
assign w47198 = pi04128 & w3115;
assign w47199 = pi07141 & w3410;
assign w47200 = pi06475 & w3486;
assign w47201 = pi02783 & w3190;
assign w47202 = pi01753 & w3548;
assign w47203 = pi07542 & w3093;
assign w47204 = pi03783 & w3424;
assign w47205 = pi02063 & w3614;
assign w47206 = pi07881 & w3229;
assign w47207 = pi02382 & w3238;
assign w47208 = pi07403 & w3430;
assign w47209 = pi07989 & w3578;
assign w47210 = pi06570 & w3344;
assign w47211 = pi04088 & w3326;
assign w47212 = pi07733 & w3106;
assign w47213 = pi07012 & w3384;
assign w47214 = pi02410 & w3620;
assign w47215 = pi07073 & w3127;
assign w47216 = pi07634 & w3446;
assign w47217 = pi03891 & w3576;
assign w47218 = pi07901 & w3342;
assign w47219 = pi07115 & w3286;
assign w47220 = pi07034 & w3506;
assign w47221 = pi07322 & w3312;
assign w47222 = pi06649 & w3288;
assign w47223 = pi04325 & w3582;
assign w47224 = pi07568 & w3516;
assign w47225 = pi02043 & w3197;
assign w47226 = pi06636 & w3550;
assign w47227 = pi04219 & w3302;
assign w47228 = pi07853 & w3188;
assign w47229 = pi06702 & w3586;
assign w47230 = pi07536 & w3125;
assign w47231 = pi06912 & w3278;
assign w47232 = pi04009 & w3494;
assign w47233 = pi07247 & w3272;
assign w47234 = pi03918 & w3348;
assign w47235 = pi04264 & w3184;
assign w47236 = pi07930 & w3316;
assign w47237 = pi07910 & w3148;
assign w47238 = pi07367 & w3374;
assign w47239 = pi02770 & w3618;
assign w47240 = pi06263 & w3086;
assign w47241 = pi07047 & w3398;
assign w47242 = pi07529 & w3596;
assign w47243 = pi07813 & w3280;
assign w47244 = pi01953 & w3322;
assign w47245 = pi04028 & w3522;
assign w47246 = pi07255 & w3376;
assign w47247 = pi03792 & w3296;
assign w47248 = pi02515 & w3368;
assign w47249 = pi08032 & w3160;
assign w47250 = pi07523 & w3352;
assign w47251 = pi01522 & w3209;
assign w47252 = pi01663 & w3192;
assign w47253 = pi07599 & w3616;
assign w47254 = pi02435 & w3194;
assign w47255 = pi03600 & w3268;
assign w47256 = pi07942 & w3324;
assign w47257 = pi04244 & w3162;
assign w47258 = pi08110 & w3408;
assign w47259 = pi07468 & w3390;
assign w47260 = pi06845 & w3227;
assign w47261 = pi02338 & w3444;
assign w47262 = pi02765 & w3169;
assign w47263 = pi06796 & w3392;
assign w47264 = pi07057 & w3234;
assign w47265 = pi09581 & w3290;
assign w47266 = pi07432 & w3458;
assign w47267 = pi07225 & w3221;
assign w47268 = pi09651 & w3574;
assign w47269 = pi07700 & w3468;
assign w47270 = pi07497 & w3270;
assign w47271 = ~w47015 & ~w47016;
assign w47272 = ~w47017 & ~w47018;
assign w47273 = ~w47019 & ~w47020;
assign w47274 = ~w47021 & ~w47022;
assign w47275 = ~w47023 & ~w47024;
assign w47276 = ~w47025 & ~w47026;
assign w47277 = ~w47027 & ~w47028;
assign w47278 = ~w47029 & ~w47030;
assign w47279 = ~w47031 & ~w47032;
assign w47280 = ~w47033 & ~w47034;
assign w47281 = ~w47035 & ~w47036;
assign w47282 = ~w47037 & ~w47038;
assign w47283 = ~w47039 & ~w47040;
assign w47284 = ~w47041 & ~w47042;
assign w47285 = ~w47043 & ~w47044;
assign w47286 = ~w47045 & ~w47046;
assign w47287 = ~w47047 & ~w47048;
assign w47288 = ~w47049 & ~w47050;
assign w47289 = ~w47051 & ~w47052;
assign w47290 = ~w47053 & ~w47054;
assign w47291 = ~w47055 & ~w47056;
assign w47292 = ~w47057 & ~w47058;
assign w47293 = ~w47059 & ~w47060;
assign w47294 = ~w47061 & ~w47062;
assign w47295 = ~w47063 & ~w47064;
assign w47296 = ~w47065 & ~w47066;
assign w47297 = ~w47067 & ~w47068;
assign w47298 = ~w47069 & ~w47070;
assign w47299 = ~w47071 & ~w47072;
assign w47300 = ~w47073 & ~w47074;
assign w47301 = ~w47075 & ~w47076;
assign w47302 = ~w47077 & ~w47078;
assign w47303 = ~w47079 & ~w47080;
assign w47304 = ~w47081 & ~w47082;
assign w47305 = ~w47083 & ~w47084;
assign w47306 = ~w47085 & ~w47086;
assign w47307 = ~w47087 & ~w47088;
assign w47308 = ~w47089 & ~w47090;
assign w47309 = ~w47091 & ~w47092;
assign w47310 = ~w47093 & ~w47094;
assign w47311 = ~w47095 & ~w47096;
assign w47312 = ~w47097 & ~w47098;
assign w47313 = ~w47099 & ~w47100;
assign w47314 = ~w47101 & ~w47102;
assign w47315 = ~w47103 & ~w47104;
assign w47316 = ~w47105 & ~w47106;
assign w47317 = ~w47107 & ~w47108;
assign w47318 = ~w47109 & ~w47110;
assign w47319 = ~w47111 & ~w47112;
assign w47320 = ~w47113 & ~w47114;
assign w47321 = ~w47115 & ~w47116;
assign w47322 = ~w47117 & ~w47118;
assign w47323 = ~w47119 & ~w47120;
assign w47324 = ~w47121 & ~w47122;
assign w47325 = ~w47123 & ~w47124;
assign w47326 = ~w47125 & ~w47126;
assign w47327 = ~w47127 & ~w47128;
assign w47328 = ~w47129 & ~w47130;
assign w47329 = ~w47131 & ~w47132;
assign w47330 = ~w47133 & ~w47134;
assign w47331 = ~w47135 & ~w47136;
assign w47332 = ~w47137 & ~w47138;
assign w47333 = ~w47139 & ~w47140;
assign w47334 = ~w47141 & ~w47142;
assign w47335 = ~w47143 & ~w47144;
assign w47336 = ~w47145 & ~w47146;
assign w47337 = ~w47147 & ~w47148;
assign w47338 = ~w47149 & ~w47150;
assign w47339 = ~w47151 & ~w47152;
assign w47340 = ~w47153 & ~w47154;
assign w47341 = ~w47155 & ~w47156;
assign w47342 = ~w47157 & ~w47158;
assign w47343 = ~w47159 & ~w47160;
assign w47344 = ~w47161 & ~w47162;
assign w47345 = ~w47163 & ~w47164;
assign w47346 = ~w47165 & ~w47166;
assign w47347 = ~w47167 & ~w47168;
assign w47348 = ~w47169 & ~w47170;
assign w47349 = ~w47171 & ~w47172;
assign w47350 = ~w47173 & ~w47174;
assign w47351 = ~w47175 & ~w47176;
assign w47352 = ~w47177 & ~w47178;
assign w47353 = ~w47179 & ~w47180;
assign w47354 = ~w47181 & ~w47182;
assign w47355 = ~w47183 & ~w47184;
assign w47356 = ~w47185 & ~w47186;
assign w47357 = ~w47187 & ~w47188;
assign w47358 = ~w47189 & ~w47190;
assign w47359 = ~w47191 & ~w47192;
assign w47360 = ~w47193 & ~w47194;
assign w47361 = ~w47195 & ~w47196;
assign w47362 = ~w47197 & ~w47198;
assign w47363 = ~w47199 & ~w47200;
assign w47364 = ~w47201 & ~w47202;
assign w47365 = ~w47203 & ~w47204;
assign w47366 = ~w47205 & ~w47206;
assign w47367 = ~w47207 & ~w47208;
assign w47368 = ~w47209 & ~w47210;
assign w47369 = ~w47211 & ~w47212;
assign w47370 = ~w47213 & ~w47214;
assign w47371 = ~w47215 & ~w47216;
assign w47372 = ~w47217 & ~w47218;
assign w47373 = ~w47219 & ~w47220;
assign w47374 = ~w47221 & ~w47222;
assign w47375 = ~w47223 & ~w47224;
assign w47376 = ~w47225 & ~w47226;
assign w47377 = ~w47227 & ~w47228;
assign w47378 = ~w47229 & ~w47230;
assign w47379 = ~w47231 & ~w47232;
assign w47380 = ~w47233 & ~w47234;
assign w47381 = ~w47235 & ~w47236;
assign w47382 = ~w47237 & ~w47238;
assign w47383 = ~w47239 & ~w47240;
assign w47384 = ~w47241 & ~w47242;
assign w47385 = ~w47243 & ~w47244;
assign w47386 = ~w47245 & ~w47246;
assign w47387 = ~w47247 & ~w47248;
assign w47388 = ~w47249 & ~w47250;
assign w47389 = ~w47251 & ~w47252;
assign w47390 = ~w47253 & ~w47254;
assign w47391 = ~w47255 & ~w47256;
assign w47392 = ~w47257 & ~w47258;
assign w47393 = ~w47259 & ~w47260;
assign w47394 = ~w47261 & ~w47262;
assign w47395 = ~w47263 & ~w47264;
assign w47396 = ~w47265 & ~w47266;
assign w47397 = ~w47267 & ~w47268;
assign w47398 = ~w47269 & ~w47270;
assign w47399 = w47397 & w47398;
assign w47400 = w47395 & w47396;
assign w47401 = w47393 & w47394;
assign w47402 = w47391 & w47392;
assign w47403 = w47389 & w47390;
assign w47404 = w47387 & w47388;
assign w47405 = w47385 & w47386;
assign w47406 = w47383 & w47384;
assign w47407 = w47381 & w47382;
assign w47408 = w47379 & w47380;
assign w47409 = w47377 & w47378;
assign w47410 = w47375 & w47376;
assign w47411 = w47373 & w47374;
assign w47412 = w47371 & w47372;
assign w47413 = w47369 & w47370;
assign w47414 = w47367 & w47368;
assign w47415 = w47365 & w47366;
assign w47416 = w47363 & w47364;
assign w47417 = w47361 & w47362;
assign w47418 = w47359 & w47360;
assign w47419 = w47357 & w47358;
assign w47420 = w47355 & w47356;
assign w47421 = w47353 & w47354;
assign w47422 = w47351 & w47352;
assign w47423 = w47349 & w47350;
assign w47424 = w47347 & w47348;
assign w47425 = w47345 & w47346;
assign w47426 = w47343 & w47344;
assign w47427 = w47341 & w47342;
assign w47428 = w47339 & w47340;
assign w47429 = w47337 & w47338;
assign w47430 = w47335 & w47336;
assign w47431 = w47333 & w47334;
assign w47432 = w47331 & w47332;
assign w47433 = w47329 & w47330;
assign w47434 = w47327 & w47328;
assign w47435 = w47325 & w47326;
assign w47436 = w47323 & w47324;
assign w47437 = w47321 & w47322;
assign w47438 = w47319 & w47320;
assign w47439 = w47317 & w47318;
assign w47440 = w47315 & w47316;
assign w47441 = w47313 & w47314;
assign w47442 = w47311 & w47312;
assign w47443 = w47309 & w47310;
assign w47444 = w47307 & w47308;
assign w47445 = w47305 & w47306;
assign w47446 = w47303 & w47304;
assign w47447 = w47301 & w47302;
assign w47448 = w47299 & w47300;
assign w47449 = w47297 & w47298;
assign w47450 = w47295 & w47296;
assign w47451 = w47293 & w47294;
assign w47452 = w47291 & w47292;
assign w47453 = w47289 & w47290;
assign w47454 = w47287 & w47288;
assign w47455 = w47285 & w47286;
assign w47456 = w47283 & w47284;
assign w47457 = w47281 & w47282;
assign w47458 = w47279 & w47280;
assign w47459 = w47277 & w47278;
assign w47460 = w47275 & w47276;
assign w47461 = w47273 & w47274;
assign w47462 = w47271 & w47272;
assign w47463 = w47461 & w47462;
assign w47464 = w47459 & w47460;
assign w47465 = w47457 & w47458;
assign w47466 = w47455 & w47456;
assign w47467 = w47453 & w47454;
assign w47468 = w47451 & w47452;
assign w47469 = w47449 & w47450;
assign w47470 = w47447 & w47448;
assign w47471 = w47445 & w47446;
assign w47472 = w47443 & w47444;
assign w47473 = w47441 & w47442;
assign w47474 = w47439 & w47440;
assign w47475 = w47437 & w47438;
assign w47476 = w47435 & w47436;
assign w47477 = w47433 & w47434;
assign w47478 = w47431 & w47432;
assign w47479 = w47429 & w47430;
assign w47480 = w47427 & w47428;
assign w47481 = w47425 & w47426;
assign w47482 = w47423 & w47424;
assign w47483 = w47421 & w47422;
assign w47484 = w47419 & w47420;
assign w47485 = w47417 & w47418;
assign w47486 = w47415 & w47416;
assign w47487 = w47413 & w47414;
assign w47488 = w47411 & w47412;
assign w47489 = w47409 & w47410;
assign w47490 = w47407 & w47408;
assign w47491 = w47405 & w47406;
assign w47492 = w47403 & w47404;
assign w47493 = w47401 & w47402;
assign w47494 = w47399 & w47400;
assign w47495 = w47493 & w47494;
assign w47496 = w47491 & w47492;
assign w47497 = w47489 & w47490;
assign w47498 = w47487 & w47488;
assign w47499 = w47485 & w47486;
assign w47500 = w47483 & w47484;
assign w47501 = w47481 & w47482;
assign w47502 = w47479 & w47480;
assign w47503 = w47477 & w47478;
assign w47504 = w47475 & w47476;
assign w47505 = w47473 & w47474;
assign w47506 = w47471 & w47472;
assign w47507 = w47469 & w47470;
assign w47508 = w47467 & w47468;
assign w47509 = w47465 & w47466;
assign w47510 = w47463 & w47464;
assign w47511 = w47509 & w47510;
assign w47512 = w47507 & w47508;
assign w47513 = w47505 & w47506;
assign w47514 = w47503 & w47504;
assign w47515 = w47501 & w47502;
assign w47516 = w47499 & w47500;
assign w47517 = w47497 & w47498;
assign w47518 = w47495 & w47496;
assign w47519 = w47517 & w47518;
assign w47520 = w47515 & w47516;
assign w47521 = w47513 & w47514;
assign w47522 = w47511 & w47512;
assign w47523 = w47521 & w47522;
assign w47524 = w47519 & w47520;
assign w47525 = w47523 & w47524;
assign w47526 = ~pi10577 & ~w47525;
assign w47527 = pi03495 & w3064;
assign w47528 = pi03210 & w3520;
assign w47529 = pi02533 & w3590;
assign w47530 = pi01869 & w3528;
assign w47531 = pi05968 & w3612;
assign w47532 = pi01599 & w3148;
assign w47533 = pi03190 & w3346;
assign w47534 = pi02144 & w3558;
assign w47535 = pi08151 & w3608;
assign w47536 = pi08142 & w3440;
assign w47537 = pi05697 & w3232;
assign w47538 = pi07271 & w3472;
assign w47539 = pi06289 & w3540;
assign w47540 = pi06152 & w3217;
assign w47541 = pi03620 & w3296;
assign w47542 = pi08102 & w3606;
assign w47543 = pi01722 & w3402;
assign w47544 = pi06437 & w3203;
assign w47545 = pi02308 & w3234;
assign w47546 = pi08183 & w3584;
assign w47547 = pi06801 & w3078;
assign w47548 = pi06204 & w3460;
assign w47549 = pi06990 & w3139;
assign w47550 = pi02276 & w3510;
assign w47551 = pi03593 & w3274;
assign w47552 = pi01904 & w3554;
assign w47553 = pi05831 & w3436;
assign w47554 = pi06760 & w3186;
assign w47555 = pi02456 & w3246;
assign w47556 = pi05788 & w3143;
assign w47557 = pi04353 & w3190;
assign w47558 = pi09529 & w3158;
assign w47559 = pi01545 & w3324;
assign w47560 = pi02278 & w3408;
assign w47561 = pi07976 & w3238;
assign w47562 = pi09730 & w3082;
assign w47563 = pi07587 & w3201;
assign w47564 = pi04439 & w3122;
assign w47565 = pi07929 & w3596;
assign w47566 = pi07389 & w3358;
assign w47567 = pi04460 & w3184;
assign w47568 = pi03155 & w3614;
assign w47569 = pi01744 & w3410;
assign w47570 = pi08085 & w3223;
assign w47571 = pi06886 & w3384;
assign w47572 = pi08203 & w3320;
assign w47573 = pi04366 & w3484;
assign w47574 = pi07343 & w3272;
assign w47575 = pi03724 & w3548;
assign w47576 = pi04070 & w3494;
assign w47577 = pi07948 & w3125;
assign w47578 = pi06530 & w3227;
assign w47579 = pi03376 & w3362;
assign w47580 = pi08071 & w3175;
assign w47581 = pi04387 & w3370;
assign w47582 = pi07252 & w3225;
assign w47583 = pi06008 & w3219;
assign w47584 = pi04466 & w3556;
assign w47585 = pi02275 & w3542;
assign w47586 = pi08177 & w3173;
assign w47587 = pi07963 & w3093;
assign w47588 = pi01818 & w3188;
assign w47589 = pi04492 & w3396;
assign w47590 = pi04414 & w3562;
assign w47591 = pi03998 & w3394;
assign w47592 = pi08209 & w3478;
assign w47593 = pi02630 & w3506;
assign w47594 = pi04117 & w3181;
assign w47595 = pi02023 & w3448;
assign w47596 = pi08196 & w3444;
assign w47597 = pi03402 & w3404;
assign w47598 = pi06971 & w3127;
assign w47599 = pi07676 & w3194;
assign w47600 = pi07357 & w3376;
assign w47601 = pi07909 & w3352;
assign w47602 = pi05986 & w3252;
assign w47603 = pi06840 & w3518;
assign w47604 = pi06270 & w3414;
assign w47605 = pi02605 & w3332;
assign w47606 = pi06716 & w3278;
assign w47607 = pi07736 & w3476;
assign w47608 = pi03991 & w3132;
assign w47609 = pi07495 & w3167;
assign w47610 = pi03552 & w3322;
assign w47611 = pi07430 & w3566;
assign w47612 = pi03626 & w3137;
assign w47613 = pi04408 & w3412;
assign w47614 = pi07439 & w3276;
assign w47615 = pi03350 & w3416;
assign w47616 = pi03933 & w3456;
assign w47617 = pi06120 & w3288;
assign w47618 = pi05744 & w3266;
assign w47619 = pi04265 & w3326;
assign w47620 = pi03633 & w3262;
assign w47621 = pi04318 & w3214;
assign w47622 = pi06964 & w3466;
assign w47623 = pi04346 & w3115;
assign w47624 = pi03873 & w3576;
assign w47625 = pi03357 & w3470;
assign w47626 = pi07032 & w3340;
assign w47627 = pi04447 & w3162;
assign w47628 = pi03278 & w3268;
assign w47629 = pi01683 & w3153;
assign w47630 = pi03264 & w3500;
assign w47631 = pi04340 & w3086;
assign w47632 = pi06178 & w3378;
assign w47633 = pi01769 & w3308;
assign w47634 = pi01970 & w3244;
assign w47635 = pi04434 & w3258;
assign w47636 = pi07655 & w3600;
assign w47637 = pi06381 & w3236;
assign w47638 = pi03607 & w3536;
assign w47639 = pi03946 & w3592;
assign w47640 = pi03977 & w3498;
assign w47641 = pi02437 & w3382;
assign w47642 = pi04473 & w3388;
assign w47643 = pi03613 & w3424;
assign w47644 = pi02591 & w3578;
assign w47645 = pi02650 & w3205;
assign w47646 = pi01876 & w3452;
assign w47647 = pi07810 & w3390;
assign w47648 = pi03164 & w3306;
assign w47649 = pi04156 & w3502;
assign w47650 = pi04453 & w3504;
assign w47651 = pi04032 & w3602;
assign w47652 = pi02622 & w3179;
assign w47653 = pi06401 & w3354;
assign w47654 = pi07456 & w3434;
assign w47655 = pi01623 & w3560;
assign w47656 = pi06788 & w3284;
assign w47657 = pi03528 & w3400;
assign w47658 = pi04379 & w3564;
assign w47659 = pi03750 & w3490;
assign w47660 = pi07621 & w3374;
assign w47661 = pi04064 & w3574;
assign w47662 = pi08222 & w3264;
assign w47663 = pi02285 & w3552;
assign w47664 = pi03880 & w3209;
assign w47665 = pi08015 & w3474;
assign w47666 = pi04030 & w3071;
assign w47667 = pi01691 & w3229;
assign w47668 = pi04479 & w3177;
assign w47669 = pi07515 & w3312;
assign w47670 = pi08038 & w3532;
assign w47671 = pi06827 & w3256;
assign w47672 = pi02599 & w3438;
assign w47673 = pi04359 & w3328;
assign w47674 = pi05892 & w3604;
assign w47675 = pi05870 & w3598;
assign w47676 = pi03519 & w3534;
assign w47677 = pi07302 & w3221;
assign w47678 = pi03240 & w3544;
assign w47679 = pi08057 & w3616;
assign w47680 = pi01517 & w3316;
assign w47681 = pi06323 & w3314;
assign w47682 = pi06507 & w3422;
assign w47683 = pi04421 & w3169;
assign w47684 = pi08190 & w3106;
assign w47685 = pi05935 & w3344;
assign w47686 = pi08124 & w3446;
assign w47687 = pi02458 & w3110;
assign w47688 = pi04292 & w3334;
assign w47689 = pi03659 & w3260;
assign w47690 = pi08229 & w3546;
assign w47691 = pi02439 & w3150;
assign w47692 = pi07999 & w3516;
assign w47693 = pi07064 & w3286;
assign w47694 = pi07329 & w3620;
assign w47695 = pi02465 & w3524;
assign w47696 = pi07131 & w3420;
assign w47697 = pi03224 & w3336;
assign w47698 = pi08307 & w3294;
assign w47699 = pi04400 & w3512;
assign w47700 = pi04043 & w3118;
assign w47701 = pi06741 & w3514;
assign w47702 = pi02535 & w3160;
assign w47703 = pi01669 & w3580;
assign w47704 = pi07176 & w3364;
assign w47705 = pi03691 & w3310;
assign w47706 = pi07603 & w3372;
assign w47707 = pi03886 & w3338;
assign w47708 = pi06335 & w3538;
assign w47709 = pi08164 & w3594;
assign w47710 = pi03184 & w3380;
assign w47711 = pi02453 & w3418;
assign w47712 = pi06389 & w3298;
assign w47713 = pi06414 & w3392;
assign w47714 = pi02627 & w3300;
assign w47715 = pi07475 & w3508;
assign w47716 = pi02088 & w3330;
assign w47717 = pi06139 & w3480;
assign w47718 = pi07704 & w3430;
assign w47719 = pi05686 & w3486;
assign w47720 = pi07151 & w3135;
assign w47721 = pi06565 & w3462;
assign w47722 = pi06486 & w3199;
assign w47723 = pi05728 & w3240;
assign w47724 = pi06550 & w3304;
assign w47725 = pi01997 & w3610;
assign w47726 = pi03796 & w3350;
assign w47727 = pi07820 & w3464;
assign w47728 = pi03917 & w3348;
assign w47729 = pi06188 & w3356;
assign w47730 = pi02104 & w3096;
assign w47731 = pi04162 & w3454;
assign w47732 = pi04393 & w3618;
assign w47733 = pi08136 & w3570;
assign w47734 = pi02518 & w3586;
assign w47735 = pi04512 & w3488;
assign w47736 = pi04505 & w3582;
assign w47737 = pi04372 & w3146;
assign w47738 = pi07784 & w3192;
assign w47739 = pi02017 & w3242;
assign w47740 = pi04246 & w3290;
assign w47741 = pi08157 & w3366;
assign w47742 = pi04499 & w3211;
assign w47743 = pi06301 & w3482;
assign w47744 = pi07723 & w3171;
assign w47745 = pi06463 & w3129;
assign w47746 = pi07850 & w3270;
assign w47747 = pi07993 & w3426;
assign w47748 = pi05955 & w3492;
assign w47749 = pi02512 & w3254;
assign w47750 = pi06087 & w3550;
assign w47751 = pi02176 & w3280;
assign w47752 = pi02733 & w3432;
assign w47753 = pi03216 & w3197;
assign w47754 = pi03574 & w3103;
assign w47755 = pi06932 & w3398;
assign w47756 = pi04077 & w3428;
assign w47757 = pi07869 & w3386;
assign w47758 = pi03763 & w3526;
assign w47759 = pi07748 & w3458;
assign w47760 = pi07794 & w3360;
assign w47761 = pi06866 & w3442;
assign w47762 = pi06102 & w3568;
assign w47763 = pi02653 & w3156;
assign w47764 = pi06584 & w3496;
assign w47765 = pi08295 & w3342;
assign w47766 = pi04485 & w3588;
assign w47767 = pi08170 & w3468;
assign w47768 = pi02083 & w3530;
assign w47769 = pi06368 & w3450;
assign w47770 = pi07003 & w3406;
assign w47771 = pi04427 & w3302;
assign w47772 = pi04103 & w3522;
assign w47773 = pi08216 & w3282;
assign w47774 = pi05851 & w3248;
assign w47775 = pi02595 & w3368;
assign w47776 = pi07564 & w3165;
assign w47777 = pi01648 & w3572;
assign w47778 = pi03489 & w3250;
assign w47779 = pi02012 & w3292;
assign w47780 = pi02032 & w3318;
assign w47781 = pi07836 & w3207;
assign w47782 = pi06160 & w3112;
assign w47783 = ~w47527 & ~w47528;
assign w47784 = ~w47529 & ~w47530;
assign w47785 = ~w47531 & ~w47532;
assign w47786 = ~w47533 & ~w47534;
assign w47787 = ~w47535 & ~w47536;
assign w47788 = ~w47537 & ~w47538;
assign w47789 = ~w47539 & ~w47540;
assign w47790 = ~w47541 & ~w47542;
assign w47791 = ~w47543 & ~w47544;
assign w47792 = ~w47545 & ~w47546;
assign w47793 = ~w47547 & ~w47548;
assign w47794 = ~w47549 & ~w47550;
assign w47795 = ~w47551 & ~w47552;
assign w47796 = ~w47553 & ~w47554;
assign w47797 = ~w47555 & ~w47556;
assign w47798 = ~w47557 & ~w47558;
assign w47799 = ~w47559 & ~w47560;
assign w47800 = ~w47561 & ~w47562;
assign w47801 = ~w47563 & ~w47564;
assign w47802 = ~w47565 & ~w47566;
assign w47803 = ~w47567 & ~w47568;
assign w47804 = ~w47569 & ~w47570;
assign w47805 = ~w47571 & ~w47572;
assign w47806 = ~w47573 & ~w47574;
assign w47807 = ~w47575 & ~w47576;
assign w47808 = ~w47577 & ~w47578;
assign w47809 = ~w47579 & ~w47580;
assign w47810 = ~w47581 & ~w47582;
assign w47811 = ~w47583 & ~w47584;
assign w47812 = ~w47585 & ~w47586;
assign w47813 = ~w47587 & ~w47588;
assign w47814 = ~w47589 & ~w47590;
assign w47815 = ~w47591 & ~w47592;
assign w47816 = ~w47593 & ~w47594;
assign w47817 = ~w47595 & ~w47596;
assign w47818 = ~w47597 & ~w47598;
assign w47819 = ~w47599 & ~w47600;
assign w47820 = ~w47601 & ~w47602;
assign w47821 = ~w47603 & ~w47604;
assign w47822 = ~w47605 & ~w47606;
assign w47823 = ~w47607 & ~w47608;
assign w47824 = ~w47609 & ~w47610;
assign w47825 = ~w47611 & ~w47612;
assign w47826 = ~w47613 & ~w47614;
assign w47827 = ~w47615 & ~w47616;
assign w47828 = ~w47617 & ~w47618;
assign w47829 = ~w47619 & ~w47620;
assign w47830 = ~w47621 & ~w47622;
assign w47831 = ~w47623 & ~w47624;
assign w47832 = ~w47625 & ~w47626;
assign w47833 = ~w47627 & ~w47628;
assign w47834 = ~w47629 & ~w47630;
assign w47835 = ~w47631 & ~w47632;
assign w47836 = ~w47633 & ~w47634;
assign w47837 = ~w47635 & ~w47636;
assign w47838 = ~w47637 & ~w47638;
assign w47839 = ~w47639 & ~w47640;
assign w47840 = ~w47641 & ~w47642;
assign w47841 = ~w47643 & ~w47644;
assign w47842 = ~w47645 & ~w47646;
assign w47843 = ~w47647 & ~w47648;
assign w47844 = ~w47649 & ~w47650;
assign w47845 = ~w47651 & ~w47652;
assign w47846 = ~w47653 & ~w47654;
assign w47847 = ~w47655 & ~w47656;
assign w47848 = ~w47657 & ~w47658;
assign w47849 = ~w47659 & ~w47660;
assign w47850 = ~w47661 & ~w47662;
assign w47851 = ~w47663 & ~w47664;
assign w47852 = ~w47665 & ~w47666;
assign w47853 = ~w47667 & ~w47668;
assign w47854 = ~w47669 & ~w47670;
assign w47855 = ~w47671 & ~w47672;
assign w47856 = ~w47673 & ~w47674;
assign w47857 = ~w47675 & ~w47676;
assign w47858 = ~w47677 & ~w47678;
assign w47859 = ~w47679 & ~w47680;
assign w47860 = ~w47681 & ~w47682;
assign w47861 = ~w47683 & ~w47684;
assign w47862 = ~w47685 & ~w47686;
assign w47863 = ~w47687 & ~w47688;
assign w47864 = ~w47689 & ~w47690;
assign w47865 = ~w47691 & ~w47692;
assign w47866 = ~w47693 & ~w47694;
assign w47867 = ~w47695 & ~w47696;
assign w47868 = ~w47697 & ~w47698;
assign w47869 = ~w47699 & ~w47700;
assign w47870 = ~w47701 & ~w47702;
assign w47871 = ~w47703 & ~w47704;
assign w47872 = ~w47705 & ~w47706;
assign w47873 = ~w47707 & ~w47708;
assign w47874 = ~w47709 & ~w47710;
assign w47875 = ~w47711 & ~w47712;
assign w47876 = ~w47713 & ~w47714;
assign w47877 = ~w47715 & ~w47716;
assign w47878 = ~w47717 & ~w47718;
assign w47879 = ~w47719 & ~w47720;
assign w47880 = ~w47721 & ~w47722;
assign w47881 = ~w47723 & ~w47724;
assign w47882 = ~w47725 & ~w47726;
assign w47883 = ~w47727 & ~w47728;
assign w47884 = ~w47729 & ~w47730;
assign w47885 = ~w47731 & ~w47732;
assign w47886 = ~w47733 & ~w47734;
assign w47887 = ~w47735 & ~w47736;
assign w47888 = ~w47737 & ~w47738;
assign w47889 = ~w47739 & ~w47740;
assign w47890 = ~w47741 & ~w47742;
assign w47891 = ~w47743 & ~w47744;
assign w47892 = ~w47745 & ~w47746;
assign w47893 = ~w47747 & ~w47748;
assign w47894 = ~w47749 & ~w47750;
assign w47895 = ~w47751 & ~w47752;
assign w47896 = ~w47753 & ~w47754;
assign w47897 = ~w47755 & ~w47756;
assign w47898 = ~w47757 & ~w47758;
assign w47899 = ~w47759 & ~w47760;
assign w47900 = ~w47761 & ~w47762;
assign w47901 = ~w47763 & ~w47764;
assign w47902 = ~w47765 & ~w47766;
assign w47903 = ~w47767 & ~w47768;
assign w47904 = ~w47769 & ~w47770;
assign w47905 = ~w47771 & ~w47772;
assign w47906 = ~w47773 & ~w47774;
assign w47907 = ~w47775 & ~w47776;
assign w47908 = ~w47777 & ~w47778;
assign w47909 = ~w47779 & ~w47780;
assign w47910 = ~w47781 & ~w47782;
assign w47911 = w47909 & w47910;
assign w47912 = w47907 & w47908;
assign w47913 = w47905 & w47906;
assign w47914 = w47903 & w47904;
assign w47915 = w47901 & w47902;
assign w47916 = w47899 & w47900;
assign w47917 = w47897 & w47898;
assign w47918 = w47895 & w47896;
assign w47919 = w47893 & w47894;
assign w47920 = w47891 & w47892;
assign w47921 = w47889 & w47890;
assign w47922 = w47887 & w47888;
assign w47923 = w47885 & w47886;
assign w47924 = w47883 & w47884;
assign w47925 = w47881 & w47882;
assign w47926 = w47879 & w47880;
assign w47927 = w47877 & w47878;
assign w47928 = w47875 & w47876;
assign w47929 = w47873 & w47874;
assign w47930 = w47871 & w47872;
assign w47931 = w47869 & w47870;
assign w47932 = w47867 & w47868;
assign w47933 = w47865 & w47866;
assign w47934 = w47863 & w47864;
assign w47935 = w47861 & w47862;
assign w47936 = w47859 & w47860;
assign w47937 = w47857 & w47858;
assign w47938 = w47855 & w47856;
assign w47939 = w47853 & w47854;
assign w47940 = w47851 & w47852;
assign w47941 = w47849 & w47850;
assign w47942 = w47847 & w47848;
assign w47943 = w47845 & w47846;
assign w47944 = w47843 & w47844;
assign w47945 = w47841 & w47842;
assign w47946 = w47839 & w47840;
assign w47947 = w47837 & w47838;
assign w47948 = w47835 & w47836;
assign w47949 = w47833 & w47834;
assign w47950 = w47831 & w47832;
assign w47951 = w47829 & w47830;
assign w47952 = w47827 & w47828;
assign w47953 = w47825 & w47826;
assign w47954 = w47823 & w47824;
assign w47955 = w47821 & w47822;
assign w47956 = w47819 & w47820;
assign w47957 = w47817 & w47818;
assign w47958 = w47815 & w47816;
assign w47959 = w47813 & w47814;
assign w47960 = w47811 & w47812;
assign w47961 = w47809 & w47810;
assign w47962 = w47807 & w47808;
assign w47963 = w47805 & w47806;
assign w47964 = w47803 & w47804;
assign w47965 = w47801 & w47802;
assign w47966 = w47799 & w47800;
assign w47967 = w47797 & w47798;
assign w47968 = w47795 & w47796;
assign w47969 = w47793 & w47794;
assign w47970 = w47791 & w47792;
assign w47971 = w47789 & w47790;
assign w47972 = w47787 & w47788;
assign w47973 = w47785 & w47786;
assign w47974 = w47783 & w47784;
assign w47975 = w47973 & w47974;
assign w47976 = w47971 & w47972;
assign w47977 = w47969 & w47970;
assign w47978 = w47967 & w47968;
assign w47979 = w47965 & w47966;
assign w47980 = w47963 & w47964;
assign w47981 = w47961 & w47962;
assign w47982 = w47959 & w47960;
assign w47983 = w47957 & w47958;
assign w47984 = w47955 & w47956;
assign w47985 = w47953 & w47954;
assign w47986 = w47951 & w47952;
assign w47987 = w47949 & w47950;
assign w47988 = w47947 & w47948;
assign w47989 = w47945 & w47946;
assign w47990 = w47943 & w47944;
assign w47991 = w47941 & w47942;
assign w47992 = w47939 & w47940;
assign w47993 = w47937 & w47938;
assign w47994 = w47935 & w47936;
assign w47995 = w47933 & w47934;
assign w47996 = w47931 & w47932;
assign w47997 = w47929 & w47930;
assign w47998 = w47927 & w47928;
assign w47999 = w47925 & w47926;
assign w48000 = w47923 & w47924;
assign w48001 = w47921 & w47922;
assign w48002 = w47919 & w47920;
assign w48003 = w47917 & w47918;
assign w48004 = w47915 & w47916;
assign w48005 = w47913 & w47914;
assign w48006 = w47911 & w47912;
assign w48007 = w48005 & w48006;
assign w48008 = w48003 & w48004;
assign w48009 = w48001 & w48002;
assign w48010 = w47999 & w48000;
assign w48011 = w47997 & w47998;
assign w48012 = w47995 & w47996;
assign w48013 = w47993 & w47994;
assign w48014 = w47991 & w47992;
assign w48015 = w47989 & w47990;
assign w48016 = w47987 & w47988;
assign w48017 = w47985 & w47986;
assign w48018 = w47983 & w47984;
assign w48019 = w47981 & w47982;
assign w48020 = w47979 & w47980;
assign w48021 = w47977 & w47978;
assign w48022 = w47975 & w47976;
assign w48023 = w48021 & w48022;
assign w48024 = w48019 & w48020;
assign w48025 = w48017 & w48018;
assign w48026 = w48015 & w48016;
assign w48027 = w48013 & w48014;
assign w48028 = w48011 & w48012;
assign w48029 = w48009 & w48010;
assign w48030 = w48007 & w48008;
assign w48031 = w48029 & w48030;
assign w48032 = w48027 & w48028;
assign w48033 = w48025 & w48026;
assign w48034 = w48023 & w48024;
assign w48035 = w48033 & w48034;
assign w48036 = w48031 & w48032;
assign w48037 = w48035 & w48036;
assign w48038 = ~pi10577 & ~w48037;
assign w48039 = pi08617 & w3314;
assign w48040 = pi09336 & w3096;
assign w48041 = pi02109 & w3438;
assign w48042 = pi09160 & w3238;
assign w48043 = pi09186 & w3532;
assign w48044 = pi01973 & w3064;
assign w48045 = pi08540 & w3528;
assign w48046 = pi09748 & w3428;
assign w48047 = pi09134 & w3352;
assign w48048 = pi09786 & w3494;
assign w48049 = pi09265 & w3173;
assign w48050 = pi09389 & w3148;
assign w48051 = pi05067 & w3582;
assign w48052 = pi01957 & w3400;
assign w48053 = pi09317 & w3546;
assign w48054 = pi08443 & w3232;
assign w48055 = pi08977 & w3276;
assign w48056 = pi01575 & w3248;
assign w48057 = pi05028 & w3556;
assign w48058 = pi01604 & w3292;
assign w48059 = pi08990 & w3508;
assign w48060 = pi02086 & w3614;
assign w48061 = pi08462 & w3143;
assign w48062 = pi09721 & w3181;
assign w48063 = pi01993 & w3330;
assign w48064 = pi04588 & w3470;
assign w48065 = pi09008 & w3165;
assign w48066 = pi08624 & w3538;
assign w48067 = pi08847 & w3572;
assign w48068 = pi01763 & w3338;
assign w48069 = pi01932 & w3296;
assign w48070 = pi09147 & w3125;
assign w48071 = pi08729 & w3278;
assign w48072 = pi09231 & w3440;
assign w48073 = pi08801 & w3300;
assign w48074 = pi04968 & w3412;
assign w48075 = pi01963 & w3322;
assign w48076 = pi08808 & w3398;
assign w48077 = pi04916 & w3190;
assign w48078 = pi01967 & w3534;
assign w48079 = pi09192 & w3616;
assign w48080 = pi08776 & w3442;
assign w48081 = pi05147 & w3482;
assign w48082 = pi04873 & w3268;
assign w48083 = pi08768 & w3518;
assign w48084 = pi09178 & w3474;
assign w48085 = pi09350 & w3188;
assign w48086 = pi04955 & w3618;
assign w48087 = pi09410 & w3324;
assign w48088 = pi09363 & w3580;
assign w48089 = pi09476 & w3418;
assign w48090 = pi08944 & w3272;
assign w48091 = pi09173 & w3516;
assign w48092 = pi09497 & w3150;
assign w48093 = pi02635 & w3554;
assign w48094 = pi09304 & w3282;
assign w48095 = pi05074 & w3112;
assign w48096 = pi09443 & w3179;
assign w48097 = pi08581 & w3378;
assign w48098 = pi08918 & w3225;
assign w48099 = pi09456 & w3368;
assign w48100 = pi08742 & w3186;
assign w48101 = pi08755 & w3078;
assign w48102 = pi08507 & w3492;
assign w48103 = pi08970 & w3566;
assign w48104 = pi05060 & w3211;
assign w48105 = pi08892 & w3364;
assign w48106 = pi09510 & w3408;
assign w48107 = pi09323 & w3542;
assign w48108 = pi08702 & w3462;
assign w48109 = pi02422 & w3578;
assign w48110 = pi09343 & w3318;
assign w48111 = pi01849 & w3610;
assign w48112 = pi08853 & w3340;
assign w48113 = pi05034 & w3388;
assign w48114 = pi02047 & w3520;
assign w48115 = pi09016 & w3201;
assign w48116 = pi08951 & w3376;
assign w48117 = pi09469 & w3524;
assign w48118 = pi01951 & w3274;
assign w48119 = pi08643 & w3298;
assign w48120 = pi08535 & w3452;
assign w48121 = pi09252 & w3594;
assign w48122 = pi05396 & w3612;
assign w48123 = pi09291 & w3320;
assign w48124 = pi09076 & w3458;
assign w48125 = pi09082 & w3192;
assign w48126 = pi09069 & w3476;
assign w48127 = pi09376 & w3560;
assign w48128 = pi09258 & w3468;
assign w48129 = pi09062 & w3171;
assign w48130 = pi08438 & w3486;
assign w48131 = pi08964 & w3448;
assign w48132 = pi01837 & w3310;
assign w48133 = pi08455 & w3266;
assign w48134 = pi09549 & w3175;
assign w48135 = pi09095 & w3390;
assign w48136 = pi09088 & w3360;
assign w48137 = pi09238 & w3608;
assign w48138 = pi08886 & w3135;
assign w48139 = pi05079 & w3242;
assign w48140 = pi08788 & w3432;
assign w48141 = pi09489 & w3110;
assign w48142 = pi04949 & w3370;
assign w48143 = pi08834 & w3139;
assign w48144 = pi02438 & w3414;
assign w48145 = pi08899 & w3156;
assign w48146 = pi04994 & w3258;
assign w48147 = pi05001 & w3122;
assign w48148 = pi04988 & w3302;
assign w48149 = pi04569 & w3197;
assign w48150 = pi08669 & w3129;
assign w48151 = pi01509 & w3118;
assign w48152 = pi01702 & w3592;
assign w48153 = pi02557 & w3217;
assign w48154 = pi08546 & w3550;
assign w48155 = pi08656 & w3392;
assign w48156 = pi04962 & w3512;
assign w48157 = pi04981 & w3169;
assign w48158 = pi09720 & w3502;
assign w48159 = pi08708 & w3496;
assign w48160 = pi02000 & w3362;
assign w48161 = pi08873 & w3410;
assign w48162 = pi08996 & w3167;
assign w48163 = pi09056 & w3430;
assign w48164 = pi09284 & w3444;
assign w48165 = pi09212 & w3606;
assign w48166 = pi02813 & w3488;
assign w48167 = pi05047 & w3588;
assign w48168 = pi08564 & w3480;
assign w48169 = pi01788 & w3350;
assign w48170 = pi08551 & w3568;
assign w48171 = pi05054 & w3396;
assign w48172 = pi08761 & w3256;
assign w48173 = pi09370 & w3229;
assign w48174 = pi01715 & w3456;
assign w48175 = pi08879 & w3420;
assign w48176 = pi09330 & w3280;
assign w48177 = pi01942 & w3536;
assign w48178 = pi01854 & w3260;
assign w48179 = pi09218 & w3446;
assign w48180 = pi09108 & w3207;
assign w48181 = pi05015 & w3504;
assign w48182 = pi09245 & w3366;
assign w48183 = pi04538 & w3346;
assign w48184 = pi08689 & w3227;
assign w48185 = pi08502 & w3344;
assign w48186 = pi09022 & w3372;
assign w48187 = pi09036 & w3600;
assign w48188 = pi08715 & w3153;
assign w48189 = pi05007 & w3162;
assign w48190 = pi01955 & w3103;
assign w48191 = pi08957 & w3358;
assign w48192 = pi08597 & w3586;
assign w48193 = pi08840 & w3406;
assign w48194 = pi01603 & w3472;
assign w48195 = pi04890 & w3334;
assign w48196 = pi08983 & w3434;
assign w48197 = pi09049 & w3590;
assign w48198 = pi04910 & w3115;
assign w48199 = pi04877 & w3290;
assign w48200 = pi08814 & w3234;
assign w48201 = pi09225 & w3570;
assign w48202 = pi05041 & w3177;
assign w48203 = pi01941 & w3424;
assign w48204 = pi02397 & w3158;
assign w48205 = pi08905 & w3205;
assign w48206 = pi09043 & w3194;
assign w48207 = pi08860 & w3286;
assign w48208 = pi09310 & w3264;
assign w48209 = pi08748 & w3284;
assign w48210 = pi04903 & w3086;
assign w48211 = pi09029 & w3374;
assign w48212 = pi09403 & w3316;
assign w48213 = pi09205 & w3223;
assign w48214 = pi08487 & w3598;
assign w48215 = pi09430 & w3602;
assign w48216 = pi09114 & w3270;
assign w48217 = pi09483 & w3246;
assign w48218 = pi08450 & w3240;
assign w48219 = pi09709 & w3454;
assign w48220 = pi04581 & w3416;
assign w48221 = pi01728 & w3348;
assign w48222 = pi08682 & w3422;
assign w48223 = pi02572 & w3312;
assign w48224 = pi08827 & w3127;
assign w48225 = pi03404 & w3252;
assign w48226 = pi08781 & w3384;
assign w48227 = pi08722 & w3082;
assign w48228 = pi08557 & w3288;
assign w48229 = pi04523 & w3306;
assign w48230 = pi01631 & w3498;
assign w48231 = pi01772 & w3209;
assign w48232 = pi09153 & w3093;
assign w48233 = pi09271 & w3584;
assign w48234 = pi08931 & w3221;
assign w48235 = pi04936 & w3146;
assign w48236 = pi01515 & w3071;
assign w48237 = pi02007 & w3336;
assign w48238 = pi09101 & w3464;
assign w48239 = pi01542 & w3394;
assign w48240 = pi02564 & w3160;
assign w48241 = pi08591 & w3460;
assign w48242 = pi01986 & w3250;
assign w48243 = pi04975 & w3562;
assign w48244 = pi09396 & w3294;
assign w48245 = pi09416 & w3332;
assign w48246 = pi04804 & w3132;
assign w48247 = pi08474 & w3436;
assign w48248 = pi09383 & w3342;
assign w48249 = pi08525 & w3219;
assign w48250 = pi01906 & w3262;
assign w48251 = pi08695 & w3304;
assign w48252 = pi01838 & w3106;
assign w48253 = pi08650 & w3354;
assign w48254 = pi04884 & w3326;
assign w48255 = pi09121 & w3386;
assign w48256 = pi08495 & w3604;
assign w48257 = pi08866 & w3552;
assign w48258 = pi08676 & w3199;
assign w48259 = pi01990 & w3530;
assign w48260 = pi05021 & w3184;
assign w48261 = pi09516 & w3510;
assign w48262 = pi09503 & w3558;
assign w48263 = pi02022 & w3500;
assign w48264 = pi08938 & w3620;
assign w48265 = pi04929 & w3484;
assign w48266 = pi08586 & w3356;
assign w48267 = pi01799 & w3526;
assign w48268 = pi04897 & w3214;
assign w48269 = pi08821 & w3466;
assign w48270 = pi01785 & w3576;
assign w48271 = pi09166 & w3426;
assign w48272 = pi08795 & w3506;
assign w48273 = pi04942 & w3564;
assign w48274 = pi09357 & w3402;
assign w48275 = pi02366 & w3574;
assign w48276 = pi04561 & w3544;
assign w48277 = pi01810 & w3548;
assign w48278 = pi09297 & w3478;
assign w48279 = pi08630 & w3450;
assign w48280 = pi09708 & w3522;
assign w48281 = pi08735 & w3514;
assign w48282 = pi08912 & w3254;
assign w48283 = pi01812 & w3490;
assign w48284 = pi02067 & w3380;
assign w48285 = pi08663 & w3203;
assign w48286 = pi01807 & w3244;
assign w48287 = pi08609 & w3540;
assign w48288 = pi09140 & w3596;
assign w48289 = pi01925 & w3137;
assign w48290 = pi09127 & w3382;
assign w48291 = pi04923 & w3328;
assign w48292 = pi08637 & w3236;
assign w48293 = pi01998 & w3404;
assign w48294 = pi01541 & w3308;
assign w48295 = ~w48039 & ~w48040;
assign w48296 = ~w48041 & ~w48042;
assign w48297 = ~w48043 & ~w48044;
assign w48298 = ~w48045 & ~w48046;
assign w48299 = ~w48047 & ~w48048;
assign w48300 = ~w48049 & ~w48050;
assign w48301 = ~w48051 & ~w48052;
assign w48302 = ~w48053 & ~w48054;
assign w48303 = ~w48055 & ~w48056;
assign w48304 = ~w48057 & ~w48058;
assign w48305 = ~w48059 & ~w48060;
assign w48306 = ~w48061 & ~w48062;
assign w48307 = ~w48063 & ~w48064;
assign w48308 = ~w48065 & ~w48066;
assign w48309 = ~w48067 & ~w48068;
assign w48310 = ~w48069 & ~w48070;
assign w48311 = ~w48071 & ~w48072;
assign w48312 = ~w48073 & ~w48074;
assign w48313 = ~w48075 & ~w48076;
assign w48314 = ~w48077 & ~w48078;
assign w48315 = ~w48079 & ~w48080;
assign w48316 = ~w48081 & ~w48082;
assign w48317 = ~w48083 & ~w48084;
assign w48318 = ~w48085 & ~w48086;
assign w48319 = ~w48087 & ~w48088;
assign w48320 = ~w48089 & ~w48090;
assign w48321 = ~w48091 & ~w48092;
assign w48322 = ~w48093 & ~w48094;
assign w48323 = ~w48095 & ~w48096;
assign w48324 = ~w48097 & ~w48098;
assign w48325 = ~w48099 & ~w48100;
assign w48326 = ~w48101 & ~w48102;
assign w48327 = ~w48103 & ~w48104;
assign w48328 = ~w48105 & ~w48106;
assign w48329 = ~w48107 & ~w48108;
assign w48330 = ~w48109 & ~w48110;
assign w48331 = ~w48111 & ~w48112;
assign w48332 = ~w48113 & ~w48114;
assign w48333 = ~w48115 & ~w48116;
assign w48334 = ~w48117 & ~w48118;
assign w48335 = ~w48119 & ~w48120;
assign w48336 = ~w48121 & ~w48122;
assign w48337 = ~w48123 & ~w48124;
assign w48338 = ~w48125 & ~w48126;
assign w48339 = ~w48127 & ~w48128;
assign w48340 = ~w48129 & ~w48130;
assign w48341 = ~w48131 & ~w48132;
assign w48342 = ~w48133 & ~w48134;
assign w48343 = ~w48135 & ~w48136;
assign w48344 = ~w48137 & ~w48138;
assign w48345 = ~w48139 & ~w48140;
assign w48346 = ~w48141 & ~w48142;
assign w48347 = ~w48143 & ~w48144;
assign w48348 = ~w48145 & ~w48146;
assign w48349 = ~w48147 & ~w48148;
assign w48350 = ~w48149 & ~w48150;
assign w48351 = ~w48151 & ~w48152;
assign w48352 = ~w48153 & ~w48154;
assign w48353 = ~w48155 & ~w48156;
assign w48354 = ~w48157 & ~w48158;
assign w48355 = ~w48159 & ~w48160;
assign w48356 = ~w48161 & ~w48162;
assign w48357 = ~w48163 & ~w48164;
assign w48358 = ~w48165 & ~w48166;
assign w48359 = ~w48167 & ~w48168;
assign w48360 = ~w48169 & ~w48170;
assign w48361 = ~w48171 & ~w48172;
assign w48362 = ~w48173 & ~w48174;
assign w48363 = ~w48175 & ~w48176;
assign w48364 = ~w48177 & ~w48178;
assign w48365 = ~w48179 & ~w48180;
assign w48366 = ~w48181 & ~w48182;
assign w48367 = ~w48183 & ~w48184;
assign w48368 = ~w48185 & ~w48186;
assign w48369 = ~w48187 & ~w48188;
assign w48370 = ~w48189 & ~w48190;
assign w48371 = ~w48191 & ~w48192;
assign w48372 = ~w48193 & ~w48194;
assign w48373 = ~w48195 & ~w48196;
assign w48374 = ~w48197 & ~w48198;
assign w48375 = ~w48199 & ~w48200;
assign w48376 = ~w48201 & ~w48202;
assign w48377 = ~w48203 & ~w48204;
assign w48378 = ~w48205 & ~w48206;
assign w48379 = ~w48207 & ~w48208;
assign w48380 = ~w48209 & ~w48210;
assign w48381 = ~w48211 & ~w48212;
assign w48382 = ~w48213 & ~w48214;
assign w48383 = ~w48215 & ~w48216;
assign w48384 = ~w48217 & ~w48218;
assign w48385 = ~w48219 & ~w48220;
assign w48386 = ~w48221 & ~w48222;
assign w48387 = ~w48223 & ~w48224;
assign w48388 = ~w48225 & ~w48226;
assign w48389 = ~w48227 & ~w48228;
assign w48390 = ~w48229 & ~w48230;
assign w48391 = ~w48231 & ~w48232;
assign w48392 = ~w48233 & ~w48234;
assign w48393 = ~w48235 & ~w48236;
assign w48394 = ~w48237 & ~w48238;
assign w48395 = ~w48239 & ~w48240;
assign w48396 = ~w48241 & ~w48242;
assign w48397 = ~w48243 & ~w48244;
assign w48398 = ~w48245 & ~w48246;
assign w48399 = ~w48247 & ~w48248;
assign w48400 = ~w48249 & ~w48250;
assign w48401 = ~w48251 & ~w48252;
assign w48402 = ~w48253 & ~w48254;
assign w48403 = ~w48255 & ~w48256;
assign w48404 = ~w48257 & ~w48258;
assign w48405 = ~w48259 & ~w48260;
assign w48406 = ~w48261 & ~w48262;
assign w48407 = ~w48263 & ~w48264;
assign w48408 = ~w48265 & ~w48266;
assign w48409 = ~w48267 & ~w48268;
assign w48410 = ~w48269 & ~w48270;
assign w48411 = ~w48271 & ~w48272;
assign w48412 = ~w48273 & ~w48274;
assign w48413 = ~w48275 & ~w48276;
assign w48414 = ~w48277 & ~w48278;
assign w48415 = ~w48279 & ~w48280;
assign w48416 = ~w48281 & ~w48282;
assign w48417 = ~w48283 & ~w48284;
assign w48418 = ~w48285 & ~w48286;
assign w48419 = ~w48287 & ~w48288;
assign w48420 = ~w48289 & ~w48290;
assign w48421 = ~w48291 & ~w48292;
assign w48422 = ~w48293 & ~w48294;
assign w48423 = w48421 & w48422;
assign w48424 = w48419 & w48420;
assign w48425 = w48417 & w48418;
assign w48426 = w48415 & w48416;
assign w48427 = w48413 & w48414;
assign w48428 = w48411 & w48412;
assign w48429 = w48409 & w48410;
assign w48430 = w48407 & w48408;
assign w48431 = w48405 & w48406;
assign w48432 = w48403 & w48404;
assign w48433 = w48401 & w48402;
assign w48434 = w48399 & w48400;
assign w48435 = w48397 & w48398;
assign w48436 = w48395 & w48396;
assign w48437 = w48393 & w48394;
assign w48438 = w48391 & w48392;
assign w48439 = w48389 & w48390;
assign w48440 = w48387 & w48388;
assign w48441 = w48385 & w48386;
assign w48442 = w48383 & w48384;
assign w48443 = w48381 & w48382;
assign w48444 = w48379 & w48380;
assign w48445 = w48377 & w48378;
assign w48446 = w48375 & w48376;
assign w48447 = w48373 & w48374;
assign w48448 = w48371 & w48372;
assign w48449 = w48369 & w48370;
assign w48450 = w48367 & w48368;
assign w48451 = w48365 & w48366;
assign w48452 = w48363 & w48364;
assign w48453 = w48361 & w48362;
assign w48454 = w48359 & w48360;
assign w48455 = w48357 & w48358;
assign w48456 = w48355 & w48356;
assign w48457 = w48353 & w48354;
assign w48458 = w48351 & w48352;
assign w48459 = w48349 & w48350;
assign w48460 = w48347 & w48348;
assign w48461 = w48345 & w48346;
assign w48462 = w48343 & w48344;
assign w48463 = w48341 & w48342;
assign w48464 = w48339 & w48340;
assign w48465 = w48337 & w48338;
assign w48466 = w48335 & w48336;
assign w48467 = w48333 & w48334;
assign w48468 = w48331 & w48332;
assign w48469 = w48329 & w48330;
assign w48470 = w48327 & w48328;
assign w48471 = w48325 & w48326;
assign w48472 = w48323 & w48324;
assign w48473 = w48321 & w48322;
assign w48474 = w48319 & w48320;
assign w48475 = w48317 & w48318;
assign w48476 = w48315 & w48316;
assign w48477 = w48313 & w48314;
assign w48478 = w48311 & w48312;
assign w48479 = w48309 & w48310;
assign w48480 = w48307 & w48308;
assign w48481 = w48305 & w48306;
assign w48482 = w48303 & w48304;
assign w48483 = w48301 & w48302;
assign w48484 = w48299 & w48300;
assign w48485 = w48297 & w48298;
assign w48486 = w48295 & w48296;
assign w48487 = w48485 & w48486;
assign w48488 = w48483 & w48484;
assign w48489 = w48481 & w48482;
assign w48490 = w48479 & w48480;
assign w48491 = w48477 & w48478;
assign w48492 = w48475 & w48476;
assign w48493 = w48473 & w48474;
assign w48494 = w48471 & w48472;
assign w48495 = w48469 & w48470;
assign w48496 = w48467 & w48468;
assign w48497 = w48465 & w48466;
assign w48498 = w48463 & w48464;
assign w48499 = w48461 & w48462;
assign w48500 = w48459 & w48460;
assign w48501 = w48457 & w48458;
assign w48502 = w48455 & w48456;
assign w48503 = w48453 & w48454;
assign w48504 = w48451 & w48452;
assign w48505 = w48449 & w48450;
assign w48506 = w48447 & w48448;
assign w48507 = w48445 & w48446;
assign w48508 = w48443 & w48444;
assign w48509 = w48441 & w48442;
assign w48510 = w48439 & w48440;
assign w48511 = w48437 & w48438;
assign w48512 = w48435 & w48436;
assign w48513 = w48433 & w48434;
assign w48514 = w48431 & w48432;
assign w48515 = w48429 & w48430;
assign w48516 = w48427 & w48428;
assign w48517 = w48425 & w48426;
assign w48518 = w48423 & w48424;
assign w48519 = w48517 & w48518;
assign w48520 = w48515 & w48516;
assign w48521 = w48513 & w48514;
assign w48522 = w48511 & w48512;
assign w48523 = w48509 & w48510;
assign w48524 = w48507 & w48508;
assign w48525 = w48505 & w48506;
assign w48526 = w48503 & w48504;
assign w48527 = w48501 & w48502;
assign w48528 = w48499 & w48500;
assign w48529 = w48497 & w48498;
assign w48530 = w48495 & w48496;
assign w48531 = w48493 & w48494;
assign w48532 = w48491 & w48492;
assign w48533 = w48489 & w48490;
assign w48534 = w48487 & w48488;
assign w48535 = w48533 & w48534;
assign w48536 = w48531 & w48532;
assign w48537 = w48529 & w48530;
assign w48538 = w48527 & w48528;
assign w48539 = w48525 & w48526;
assign w48540 = w48523 & w48524;
assign w48541 = w48521 & w48522;
assign w48542 = w48519 & w48520;
assign w48543 = w48541 & w48542;
assign w48544 = w48539 & w48540;
assign w48545 = w48537 & w48538;
assign w48546 = w48535 & w48536;
assign w48547 = w48545 & w48546;
assign w48548 = w48543 & w48544;
assign w48549 = w48547 & w48548;
assign w48550 = ~pi10577 & ~w48549;
assign w48551 = pi04917 & w3190;
assign w48552 = pi09009 & w3165;
assign w48553 = pi04524 & w3306;
assign w48554 = pi08592 & w3460;
assign w48555 = pi08576 & w3112;
assign w48556 = pi09351 & w3188;
assign w48557 = pi08867 & w3552;
assign w48558 = pi04832 & w3574;
assign w48559 = pi09023 & w3372;
assign w48560 = pi05348 & w3378;
assign w48561 = pi09232 & w3440;
assign w48562 = pi04725 & w3244;
assign w48563 = pi02501 & w3356;
assign w48564 = pi04963 & w3512;
assign w48565 = pi08657 & w3392;
assign w48566 = pi04517 & w3614;
assign w48567 = pi05022 & w3184;
assign w48568 = pi02561 & w3276;
assign w48569 = pi02542 & w3135;
assign w48570 = pi04825 & w3118;
assign w48571 = pi05042 & w3177;
assign w48572 = pi08789 & w3432;
assign w48573 = pi09324 & w3542;
assign w48574 = pi01555 & w3572;
assign w48575 = pi08971 & w3566;
assign w48576 = pi04858 & w3181;
assign w48577 = pi04989 & w3302;
assign w48578 = pi08638 & w3236;
assign w48579 = pi08854 & w3340;
assign w48580 = pi09199 & w3175;
assign w48581 = pi02331 & w3173;
assign w48582 = pi04878 & w3290;
assign w48583 = pi01525 & w3620;
assign w48584 = pi08984 & w3434;
assign w48585 = pi02560 & w3318;
assign w48586 = pi02335 & w3608;
assign w48587 = pi08503 & w3219;
assign w48588 = pi09444 & w3179;
assign w48589 = pi01858 & w3374;
assign w48590 = pi08736 & w3514;
assign w48591 = pi04539 & w3346;
assign w48592 = pi04885 & w3326;
assign w48593 = pi08696 & w3304;
assign w48594 = pi05029 & w3556;
assign w48595 = pi04562 & w3544;
assign w48596 = pi09272 & w3584;
assign w48597 = pi04891 & w3334;
assign w48598 = pi08565 & w3480;
assign w48599 = pi08677 & w3199;
assign w48600 = pi04851 & w3522;
assign w48601 = pi01571 & w3402;
assign w48602 = pi04797 & w3498;
assign w48603 = pi04666 & w3536;
assign w48604 = pi04757 & w3576;
assign w48605 = pi08463 & w3143;
assign w48606 = pi01813 & w3398;
assign w48607 = pi09259 & w3468;
assign w48608 = pi01949 & w3352;
assign w48609 = pi04653 & w3103;
assign w48610 = pi09364 & w3580;
assign w48611 = pi04805 & w3132;
assign w48612 = pi08893 & w3364;
assign w48613 = pi02446 & w3518;
assign w48614 = pi04930 & w3484;
assign w48615 = pi04937 & w3146;
assign w48616 = pi04550 & w3197;
assign w48617 = pi04982 & w3169;
assign w48618 = pi02543 & w3238;
assign w48619 = pi04898 & w3214;
assign w48620 = pi08514 & w3612;
assign w48621 = pi09517 & w3510;
assign w48622 = pi04614 & w3530;
assign w48623 = pi09450 & w3438;
assign w48624 = pi04589 & w3470;
assign w48625 = pi02485 & w3516;
assign w48626 = pi09463 & w3160;
assign w48627 = pi08618 & w3314;
assign w48628 = pi09404 & w3316;
assign w48629 = pi09390 & w3148;
assign w48630 = pi08716 & w3153;
assign w48631 = pi04943 & w3564;
assign w48632 = pi04530 & w3380;
assign w48633 = pi08958 & w3358;
assign w48634 = pi01931 & w3254;
assign w48635 = pi09285 & w3444;
assign w48636 = pi09457 & w3368;
assign w48637 = pi02244 & w3482;
assign w48638 = pi08468 & w3308;
assign w48639 = pi08520 & w3252;
assign w48640 = pi09377 & w3560;
assign w48641 = pi08945 & w3272;
assign w48642 = pi04568 & w3500;
assign w48643 = pi04660 & w3274;
assign w48644 = pi04545 & w3520;
assign w48645 = pi04595 & w3362;
assign w48646 = pi01652 & w3282;
assign w48647 = pi09498 & w3150;
assign w48648 = pi08723 & w3082;
assign w48649 = pi08775 & w3442;
assign w48650 = pi08530 & w3554;
assign w48651 = pi04640 & w3400;
assign w48652 = pi09311 & w3264;
assign w48653 = pi09154 & w3093;
assign w48654 = pi08481 & w3248;
assign w48655 = pi09246 & w3366;
assign w48656 = pi09477 & w3418;
assign w48657 = pi09128 & w3382;
assign w48658 = pi08802 & w3300;
assign w48659 = pi01601 & w3203;
assign w48660 = pi04718 & w3310;
assign w48661 = pi09417 & w3332;
assign w48662 = pi04791 & w3592;
assign w48663 = pi02474 & w3186;
assign w48664 = pi08437 & w3486;
assign w48665 = pi02544 & w3386;
assign w48666 = pi09484 & w3246;
assign w48667 = pi08598 & w3586;
assign w48668 = pi04556 & w3336;
assign w48669 = pi04811 & w3394;
assign w48670 = pi08841 & w3406;
assign w48671 = pi04744 & w3526;
assign w48672 = pi04705 & w3260;
assign w48673 = pi02594 & w3278;
assign w48674 = pi09089 & w3360;
assign w48675 = pi08644 & w3298;
assign w48676 = pi04838 & w3494;
assign w48677 = pi04699 & w3292;
assign w48678 = pi08651 & w3354;
assign w48679 = pi01561 & w3139;
assign w48680 = pi04686 & w3137;
assign w48681 = pi04627 & w3064;
assign w48682 = pi05055 & w3396;
assign w48683 = pi08603 & w3414;
assign w48684 = pi08690 & w3227;
assign w48685 = pi02582 & w3410;
assign w48686 = pi04976 & w3562;
assign w48687 = pi04764 & w3209;
assign w48688 = pi04712 & w3610;
assign w48689 = pi05008 & w3162;
assign w48690 = pi04995 & w3258;
assign w48691 = pi05035 & w3388;
assign w48692 = pi08709 & w3496;
assign w48693 = pi04673 & w3424;
assign w48694 = pi04574 & w3268;
assign w48695 = pi08919 & w3225;
assign w48696 = pi08558 & w3288;
assign w48697 = pi04731 & w3548;
assign w48698 = pi08932 & w3221;
assign w48699 = pi02479 & w3342;
assign w48700 = pi01725 & w3546;
assign w48701 = pi01909 & w3194;
assign w48702 = pi08631 & w3450;
assign w48703 = pi08828 & w3127;
assign w48704 = pi08547 & w3550;
assign w48705 = pi09504 & w3558;
assign w48706 = pi09037 & w3600;
assign w48707 = pi09337 & w3096;
assign w48708 = pi08488 & w3598;
assign w48709 = pi04771 & w3338;
assign w48710 = pi01583 & w3376;
assign w48711 = pi04679 & w3296;
assign w48712 = pi04608 & w3330;
assign w48713 = pi08496 & w3604;
assign w48714 = pi09278 & w3106;
assign w48715 = pi04864 & w3502;
assign w48716 = pi07569 & w3606;
assign w48717 = pi08925 & w3472;
assign w48718 = pi02541 & w3201;
assign w48719 = pi05712 & w3192;
assign w48720 = pi04911 & w3115;
assign w48721 = pi02606 & w3452;
assign w48722 = pi04818 & w3071;
assign w48723 = pi08749 & w3284;
assign w48724 = pi04871 & w3454;
assign w48725 = pi09298 & w3478;
assign w48726 = pi09470 & w3524;
assign w48727 = pi02587 & w3532;
assign w48728 = pi04969 & w3412;
assign w48729 = pi02470 & w3078;
assign w48730 = pi01911 & w3506;
assign w48731 = pi08451 & w3240;
assign w48732 = pi04738 & w3490;
assign w48733 = pi04784 & w3456;
assign w48734 = pi02814 & w3488;
assign w48735 = pi08880 & w3420;
assign w48736 = pi09206 & w3223;
assign w48737 = pi09511 & w3408;
assign w48738 = pi08683 & w3422;
assign w48739 = pi08475 & w3436;
assign w48740 = pi04845 & w3428;
assign w48741 = pi08542 & w3528;
assign w48742 = pi01798 & w3430;
assign w48743 = pi04621 & w3250;
assign w48744 = pi04904 & w3086;
assign w48745 = pi04582 & w3416;
assign w48746 = pi09075 & w3458;
assign w48747 = pi09141 & w3596;
assign w48748 = pi09193 & w3616;
assign w48749 = pi09424 & w3158;
assign w48750 = pi01524 & w3156;
assign w48751 = pi05002 & w3122;
assign w48752 = pi05068 & w3582;
assign w48753 = pi04692 & w3262;
assign w48754 = pi08552 & w3568;
assign w48755 = pi05791 & w3286;
assign w48756 = pi08670 & w3129;
assign w48757 = pi07650 & w3217;
assign w48758 = pi09437 & w3578;
assign w48759 = pi05061 & w3211;
assign w48760 = pi02610 & w3390;
assign w48761 = pi01529 & w3229;
assign w48762 = pi01519 & w3280;
assign w48763 = pi02332 & w3594;
assign w48764 = pi09102 & w3464;
assign w48765 = pi01598 & w3466;
assign w48766 = pi01685 & w3320;
assign w48767 = pi08444 & w3232;
assign w48768 = pi01910 & w3540;
assign w48769 = pi05048 & w3588;
assign w48770 = pi08762 & w3256;
assign w48771 = pi09050 & w3590;
assign w48772 = pi08625 & w3538;
assign w48773 = pi08815 & w3234;
assign w48774 = pi01558 & w3476;
assign w48775 = pi04601 & w3404;
assign w48776 = pi09179 & w3474;
assign w48777 = pi01550 & w3448;
assign w48778 = pi04956 & w3618;
assign w48779 = pi02586 & w3294;
assign w48780 = pi08906 & w3205;
assign w48781 = pi08703 & w3462;
assign w48782 = pi02289 & w3570;
assign w48783 = pi02510 & w3324;
assign w48784 = pi09219 & w3446;
assign w48785 = pi09167 & w3426;
assign w48786 = pi09431 & w3602;
assign w48787 = pi08782 & w3384;
assign w48788 = pi02741 & w3242;
assign w48789 = pi09063 & w3171;
assign w48790 = pi04950 & w3370;
assign w48791 = pi04751 & w3350;
assign w48792 = pi09490 & w3110;
assign w48793 = pi08997 & w3167;
assign w48794 = pi02609 & w3207;
assign w48795 = pi09756 & w3125;
assign w48796 = pi04924 & w3328;
assign w48797 = pi02597 & w3508;
assign w48798 = pi09115 & w3270;
assign w48799 = pi02255 & w3344;
assign w48800 = pi08508 & w3492;
assign w48801 = pi05016 & w3504;
assign w48802 = pi04647 & w3322;
assign w48803 = pi09003 & w3312;
assign w48804 = pi04778 & w3348;
assign w48805 = pi04634 & w3534;
assign w48806 = pi08456 & w3266;
assign w48807 = ~w48551 & ~w48552;
assign w48808 = ~w48553 & ~w48554;
assign w48809 = ~w48555 & ~w48556;
assign w48810 = ~w48557 & ~w48558;
assign w48811 = ~w48559 & ~w48560;
assign w48812 = ~w48561 & ~w48562;
assign w48813 = ~w48563 & ~w48564;
assign w48814 = ~w48565 & ~w48566;
assign w48815 = ~w48567 & ~w48568;
assign w48816 = ~w48569 & ~w48570;
assign w48817 = ~w48571 & ~w48572;
assign w48818 = ~w48573 & ~w48574;
assign w48819 = ~w48575 & ~w48576;
assign w48820 = ~w48577 & ~w48578;
assign w48821 = ~w48579 & ~w48580;
assign w48822 = ~w48581 & ~w48582;
assign w48823 = ~w48583 & ~w48584;
assign w48824 = ~w48585 & ~w48586;
assign w48825 = ~w48587 & ~w48588;
assign w48826 = ~w48589 & ~w48590;
assign w48827 = ~w48591 & ~w48592;
assign w48828 = ~w48593 & ~w48594;
assign w48829 = ~w48595 & ~w48596;
assign w48830 = ~w48597 & ~w48598;
assign w48831 = ~w48599 & ~w48600;
assign w48832 = ~w48601 & ~w48602;
assign w48833 = ~w48603 & ~w48604;
assign w48834 = ~w48605 & ~w48606;
assign w48835 = ~w48607 & ~w48608;
assign w48836 = ~w48609 & ~w48610;
assign w48837 = ~w48611 & ~w48612;
assign w48838 = ~w48613 & ~w48614;
assign w48839 = ~w48615 & ~w48616;
assign w48840 = ~w48617 & ~w48618;
assign w48841 = ~w48619 & ~w48620;
assign w48842 = ~w48621 & ~w48622;
assign w48843 = ~w48623 & ~w48624;
assign w48844 = ~w48625 & ~w48626;
assign w48845 = ~w48627 & ~w48628;
assign w48846 = ~w48629 & ~w48630;
assign w48847 = ~w48631 & ~w48632;
assign w48848 = ~w48633 & ~w48634;
assign w48849 = ~w48635 & ~w48636;
assign w48850 = ~w48637 & ~w48638;
assign w48851 = ~w48639 & ~w48640;
assign w48852 = ~w48641 & ~w48642;
assign w48853 = ~w48643 & ~w48644;
assign w48854 = ~w48645 & ~w48646;
assign w48855 = ~w48647 & ~w48648;
assign w48856 = ~w48649 & ~w48650;
assign w48857 = ~w48651 & ~w48652;
assign w48858 = ~w48653 & ~w48654;
assign w48859 = ~w48655 & ~w48656;
assign w48860 = ~w48657 & ~w48658;
assign w48861 = ~w48659 & ~w48660;
assign w48862 = ~w48661 & ~w48662;
assign w48863 = ~w48663 & ~w48664;
assign w48864 = ~w48665 & ~w48666;
assign w48865 = ~w48667 & ~w48668;
assign w48866 = ~w48669 & ~w48670;
assign w48867 = ~w48671 & ~w48672;
assign w48868 = ~w48673 & ~w48674;
assign w48869 = ~w48675 & ~w48676;
assign w48870 = ~w48677 & ~w48678;
assign w48871 = ~w48679 & ~w48680;
assign w48872 = ~w48681 & ~w48682;
assign w48873 = ~w48683 & ~w48684;
assign w48874 = ~w48685 & ~w48686;
assign w48875 = ~w48687 & ~w48688;
assign w48876 = ~w48689 & ~w48690;
assign w48877 = ~w48691 & ~w48692;
assign w48878 = ~w48693 & ~w48694;
assign w48879 = ~w48695 & ~w48696;
assign w48880 = ~w48697 & ~w48698;
assign w48881 = ~w48699 & ~w48700;
assign w48882 = ~w48701 & ~w48702;
assign w48883 = ~w48703 & ~w48704;
assign w48884 = ~w48705 & ~w48706;
assign w48885 = ~w48707 & ~w48708;
assign w48886 = ~w48709 & ~w48710;
assign w48887 = ~w48711 & ~w48712;
assign w48888 = ~w48713 & ~w48714;
assign w48889 = ~w48715 & ~w48716;
assign w48890 = ~w48717 & ~w48718;
assign w48891 = ~w48719 & ~w48720;
assign w48892 = ~w48721 & ~w48722;
assign w48893 = ~w48723 & ~w48724;
assign w48894 = ~w48725 & ~w48726;
assign w48895 = ~w48727 & ~w48728;
assign w48896 = ~w48729 & ~w48730;
assign w48897 = ~w48731 & ~w48732;
assign w48898 = ~w48733 & ~w48734;
assign w48899 = ~w48735 & ~w48736;
assign w48900 = ~w48737 & ~w48738;
assign w48901 = ~w48739 & ~w48740;
assign w48902 = ~w48741 & ~w48742;
assign w48903 = ~w48743 & ~w48744;
assign w48904 = ~w48745 & ~w48746;
assign w48905 = ~w48747 & ~w48748;
assign w48906 = ~w48749 & ~w48750;
assign w48907 = ~w48751 & ~w48752;
assign w48908 = ~w48753 & ~w48754;
assign w48909 = ~w48755 & ~w48756;
assign w48910 = ~w48757 & ~w48758;
assign w48911 = ~w48759 & ~w48760;
assign w48912 = ~w48761 & ~w48762;
assign w48913 = ~w48763 & ~w48764;
assign w48914 = ~w48765 & ~w48766;
assign w48915 = ~w48767 & ~w48768;
assign w48916 = ~w48769 & ~w48770;
assign w48917 = ~w48771 & ~w48772;
assign w48918 = ~w48773 & ~w48774;
assign w48919 = ~w48775 & ~w48776;
assign w48920 = ~w48777 & ~w48778;
assign w48921 = ~w48779 & ~w48780;
assign w48922 = ~w48781 & ~w48782;
assign w48923 = ~w48783 & ~w48784;
assign w48924 = ~w48785 & ~w48786;
assign w48925 = ~w48787 & ~w48788;
assign w48926 = ~w48789 & ~w48790;
assign w48927 = ~w48791 & ~w48792;
assign w48928 = ~w48793 & ~w48794;
assign w48929 = ~w48795 & ~w48796;
assign w48930 = ~w48797 & ~w48798;
assign w48931 = ~w48799 & ~w48800;
assign w48932 = ~w48801 & ~w48802;
assign w48933 = ~w48803 & ~w48804;
assign w48934 = ~w48805 & ~w48806;
assign w48935 = w48933 & w48934;
assign w48936 = w48931 & w48932;
assign w48937 = w48929 & w48930;
assign w48938 = w48927 & w48928;
assign w48939 = w48925 & w48926;
assign w48940 = w48923 & w48924;
assign w48941 = w48921 & w48922;
assign w48942 = w48919 & w48920;
assign w48943 = w48917 & w48918;
assign w48944 = w48915 & w48916;
assign w48945 = w48913 & w48914;
assign w48946 = w48911 & w48912;
assign w48947 = w48909 & w48910;
assign w48948 = w48907 & w48908;
assign w48949 = w48905 & w48906;
assign w48950 = w48903 & w48904;
assign w48951 = w48901 & w48902;
assign w48952 = w48899 & w48900;
assign w48953 = w48897 & w48898;
assign w48954 = w48895 & w48896;
assign w48955 = w48893 & w48894;
assign w48956 = w48891 & w48892;
assign w48957 = w48889 & w48890;
assign w48958 = w48887 & w48888;
assign w48959 = w48885 & w48886;
assign w48960 = w48883 & w48884;
assign w48961 = w48881 & w48882;
assign w48962 = w48879 & w48880;
assign w48963 = w48877 & w48878;
assign w48964 = w48875 & w48876;
assign w48965 = w48873 & w48874;
assign w48966 = w48871 & w48872;
assign w48967 = w48869 & w48870;
assign w48968 = w48867 & w48868;
assign w48969 = w48865 & w48866;
assign w48970 = w48863 & w48864;
assign w48971 = w48861 & w48862;
assign w48972 = w48859 & w48860;
assign w48973 = w48857 & w48858;
assign w48974 = w48855 & w48856;
assign w48975 = w48853 & w48854;
assign w48976 = w48851 & w48852;
assign w48977 = w48849 & w48850;
assign w48978 = w48847 & w48848;
assign w48979 = w48845 & w48846;
assign w48980 = w48843 & w48844;
assign w48981 = w48841 & w48842;
assign w48982 = w48839 & w48840;
assign w48983 = w48837 & w48838;
assign w48984 = w48835 & w48836;
assign w48985 = w48833 & w48834;
assign w48986 = w48831 & w48832;
assign w48987 = w48829 & w48830;
assign w48988 = w48827 & w48828;
assign w48989 = w48825 & w48826;
assign w48990 = w48823 & w48824;
assign w48991 = w48821 & w48822;
assign w48992 = w48819 & w48820;
assign w48993 = w48817 & w48818;
assign w48994 = w48815 & w48816;
assign w48995 = w48813 & w48814;
assign w48996 = w48811 & w48812;
assign w48997 = w48809 & w48810;
assign w48998 = w48807 & w48808;
assign w48999 = w48997 & w48998;
assign w49000 = w48995 & w48996;
assign w49001 = w48993 & w48994;
assign w49002 = w48991 & w48992;
assign w49003 = w48989 & w48990;
assign w49004 = w48987 & w48988;
assign w49005 = w48985 & w48986;
assign w49006 = w48983 & w48984;
assign w49007 = w48981 & w48982;
assign w49008 = w48979 & w48980;
assign w49009 = w48977 & w48978;
assign w49010 = w48975 & w48976;
assign w49011 = w48973 & w48974;
assign w49012 = w48971 & w48972;
assign w49013 = w48969 & w48970;
assign w49014 = w48967 & w48968;
assign w49015 = w48965 & w48966;
assign w49016 = w48963 & w48964;
assign w49017 = w48961 & w48962;
assign w49018 = w48959 & w48960;
assign w49019 = w48957 & w48958;
assign w49020 = w48955 & w48956;
assign w49021 = w48953 & w48954;
assign w49022 = w48951 & w48952;
assign w49023 = w48949 & w48950;
assign w49024 = w48947 & w48948;
assign w49025 = w48945 & w48946;
assign w49026 = w48943 & w48944;
assign w49027 = w48941 & w48942;
assign w49028 = w48939 & w48940;
assign w49029 = w48937 & w48938;
assign w49030 = w48935 & w48936;
assign w49031 = w49029 & w49030;
assign w49032 = w49027 & w49028;
assign w49033 = w49025 & w49026;
assign w49034 = w49023 & w49024;
assign w49035 = w49021 & w49022;
assign w49036 = w49019 & w49020;
assign w49037 = w49017 & w49018;
assign w49038 = w49015 & w49016;
assign w49039 = w49013 & w49014;
assign w49040 = w49011 & w49012;
assign w49041 = w49009 & w49010;
assign w49042 = w49007 & w49008;
assign w49043 = w49005 & w49006;
assign w49044 = w49003 & w49004;
assign w49045 = w49001 & w49002;
assign w49046 = w48999 & w49000;
assign w49047 = w49045 & w49046;
assign w49048 = w49043 & w49044;
assign w49049 = w49041 & w49042;
assign w49050 = w49039 & w49040;
assign w49051 = w49037 & w49038;
assign w49052 = w49035 & w49036;
assign w49053 = w49033 & w49034;
assign w49054 = w49031 & w49032;
assign w49055 = w49053 & w49054;
assign w49056 = w49051 & w49052;
assign w49057 = w49049 & w49050;
assign w49058 = w49047 & w49048;
assign w49059 = w49057 & w49058;
assign w49060 = w49055 & w49056;
assign w49061 = w49059 & w49060;
assign w49062 = ~pi10577 & ~w49061;
assign w49063 = pi08141 & w3440;
assign w49064 = pi08189 & w3106;
assign w49065 = pi06203 & w3460;
assign w49066 = pi08163 & w3594;
assign w49067 = pi03885 & w3338;
assign w49068 = pi03263 & w3500;
assign w49069 = pi02492 & w3430;
assign w49070 = pi08255 & w3318;
assign w49071 = pi04394 & w3618;
assign w49072 = pi06413 & w3392;
assign w49073 = pi08360 & w3438;
assign w49074 = pi07847 & w3270;
assign w49075 = pi07974 & w3238;
assign w49076 = pi08379 & w3524;
assign w49077 = pi07148 & w3135;
assign w49078 = pi06387 & w3298;
assign w49079 = pi07340 & w3272;
assign w49080 = pi06305 & w3482;
assign w49081 = pi06461 & w3129;
assign w49082 = pi08176 & w3173;
assign w49083 = pi06891 & w3432;
assign w49084 = pi09563 & w3620;
assign w49085 = pi04365 & w3484;
assign w49086 = pi04478 & w3177;
assign w49087 = pi08294 & w3342;
assign w49088 = pi08202 & w3320;
assign w49089 = pi07907 & w3352;
assign w49090 = pi07002 & w3406;
assign w49091 = pi04407 & w3412;
assign w49092 = pi04076 & w3428;
assign w49093 = pi06738 & w3514;
assign w49094 = pi05849 & w3248;
assign w49095 = pi03932 & w3456;
assign w49096 = pi06549 & w3304;
assign w49097 = pi04339 & w3086;
assign w49098 = pi06787 & w3284;
assign w49099 = pi06286 & w3540;
assign w49100 = pi06185 & w3356;
assign w49101 = pi09688 & w3604;
assign w49102 = pi04380 & w3564;
assign w49103 = pi04161 & w3454;
assign w49104 = pi04243 & w3290;
assign w49105 = pi06266 & w3414;
assign w49106 = pi05830 & w3436;
assign w49107 = pi04317 & w3214;
assign w49108 = pi04426 & w3302;
assign w49109 = pi07987 & w3426;
assign w49110 = pi07952 & w3125;
assign w49111 = pi08120 & w3446;
assign w49112 = pi05983 & w3252;
assign w49113 = pi04498 & w3211;
assign w49114 = pi08352 & w3179;
assign w49115 = pi02208 & w3346;
assign w49116 = pi06099 & w3568;
assign w49117 = pi03239 & w3544;
assign w49118 = pi04352 & w3190;
assign w49119 = pi01635 & w3472;
assign w49120 = pi06482 & w3199;
assign w49121 = pi06885 & w3384;
assign w49122 = pi08235 & w3542;
assign w49123 = pi03275 & w3268;
assign w49124 = pi07408 & w3448;
assign w49125 = pi08320 & w3324;
assign w49126 = pi05967 & w3612;
assign w49127 = pi08156 & w3366;
assign w49128 = pi03209 & w3520;
assign w49129 = pi08339 & w3602;
assign w49130 = pi08365 & w3368;
assign w49131 = pi04116 & w3181;
assign w49132 = pi08399 & w3110;
assign w49133 = pi07175 & w3364;
assign w49134 = pi03673 & w3610;
assign w49135 = pi07867 & w3386;
assign w49136 = pi07128 & w3420;
assign w49137 = pi03183 & w3380;
assign w49138 = pi08221 & w3264;
assign w49139 = pi06930 & w3398;
assign w49140 = pi05789 & w3143;
assign w49141 = pi04465 & w3556;
assign w49142 = pi06059 & w3452;
assign w49143 = pi04491 & w3396;
assign w49144 = pi08333 & w3158;
assign w49145 = pi08169 & w3468;
assign w49146 = pi04446 & w3162;
assign w49147 = pi07438 & w3276;
assign w49148 = pi01642 & w3372;
assign w49149 = pi03619 & w3296;
assign w49150 = pi09794 & w3340;
assign w49151 = pi02061 & w3534;
assign w49152 = pi08300 & w3148;
assign w49153 = pi08215 & w3282;
assign w49154 = pi07107 & w3552;
assign w49155 = pi01578 & w3294;
assign w49156 = pi07833 & w3207;
assign w49157 = pi03494 & w3064;
assign w49158 = pi01493 & w3348;
assign w49159 = pi04452 & w3504;
assign w49160 = pi04102 & w3522;
assign w49161 = pi08195 & w3444;
assign w49162 = pi03401 & w3404;
assign w49163 = pi03713 & w3244;
assign w49164 = pi07217 & w3205;
assign w49165 = pi05934 & w3344;
assign w49166 = pi04440 & w3122;
assign w49167 = pi08431 & w3242;
assign w49168 = pi07512 & w3312;
assign w49169 = pi08134 & w3570;
assign w49170 = pi07453 & w3434;
assign w49171 = pi06119 & w3288;
assign w49172 = pi01719 & w3606;
assign w49173 = pi03872 & w3576;
assign w49174 = pi06322 & w3314;
assign w49175 = pi06380 & w3236;
assign w49176 = pi03879 & w3209;
assign w49177 = pi03349 & w3416;
assign w49178 = pi06826 & w3256;
assign w49179 = pi06086 & w3550;
assign w49180 = pi08425 & w3510;
assign w49181 = pi08346 & w3578;
assign w49182 = pi04472 & w3388;
assign w49183 = pi09614 & w3118;
assign w49184 = pi07244 & w3225;
assign w49185 = pi04069 & w3494;
assign w49186 = pi06839 & w3518;
assign w49187 = pi03456 & w3530;
assign w49188 = pi07305 & w3221;
assign w49189 = pi07387 & w3358;
assign w49190 = pi06400 & w3354;
assign w49191 = pi08018 & w3474;
assign w49192 = pi07741 & w3458;
assign w49193 = pi08268 & w3402;
assign w49194 = pi03356 & w3470;
assign w49195 = pi08150 & w3608;
assign w49196 = pi07927 & w3596;
assign w49197 = pi04027 & w3071;
assign w49198 = pi08070 & w3175;
assign w49199 = pi07204 & w3156;
assign w49200 = pi02794 & w3516;
assign w49201 = pi03975 & w3498;
assign w49202 = pi03527 & w3400;
assign w49203 = pi04413 & w3562;
assign w49204 = pi04371 & w3146;
assign w49205 = pi07780 & w3192;
assign w49206 = pi08326 & w3332;
assign w49207 = pi02373 & w3278;
assign w49208 = pi04263 & w3326;
assign w49209 = pi05740 & w3266;
assign w49210 = pi03990 & w3132;
assign w49211 = pi03749 & w3490;
assign w49212 = pi06159 & w3112;
assign w49213 = pi04420 & w3169;
assign w49214 = pi08418 & w3408;
assign w49215 = pi09686 & w3286;
assign w49216 = pi05684 & w3486;
assign w49217 = pi06800 & w3078;
assign w49218 = pi03658 & w3260;
assign w49219 = pi03488 & w3250;
assign w49220 = pi05869 & w3598;
assign w49221 = pi09767 & w3203;
assign w49222 = pi03409 & w3330;
assign w49223 = pi06073 & w3528;
assign w49224 = pi07120 & w3410;
assign w49225 = pi04063 & w3574;
assign w49226 = pi03373 & w3362;
assign w49227 = pi03550 & w3322;
assign w49228 = pi07654 & w3600;
assign w49229 = pi07819 & w3464;
assign w49230 = pi05954 & w3492;
assign w49231 = pi07673 & w3194;
assign w49232 = pi02223 & w3240;
assign w49233 = pi02379 & w3476;
assign w49234 = pi06336 & w3538;
assign w49235 = pi04386 & w3370;
assign w49236 = pi08037 & w3532;
assign w49237 = pi06177 & w3378;
assign w49238 = pi07230 & w3254;
assign w49239 = pi08313 & w3316;
assign w49240 = pi06366 & w3450;
assign w49241 = pi07807 & w3390;
assign w49242 = pi03690 & w3310;
assign w49243 = pi08208 & w3478;
assign w49244 = pi02361 & w3232;
assign w49245 = pi04459 & w3184;
assign w49246 = pi08386 & w3418;
assign w49247 = pi02229 & w3306;
assign w49248 = pi08392 & w3246;
assign w49249 = pi08287 & w3560;
assign w49250 = pi06917 & w3300;
assign w49251 = pi04358 & w3328;
assign w49252 = pi04345 & w3115;
assign w49253 = pi07016 & w3572;
assign w49254 = pi02202 & w3197;
assign w49255 = pi08261 & w3188;
assign w49256 = pi06581 & w3496;
assign w49257 = pi07961 & w3093;
assign w49258 = pi03762 & w3526;
assign w49259 = pi08082 & w3223;
assign w49260 = pi08373 & w3160;
assign w49261 = pi03573 & w3103;
assign w49262 = pi03793 & w3350;
assign w49263 = pi06865 & w3442;
assign w49264 = pi07427 & w3566;
assign w49265 = pi03625 & w3137;
assign w49266 = pi07354 & w3376;
assign w49267 = pi06151 & w3217;
assign w49268 = pi07473 & w3508;
assign w49269 = pi04155 & w3502;
assign w49270 = pi03997 & w3394;
assign w49271 = pi07888 & w3382;
assign w49272 = pi03153 & w3614;
assign w49273 = pi08242 & w3280;
assign w49274 = pi08274 & w3580;
assign w49275 = pi06601 & w3153;
assign w49276 = pi06963 & w3466;
assign w49277 = pi02444 & w3171;
assign w49278 = pi06970 & w3127;
assign w49279 = pi06038 & w3554;
assign w49280 = pi01859 & w3186;
assign w49281 = pi08182 & w3584;
assign w49282 = pi01611 & w3374;
assign w49283 = pi06003 & w3219;
assign w49284 = pi07793 & w3360;
assign w49285 = pi07591 & w3201;
assign w49286 = pi03612 & w3424;
assign w49287 = pi06219 & w3586;
assign w49288 = pi07683 & w3590;
assign w49289 = pi06904 & w3506;
assign w49290 = pi04399 & w3512;
assign w49291 = pi08228 & w3546;
assign w49292 = pi06528 & w3227;
assign w49293 = pi03632 & w3262;
assign w49294 = pi03591 & w3274;
assign w49295 = pi08405 & w3150;
assign w49296 = pi04433 & w3258;
assign w49297 = pi04511 & w3488;
assign w49298 = pi06564 & w3462;
assign w49299 = pi08248 & w3096;
assign w49300 = pi06138 & w3480;
assign w49301 = pi07559 & w3165;
assign w49302 = pi07492 & w3167;
assign w49303 = pi06506 & w3422;
assign w49304 = pi08281 & w3229;
assign w49305 = pi05809 & w3308;
assign w49306 = pi06989 & w3139;
assign w49307 = pi06688 & w3082;
assign w49308 = pi04504 & w3582;
assign w49309 = pi03945 & w3592;
assign w49310 = pi08054 & w3616;
assign w49311 = pi08410 & w3558;
assign w49312 = pi03223 & w3336;
assign w49313 = pi04290 & w3334;
assign w49314 = pi03640 & w3292;
assign w49315 = pi03606 & w3536;
assign w49316 = pi06943 & w3234;
assign w49317 = pi03723 & w3548;
assign w49318 = pi04486 & w3588;
assign w49319 = ~w49063 & ~w49064;
assign w49320 = ~w49065 & ~w49066;
assign w49321 = ~w49067 & ~w49068;
assign w49322 = ~w49069 & ~w49070;
assign w49323 = ~w49071 & ~w49072;
assign w49324 = ~w49073 & ~w49074;
assign w49325 = ~w49075 & ~w49076;
assign w49326 = ~w49077 & ~w49078;
assign w49327 = ~w49079 & ~w49080;
assign w49328 = ~w49081 & ~w49082;
assign w49329 = ~w49083 & ~w49084;
assign w49330 = ~w49085 & ~w49086;
assign w49331 = ~w49087 & ~w49088;
assign w49332 = ~w49089 & ~w49090;
assign w49333 = ~w49091 & ~w49092;
assign w49334 = ~w49093 & ~w49094;
assign w49335 = ~w49095 & ~w49096;
assign w49336 = ~w49097 & ~w49098;
assign w49337 = ~w49099 & ~w49100;
assign w49338 = ~w49101 & ~w49102;
assign w49339 = ~w49103 & ~w49104;
assign w49340 = ~w49105 & ~w49106;
assign w49341 = ~w49107 & ~w49108;
assign w49342 = ~w49109 & ~w49110;
assign w49343 = ~w49111 & ~w49112;
assign w49344 = ~w49113 & ~w49114;
assign w49345 = ~w49115 & ~w49116;
assign w49346 = ~w49117 & ~w49118;
assign w49347 = ~w49119 & ~w49120;
assign w49348 = ~w49121 & ~w49122;
assign w49349 = ~w49123 & ~w49124;
assign w49350 = ~w49125 & ~w49126;
assign w49351 = ~w49127 & ~w49128;
assign w49352 = ~w49129 & ~w49130;
assign w49353 = ~w49131 & ~w49132;
assign w49354 = ~w49133 & ~w49134;
assign w49355 = ~w49135 & ~w49136;
assign w49356 = ~w49137 & ~w49138;
assign w49357 = ~w49139 & ~w49140;
assign w49358 = ~w49141 & ~w49142;
assign w49359 = ~w49143 & ~w49144;
assign w49360 = ~w49145 & ~w49146;
assign w49361 = ~w49147 & ~w49148;
assign w49362 = ~w49149 & ~w49150;
assign w49363 = ~w49151 & ~w49152;
assign w49364 = ~w49153 & ~w49154;
assign w49365 = ~w49155 & ~w49156;
assign w49366 = ~w49157 & ~w49158;
assign w49367 = ~w49159 & ~w49160;
assign w49368 = ~w49161 & ~w49162;
assign w49369 = ~w49163 & ~w49164;
assign w49370 = ~w49165 & ~w49166;
assign w49371 = ~w49167 & ~w49168;
assign w49372 = ~w49169 & ~w49170;
assign w49373 = ~w49171 & ~w49172;
assign w49374 = ~w49173 & ~w49174;
assign w49375 = ~w49175 & ~w49176;
assign w49376 = ~w49177 & ~w49178;
assign w49377 = ~w49179 & ~w49180;
assign w49378 = ~w49181 & ~w49182;
assign w49379 = ~w49183 & ~w49184;
assign w49380 = ~w49185 & ~w49186;
assign w49381 = ~w49187 & ~w49188;
assign w49382 = ~w49189 & ~w49190;
assign w49383 = ~w49191 & ~w49192;
assign w49384 = ~w49193 & ~w49194;
assign w49385 = ~w49195 & ~w49196;
assign w49386 = ~w49197 & ~w49198;
assign w49387 = ~w49199 & ~w49200;
assign w49388 = ~w49201 & ~w49202;
assign w49389 = ~w49203 & ~w49204;
assign w49390 = ~w49205 & ~w49206;
assign w49391 = ~w49207 & ~w49208;
assign w49392 = ~w49209 & ~w49210;
assign w49393 = ~w49211 & ~w49212;
assign w49394 = ~w49213 & ~w49214;
assign w49395 = ~w49215 & ~w49216;
assign w49396 = ~w49217 & ~w49218;
assign w49397 = ~w49219 & ~w49220;
assign w49398 = ~w49221 & ~w49222;
assign w49399 = ~w49223 & ~w49224;
assign w49400 = ~w49225 & ~w49226;
assign w49401 = ~w49227 & ~w49228;
assign w49402 = ~w49229 & ~w49230;
assign w49403 = ~w49231 & ~w49232;
assign w49404 = ~w49233 & ~w49234;
assign w49405 = ~w49235 & ~w49236;
assign w49406 = ~w49237 & ~w49238;
assign w49407 = ~w49239 & ~w49240;
assign w49408 = ~w49241 & ~w49242;
assign w49409 = ~w49243 & ~w49244;
assign w49410 = ~w49245 & ~w49246;
assign w49411 = ~w49247 & ~w49248;
assign w49412 = ~w49249 & ~w49250;
assign w49413 = ~w49251 & ~w49252;
assign w49414 = ~w49253 & ~w49254;
assign w49415 = ~w49255 & ~w49256;
assign w49416 = ~w49257 & ~w49258;
assign w49417 = ~w49259 & ~w49260;
assign w49418 = ~w49261 & ~w49262;
assign w49419 = ~w49263 & ~w49264;
assign w49420 = ~w49265 & ~w49266;
assign w49421 = ~w49267 & ~w49268;
assign w49422 = ~w49269 & ~w49270;
assign w49423 = ~w49271 & ~w49272;
assign w49424 = ~w49273 & ~w49274;
assign w49425 = ~w49275 & ~w49276;
assign w49426 = ~w49277 & ~w49278;
assign w49427 = ~w49279 & ~w49280;
assign w49428 = ~w49281 & ~w49282;
assign w49429 = ~w49283 & ~w49284;
assign w49430 = ~w49285 & ~w49286;
assign w49431 = ~w49287 & ~w49288;
assign w49432 = ~w49289 & ~w49290;
assign w49433 = ~w49291 & ~w49292;
assign w49434 = ~w49293 & ~w49294;
assign w49435 = ~w49295 & ~w49296;
assign w49436 = ~w49297 & ~w49298;
assign w49437 = ~w49299 & ~w49300;
assign w49438 = ~w49301 & ~w49302;
assign w49439 = ~w49303 & ~w49304;
assign w49440 = ~w49305 & ~w49306;
assign w49441 = ~w49307 & ~w49308;
assign w49442 = ~w49309 & ~w49310;
assign w49443 = ~w49311 & ~w49312;
assign w49444 = ~w49313 & ~w49314;
assign w49445 = ~w49315 & ~w49316;
assign w49446 = ~w49317 & ~w49318;
assign w49447 = w49445 & w49446;
assign w49448 = w49443 & w49444;
assign w49449 = w49441 & w49442;
assign w49450 = w49439 & w49440;
assign w49451 = w49437 & w49438;
assign w49452 = w49435 & w49436;
assign w49453 = w49433 & w49434;
assign w49454 = w49431 & w49432;
assign w49455 = w49429 & w49430;
assign w49456 = w49427 & w49428;
assign w49457 = w49425 & w49426;
assign w49458 = w49423 & w49424;
assign w49459 = w49421 & w49422;
assign w49460 = w49419 & w49420;
assign w49461 = w49417 & w49418;
assign w49462 = w49415 & w49416;
assign w49463 = w49413 & w49414;
assign w49464 = w49411 & w49412;
assign w49465 = w49409 & w49410;
assign w49466 = w49407 & w49408;
assign w49467 = w49405 & w49406;
assign w49468 = w49403 & w49404;
assign w49469 = w49401 & w49402;
assign w49470 = w49399 & w49400;
assign w49471 = w49397 & w49398;
assign w49472 = w49395 & w49396;
assign w49473 = w49393 & w49394;
assign w49474 = w49391 & w49392;
assign w49475 = w49389 & w49390;
assign w49476 = w49387 & w49388;
assign w49477 = w49385 & w49386;
assign w49478 = w49383 & w49384;
assign w49479 = w49381 & w49382;
assign w49480 = w49379 & w49380;
assign w49481 = w49377 & w49378;
assign w49482 = w49375 & w49376;
assign w49483 = w49373 & w49374;
assign w49484 = w49371 & w49372;
assign w49485 = w49369 & w49370;
assign w49486 = w49367 & w49368;
assign w49487 = w49365 & w49366;
assign w49488 = w49363 & w49364;
assign w49489 = w49361 & w49362;
assign w49490 = w49359 & w49360;
assign w49491 = w49357 & w49358;
assign w49492 = w49355 & w49356;
assign w49493 = w49353 & w49354;
assign w49494 = w49351 & w49352;
assign w49495 = w49349 & w49350;
assign w49496 = w49347 & w49348;
assign w49497 = w49345 & w49346;
assign w49498 = w49343 & w49344;
assign w49499 = w49341 & w49342;
assign w49500 = w49339 & w49340;
assign w49501 = w49337 & w49338;
assign w49502 = w49335 & w49336;
assign w49503 = w49333 & w49334;
assign w49504 = w49331 & w49332;
assign w49505 = w49329 & w49330;
assign w49506 = w49327 & w49328;
assign w49507 = w49325 & w49326;
assign w49508 = w49323 & w49324;
assign w49509 = w49321 & w49322;
assign w49510 = w49319 & w49320;
assign w49511 = w49509 & w49510;
assign w49512 = w49507 & w49508;
assign w49513 = w49505 & w49506;
assign w49514 = w49503 & w49504;
assign w49515 = w49501 & w49502;
assign w49516 = w49499 & w49500;
assign w49517 = w49497 & w49498;
assign w49518 = w49495 & w49496;
assign w49519 = w49493 & w49494;
assign w49520 = w49491 & w49492;
assign w49521 = w49489 & w49490;
assign w49522 = w49487 & w49488;
assign w49523 = w49485 & w49486;
assign w49524 = w49483 & w49484;
assign w49525 = w49481 & w49482;
assign w49526 = w49479 & w49480;
assign w49527 = w49477 & w49478;
assign w49528 = w49475 & w49476;
assign w49529 = w49473 & w49474;
assign w49530 = w49471 & w49472;
assign w49531 = w49469 & w49470;
assign w49532 = w49467 & w49468;
assign w49533 = w49465 & w49466;
assign w49534 = w49463 & w49464;
assign w49535 = w49461 & w49462;
assign w49536 = w49459 & w49460;
assign w49537 = w49457 & w49458;
assign w49538 = w49455 & w49456;
assign w49539 = w49453 & w49454;
assign w49540 = w49451 & w49452;
assign w49541 = w49449 & w49450;
assign w49542 = w49447 & w49448;
assign w49543 = w49541 & w49542;
assign w49544 = w49539 & w49540;
assign w49545 = w49537 & w49538;
assign w49546 = w49535 & w49536;
assign w49547 = w49533 & w49534;
assign w49548 = w49531 & w49532;
assign w49549 = w49529 & w49530;
assign w49550 = w49527 & w49528;
assign w49551 = w49525 & w49526;
assign w49552 = w49523 & w49524;
assign w49553 = w49521 & w49522;
assign w49554 = w49519 & w49520;
assign w49555 = w49517 & w49518;
assign w49556 = w49515 & w49516;
assign w49557 = w49513 & w49514;
assign w49558 = w49511 & w49512;
assign w49559 = w49557 & w49558;
assign w49560 = w49555 & w49556;
assign w49561 = w49553 & w49554;
assign w49562 = w49551 & w49552;
assign w49563 = w49549 & w49550;
assign w49564 = w49547 & w49548;
assign w49565 = w49545 & w49546;
assign w49566 = w49543 & w49544;
assign w49567 = w49565 & w49566;
assign w49568 = w49563 & w49564;
assign w49569 = w49561 & w49562;
assign w49570 = w49559 & w49560;
assign w49571 = w49569 & w49570;
assign w49572 = w49567 & w49568;
assign w49573 = w49571 & w49572;
assign w49574 = ~pi10577 & ~w49573;
assign w49575 = pi09369 & w3229;
assign w49576 = pi02746 & w3582;
assign w49577 = pi04607 & w3330;
assign w49578 = pi04691 & w3262;
assign w49579 = pi09048 & w3590;
assign w49580 = pi08707 & w3496;
assign w49581 = pi02574 & w3480;
assign w49582 = pi09074 & w3458;
assign w49583 = pi09230 & w3440;
assign w49584 = pi04704 & w3260;
assign w49585 = pi09061 & w3171;
assign w49586 = pi04613 & w3530;
assign w49587 = pi08570 & w3217;
assign w49588 = pi04672 & w3424;
assign w49589 = pi04810 & w3394;
assign w49590 = pi08655 & w3392;
assign w49591 = pi04522 & w3306;
assign w49592 = pi08989 & w3508;
assign w49593 = pi09382 & w3342;
assign w49594 = pi09482 & w3246;
assign w49595 = pi02751 & w3396;
assign w49596 = pi08885 & w3135;
assign w49597 = pi04626 & w3064;
assign w49598 = pi02748 & w3211;
assign w49599 = pi08937 & w3620;
assign w49600 = pi04750 & w3350;
assign w49601 = pi09244 & w3366;
assign w49602 = pi09641 & w3370;
assign w49603 = pi04600 & w3404;
assign w49604 = pi08956 & w3358;
assign w49605 = pi08741 & w3186;
assign w49606 = pi02494 & w3460;
assign w49607 = pi08898 & w3156;
assign w49608 = pi08524 & w3219;
assign w49609 = pi08872 & w3410;
assign w49610 = pi08636 & w3236;
assign w49611 = pi09349 & w3188;
assign w49612 = pi09640 & w3564;
assign w49613 = pi08826 & w3127;
assign w49614 = pi04537 & w3346;
assign w49615 = pi02754 & w3588;
assign w49616 = pi08800 & w3300;
assign w49617 = pi09028 & w3374;
assign w49618 = pi08580 & w3378;
assign w49619 = pi04543 & w3520;
assign w49620 = pi09146 & w3125;
assign w49621 = pi08904 & w3205;
assign w49622 = pi04844 & w3428;
assign w49623 = pi08461 & w3143;
assign w49624 = pi08943 & w3272;
assign w49625 = pi09362 & w3580;
assign w49626 = pi09462 & w3160;
assign w49627 = pi09375 & w3560;
assign w49628 = pi09707 & w3326;
assign w49629 = pi09436 & w3578;
assign w49630 = pi08721 & w3082;
assign w49631 = pi04737 & w3490;
assign w49632 = pi01940 & w3482;
assign w49633 = pi09197 & w3175;
assign w49634 = pi09152 & w3093;
assign w49635 = pi08747 & w3284;
assign w49636 = pi01734 & w3266;
assign w49637 = pi09100 & w3464;
assign w49638 = pi08602 & w3414;
assign w49639 = pi09575 & w3122;
assign w49640 = pi08976 & w3276;
assign w49641 = pi04516 & w3614;
assign w49642 = pi04756 & w3576;
assign w49643 = pi09356 & w3402;
assign w49644 = pi09002 & w3312;
assign w49645 = pi08436 & w3486;
assign w49646 = pi02049 & w3232;
assign w49647 = pi09711 & w3290;
assign w49648 = pi08668 & w3129;
assign w49649 = pi01943 & w3538;
assign w49650 = pi09094 & w3390;
assign w49651 = pi09696 & w3214;
assign w49652 = pi09087 & w3360;
assign w49653 = pi08734 & w3514;
assign w49654 = pi08969 & w3566;
assign w49655 = pi09342 & w3318;
assign w49656 = pi04685 & w3137;
assign w49657 = pi09442 & w3179;
assign w49658 = pi01593 & w3418;
assign w49659 = pi09678 & w3190;
assign w49660 = pi08575 & w3112;
assign w49661 = pi04730 & w3548;
assign w49662 = pi09107 & w3207;
assign w49663 = pi09335 & w3096;
assign w49664 = pi04567 & w3500;
assign w49665 = pi08675 & w3199;
assign w49666 = pi05322 & w3550;
assign w49667 = pi09021 & w3372;
assign w49668 = pi08891 & w3364;
assign w49669 = pi04639 & w3400;
assign w49670 = pi01777 & w3568;
assign w49671 = pi08519 & w3252;
assign w49672 = pi04633 & w3534;
assign w49673 = pi04783 & w3456;
assign w49674 = pi04678 & w3296;
assign w49675 = pi09538 & w3556;
assign w49676 = pi09264 & w3173;
assign w49677 = pi09217 & w3446;
assign w49678 = pi04863 & w3502;
assign w49679 = pi09515 & w3510;
assign w49680 = pi05922 & w3492;
assign w49681 = pi08865 & w3552;
assign w49682 = pi09689 & w3086;
assign w49683 = pi08917 & w3225;
assign w49684 = pi04790 & w3592;
assign w49685 = pi09224 & w3570;
assign w49686 = pi08780 & w3384;
assign w49687 = pi08852 & w3340;
assign w49688 = pi04717 & w3310;
assign w49689 = pi04594 & w3362;
assign w49690 = pi04777 & w3348;
assign w49691 = pi09578 & w3258;
assign w49692 = pi09211 & w3606;
assign w49693 = pi09068 & w3476;
assign w49694 = pi09015 & w3201;
assign w49695 = pi09597 & w3169;
assign w49696 = pi09257 & w3468;
assign w49697 = pi04796 & w3498;
assign w49698 = pi09757 & w3452;
assign w49699 = pi04620 & w3250;
assign w49700 = pi04659 & w3274;
assign w49701 = pi08833 & w3139;
assign w49702 = pi08556 & w3288;
assign w49703 = pi04857 & w3181;
assign w49704 = pi08963 & w3448;
assign w49705 = pi05078 & w3242;
assign w49706 = pi09126 & w3382;
assign w49707 = pi08529 & w3554;
assign w49708 = pi04823 & w3118;
assign w49709 = pi08701 & w3462;
assign w49710 = pi09165 & w3426;
assign w49711 = pi08760 & w3256;
assign w49712 = pi09496 & w3150;
assign w49713 = pi09388 & w3148;
assign w49714 = pi09402 & w3316;
assign w49715 = pi04763 & w3209;
assign w49716 = pi09667 & w3115;
assign w49717 = pi03901 & w3177;
assign w49718 = pi08754 & w3078;
assign w49719 = pi09042 & w3194;
assign w49720 = pi09303 & w3282;
assign w49721 = pi09322 & w3542;
assign w49722 = pi08480 & w3248;
assign w49723 = pi09316 & w3546;
assign w49724 = pi09637 & w3618;
assign w49725 = pi09670 & w3328;
assign w49726 = pi02569 & w3110;
assign w49727 = pi02013 & w3268;
assign w49728 = pi04646 & w3322;
assign w49729 = pi09296 & w3478;
assign w49730 = pi09204 & w3223;
assign w49731 = pi09527 & w3388;
assign w49732 = pi08585 & w3356;
assign w49733 = pi09590 & w3302;
assign w49734 = pi09270 & w3584;
assign w49735 = pi04870 & w3454;
assign w49736 = pi04837 & w3494;
assign w49737 = pi08794 & w3506;
assign w49738 = pi09455 & w3368;
assign w49739 = pi09657 & w3146;
assign w49740 = pi08924 & w3472;
assign w49741 = pi09290 & w3320;
assign w49742 = pi04711 & w3610;
assign w49743 = pi04698 & w3292;
assign w49744 = pi08473 & w3436;
assign w49745 = pi09567 & w3162;
assign w49746 = pi09661 & w3484;
assign w49747 = pi02002 & w3470;
assign w49748 = pi09283 & w3444;
assign w49749 = pi08807 & w3398;
assign w49750 = pi04817 & w3071;
assign w49751 = pi09502 & w3558;
assign w49752 = pi08911 & w3254;
assign w49753 = pi04850 & w3522;
assign w49754 = pi08486 & w3598;
assign w49755 = pi02742 & w3488;
assign w49756 = pi09177 & w3474;
assign w49757 = pi05014 & w3504;
assign w49758 = pi08629 & w3450;
assign w49759 = pi08813 & w3234;
assign w49760 = pi09133 & w3352;
assign w49761 = pi09007 & w3165;
assign w49762 = pi08494 & w3604;
assign w49763 = pi08787 & w3432;
assign w49764 = pi09704 & w3334;
assign w49765 = pi08714 & w3153;
assign w49766 = pi04555 & w3336;
assign w49767 = pi08846 & w3572;
assign w49768 = pi09611 & w3562;
assign w49769 = pi01672 & w3308;
assign w49770 = pi09429 & w3602;
assign w49771 = pi04529 & w3380;
assign w49772 = pi07679 & w3528;
assign w49773 = pi08774 & w3442;
assign w49774 = pi09139 & w3596;
assign w49775 = pi08501 & w3344;
assign w49776 = pi04831 & w3574;
assign w49777 = pi09627 & w3512;
assign w49778 = pi04549 & w3197;
assign w49779 = pi08995 & w3167;
assign w49780 = pi09449 & w3438;
assign w49781 = pi08820 & w3466;
assign w49782 = pi08513 & w3612;
assign w49783 = pi08681 & w3422;
assign w49784 = pi09423 & w3158;
assign w49785 = pi09120 & w3386;
assign w49786 = pi08608 & w3540;
assign w49787 = pi09309 & w3264;
assign w49788 = pi04665 & w3536;
assign w49789 = pi02031 & w3544;
assign w49790 = pi08449 & w3240;
assign w49791 = pi02009 & w3416;
assign w49792 = pi09509 & w3408;
assign w49793 = pi08694 & w3304;
assign w49794 = pi04743 & w3526;
assign w49795 = pi08642 & w3298;
assign w49796 = pi04652 & w3103;
assign w49797 = pi09277 & w3106;
assign w49798 = pi09415 & w3332;
assign w49799 = pi09113 & w3270;
assign w49800 = pi08688 & w3227;
assign w49801 = pi08839 & w3406;
assign w49802 = pi09409 & w3324;
assign w49803 = pi08950 & w3376;
assign w49804 = pi09468 & w3524;
assign w49805 = pi09081 & w3192;
assign w49806 = pi09191 & w3616;
assign w49807 = pi09237 & w3608;
assign w49808 = pi08728 & w3278;
assign w49809 = pi08930 & w3221;
assign w49810 = pi09616 & w3412;
assign w49811 = pi08878 & w3420;
assign w49812 = pi09526 & w3184;
assign w49813 = pi09159 & w3238;
assign w49814 = pi09329 & w3280;
assign w49815 = pi09172 & w3516;
assign w49816 = pi08616 & w3314;
assign w49817 = pi09035 & w3600;
assign w49818 = pi08859 & w3286;
assign w49819 = pi09185 & w3532;
assign w49820 = pi09395 & w3294;
assign w49821 = pi09055 & w3430;
assign w49822 = pi04803 & w3132;
assign w49823 = pi08982 & w3434;
assign w49824 = pi08649 & w3354;
assign w49825 = pi09251 & w3594;
assign w49826 = pi08767 & w3518;
assign w49827 = pi05326 & w3586;
assign w49828 = pi04724 & w3244;
assign w49829 = pi08662 & w3203;
assign w49830 = pi04769 & w3338;
assign w49831 = ~w49575 & ~w49576;
assign w49832 = ~w49577 & ~w49578;
assign w49833 = ~w49579 & ~w49580;
assign w49834 = ~w49581 & ~w49582;
assign w49835 = ~w49583 & ~w49584;
assign w49836 = ~w49585 & ~w49586;
assign w49837 = ~w49587 & ~w49588;
assign w49838 = ~w49589 & ~w49590;
assign w49839 = ~w49591 & ~w49592;
assign w49840 = ~w49593 & ~w49594;
assign w49841 = ~w49595 & ~w49596;
assign w49842 = ~w49597 & ~w49598;
assign w49843 = ~w49599 & ~w49600;
assign w49844 = ~w49601 & ~w49602;
assign w49845 = ~w49603 & ~w49604;
assign w49846 = ~w49605 & ~w49606;
assign w49847 = ~w49607 & ~w49608;
assign w49848 = ~w49609 & ~w49610;
assign w49849 = ~w49611 & ~w49612;
assign w49850 = ~w49613 & ~w49614;
assign w49851 = ~w49615 & ~w49616;
assign w49852 = ~w49617 & ~w49618;
assign w49853 = ~w49619 & ~w49620;
assign w49854 = ~w49621 & ~w49622;
assign w49855 = ~w49623 & ~w49624;
assign w49856 = ~w49625 & ~w49626;
assign w49857 = ~w49627 & ~w49628;
assign w49858 = ~w49629 & ~w49630;
assign w49859 = ~w49631 & ~w49632;
assign w49860 = ~w49633 & ~w49634;
assign w49861 = ~w49635 & ~w49636;
assign w49862 = ~w49637 & ~w49638;
assign w49863 = ~w49639 & ~w49640;
assign w49864 = ~w49641 & ~w49642;
assign w49865 = ~w49643 & ~w49644;
assign w49866 = ~w49645 & ~w49646;
assign w49867 = ~w49647 & ~w49648;
assign w49868 = ~w49649 & ~w49650;
assign w49869 = ~w49651 & ~w49652;
assign w49870 = ~w49653 & ~w49654;
assign w49871 = ~w49655 & ~w49656;
assign w49872 = ~w49657 & ~w49658;
assign w49873 = ~w49659 & ~w49660;
assign w49874 = ~w49661 & ~w49662;
assign w49875 = ~w49663 & ~w49664;
assign w49876 = ~w49665 & ~w49666;
assign w49877 = ~w49667 & ~w49668;
assign w49878 = ~w49669 & ~w49670;
assign w49879 = ~w49671 & ~w49672;
assign w49880 = ~w49673 & ~w49674;
assign w49881 = ~w49675 & ~w49676;
assign w49882 = ~w49677 & ~w49678;
assign w49883 = ~w49679 & ~w49680;
assign w49884 = ~w49681 & ~w49682;
assign w49885 = ~w49683 & ~w49684;
assign w49886 = ~w49685 & ~w49686;
assign w49887 = ~w49687 & ~w49688;
assign w49888 = ~w49689 & ~w49690;
assign w49889 = ~w49691 & ~w49692;
assign w49890 = ~w49693 & ~w49694;
assign w49891 = ~w49695 & ~w49696;
assign w49892 = ~w49697 & ~w49698;
assign w49893 = ~w49699 & ~w49700;
assign w49894 = ~w49701 & ~w49702;
assign w49895 = ~w49703 & ~w49704;
assign w49896 = ~w49705 & ~w49706;
assign w49897 = ~w49707 & ~w49708;
assign w49898 = ~w49709 & ~w49710;
assign w49899 = ~w49711 & ~w49712;
assign w49900 = ~w49713 & ~w49714;
assign w49901 = ~w49715 & ~w49716;
assign w49902 = ~w49717 & ~w49718;
assign w49903 = ~w49719 & ~w49720;
assign w49904 = ~w49721 & ~w49722;
assign w49905 = ~w49723 & ~w49724;
assign w49906 = ~w49725 & ~w49726;
assign w49907 = ~w49727 & ~w49728;
assign w49908 = ~w49729 & ~w49730;
assign w49909 = ~w49731 & ~w49732;
assign w49910 = ~w49733 & ~w49734;
assign w49911 = ~w49735 & ~w49736;
assign w49912 = ~w49737 & ~w49738;
assign w49913 = ~w49739 & ~w49740;
assign w49914 = ~w49741 & ~w49742;
assign w49915 = ~w49743 & ~w49744;
assign w49916 = ~w49745 & ~w49746;
assign w49917 = ~w49747 & ~w49748;
assign w49918 = ~w49749 & ~w49750;
assign w49919 = ~w49751 & ~w49752;
assign w49920 = ~w49753 & ~w49754;
assign w49921 = ~w49755 & ~w49756;
assign w49922 = ~w49757 & ~w49758;
assign w49923 = ~w49759 & ~w49760;
assign w49924 = ~w49761 & ~w49762;
assign w49925 = ~w49763 & ~w49764;
assign w49926 = ~w49765 & ~w49766;
assign w49927 = ~w49767 & ~w49768;
assign w49928 = ~w49769 & ~w49770;
assign w49929 = ~w49771 & ~w49772;
assign w49930 = ~w49773 & ~w49774;
assign w49931 = ~w49775 & ~w49776;
assign w49932 = ~w49777 & ~w49778;
assign w49933 = ~w49779 & ~w49780;
assign w49934 = ~w49781 & ~w49782;
assign w49935 = ~w49783 & ~w49784;
assign w49936 = ~w49785 & ~w49786;
assign w49937 = ~w49787 & ~w49788;
assign w49938 = ~w49789 & ~w49790;
assign w49939 = ~w49791 & ~w49792;
assign w49940 = ~w49793 & ~w49794;
assign w49941 = ~w49795 & ~w49796;
assign w49942 = ~w49797 & ~w49798;
assign w49943 = ~w49799 & ~w49800;
assign w49944 = ~w49801 & ~w49802;
assign w49945 = ~w49803 & ~w49804;
assign w49946 = ~w49805 & ~w49806;
assign w49947 = ~w49807 & ~w49808;
assign w49948 = ~w49809 & ~w49810;
assign w49949 = ~w49811 & ~w49812;
assign w49950 = ~w49813 & ~w49814;
assign w49951 = ~w49815 & ~w49816;
assign w49952 = ~w49817 & ~w49818;
assign w49953 = ~w49819 & ~w49820;
assign w49954 = ~w49821 & ~w49822;
assign w49955 = ~w49823 & ~w49824;
assign w49956 = ~w49825 & ~w49826;
assign w49957 = ~w49827 & ~w49828;
assign w49958 = ~w49829 & ~w49830;
assign w49959 = w49957 & w49958;
assign w49960 = w49955 & w49956;
assign w49961 = w49953 & w49954;
assign w49962 = w49951 & w49952;
assign w49963 = w49949 & w49950;
assign w49964 = w49947 & w49948;
assign w49965 = w49945 & w49946;
assign w49966 = w49943 & w49944;
assign w49967 = w49941 & w49942;
assign w49968 = w49939 & w49940;
assign w49969 = w49937 & w49938;
assign w49970 = w49935 & w49936;
assign w49971 = w49933 & w49934;
assign w49972 = w49931 & w49932;
assign w49973 = w49929 & w49930;
assign w49974 = w49927 & w49928;
assign w49975 = w49925 & w49926;
assign w49976 = w49923 & w49924;
assign w49977 = w49921 & w49922;
assign w49978 = w49919 & w49920;
assign w49979 = w49917 & w49918;
assign w49980 = w49915 & w49916;
assign w49981 = w49913 & w49914;
assign w49982 = w49911 & w49912;
assign w49983 = w49909 & w49910;
assign w49984 = w49907 & w49908;
assign w49985 = w49905 & w49906;
assign w49986 = w49903 & w49904;
assign w49987 = w49901 & w49902;
assign w49988 = w49899 & w49900;
assign w49989 = w49897 & w49898;
assign w49990 = w49895 & w49896;
assign w49991 = w49893 & w49894;
assign w49992 = w49891 & w49892;
assign w49993 = w49889 & w49890;
assign w49994 = w49887 & w49888;
assign w49995 = w49885 & w49886;
assign w49996 = w49883 & w49884;
assign w49997 = w49881 & w49882;
assign w49998 = w49879 & w49880;
assign w49999 = w49877 & w49878;
assign w50000 = w49875 & w49876;
assign w50001 = w49873 & w49874;
assign w50002 = w49871 & w49872;
assign w50003 = w49869 & w49870;
assign w50004 = w49867 & w49868;
assign w50005 = w49865 & w49866;
assign w50006 = w49863 & w49864;
assign w50007 = w49861 & w49862;
assign w50008 = w49859 & w49860;
assign w50009 = w49857 & w49858;
assign w50010 = w49855 & w49856;
assign w50011 = w49853 & w49854;
assign w50012 = w49851 & w49852;
assign w50013 = w49849 & w49850;
assign w50014 = w49847 & w49848;
assign w50015 = w49845 & w49846;
assign w50016 = w49843 & w49844;
assign w50017 = w49841 & w49842;
assign w50018 = w49839 & w49840;
assign w50019 = w49837 & w49838;
assign w50020 = w49835 & w49836;
assign w50021 = w49833 & w49834;
assign w50022 = w49831 & w49832;
assign w50023 = w50021 & w50022;
assign w50024 = w50019 & w50020;
assign w50025 = w50017 & w50018;
assign w50026 = w50015 & w50016;
assign w50027 = w50013 & w50014;
assign w50028 = w50011 & w50012;
assign w50029 = w50009 & w50010;
assign w50030 = w50007 & w50008;
assign w50031 = w50005 & w50006;
assign w50032 = w50003 & w50004;
assign w50033 = w50001 & w50002;
assign w50034 = w49999 & w50000;
assign w50035 = w49997 & w49998;
assign w50036 = w49995 & w49996;
assign w50037 = w49993 & w49994;
assign w50038 = w49991 & w49992;
assign w50039 = w49989 & w49990;
assign w50040 = w49987 & w49988;
assign w50041 = w49985 & w49986;
assign w50042 = w49983 & w49984;
assign w50043 = w49981 & w49982;
assign w50044 = w49979 & w49980;
assign w50045 = w49977 & w49978;
assign w50046 = w49975 & w49976;
assign w50047 = w49973 & w49974;
assign w50048 = w49971 & w49972;
assign w50049 = w49969 & w49970;
assign w50050 = w49967 & w49968;
assign w50051 = w49965 & w49966;
assign w50052 = w49963 & w49964;
assign w50053 = w49961 & w49962;
assign w50054 = w49959 & w49960;
assign w50055 = w50053 & w50054;
assign w50056 = w50051 & w50052;
assign w50057 = w50049 & w50050;
assign w50058 = w50047 & w50048;
assign w50059 = w50045 & w50046;
assign w50060 = w50043 & w50044;
assign w50061 = w50041 & w50042;
assign w50062 = w50039 & w50040;
assign w50063 = w50037 & w50038;
assign w50064 = w50035 & w50036;
assign w50065 = w50033 & w50034;
assign w50066 = w50031 & w50032;
assign w50067 = w50029 & w50030;
assign w50068 = w50027 & w50028;
assign w50069 = w50025 & w50026;
assign w50070 = w50023 & w50024;
assign w50071 = w50069 & w50070;
assign w50072 = w50067 & w50068;
assign w50073 = w50065 & w50066;
assign w50074 = w50063 & w50064;
assign w50075 = w50061 & w50062;
assign w50076 = w50059 & w50060;
assign w50077 = w50057 & w50058;
assign w50078 = w50055 & w50056;
assign w50079 = w50077 & w50078;
assign w50080 = w50075 & w50076;
assign w50081 = w50073 & w50074;
assign w50082 = w50071 & w50072;
assign w50083 = w50081 & w50082;
assign w50084 = w50079 & w50080;
assign w50085 = w50083 & w50084;
assign w50086 = ~pi10577 & ~w50085;
assign w50087 = pi03670 & w3610;
assign w50088 = pi04419 & w3169;
assign w50089 = pi01855 & w3350;
assign w50090 = pi03748 & w3490;
assign w50091 = pi06334 & w3538;
assign w50092 = pi07866 & w3386;
assign w50093 = pi08069 & w3175;
assign w50094 = pi02138 & w3177;
assign w50095 = pi07596 & w3372;
assign w50096 = pi05805 & w3308;
assign w50097 = pi05696 & w3232;
assign w50098 = pi09594 & w3494;
assign w50099 = pi08332 & w3158;
assign w50100 = pi05867 & w3598;
assign w50101 = pi03514 & w3534;
assign w50102 = pi03605 & w3536;
assign w50103 = pi07424 & w3566;
assign w50104 = pi09790 & w3238;
assign w50105 = pi07804 & w3390;
assign w50106 = pi03526 & w3400;
assign w50107 = pi02156 & w3556;
assign w50108 = pi02133 & w3416;
assign w50109 = pi06084 & w3550;
assign w50110 = pi07682 & w3590;
assign w50111 = pi03618 & w3296;
assign w50112 = pi08345 & w3578;
assign w50113 = pi03215 & w3197;
assign w50114 = pi08207 & w3478;
assign w50115 = pi06432 & w3203;
assign w50116 = pi01982 & w3396;
assign w50117 = pi08162 & w3594;
assign w50118 = pi02068 & w3064;
assign w50119 = pi04241 & w3290;
assign w50120 = pi03408 & w3330;
assign w50121 = pi04115 & w3181;
assign w50122 = pi07173 & w3364;
assign w50123 = pi08155 & w3366;
assign w50124 = pi06176 & w3378;
assign w50125 = pi05887 & w3604;
assign w50126 = pi06300 & w3482;
assign w50127 = pi02110 & w3404;
assign w50128 = pi08391 & w3246;
assign w50129 = pi02245 & w3370;
assign w50130 = pi06961 & w3466;
assign w50131 = pi03355 & w3470;
assign w50132 = pi02298 & w3414;
assign w50133 = pi06460 & w3129;
assign w50134 = pi05953 & w3492;
assign w50135 = pi03878 & w3209;
assign w50136 = pi07450 & w3434;
assign w50137 = pi08254 & w3318;
assign w50138 = pi03657 & w3260;
assign w50139 = pi06799 & w3078;
assign w50140 = pi07264 & w3472;
assign w50141 = pi08280 & w3229;
assign w50142 = pi08201 & w3320;
assign w50143 = pi04062 & w3574;
assign w50144 = pi06734 & w3514;
assign w50145 = pi01646 & w3135;
assign w50146 = pi07405 & w3448;
assign w50147 = pi04445 & w3162;
assign w50148 = pi03182 & w3380;
assign w50149 = pi06505 & w3422;
assign w50150 = pi03711 & w3244;
assign w50151 = pi02184 & w3122;
assign w50152 = pi07349 & w3376;
assign w50153 = pi07556 & w3165;
assign w50154 = pi03973 & w3498;
assign w50155 = pi08417 & w3408;
assign w50156 = pi06097 & w3568;
assign w50157 = pi06000 & w3219;
assign w50158 = pi07924 & w3596;
assign w50159 = pi04510 & w3488;
assign w50160 = pi06884 & w3384;
assign w50161 = pi04497 & w3211;
assign w50162 = pi02205 & w3302;
assign w50163 = pi08293 & w3342;
assign w50164 = pi08099 & w3606;
assign w50165 = pi08319 & w3324;
assign w50166 = pi07885 & w3382;
assign w50167 = pi01688 & w3153;
assign w50168 = pi06929 & w3398;
assign w50169 = pi02368 & w3458;
assign w50170 = pi04471 & w3388;
assign w50171 = pi05736 & w3266;
assign w50172 = pi08372 & w3160;
assign w50173 = pi08052 & w3616;
assign w50174 = pi04351 & w3190;
assign w50175 = pi08325 & w3332;
assign w50176 = pi07845 & w3270;
assign w50177 = pi08168 & w3468;
assign w50178 = pi08424 & w3510;
assign w50179 = pi08181 & w3584;
assign w50180 = pi02021 & w3424;
assign w50181 = pi07731 & w3476;
assign w50182 = pi03912 & w3348;
assign w50183 = pi08175 & w3173;
assign w50184 = pi01696 & w3576;
assign w50185 = pi08430 & w3242;
assign w50186 = pi08398 & w3110;
assign w50187 = pi06838 & w3518;
assign w50188 = pi08129 & w3570;
assign w50189 = pi02020 & w3137;
assign w50190 = pi08359 & w3438;
assign w50191 = pi08214 & w3282;
assign w50192 = pi07616 & w3374;
assign w50193 = pi07998 & w3516;
assign w50194 = pi04432 & w3258;
assign w50195 = pi02236 & w3512;
assign w50196 = pi01706 & w3276;
assign w50197 = pi06631 & w3272;
assign w50198 = pi04075 & w3428;
assign w50199 = pi02242 & w3328;
assign w50200 = pi03944 & w3592;
assign w50201 = pi01991 & w3310;
assign w50202 = pi02776 & w3454;
assign w50203 = pi07470 & w3508;
assign w50204 = pi08079 & w3223;
assign w50205 = pi02173 & w3504;
assign w50206 = pi01897 & w3304;
assign w50207 = pi02203 & w3520;
assign w50208 = pi07509 & w3312;
assign w50209 = pi07015 & w3572;
assign w50210 = pi03222 & w3336;
assign w50211 = pi06412 & w3392;
assign w50212 = pi08188 & w3106;
assign w50213 = pi08385 & w3418;
assign w50214 = pi04154 & w3502;
assign w50215 = pi01636 & w3256;
assign w50216 = pi03589 & w3274;
assign w50217 = pi03931 & w3456;
assign w50218 = pi04041 & w3118;
assign w50219 = pi07830 & w3207;
assign w50220 = pi08234 & w3542;
assign w50221 = pi08227 & w3546;
assign w50222 = pi07126 & w3420;
assign w50223 = pi06399 & w3354;
assign w50224 = pi02300 & w3227;
assign w50225 = pi06987 & w3139;
assign w50226 = pi08412 & w3558;
assign w50227 = pi08149 & w3608;
assign w50228 = pi05682 & w3486;
assign w50229 = pi07818 & w3464;
assign w50230 = pi02347 & w3586;
assign w50231 = pi03722 & w3548;
assign w50232 = pi06321 & w3314;
assign w50233 = pi06968 & w3127;
assign w50234 = pi09736 & w3286;
assign w50235 = pi06157 & w3112;
assign w50236 = pi06055 & w3452;
assign w50237 = pi06864 & w3442;
assign w50238 = pi03996 & w3394;
assign w50239 = pi07203 & w3156;
assign w50240 = pi08013 & w3474;
assign w50241 = pi01629 & w3093;
assign w50242 = pi07489 & w3167;
assign w50243 = pi07328 & w3620;
assign w50244 = pi07249 & w3225;
assign w50245 = pi06708 & w3278;
assign w50246 = pi06942 & w3234;
assign w50247 = pi02445 & w3532;
assign w50248 = pi02080 & w3530;
assign w50249 = pi08338 & w3602;
assign w50250 = pi05826 & w3436;
assign w50251 = pi03272 & w3268;
assign w50252 = pi07779 & w3192;
assign w50253 = pi06377 & w3236;
assign w50254 = pi08286 & w3560;
assign w50255 = pi08122 & w3446;
assign w50256 = pi04364 & w3484;
assign w50257 = pi06072 & w3528;
assign w50258 = pi03487 & w3250;
assign w50259 = pi08404 & w3150;
assign w50260 = pi08267 & w3402;
assign w50261 = pi02520 & w3194;
assign w50262 = pi07718 & w3171;
assign w50263 = pi08364 & w3368;
assign w50264 = pi01808 & w3496;
assign w50265 = pi09671 & w3132;
assign w50266 = pi01784 & w3288;
assign w50267 = pi04101 & w3522;
assign w50268 = pi03631 & w3262;
assign w50269 = pi08299 & w3148;
assign w50270 = pi07385 & w3358;
assign w50271 = pi02039 & w3103;
assign w50272 = pi08194 & w3444;
assign w50273 = pi05724 & w3240;
assign w50274 = pi07000 & w3406;
assign w50275 = pi06786 & w3284;
assign w50276 = pi07106 & w3552;
assign w50277 = pi07229 & w3254;
assign w50278 = pi08260 & w3188;
assign w50279 = pi04289 & w3334;
assign w50280 = pi02010 & w3292;
assign w50281 = pi07296 & w3221;
assign w50282 = pi06183 & w3356;
assign w50283 = pi06150 & w3217;
assign w50284 = pi08312 & w3316;
assign w50285 = pi03262 & w3500;
assign w50286 = pi02125 & w3362;
assign w50287 = pi08273 & w3580;
assign w50288 = pi05933 & w3344;
assign w50289 = pi08351 & w3179;
assign w50290 = pi04458 & w3184;
assign w50291 = pi07216 & w3205;
assign w50292 = pi04484 & w3588;
assign w50293 = pi03163 & w3306;
assign w50294 = pi04406 & w3412;
assign w50295 = pi06480 & w3199;
assign w50296 = pi06916 & w3300;
assign w50297 = pi05981 & w3252;
assign w50298 = pi08247 & w3096;
assign w50299 = pi02237 & w3614;
assign w50300 = pi06385 & w3298;
assign w50301 = pi04026 & w3071;
assign w50302 = pi06754 & w3186;
assign w50303 = pi08377 & w3524;
assign w50304 = pi08220 & w3264;
assign w50305 = pi08306 & w3294;
assign w50306 = pi03548 & w3322;
assign w50307 = pi06202 & w3460;
assign w50308 = pi06890 & w3432;
assign w50309 = pi04338 & w3086;
assign w50310 = pi03189 & w3346;
assign w50311 = pi07946 & w3125;
assign w50312 = pi07026 & w3340;
assign w50313 = pi06903 & w3506;
assign w50314 = pi06563 & w3462;
assign w50315 = pi02562 & w3426;
assign w50316 = pi06367 & w3450;
assign w50317 = pi01622 & w3338;
assign w50318 = pi02222 & w3562;
assign w50319 = pi07697 & w3430;
assign w50320 = pi05847 & w3248;
assign w50321 = pi02364 & w3115;
assign w50322 = pi07119 & w3410;
assign w50323 = pi07905 & w3352;
assign w50324 = pi07651 & w3600;
assign w50325 = pi05785 & w3143;
assign w50326 = pi04315 & w3214;
assign w50327 = pi02259 & w3146;
assign w50328 = pi04261 & w3326;
assign w50329 = pi01731 & w3201;
assign w50330 = pi03761 & w3526;
assign w50331 = pi04392 & w3618;
assign w50332 = pi05966 & w3612;
assign w50333 = pi08241 & w3280;
assign w50334 = pi02094 & w3582;
assign w50335 = pi07792 & w3360;
assign w50336 = pi06137 & w3480;
assign w50337 = pi01516 & w3440;
assign w50338 = pi02311 & w3540;
assign w50339 = pi06035 & w3554;
assign w50340 = pi06695 & w3082;
assign w50341 = pi04378 & w3564;
assign w50342 = pi03237 & w3544;
assign w50343 = ~w50087 & ~w50088;
assign w50344 = ~w50089 & ~w50090;
assign w50345 = ~w50091 & ~w50092;
assign w50346 = ~w50093 & ~w50094;
assign w50347 = ~w50095 & ~w50096;
assign w50348 = ~w50097 & ~w50098;
assign w50349 = ~w50099 & ~w50100;
assign w50350 = ~w50101 & ~w50102;
assign w50351 = ~w50103 & ~w50104;
assign w50352 = ~w50105 & ~w50106;
assign w50353 = ~w50107 & ~w50108;
assign w50354 = ~w50109 & ~w50110;
assign w50355 = ~w50111 & ~w50112;
assign w50356 = ~w50113 & ~w50114;
assign w50357 = ~w50115 & ~w50116;
assign w50358 = ~w50117 & ~w50118;
assign w50359 = ~w50119 & ~w50120;
assign w50360 = ~w50121 & ~w50122;
assign w50361 = ~w50123 & ~w50124;
assign w50362 = ~w50125 & ~w50126;
assign w50363 = ~w50127 & ~w50128;
assign w50364 = ~w50129 & ~w50130;
assign w50365 = ~w50131 & ~w50132;
assign w50366 = ~w50133 & ~w50134;
assign w50367 = ~w50135 & ~w50136;
assign w50368 = ~w50137 & ~w50138;
assign w50369 = ~w50139 & ~w50140;
assign w50370 = ~w50141 & ~w50142;
assign w50371 = ~w50143 & ~w50144;
assign w50372 = ~w50145 & ~w50146;
assign w50373 = ~w50147 & ~w50148;
assign w50374 = ~w50149 & ~w50150;
assign w50375 = ~w50151 & ~w50152;
assign w50376 = ~w50153 & ~w50154;
assign w50377 = ~w50155 & ~w50156;
assign w50378 = ~w50157 & ~w50158;
assign w50379 = ~w50159 & ~w50160;
assign w50380 = ~w50161 & ~w50162;
assign w50381 = ~w50163 & ~w50164;
assign w50382 = ~w50165 & ~w50166;
assign w50383 = ~w50167 & ~w50168;
assign w50384 = ~w50169 & ~w50170;
assign w50385 = ~w50171 & ~w50172;
assign w50386 = ~w50173 & ~w50174;
assign w50387 = ~w50175 & ~w50176;
assign w50388 = ~w50177 & ~w50178;
assign w50389 = ~w50179 & ~w50180;
assign w50390 = ~w50181 & ~w50182;
assign w50391 = ~w50183 & ~w50184;
assign w50392 = ~w50185 & ~w50186;
assign w50393 = ~w50187 & ~w50188;
assign w50394 = ~w50189 & ~w50190;
assign w50395 = ~w50191 & ~w50192;
assign w50396 = ~w50193 & ~w50194;
assign w50397 = ~w50195 & ~w50196;
assign w50398 = ~w50197 & ~w50198;
assign w50399 = ~w50199 & ~w50200;
assign w50400 = ~w50201 & ~w50202;
assign w50401 = ~w50203 & ~w50204;
assign w50402 = ~w50205 & ~w50206;
assign w50403 = ~w50207 & ~w50208;
assign w50404 = ~w50209 & ~w50210;
assign w50405 = ~w50211 & ~w50212;
assign w50406 = ~w50213 & ~w50214;
assign w50407 = ~w50215 & ~w50216;
assign w50408 = ~w50217 & ~w50218;
assign w50409 = ~w50219 & ~w50220;
assign w50410 = ~w50221 & ~w50222;
assign w50411 = ~w50223 & ~w50224;
assign w50412 = ~w50225 & ~w50226;
assign w50413 = ~w50227 & ~w50228;
assign w50414 = ~w50229 & ~w50230;
assign w50415 = ~w50231 & ~w50232;
assign w50416 = ~w50233 & ~w50234;
assign w50417 = ~w50235 & ~w50236;
assign w50418 = ~w50237 & ~w50238;
assign w50419 = ~w50239 & ~w50240;
assign w50420 = ~w50241 & ~w50242;
assign w50421 = ~w50243 & ~w50244;
assign w50422 = ~w50245 & ~w50246;
assign w50423 = ~w50247 & ~w50248;
assign w50424 = ~w50249 & ~w50250;
assign w50425 = ~w50251 & ~w50252;
assign w50426 = ~w50253 & ~w50254;
assign w50427 = ~w50255 & ~w50256;
assign w50428 = ~w50257 & ~w50258;
assign w50429 = ~w50259 & ~w50260;
assign w50430 = ~w50261 & ~w50262;
assign w50431 = ~w50263 & ~w50264;
assign w50432 = ~w50265 & ~w50266;
assign w50433 = ~w50267 & ~w50268;
assign w50434 = ~w50269 & ~w50270;
assign w50435 = ~w50271 & ~w50272;
assign w50436 = ~w50273 & ~w50274;
assign w50437 = ~w50275 & ~w50276;
assign w50438 = ~w50277 & ~w50278;
assign w50439 = ~w50279 & ~w50280;
assign w50440 = ~w50281 & ~w50282;
assign w50441 = ~w50283 & ~w50284;
assign w50442 = ~w50285 & ~w50286;
assign w50443 = ~w50287 & ~w50288;
assign w50444 = ~w50289 & ~w50290;
assign w50445 = ~w50291 & ~w50292;
assign w50446 = ~w50293 & ~w50294;
assign w50447 = ~w50295 & ~w50296;
assign w50448 = ~w50297 & ~w50298;
assign w50449 = ~w50299 & ~w50300;
assign w50450 = ~w50301 & ~w50302;
assign w50451 = ~w50303 & ~w50304;
assign w50452 = ~w50305 & ~w50306;
assign w50453 = ~w50307 & ~w50308;
assign w50454 = ~w50309 & ~w50310;
assign w50455 = ~w50311 & ~w50312;
assign w50456 = ~w50313 & ~w50314;
assign w50457 = ~w50315 & ~w50316;
assign w50458 = ~w50317 & ~w50318;
assign w50459 = ~w50319 & ~w50320;
assign w50460 = ~w50321 & ~w50322;
assign w50461 = ~w50323 & ~w50324;
assign w50462 = ~w50325 & ~w50326;
assign w50463 = ~w50327 & ~w50328;
assign w50464 = ~w50329 & ~w50330;
assign w50465 = ~w50331 & ~w50332;
assign w50466 = ~w50333 & ~w50334;
assign w50467 = ~w50335 & ~w50336;
assign w50468 = ~w50337 & ~w50338;
assign w50469 = ~w50339 & ~w50340;
assign w50470 = ~w50341 & ~w50342;
assign w50471 = w50469 & w50470;
assign w50472 = w50467 & w50468;
assign w50473 = w50465 & w50466;
assign w50474 = w50463 & w50464;
assign w50475 = w50461 & w50462;
assign w50476 = w50459 & w50460;
assign w50477 = w50457 & w50458;
assign w50478 = w50455 & w50456;
assign w50479 = w50453 & w50454;
assign w50480 = w50451 & w50452;
assign w50481 = w50449 & w50450;
assign w50482 = w50447 & w50448;
assign w50483 = w50445 & w50446;
assign w50484 = w50443 & w50444;
assign w50485 = w50441 & w50442;
assign w50486 = w50439 & w50440;
assign w50487 = w50437 & w50438;
assign w50488 = w50435 & w50436;
assign w50489 = w50433 & w50434;
assign w50490 = w50431 & w50432;
assign w50491 = w50429 & w50430;
assign w50492 = w50427 & w50428;
assign w50493 = w50425 & w50426;
assign w50494 = w50423 & w50424;
assign w50495 = w50421 & w50422;
assign w50496 = w50419 & w50420;
assign w50497 = w50417 & w50418;
assign w50498 = w50415 & w50416;
assign w50499 = w50413 & w50414;
assign w50500 = w50411 & w50412;
assign w50501 = w50409 & w50410;
assign w50502 = w50407 & w50408;
assign w50503 = w50405 & w50406;
assign w50504 = w50403 & w50404;
assign w50505 = w50401 & w50402;
assign w50506 = w50399 & w50400;
assign w50507 = w50397 & w50398;
assign w50508 = w50395 & w50396;
assign w50509 = w50393 & w50394;
assign w50510 = w50391 & w50392;
assign w50511 = w50389 & w50390;
assign w50512 = w50387 & w50388;
assign w50513 = w50385 & w50386;
assign w50514 = w50383 & w50384;
assign w50515 = w50381 & w50382;
assign w50516 = w50379 & w50380;
assign w50517 = w50377 & w50378;
assign w50518 = w50375 & w50376;
assign w50519 = w50373 & w50374;
assign w50520 = w50371 & w50372;
assign w50521 = w50369 & w50370;
assign w50522 = w50367 & w50368;
assign w50523 = w50365 & w50366;
assign w50524 = w50363 & w50364;
assign w50525 = w50361 & w50362;
assign w50526 = w50359 & w50360;
assign w50527 = w50357 & w50358;
assign w50528 = w50355 & w50356;
assign w50529 = w50353 & w50354;
assign w50530 = w50351 & w50352;
assign w50531 = w50349 & w50350;
assign w50532 = w50347 & w50348;
assign w50533 = w50345 & w50346;
assign w50534 = w50343 & w50344;
assign w50535 = w50533 & w50534;
assign w50536 = w50531 & w50532;
assign w50537 = w50529 & w50530;
assign w50538 = w50527 & w50528;
assign w50539 = w50525 & w50526;
assign w50540 = w50523 & w50524;
assign w50541 = w50521 & w50522;
assign w50542 = w50519 & w50520;
assign w50543 = w50517 & w50518;
assign w50544 = w50515 & w50516;
assign w50545 = w50513 & w50514;
assign w50546 = w50511 & w50512;
assign w50547 = w50509 & w50510;
assign w50548 = w50507 & w50508;
assign w50549 = w50505 & w50506;
assign w50550 = w50503 & w50504;
assign w50551 = w50501 & w50502;
assign w50552 = w50499 & w50500;
assign w50553 = w50497 & w50498;
assign w50554 = w50495 & w50496;
assign w50555 = w50493 & w50494;
assign w50556 = w50491 & w50492;
assign w50557 = w50489 & w50490;
assign w50558 = w50487 & w50488;
assign w50559 = w50485 & w50486;
assign w50560 = w50483 & w50484;
assign w50561 = w50481 & w50482;
assign w50562 = w50479 & w50480;
assign w50563 = w50477 & w50478;
assign w50564 = w50475 & w50476;
assign w50565 = w50473 & w50474;
assign w50566 = w50471 & w50472;
assign w50567 = w50565 & w50566;
assign w50568 = w50563 & w50564;
assign w50569 = w50561 & w50562;
assign w50570 = w50559 & w50560;
assign w50571 = w50557 & w50558;
assign w50572 = w50555 & w50556;
assign w50573 = w50553 & w50554;
assign w50574 = w50551 & w50552;
assign w50575 = w50549 & w50550;
assign w50576 = w50547 & w50548;
assign w50577 = w50545 & w50546;
assign w50578 = w50543 & w50544;
assign w50579 = w50541 & w50542;
assign w50580 = w50539 & w50540;
assign w50581 = w50537 & w50538;
assign w50582 = w50535 & w50536;
assign w50583 = w50581 & w50582;
assign w50584 = w50579 & w50580;
assign w50585 = w50577 & w50578;
assign w50586 = w50575 & w50576;
assign w50587 = w50573 & w50574;
assign w50588 = w50571 & w50572;
assign w50589 = w50569 & w50570;
assign w50590 = w50567 & w50568;
assign w50591 = w50589 & w50590;
assign w50592 = w50587 & w50588;
assign w50593 = w50585 & w50586;
assign w50594 = w50583 & w50584;
assign w50595 = w50593 & w50594;
assign w50596 = w50591 & w50592;
assign w50597 = w50595 & w50596;
assign w50598 = ~pi10577 & ~w50597;
assign w50599 = pi08219 & w3264;
assign w50600 = pi02131 & w3096;
assign w50601 = pi07969 & w3238;
assign w50602 = pi04482 & w3588;
assign w50603 = pi02488 & w3612;
assign w50604 = pi07551 & w3165;
assign w50605 = pi07727 & w3476;
assign w50606 = pi06181 & w3356;
assign w50607 = pi02537 & w3590;
assign w50608 = pi06824 & w3256;
assign w50609 = pi01778 & w3078;
assign w50610 = pi02534 & w3254;
assign w50611 = pi06752 & w3186;
assign w50612 = pi03233 & w3544;
assign w50613 = pi06111 & w3288;
assign w50614 = pi08383 & w3418;
assign w50615 = pi03629 & w3262;
assign w50616 = pi07613 & w3374;
assign w50617 = pi03603 & w3536;
assign w50618 = pi01689 & w3434;
assign w50619 = pi01829 & w3606;
assign w50620 = pi03883 & w3338;
assign w50621 = pi07940 & w3125;
assign w50622 = pi04060 & w3574;
assign w50623 = pi04375 & w3564;
assign w50624 = pi06595 & w3153;
assign w50625 = pi08154 & w3366;
assign w50626 = pi06155 & w3112;
assign w50627 = pi05881 & w3604;
assign w50628 = pi06359 & w3450;
assign w50629 = pi04336 & w3086;
assign w50630 = pi03213 & w3197;
assign w50631 = pi06575 & w3496;
assign w50632 = pi06683 & w3082;
assign w50633 = pi08291 & w3342;
assign w50634 = pi04362 & w3484;
assign w50635 = pi06882 & w3384;
assign w50636 = pi07693 & w3430;
assign w50637 = pi04256 & w3326;
assign w50638 = pi02040 & w3103;
assign w50639 = pi06083 & w3550;
assign w50640 = pi03353 & w3470;
assign w50641 = pi08193 & w3444;
assign w50642 = pi03161 & w3306;
assign w50643 = pi06212 & w3586;
assign w50644 = pi07326 & w3620;
assign w50645 = pi08240 & w3280;
assign w50646 = pi04349 & w3190;
assign w50647 = pi08127 & w3570;
assign w50648 = pi03688 & w3310;
assign w50649 = pi03480 & w3250;
assign w50650 = pi06901 & w3506;
assign w50651 = pi02025 & w3448;
assign w50652 = pi07239 & w3225;
assign w50653 = pi07996 & w3516;
assign w50654 = pi06031 & w3554;
assign w50655 = pi07778 & w3192;
assign w50656 = pi06994 & w3406;
assign w50657 = pi05694 & w3232;
assign w50658 = pi04411 & w3562;
assign w50659 = pi04023 & w3071;
assign w50660 = pi01720 & w3580;
assign w50661 = pi07843 & w3270;
assign w50662 = pi03988 & w3132;
assign w50663 = pi04037 & w3118;
assign w50664 = pi03655 & w3260;
assign w50665 = pi03910 & w3348;
assign w50666 = pi03508 & w3534;
assign w50667 = pi06928 & w3398;
assign w50668 = pi06473 & w3199;
assign w50669 = pi03399 & w3404;
assign w50670 = pi03260 & w3500;
assign w50671 = pi06915 & w3300;
assign w50672 = pi03759 & w3526;
assign w50673 = pi08206 & w3478;
assign w50674 = pi03347 & w3416;
assign w50675 = pi07899 & w3352;
assign w50676 = pi08357 & w3438;
assign w50677 = pi04237 & w3290;
assign w50678 = pi03784 & w3350;
assign w50679 = pi06521 & w3227;
assign w50680 = pi06200 & w3460;
assign w50681 = pi04404 & w3412;
assign w50682 = pi01597 & w3148;
assign w50683 = pi08343 & w3578;
assign w50684 = pi07008 & w3572;
assign w50685 = pi04067 & w3494;
assign w50686 = pi02286 & w3596;
assign w50687 = pi02310 & w3552;
assign w50688 = pi07505 & w3312;
assign w50689 = pi07339 & w3272;
assign w50690 = pi07436 & w3276;
assign w50691 = pi08075 & w3223;
assign w50692 = pi03268 & w3268;
assign w50693 = pi06091 & w3568;
assign w50694 = pi01661 & w3560;
assign w50695 = pi06981 & w3139;
assign w50696 = pi06835 & w3518;
assign w50697 = pi03636 & w3292;
assign w50698 = pi07140 & w3135;
assign w50699 = pi04097 & w3522;
assign w50700 = pi07379 & w3358;
assign w50701 = pi09542 & w3344;
assign w50702 = pi07799 & w3390;
assign w50703 = pi08369 & w3160;
assign w50704 = pi08180 & w3584;
assign w50705 = pi04430 & w3258;
assign w50706 = pi08336 & w3602;
assign w50707 = pi06967 & w3127;
assign w50708 = pi07982 & w3426;
assign w50709 = pi02425 & w3382;
assign w50710 = pi05823 & w3436;
assign w50711 = pi07858 & w3386;
assign w50712 = pi08114 & w3446;
assign w50713 = pi03746 & w3490;
assign w50714 = pi03187 & w3346;
assign w50715 = pi05676 & w3486;
assign w50716 = pi09755 & w3378;
assign w50717 = pi08147 & w3608;
assign w50718 = pi03994 & w3394;
assign w50719 = pi06561 & w3462;
assign w50720 = pi07817 & w3464;
assign w50721 = pi07169 & w3364;
assign w50722 = pi04489 & w3396;
assign w50723 = pi02450 & w3150;
assign w50724 = pi01533 & w3332;
assign w50725 = pi06889 & w3432;
assign w50726 = pi07214 & w3205;
assign w50727 = pi08278 & w3229;
assign w50728 = pi07712 & w3171;
assign w50729 = pi07201 & w3156;
assign w50730 = pi06384 & w3298;
assign w50731 = pi04152 & w3502;
assign w50732 = pi07294 & w3221;
assign w50733 = pi04397 & w3512;
assign w50734 = pi06050 & w3452;
assign w50735 = pi04389 & w3618;
assign w50736 = pi01789 & w3284;
assign w50737 = pi03545 & w3322;
assign w50738 = pi07593 & w3372;
assign w50739 = pi06071 & w3528;
assign w50740 = pi03969 & w3498;
assign w50741 = pi01535 & w3188;
assign w50742 = pi04113 & w3181;
assign w50743 = pi03610 & w3424;
assign w50744 = pi08252 & w3318;
assign w50745 = pi06279 & w3540;
assign w50746 = pi08317 & w3324;
assign w50747 = pi08411 & w3558;
assign w50748 = pi07791 & w3360;
assign w50749 = pi04469 & w3388;
assign w50750 = pi03585 & w3274;
assign w50751 = pi08212 & w3282;
assign w50752 = pi08186 & w3106;
assign w50753 = pi06941 & w3234;
assign w50754 = pi06457 & w3129;
assign w50755 = pi02196 & w3242;
assign w50756 = pi07738 & w3458;
assign w50757 = pi01569 & w3316;
assign w50758 = pi06955 & w3466;
assign w50759 = pi03367 & w3362;
assign w50760 = pi03452 & w3530;
assign w50761 = pi04508 & w3488;
assign w50762 = pi04456 & w3184;
assign w50763 = pi07665 & w3194;
assign w50764 = pi03220 & w3336;
assign w50765 = pi04437 & w3122;
assign w50766 = pi09699 & w3508;
assign w50767 = pi03876 & w3209;
assign w50768 = pi03406 & w3330;
assign w50769 = pi07347 & w3376;
assign w50770 = pi03180 & w3380;
assign w50771 = pi02460 & w3246;
assign w50772 = pi05997 & w3219;
assign w50773 = pi05780 & w3143;
assign w50774 = pi06258 & w3414;
assign w50775 = pi03623 & w3137;
assign w50776 = pi06374 & w3236;
assign w50777 = pi03492 & w3064;
assign w50778 = pi03720 & w3548;
assign w50779 = pi06503 & w3422;
assign w50780 = pi08422 & w3510;
assign w50781 = pi09548 & w3203;
assign w50782 = pi02159 & w3408;
assign w50783 = pi03668 & w3610;
assign w50784 = pi07580 & w3201;
assign w50785 = pi03524 & w3400;
assign w50786 = pi06319 & w3314;
assign w50787 = pi05801 & w3308;
assign w50788 = pi08035 & w3532;
assign w50789 = pi01852 & w3420;
assign w50790 = pi06861 & w3442;
assign w50791 = pi04284 & w3334;
assign w50792 = pi03942 & w3592;
assign w50793 = pi06130 & w3480;
assign w50794 = pi08067 & w3175;
assign w50795 = pi06145 & w3217;
assign w50796 = pi03148 & w3614;
assign w50797 = pi04310 & w3214;
assign w50798 = pi04073 & w3428;
assign w50799 = pi05734 & w3266;
assign w50800 = pi08160 & w3594;
assign w50801 = pi06733 & w3514;
assign w50802 = pi08167 & w3468;
assign w50803 = pi07486 & w3167;
assign w50804 = pi08173 & w3173;
assign w50805 = pi06410 & w3392;
assign w50806 = pi08199 & w3320;
assign w50807 = pi07114 & w3410;
assign w50808 = pi08048 & w3616;
assign w50809 = pi02637 & w3474;
assign w50810 = pi02602 & w3368;
assign w50811 = pi08349 & w3179;
assign w50812 = pi05952 & w3492;
assign w50813 = pi02419 & w3252;
assign w50814 = pi04451 & w3504;
assign w50815 = pi04159 & w3454;
assign w50816 = pi07261 & w3472;
assign w50817 = pi01887 & w3482;
assign w50818 = pi04495 & w3211;
assign w50819 = pi03870 & w3576;
assign w50820 = pi04443 & w3162;
assign w50821 = pi04502 & w3582;
assign w50822 = pi09734 & w3286;
assign w50823 = pi09751 & w3456;
assign w50824 = pi06397 & w3354;
assign w50825 = pi05842 & w3248;
assign w50826 = pi07021 & w3340;
assign w50827 = pi08330 & w3158;
assign w50828 = pi04424 & w3302;
assign w50829 = pi08265 & w3402;
assign w50830 = pi01621 & w3093;
assign w50831 = pi08225 & w3546;
assign w50832 = pi06332 & w3538;
assign w50833 = pi04356 & w3328;
assign w50834 = pi04463 & w3556;
assign w50835 = pi05860 & w3598;
assign w50836 = pi03707 & w3244;
assign w50837 = pi02536 & w3524;
assign w50838 = pi08397 & w3110;
assign w50839 = pi02279 & w3542;
assign w50840 = pi07827 & w3207;
assign w50841 = pi04343 & w3115;
assign w50842 = pi04369 & w3146;
assign w50843 = pi06540 & w3304;
assign w50844 = pi04476 & w3177;
assign w50845 = pi06707 & w3278;
assign w50846 = pi08139 & w3440;
assign w50847 = pi07420 & w3566;
assign w50848 = pi04384 & w3370;
assign w50849 = pi04417 & w3169;
assign w50850 = pi03616 & w3296;
assign w50851 = pi08304 & w3294;
assign w50852 = pi03201 & w3520;
assign w50853 = pi05721 & w3240;
assign w50854 = pi09576 & w3600;
assign w50855 = ~w50599 & ~w50600;
assign w50856 = ~w50601 & ~w50602;
assign w50857 = ~w50603 & ~w50604;
assign w50858 = ~w50605 & ~w50606;
assign w50859 = ~w50607 & ~w50608;
assign w50860 = ~w50609 & ~w50610;
assign w50861 = ~w50611 & ~w50612;
assign w50862 = ~w50613 & ~w50614;
assign w50863 = ~w50615 & ~w50616;
assign w50864 = ~w50617 & ~w50618;
assign w50865 = ~w50619 & ~w50620;
assign w50866 = ~w50621 & ~w50622;
assign w50867 = ~w50623 & ~w50624;
assign w50868 = ~w50625 & ~w50626;
assign w50869 = ~w50627 & ~w50628;
assign w50870 = ~w50629 & ~w50630;
assign w50871 = ~w50631 & ~w50632;
assign w50872 = ~w50633 & ~w50634;
assign w50873 = ~w50635 & ~w50636;
assign w50874 = ~w50637 & ~w50638;
assign w50875 = ~w50639 & ~w50640;
assign w50876 = ~w50641 & ~w50642;
assign w50877 = ~w50643 & ~w50644;
assign w50878 = ~w50645 & ~w50646;
assign w50879 = ~w50647 & ~w50648;
assign w50880 = ~w50649 & ~w50650;
assign w50881 = ~w50651 & ~w50652;
assign w50882 = ~w50653 & ~w50654;
assign w50883 = ~w50655 & ~w50656;
assign w50884 = ~w50657 & ~w50658;
assign w50885 = ~w50659 & ~w50660;
assign w50886 = ~w50661 & ~w50662;
assign w50887 = ~w50663 & ~w50664;
assign w50888 = ~w50665 & ~w50666;
assign w50889 = ~w50667 & ~w50668;
assign w50890 = ~w50669 & ~w50670;
assign w50891 = ~w50671 & ~w50672;
assign w50892 = ~w50673 & ~w50674;
assign w50893 = ~w50675 & ~w50676;
assign w50894 = ~w50677 & ~w50678;
assign w50895 = ~w50679 & ~w50680;
assign w50896 = ~w50681 & ~w50682;
assign w50897 = ~w50683 & ~w50684;
assign w50898 = ~w50685 & ~w50686;
assign w50899 = ~w50687 & ~w50688;
assign w50900 = ~w50689 & ~w50690;
assign w50901 = ~w50691 & ~w50692;
assign w50902 = ~w50693 & ~w50694;
assign w50903 = ~w50695 & ~w50696;
assign w50904 = ~w50697 & ~w50698;
assign w50905 = ~w50699 & ~w50700;
assign w50906 = ~w50701 & ~w50702;
assign w50907 = ~w50703 & ~w50704;
assign w50908 = ~w50705 & ~w50706;
assign w50909 = ~w50707 & ~w50708;
assign w50910 = ~w50709 & ~w50710;
assign w50911 = ~w50711 & ~w50712;
assign w50912 = ~w50713 & ~w50714;
assign w50913 = ~w50715 & ~w50716;
assign w50914 = ~w50717 & ~w50718;
assign w50915 = ~w50719 & ~w50720;
assign w50916 = ~w50721 & ~w50722;
assign w50917 = ~w50723 & ~w50724;
assign w50918 = ~w50725 & ~w50726;
assign w50919 = ~w50727 & ~w50728;
assign w50920 = ~w50729 & ~w50730;
assign w50921 = ~w50731 & ~w50732;
assign w50922 = ~w50733 & ~w50734;
assign w50923 = ~w50735 & ~w50736;
assign w50924 = ~w50737 & ~w50738;
assign w50925 = ~w50739 & ~w50740;
assign w50926 = ~w50741 & ~w50742;
assign w50927 = ~w50743 & ~w50744;
assign w50928 = ~w50745 & ~w50746;
assign w50929 = ~w50747 & ~w50748;
assign w50930 = ~w50749 & ~w50750;
assign w50931 = ~w50751 & ~w50752;
assign w50932 = ~w50753 & ~w50754;
assign w50933 = ~w50755 & ~w50756;
assign w50934 = ~w50757 & ~w50758;
assign w50935 = ~w50759 & ~w50760;
assign w50936 = ~w50761 & ~w50762;
assign w50937 = ~w50763 & ~w50764;
assign w50938 = ~w50765 & ~w50766;
assign w50939 = ~w50767 & ~w50768;
assign w50940 = ~w50769 & ~w50770;
assign w50941 = ~w50771 & ~w50772;
assign w50942 = ~w50773 & ~w50774;
assign w50943 = ~w50775 & ~w50776;
assign w50944 = ~w50777 & ~w50778;
assign w50945 = ~w50779 & ~w50780;
assign w50946 = ~w50781 & ~w50782;
assign w50947 = ~w50783 & ~w50784;
assign w50948 = ~w50785 & ~w50786;
assign w50949 = ~w50787 & ~w50788;
assign w50950 = ~w50789 & ~w50790;
assign w50951 = ~w50791 & ~w50792;
assign w50952 = ~w50793 & ~w50794;
assign w50953 = ~w50795 & ~w50796;
assign w50954 = ~w50797 & ~w50798;
assign w50955 = ~w50799 & ~w50800;
assign w50956 = ~w50801 & ~w50802;
assign w50957 = ~w50803 & ~w50804;
assign w50958 = ~w50805 & ~w50806;
assign w50959 = ~w50807 & ~w50808;
assign w50960 = ~w50809 & ~w50810;
assign w50961 = ~w50811 & ~w50812;
assign w50962 = ~w50813 & ~w50814;
assign w50963 = ~w50815 & ~w50816;
assign w50964 = ~w50817 & ~w50818;
assign w50965 = ~w50819 & ~w50820;
assign w50966 = ~w50821 & ~w50822;
assign w50967 = ~w50823 & ~w50824;
assign w50968 = ~w50825 & ~w50826;
assign w50969 = ~w50827 & ~w50828;
assign w50970 = ~w50829 & ~w50830;
assign w50971 = ~w50831 & ~w50832;
assign w50972 = ~w50833 & ~w50834;
assign w50973 = ~w50835 & ~w50836;
assign w50974 = ~w50837 & ~w50838;
assign w50975 = ~w50839 & ~w50840;
assign w50976 = ~w50841 & ~w50842;
assign w50977 = ~w50843 & ~w50844;
assign w50978 = ~w50845 & ~w50846;
assign w50979 = ~w50847 & ~w50848;
assign w50980 = ~w50849 & ~w50850;
assign w50981 = ~w50851 & ~w50852;
assign w50982 = ~w50853 & ~w50854;
assign w50983 = w50981 & w50982;
assign w50984 = w50979 & w50980;
assign w50985 = w50977 & w50978;
assign w50986 = w50975 & w50976;
assign w50987 = w50973 & w50974;
assign w50988 = w50971 & w50972;
assign w50989 = w50969 & w50970;
assign w50990 = w50967 & w50968;
assign w50991 = w50965 & w50966;
assign w50992 = w50963 & w50964;
assign w50993 = w50961 & w50962;
assign w50994 = w50959 & w50960;
assign w50995 = w50957 & w50958;
assign w50996 = w50955 & w50956;
assign w50997 = w50953 & w50954;
assign w50998 = w50951 & w50952;
assign w50999 = w50949 & w50950;
assign w51000 = w50947 & w50948;
assign w51001 = w50945 & w50946;
assign w51002 = w50943 & w50944;
assign w51003 = w50941 & w50942;
assign w51004 = w50939 & w50940;
assign w51005 = w50937 & w50938;
assign w51006 = w50935 & w50936;
assign w51007 = w50933 & w50934;
assign w51008 = w50931 & w50932;
assign w51009 = w50929 & w50930;
assign w51010 = w50927 & w50928;
assign w51011 = w50925 & w50926;
assign w51012 = w50923 & w50924;
assign w51013 = w50921 & w50922;
assign w51014 = w50919 & w50920;
assign w51015 = w50917 & w50918;
assign w51016 = w50915 & w50916;
assign w51017 = w50913 & w50914;
assign w51018 = w50911 & w50912;
assign w51019 = w50909 & w50910;
assign w51020 = w50907 & w50908;
assign w51021 = w50905 & w50906;
assign w51022 = w50903 & w50904;
assign w51023 = w50901 & w50902;
assign w51024 = w50899 & w50900;
assign w51025 = w50897 & w50898;
assign w51026 = w50895 & w50896;
assign w51027 = w50893 & w50894;
assign w51028 = w50891 & w50892;
assign w51029 = w50889 & w50890;
assign w51030 = w50887 & w50888;
assign w51031 = w50885 & w50886;
assign w51032 = w50883 & w50884;
assign w51033 = w50881 & w50882;
assign w51034 = w50879 & w50880;
assign w51035 = w50877 & w50878;
assign w51036 = w50875 & w50876;
assign w51037 = w50873 & w50874;
assign w51038 = w50871 & w50872;
assign w51039 = w50869 & w50870;
assign w51040 = w50867 & w50868;
assign w51041 = w50865 & w50866;
assign w51042 = w50863 & w50864;
assign w51043 = w50861 & w50862;
assign w51044 = w50859 & w50860;
assign w51045 = w50857 & w50858;
assign w51046 = w50855 & w50856;
assign w51047 = w51045 & w51046;
assign w51048 = w51043 & w51044;
assign w51049 = w51041 & w51042;
assign w51050 = w51039 & w51040;
assign w51051 = w51037 & w51038;
assign w51052 = w51035 & w51036;
assign w51053 = w51033 & w51034;
assign w51054 = w51031 & w51032;
assign w51055 = w51029 & w51030;
assign w51056 = w51027 & w51028;
assign w51057 = w51025 & w51026;
assign w51058 = w51023 & w51024;
assign w51059 = w51021 & w51022;
assign w51060 = w51019 & w51020;
assign w51061 = w51017 & w51018;
assign w51062 = w51015 & w51016;
assign w51063 = w51013 & w51014;
assign w51064 = w51011 & w51012;
assign w51065 = w51009 & w51010;
assign w51066 = w51007 & w51008;
assign w51067 = w51005 & w51006;
assign w51068 = w51003 & w51004;
assign w51069 = w51001 & w51002;
assign w51070 = w50999 & w51000;
assign w51071 = w50997 & w50998;
assign w51072 = w50995 & w50996;
assign w51073 = w50993 & w50994;
assign w51074 = w50991 & w50992;
assign w51075 = w50989 & w50990;
assign w51076 = w50987 & w50988;
assign w51077 = w50985 & w50986;
assign w51078 = w50983 & w50984;
assign w51079 = w51077 & w51078;
assign w51080 = w51075 & w51076;
assign w51081 = w51073 & w51074;
assign w51082 = w51071 & w51072;
assign w51083 = w51069 & w51070;
assign w51084 = w51067 & w51068;
assign w51085 = w51065 & w51066;
assign w51086 = w51063 & w51064;
assign w51087 = w51061 & w51062;
assign w51088 = w51059 & w51060;
assign w51089 = w51057 & w51058;
assign w51090 = w51055 & w51056;
assign w51091 = w51053 & w51054;
assign w51092 = w51051 & w51052;
assign w51093 = w51049 & w51050;
assign w51094 = w51047 & w51048;
assign w51095 = w51093 & w51094;
assign w51096 = w51091 & w51092;
assign w51097 = w51089 & w51090;
assign w51098 = w51087 & w51088;
assign w51099 = w51085 & w51086;
assign w51100 = w51083 & w51084;
assign w51101 = w51081 & w51082;
assign w51102 = w51079 & w51080;
assign w51103 = w51101 & w51102;
assign w51104 = w51099 & w51100;
assign w51105 = w51097 & w51098;
assign w51106 = w51095 & w51096;
assign w51107 = w51105 & w51106;
assign w51108 = w51103 & w51104;
assign w51109 = w51107 & w51108;
assign w51110 = ~pi10577 & ~w51109;
assign w51111 = pi09368 & w3229;
assign w51112 = pi09086 & w3360;
assign w51113 = pi05006 & w3162;
assign w51114 = pi04822 & w3118;
assign w51115 = pi09132 & w3352;
assign w51116 = pi05000 & w3122;
assign w51117 = pi04776 & w3348;
assign w51118 = pi09216 & w3446;
assign w51119 = pi08845 & w3572;
assign w51120 = pi08485 & w3598;
assign w51121 = pi05033 & w3388;
assign w51122 = pi09408 & w3324;
assign w51123 = pi04690 & w3262;
assign w51124 = pi08923 & w3472;
assign w51125 = pi04684 & w3137;
assign w51126 = pi08949 & w3376;
assign w51127 = pi09302 & w3282;
assign w51128 = pi08825 & w3127;
assign w51129 = pi08806 & w3398;
assign w51130 = pi09269 & w3584;
assign w51131 = pi09441 & w3179;
assign w51132 = pi02037 & w3336;
assign w51133 = pi09488 & w3110;
assign w51134 = pi05013 & w3504;
assign w51135 = pi04795 & w3498;
assign w51136 = pi02477 & w3586;
assign w51137 = pi09328 & w3280;
assign w51138 = pi04789 & w3592;
assign w51139 = pi08601 & w3414;
assign w51140 = pi08812 & w3234;
assign w51141 = pi09047 & w3590;
assign w51142 = pi04749 & w3350;
assign w51143 = pi09435 & w3578;
assign w51144 = pi01568 & w3422;
assign w51145 = pi04560 & w3544;
assign w51146 = pi04935 & w3146;
assign w51147 = pi05027 & w3556;
assign w51148 = pi09414 & w3332;
assign w51149 = pi09125 & w3382;
assign w51150 = pi08759 & w3256;
assign w51151 = pi08753 & w3078;
assign w51152 = pi09448 & w3438;
assign w51153 = pi04566 & w3500;
assign w51154 = pi09145 & w3125;
assign w51155 = pi09348 & w3188;
assign w51156 = pi08448 & w3240;
assign w51157 = pi09355 & w3402;
assign w51158 = pi09073 & w3458;
assign w51159 = pi04954 & w3618;
assign w51160 = pi04619 & w3250;
assign w51161 = pi04703 & w3260;
assign w51162 = pi04824 & w3153;
assign w51163 = pi01559 & w3227;
assign w51164 = pi05020 & w3184;
assign w51165 = pi08733 & w3514;
assign w51166 = pi04645 & w3322;
assign w51167 = pi04836 & w3494;
assign w51168 = pi04987 & w3302;
assign w51169 = pi09099 & w3464;
assign w51170 = pi04638 & w3400;
assign w51171 = pi05072 & w3488;
assign w51172 = pi08942 & w3272;
assign w51173 = pi09138 & w3596;
assign w51174 = pi08623 & w3538;
assign w51175 = pi09308 & w3264;
assign w51176 = pi04521 & w3306;
assign w51177 = pi04980 & w3169;
assign w51178 = pi07269 & w3554;
assign w51179 = pi09041 & w3194;
assign w51180 = pi09374 & w3560;
assign w51181 = pi05046 & w3588;
assign w51182 = pi09334 & w3096;
assign w51183 = pi04974 & w3562;
assign w51184 = pi04716 & w3310;
assign w51185 = pi08574 & w3112;
assign w51186 = pi09011 & w3165;
assign w51187 = pi09747 & w3474;
assign w51188 = pi05472 & w3540;
assign w51189 = pi04729 & w3548;
assign w51190 = pi05059 & w3211;
assign w51191 = pi09295 & w3478;
assign w51192 = pi02429 & w3510;
assign w51193 = pi08864 & w3552;
assign w51194 = pi04869 & w3454;
assign w51195 = pi09341 & w3318;
assign w51196 = pi04593 & w3362;
assign w51197 = pi08442 & w3232;
assign w51198 = pi09475 & w3418;
assign w51199 = pi04856 & w3181;
assign w51200 = pi09151 & w3093;
assign w51201 = pi09060 & w3171;
assign w51202 = pi09508 & w3408;
assign w51203 = pi09401 & w3316;
assign w51204 = pi08766 & w3518;
assign w51205 = pi04528 & w3380;
assign w51206 = pi04802 & w3132;
assign w51207 = pi05174 & w3288;
assign w51208 = pi01537 & w3462;
assign w51209 = pi08727 & w3278;
assign w51210 = pi09428 & w3602;
assign w51211 = pi04736 & w3490;
assign w51212 = pi09223 & w3570;
assign w51213 = pi08916 & w3225;
assign w51214 = pi09001 & w3312;
assign w51215 = pi09093 & w3390;
assign w51216 = pi04889 & w3334;
assign w51217 = pi08435 & w3486;
assign w51218 = pi04576 & w3197;
assign w51219 = pi08890 & w3364;
assign w51220 = pi04941 & w3564;
assign w51221 = pi01922 & w3384;
assign w51222 = pi01698 & w3392;
assign w51223 = pi09263 & w3173;
assign w51224 = pi04755 & w3576;
assign w51225 = pi04849 & w3522;
assign w51226 = pi08569 & w3217;
assign w51227 = pi09256 & w3468;
assign w51228 = pi08871 & w3410;
assign w51229 = pi02598 & w3550;
assign w51230 = pi08877 & w3420;
assign w51231 = pi04697 & w3292;
assign w51232 = pi09171 & w3516;
assign w51233 = pi08858 & w3286;
assign w51234 = pi04544 & w3520;
assign w51235 = pi09361 & w3580;
assign w51236 = pi09454 & w3368;
assign w51237 = pi09321 & w3542;
assign w51238 = pi08472 & w3436;
assign w51239 = pi08579 & w3378;
assign w51240 = pi09387 & w3148;
assign w51241 = pi08746 & w3284;
assign w51242 = pi09210 & w3606;
assign w51243 = pi08962 & w3448;
assign w51244 = pi01590 & w3129;
assign w51245 = pi08500 & w3344;
assign w51246 = pi08460 & w3143;
assign w51247 = pi04723 & w3244;
assign w51248 = pi08929 & w3221;
assign w51249 = pi09184 & w3532;
assign w51250 = pi08590 & w3460;
assign w51251 = pi09381 & w3342;
assign w51252 = pi01510 & w3236;
assign w51253 = pi09394 & w3294;
assign w51254 = pi09027 & w3374;
assign w51255 = pi09494 & w3150;
assign w51256 = pi04993 & w3258;
assign w51257 = pi08936 & w3620;
assign w51258 = pi04843 & w3428;
assign w51259 = pi05053 & w3396;
assign w51260 = pi09158 & w3238;
assign w51261 = pi08838 & w3406;
assign w51262 = pi04625 & w3064;
assign w51263 = pi09164 & w3426;
assign w51264 = pi01572 & w3558;
assign w51265 = pi04742 & w3526;
assign w51266 = pi01885 & w3314;
assign w51267 = pi08478 & w3248;
assign w51268 = pi04536 & w3346;
assign w51269 = pi08981 & w3434;
assign w51270 = pi08550 & w3568;
assign w51271 = pi09250 & w3594;
assign w51272 = pi04816 & w3071;
assign w51273 = pi09236 & w3608;
assign w51274 = pi01539 & w3604;
assign w51275 = pi02963 & w3470;
assign w51276 = pi09080 & w3192;
assign w51277 = pi08851 & w3340;
assign w51278 = pi01834 & w3298;
assign w51279 = pi04651 & w3103;
assign w51280 = pi04928 & w3484;
assign w51281 = pi09034 & w3600;
assign w51282 = pi08740 & w3186;
assign w51283 = pi08799 & w3300;
assign w51284 = pi01694 & w3203;
assign w51285 = pi09243 & w3366;
assign w51286 = pi04915 & w3190;
assign w51287 = pi04967 & w3412;
assign w51288 = pi08994 & w3167;
assign w51289 = pi08988 & w3508;
assign w51290 = pi04909 & w3115;
assign w51291 = pi04599 & w3404;
assign w51292 = pi04876 & w3290;
assign w51293 = pi09481 & w3246;
assign w51294 = pi08457 & w3266;
assign w51295 = pi08467 & w3308;
assign w51296 = pi05040 & w3177;
assign w51297 = pi04862 & w3502;
assign w51298 = pi09461 & w3160;
assign w51299 = pi04922 & w3328;
assign w51300 = pi08910 & w3254;
assign w51301 = pi08612 & w3482;
assign w51302 = pi04573 & w3268;
assign w51303 = pi09020 & w3372;
assign w51304 = pi09422 & w3158;
assign w51305 = pi09276 & w3106;
assign w51306 = pi04710 & w3610;
assign w51307 = pi08955 & w3358;
assign w51308 = pi09067 & w3476;
assign w51309 = pi08512 & w3612;
assign w51310 = pi09783 & w3496;
assign w51311 = pi08534 & w3452;
assign w51312 = pi04883 & w3326;
assign w51313 = pi01591 & w3199;
assign w51314 = pi08773 & w3442;
assign w51315 = pi04580 & w3416;
assign w51316 = pi08884 & w3135;
assign w51317 = pi09289 & w3320;
assign w51318 = pi04782 & w3456;
assign w51319 = pi04902 & w3086;
assign w51320 = pi04768 & w3338;
assign w51321 = pi09229 & w3440;
assign w51322 = pi08518 & w3252;
assign w51323 = pi08720 & w3082;
assign w51324 = pi09282 & w3444;
assign w51325 = pi08903 & w3205;
assign w51326 = pi08832 & w3139;
assign w51327 = pi04961 & w3512;
assign w51328 = pi08897 & w3156;
assign w51329 = pi08561 & w3480;
assign w51330 = pi04606 & w3330;
assign w51331 = pi04612 & w3530;
assign w51332 = pi09106 & w3207;
assign w51333 = pi08793 & w3506;
assign w51334 = pi08975 & w3276;
assign w51335 = pi01735 & w3354;
assign w51336 = pi09014 & w3201;
assign w51337 = pi02482 & w3175;
assign w51338 = pi09315 & w3546;
assign w51339 = pi04632 & w3534;
assign w51340 = pi05066 & w3582;
assign w51341 = pi04515 & w3614;
assign w51342 = pi09203 & w3223;
assign w51343 = pi04896 & w3214;
assign w51344 = pi01553 & w3304;
assign w51345 = pi09190 & w3616;
assign w51346 = pi08539 & w3528;
assign w51347 = pi05366 & w3356;
assign w51348 = pi04762 & w3209;
assign w51349 = pi09112 & w3270;
assign w51350 = pi04677 & w3296;
assign w51351 = pi09054 & w3430;
assign w51352 = pi08968 & w3566;
assign w51353 = pi08506 & w3492;
assign w51354 = pi05077 & w3242;
assign w51355 = pi08819 & w3466;
assign w51356 = pi01908 & w3450;
assign w51357 = pi08523 & w3219;
assign w51358 = pi04948 & w3370;
assign w51359 = pi04809 & w3394;
assign w51360 = pi09467 & w3524;
assign w51361 = pi04664 & w3536;
assign w51362 = pi09119 & w3386;
assign w51363 = pi04658 & w3274;
assign w51364 = pi04830 & w3574;
assign w51365 = pi04671 & w3424;
assign w51366 = pi08786 & w3432;
assign w51367 = ~w51111 & ~w51112;
assign w51368 = ~w51113 & ~w51114;
assign w51369 = ~w51115 & ~w51116;
assign w51370 = ~w51117 & ~w51118;
assign w51371 = ~w51119 & ~w51120;
assign w51372 = ~w51121 & ~w51122;
assign w51373 = ~w51123 & ~w51124;
assign w51374 = ~w51125 & ~w51126;
assign w51375 = ~w51127 & ~w51128;
assign w51376 = ~w51129 & ~w51130;
assign w51377 = ~w51131 & ~w51132;
assign w51378 = ~w51133 & ~w51134;
assign w51379 = ~w51135 & ~w51136;
assign w51380 = ~w51137 & ~w51138;
assign w51381 = ~w51139 & ~w51140;
assign w51382 = ~w51141 & ~w51142;
assign w51383 = ~w51143 & ~w51144;
assign w51384 = ~w51145 & ~w51146;
assign w51385 = ~w51147 & ~w51148;
assign w51386 = ~w51149 & ~w51150;
assign w51387 = ~w51151 & ~w51152;
assign w51388 = ~w51153 & ~w51154;
assign w51389 = ~w51155 & ~w51156;
assign w51390 = ~w51157 & ~w51158;
assign w51391 = ~w51159 & ~w51160;
assign w51392 = ~w51161 & ~w51162;
assign w51393 = ~w51163 & ~w51164;
assign w51394 = ~w51165 & ~w51166;
assign w51395 = ~w51167 & ~w51168;
assign w51396 = ~w51169 & ~w51170;
assign w51397 = ~w51171 & ~w51172;
assign w51398 = ~w51173 & ~w51174;
assign w51399 = ~w51175 & ~w51176;
assign w51400 = ~w51177 & ~w51178;
assign w51401 = ~w51179 & ~w51180;
assign w51402 = ~w51181 & ~w51182;
assign w51403 = ~w51183 & ~w51184;
assign w51404 = ~w51185 & ~w51186;
assign w51405 = ~w51187 & ~w51188;
assign w51406 = ~w51189 & ~w51190;
assign w51407 = ~w51191 & ~w51192;
assign w51408 = ~w51193 & ~w51194;
assign w51409 = ~w51195 & ~w51196;
assign w51410 = ~w51197 & ~w51198;
assign w51411 = ~w51199 & ~w51200;
assign w51412 = ~w51201 & ~w51202;
assign w51413 = ~w51203 & ~w51204;
assign w51414 = ~w51205 & ~w51206;
assign w51415 = ~w51207 & ~w51208;
assign w51416 = ~w51209 & ~w51210;
assign w51417 = ~w51211 & ~w51212;
assign w51418 = ~w51213 & ~w51214;
assign w51419 = ~w51215 & ~w51216;
assign w51420 = ~w51217 & ~w51218;
assign w51421 = ~w51219 & ~w51220;
assign w51422 = ~w51221 & ~w51222;
assign w51423 = ~w51223 & ~w51224;
assign w51424 = ~w51225 & ~w51226;
assign w51425 = ~w51227 & ~w51228;
assign w51426 = ~w51229 & ~w51230;
assign w51427 = ~w51231 & ~w51232;
assign w51428 = ~w51233 & ~w51234;
assign w51429 = ~w51235 & ~w51236;
assign w51430 = ~w51237 & ~w51238;
assign w51431 = ~w51239 & ~w51240;
assign w51432 = ~w51241 & ~w51242;
assign w51433 = ~w51243 & ~w51244;
assign w51434 = ~w51245 & ~w51246;
assign w51435 = ~w51247 & ~w51248;
assign w51436 = ~w51249 & ~w51250;
assign w51437 = ~w51251 & ~w51252;
assign w51438 = ~w51253 & ~w51254;
assign w51439 = ~w51255 & ~w51256;
assign w51440 = ~w51257 & ~w51258;
assign w51441 = ~w51259 & ~w51260;
assign w51442 = ~w51261 & ~w51262;
assign w51443 = ~w51263 & ~w51264;
assign w51444 = ~w51265 & ~w51266;
assign w51445 = ~w51267 & ~w51268;
assign w51446 = ~w51269 & ~w51270;
assign w51447 = ~w51271 & ~w51272;
assign w51448 = ~w51273 & ~w51274;
assign w51449 = ~w51275 & ~w51276;
assign w51450 = ~w51277 & ~w51278;
assign w51451 = ~w51279 & ~w51280;
assign w51452 = ~w51281 & ~w51282;
assign w51453 = ~w51283 & ~w51284;
assign w51454 = ~w51285 & ~w51286;
assign w51455 = ~w51287 & ~w51288;
assign w51456 = ~w51289 & ~w51290;
assign w51457 = ~w51291 & ~w51292;
assign w51458 = ~w51293 & ~w51294;
assign w51459 = ~w51295 & ~w51296;
assign w51460 = ~w51297 & ~w51298;
assign w51461 = ~w51299 & ~w51300;
assign w51462 = ~w51301 & ~w51302;
assign w51463 = ~w51303 & ~w51304;
assign w51464 = ~w51305 & ~w51306;
assign w51465 = ~w51307 & ~w51308;
assign w51466 = ~w51309 & ~w51310;
assign w51467 = ~w51311 & ~w51312;
assign w51468 = ~w51313 & ~w51314;
assign w51469 = ~w51315 & ~w51316;
assign w51470 = ~w51317 & ~w51318;
assign w51471 = ~w51319 & ~w51320;
assign w51472 = ~w51321 & ~w51322;
assign w51473 = ~w51323 & ~w51324;
assign w51474 = ~w51325 & ~w51326;
assign w51475 = ~w51327 & ~w51328;
assign w51476 = ~w51329 & ~w51330;
assign w51477 = ~w51331 & ~w51332;
assign w51478 = ~w51333 & ~w51334;
assign w51479 = ~w51335 & ~w51336;
assign w51480 = ~w51337 & ~w51338;
assign w51481 = ~w51339 & ~w51340;
assign w51482 = ~w51341 & ~w51342;
assign w51483 = ~w51343 & ~w51344;
assign w51484 = ~w51345 & ~w51346;
assign w51485 = ~w51347 & ~w51348;
assign w51486 = ~w51349 & ~w51350;
assign w51487 = ~w51351 & ~w51352;
assign w51488 = ~w51353 & ~w51354;
assign w51489 = ~w51355 & ~w51356;
assign w51490 = ~w51357 & ~w51358;
assign w51491 = ~w51359 & ~w51360;
assign w51492 = ~w51361 & ~w51362;
assign w51493 = ~w51363 & ~w51364;
assign w51494 = ~w51365 & ~w51366;
assign w51495 = w51493 & w51494;
assign w51496 = w51491 & w51492;
assign w51497 = w51489 & w51490;
assign w51498 = w51487 & w51488;
assign w51499 = w51485 & w51486;
assign w51500 = w51483 & w51484;
assign w51501 = w51481 & w51482;
assign w51502 = w51479 & w51480;
assign w51503 = w51477 & w51478;
assign w51504 = w51475 & w51476;
assign w51505 = w51473 & w51474;
assign w51506 = w51471 & w51472;
assign w51507 = w51469 & w51470;
assign w51508 = w51467 & w51468;
assign w51509 = w51465 & w51466;
assign w51510 = w51463 & w51464;
assign w51511 = w51461 & w51462;
assign w51512 = w51459 & w51460;
assign w51513 = w51457 & w51458;
assign w51514 = w51455 & w51456;
assign w51515 = w51453 & w51454;
assign w51516 = w51451 & w51452;
assign w51517 = w51449 & w51450;
assign w51518 = w51447 & w51448;
assign w51519 = w51445 & w51446;
assign w51520 = w51443 & w51444;
assign w51521 = w51441 & w51442;
assign w51522 = w51439 & w51440;
assign w51523 = w51437 & w51438;
assign w51524 = w51435 & w51436;
assign w51525 = w51433 & w51434;
assign w51526 = w51431 & w51432;
assign w51527 = w51429 & w51430;
assign w51528 = w51427 & w51428;
assign w51529 = w51425 & w51426;
assign w51530 = w51423 & w51424;
assign w51531 = w51421 & w51422;
assign w51532 = w51419 & w51420;
assign w51533 = w51417 & w51418;
assign w51534 = w51415 & w51416;
assign w51535 = w51413 & w51414;
assign w51536 = w51411 & w51412;
assign w51537 = w51409 & w51410;
assign w51538 = w51407 & w51408;
assign w51539 = w51405 & w51406;
assign w51540 = w51403 & w51404;
assign w51541 = w51401 & w51402;
assign w51542 = w51399 & w51400;
assign w51543 = w51397 & w51398;
assign w51544 = w51395 & w51396;
assign w51545 = w51393 & w51394;
assign w51546 = w51391 & w51392;
assign w51547 = w51389 & w51390;
assign w51548 = w51387 & w51388;
assign w51549 = w51385 & w51386;
assign w51550 = w51383 & w51384;
assign w51551 = w51381 & w51382;
assign w51552 = w51379 & w51380;
assign w51553 = w51377 & w51378;
assign w51554 = w51375 & w51376;
assign w51555 = w51373 & w51374;
assign w51556 = w51371 & w51372;
assign w51557 = w51369 & w51370;
assign w51558 = w51367 & w51368;
assign w51559 = w51557 & w51558;
assign w51560 = w51555 & w51556;
assign w51561 = w51553 & w51554;
assign w51562 = w51551 & w51552;
assign w51563 = w51549 & w51550;
assign w51564 = w51547 & w51548;
assign w51565 = w51545 & w51546;
assign w51566 = w51543 & w51544;
assign w51567 = w51541 & w51542;
assign w51568 = w51539 & w51540;
assign w51569 = w51537 & w51538;
assign w51570 = w51535 & w51536;
assign w51571 = w51533 & w51534;
assign w51572 = w51531 & w51532;
assign w51573 = w51529 & w51530;
assign w51574 = w51527 & w51528;
assign w51575 = w51525 & w51526;
assign w51576 = w51523 & w51524;
assign w51577 = w51521 & w51522;
assign w51578 = w51519 & w51520;
assign w51579 = w51517 & w51518;
assign w51580 = w51515 & w51516;
assign w51581 = w51513 & w51514;
assign w51582 = w51511 & w51512;
assign w51583 = w51509 & w51510;
assign w51584 = w51507 & w51508;
assign w51585 = w51505 & w51506;
assign w51586 = w51503 & w51504;
assign w51587 = w51501 & w51502;
assign w51588 = w51499 & w51500;
assign w51589 = w51497 & w51498;
assign w51590 = w51495 & w51496;
assign w51591 = w51589 & w51590;
assign w51592 = w51587 & w51588;
assign w51593 = w51585 & w51586;
assign w51594 = w51583 & w51584;
assign w51595 = w51581 & w51582;
assign w51596 = w51579 & w51580;
assign w51597 = w51577 & w51578;
assign w51598 = w51575 & w51576;
assign w51599 = w51573 & w51574;
assign w51600 = w51571 & w51572;
assign w51601 = w51569 & w51570;
assign w51602 = w51567 & w51568;
assign w51603 = w51565 & w51566;
assign w51604 = w51563 & w51564;
assign w51605 = w51561 & w51562;
assign w51606 = w51559 & w51560;
assign w51607 = w51605 & w51606;
assign w51608 = w51603 & w51604;
assign w51609 = w51601 & w51602;
assign w51610 = w51599 & w51600;
assign w51611 = w51597 & w51598;
assign w51612 = w51595 & w51596;
assign w51613 = w51593 & w51594;
assign w51614 = w51591 & w51592;
assign w51615 = w51613 & w51614;
assign w51616 = w51611 & w51612;
assign w51617 = w51609 & w51610;
assign w51618 = w51607 & w51608;
assign w51619 = w51617 & w51618;
assign w51620 = w51615 & w51616;
assign w51621 = w51619 & w51620;
assign w51622 = ~pi10577 & ~w51621;
assign w51623 = pi04719 & w3310;
assign w51624 = pi02815 & w3488;
assign w51625 = pi09207 & w3223;
assign w51626 = pi08920 & w3225;
assign w51627 = pi09253 & w3594;
assign w51628 = pi09051 & w3590;
assign w51629 = pi09266 & w3173;
assign w51630 = pi08509 & w3492;
assign w51631 = pi04798 & w3498;
assign w51632 = pi04654 & w3103;
assign w51633 = pi09044 & w3194;
assign w51634 = pi03246 & w3153;
assign w51635 = pi08965 & w3448;
assign w51636 = pi04693 & w3262;
assign w51637 = pi04726 & w3244;
assign w51638 = pi09438 & w3578;
assign w51639 = pi08939 & w3620;
assign w51640 = pi04713 & w3610;
assign w51641 = pi08894 & w3364;
assign w51642 = pi08842 & w3406;
assign w51643 = pi08998 & w3167;
assign w51644 = pi08972 & w3566;
assign w51645 = pi04518 & w3614;
assign w51646 = pi09273 & w3584;
assign w51647 = pi09103 & w3464;
assign w51648 = pi09365 & w3580;
assign w51649 = pi08881 & w3420;
assign w51650 = pi09331 & w3280;
assign w51651 = pi01540 & w3150;
assign w51652 = pi09122 & w3386;
assign w51653 = pi08684 & w3422;
assign w51654 = pi09180 & w3474;
assign w51655 = pi04551 & w3197;
assign w51656 = pi08887 & w3135;
assign w51657 = pi09239 & w3608;
assign w51658 = pi04819 & w3071;
assign w51659 = pi09017 & w3201;
assign w51660 = pi04732 & w3548;
assign w51661 = pi08582 & w3378;
assign w51662 = pi09142 & w3596;
assign w51663 = pi04531 & w3380;
assign w51664 = pi04765 & w3209;
assign w51665 = pi05017 & w3504;
assign w51666 = pi08743 & w3186;
assign w51667 = pi09425 & w3158;
assign w51668 = pi04990 & w3302;
assign w51669 = pi08521 & w3252;
assign w51670 = pi08763 & w3256;
assign w51671 = pi08724 & w3082;
assign w51672 = pi09305 & w3282;
assign w51673 = pi08671 & w3129;
assign w51674 = pi08469 & w3308;
assign w51675 = pi09312 & w3264;
assign w51676 = pi01587 & w3199;
assign w51677 = pi09397 & w3294;
assign w51678 = pi09030 & w3374;
assign w51679 = pi04641 & w3400;
assign w51680 = pi04596 & w3362;
assign w51681 = pi09168 & w3426;
assign w51682 = pi04575 & w3268;
assign w51683 = pi02575 & w3288;
assign w51684 = pi04667 & w3536;
assign w51685 = pi04525 & w3306;
assign w51686 = pi08526 & w3219;
assign w51687 = pi07994 & w3540;
assign w51688 = pi05056 & w3396;
assign w51689 = pi09478 & w3418;
assign w51690 = pi05009 & w3162;
assign w51691 = pi04583 & w3416;
assign w51692 = pi05062 & w3211;
assign w51693 = pi04602 & w3404;
assign w51694 = pi08476 & w3436;
assign w51695 = pi04886 & w3326;
assign w51696 = pi08790 & w3432;
assign w51697 = pi09384 & w3342;
assign w51698 = pi08572 & w3217;
assign w51699 = pi09344 & w3318;
assign w51700 = pi09772 & w3344;
assign w51701 = pi09292 & w3320;
assign w51702 = pi09194 & w3616;
assign w51703 = pi08809 & w3398;
assign w51704 = pi04812 & w3394;
assign w51705 = pi04772 & w3338;
assign w51706 = pi09174 & w3516;
assign w51707 = pi09299 & w3478;
assign w51708 = pi09485 & w3246;
assign w51709 = pi04609 & w3330;
assign w51710 = pi08489 & w3598;
assign w51711 = pi08777 & w3442;
assign w51712 = pi08613 & w3482;
assign w51713 = pi08868 & w3552;
assign w51714 = pi08816 & w3234;
assign w51715 = pi09116 & w3270;
assign w51716 = pi09432 & w3602;
assign w51717 = pi04879 & w3290;
assign w51718 = pi05023 & w3184;
assign w51719 = pi04983 & w3169;
assign w51720 = pi04622 & w3250;
assign w51721 = pi08861 & w3286;
assign w51722 = pi09378 & w3560;
assign w51723 = pi09418 & w3332;
assign w51724 = pi05049 & w3588;
assign w51725 = pi04540 & w3346;
assign w51726 = pi08829 & w3127;
assign w51727 = pi04918 & w3190;
assign w51728 = pi04846 & w3428;
assign w51729 = pi09187 & w3532;
assign w51730 = pi09200 & w3175;
assign w51731 = pi01730 & w3266;
assign w51732 = pi04839 & w3494;
assign w51733 = pi04674 & w3424;
assign w51734 = pi09090 & w3360;
assign w51735 = pi09004 & w3312;
assign w51736 = pi09286 & w3444;
assign w51737 = pi08933 & w3221;
assign w51738 = pi04925 & w3328;
assign w51739 = pi08978 & w3276;
assign w51740 = pi08756 & w3078;
assign w51741 = pi08959 & w3358;
assign w51742 = pi09155 & w3093;
assign w51743 = pi04852 & w3522;
assign w51744 = pi09096 & w3390;
assign w51745 = pi01815 & w3236;
assign w51746 = pi04758 & w3576;
assign w51747 = pi08913 & w3254;
assign w51748 = pi04833 & w3574;
assign w51749 = pi08991 & w3508;
assign w51750 = pi08737 & w3514;
assign w51751 = pi08553 & w3568;
assign w51752 = pi08803 & w3300;
assign w51753 = pi09464 & w3160;
assign w51754 = pi04905 & w3086;
assign w51755 = pi05030 & w3556;
assign w51756 = pi04785 & w3456;
assign w51757 = pi09226 & w3570;
assign w51758 = pi04912 & w3115;
assign w51759 = pi04865 & w3502;
assign w51760 = pi08730 & w3278;
assign w51761 = pi08710 & w3496;
assign w51762 = pi09371 & w3229;
assign w51763 = pi08946 & w3272;
assign w51764 = pi09352 & w3188;
assign w51765 = pi09161 & w3238;
assign w51766 = pi01552 & w3586;
assign w51767 = pi09411 & w3324;
assign w51768 = pi09010 & w3165;
assign w51769 = pi04570 & w3500;
assign w51770 = pi04957 & w3618;
assign w51771 = pi09391 & w3148;
assign w51772 = pi01547 & w3558;
assign w51773 = pi04826 & w3118;
assign w51774 = pi08848 & w3572;
assign w51775 = pi09458 & w3368;
assign w51776 = pi01718 & w3240;
assign w51777 = pi01536 & w3604;
assign w51778 = pi09318 & w3546;
assign w51779 = pi04680 & w3296;
assign w51780 = pi05036 & w3388;
assign w51781 = pi08587 & w3356;
assign w51782 = pi09445 & w3179;
assign w51783 = pi04706 & w3260;
assign w51784 = pi08952 & w3376;
assign w51785 = pi04899 & w3214;
assign w51786 = pi04739 & w3490;
assign w51787 = pi08604 & w3414;
assign w51788 = pi09451 & w3438;
assign w51789 = pi04635 & w3534;
assign w51790 = pi09279 & w3106;
assign w51791 = pi09220 & w3446;
assign w51792 = pi08697 & w3304;
assign w51793 = pi02078 & w3486;
assign w51794 = pi09213 & w3606;
assign w51795 = pi04806 & w3132;
assign w51796 = pi04700 & w3292;
assign w51797 = pi01526 & w3227;
assign w51798 = pi04892 & w3334;
assign w51799 = pi09471 & w3524;
assign w51800 = pi08822 & w3466;
assign w51801 = pi04964 & w3512;
assign w51802 = pi08985 & w3434;
assign w51803 = pi08907 & w3205;
assign w51804 = pi02442 & w3510;
assign w51805 = pi04745 & w3526;
assign w51806 = pi09070 & w3476;
assign w51807 = pi08515 & w3612;
assign w51808 = pi09247 & w3366;
assign w51809 = pi09472 & w3112;
assign w51810 = pi08632 & w3450;
assign w51811 = pi09077 & w3458;
assign w51812 = pi04557 & w3336;
assign w51813 = pi09233 & w3440;
assign w51814 = pi08619 & w3314;
assign w51815 = pi08926 & w3472;
assign w51816 = pi08750 & w3284;
assign w51817 = pi08900 & w3156;
assign w51818 = pi04931 & w3484;
assign w51819 = pi08593 & w3460;
assign w51820 = pi08664 & w3203;
assign w51821 = pi08855 & w3340;
assign w51822 = pi04779 & w3348;
assign w51823 = pi09135 & w3352;
assign w51824 = pi09260 & w3468;
assign w51825 = pi08482 & w3248;
assign w51826 = pi04752 & w3350;
assign w51827 = pi04970 & w3412;
assign w51828 = pi09064 & w3171;
assign w51829 = pi09083 & w3192;
assign w51830 = pi08658 & w3392;
assign w51831 = pi02601 & w3528;
assign w51832 = pi01530 & w3462;
assign w51833 = pi05043 & w3177;
assign w51834 = pi08531 & w3554;
assign w51835 = pi09057 & w3430;
assign w51836 = pi04938 & w3146;
assign w51837 = pi08645 & w3298;
assign w51838 = pi09038 & w3600;
assign w51839 = pi08874 & w3410;
assign w51840 = pi08769 & w3518;
assign w51841 = pi04546 & w3520;
assign w51842 = pi09405 & w3316;
assign w51843 = pi09491 & w3110;
assign w51844 = pi05003 & w3122;
assign w51845 = pi09540 & w3408;
assign w51846 = pi04590 & w3470;
assign w51847 = pi08548 & w3550;
assign w51848 = pi08835 & w3139;
assign w51849 = pi04615 & w3530;
assign w51850 = pi08566 & w3480;
assign w51851 = pi01914 & w3232;
assign w51852 = pi04792 & w3592;
assign w51853 = pi04628 & w3064;
assign w51854 = pi04872 & w3454;
assign w51855 = pi09325 & w3542;
assign w51856 = pi04951 & w3370;
assign w51857 = pi09129 & w3382;
assign w51858 = pi09109 & w3207;
assign w51859 = pi04977 & w3562;
assign w51860 = pi09338 & w3096;
assign w51861 = pi08796 & w3506;
assign w51862 = pi05069 & w3582;
assign w51863 = pi04687 & w3137;
assign w51864 = pi04648 & w3322;
assign w51865 = pi09024 & w3372;
assign w51866 = pi04944 & w3564;
assign w51867 = pi01959 & w3384;
assign w51868 = pi01930 & w3538;
assign w51869 = pi01721 & w3354;
assign w51870 = pi09148 & w3125;
assign w51871 = pi08536 & w3452;
assign w51872 = pi08464 & w3143;
assign w51873 = pi04996 & w3258;
assign w51874 = pi04563 & w3544;
assign w51875 = pi04661 & w3274;
assign w51876 = pi09358 & w3402;
assign w51877 = pi05080 & w3242;
assign w51878 = pi04859 & w3181;
assign w51879 = ~w51623 & ~w51624;
assign w51880 = ~w51625 & ~w51626;
assign w51881 = ~w51627 & ~w51628;
assign w51882 = ~w51629 & ~w51630;
assign w51883 = ~w51631 & ~w51632;
assign w51884 = ~w51633 & ~w51634;
assign w51885 = ~w51635 & ~w51636;
assign w51886 = ~w51637 & ~w51638;
assign w51887 = ~w51639 & ~w51640;
assign w51888 = ~w51641 & ~w51642;
assign w51889 = ~w51643 & ~w51644;
assign w51890 = ~w51645 & ~w51646;
assign w51891 = ~w51647 & ~w51648;
assign w51892 = ~w51649 & ~w51650;
assign w51893 = ~w51651 & ~w51652;
assign w51894 = ~w51653 & ~w51654;
assign w51895 = ~w51655 & ~w51656;
assign w51896 = ~w51657 & ~w51658;
assign w51897 = ~w51659 & ~w51660;
assign w51898 = ~w51661 & ~w51662;
assign w51899 = ~w51663 & ~w51664;
assign w51900 = ~w51665 & ~w51666;
assign w51901 = ~w51667 & ~w51668;
assign w51902 = ~w51669 & ~w51670;
assign w51903 = ~w51671 & ~w51672;
assign w51904 = ~w51673 & ~w51674;
assign w51905 = ~w51675 & ~w51676;
assign w51906 = ~w51677 & ~w51678;
assign w51907 = ~w51679 & ~w51680;
assign w51908 = ~w51681 & ~w51682;
assign w51909 = ~w51683 & ~w51684;
assign w51910 = ~w51685 & ~w51686;
assign w51911 = ~w51687 & ~w51688;
assign w51912 = ~w51689 & ~w51690;
assign w51913 = ~w51691 & ~w51692;
assign w51914 = ~w51693 & ~w51694;
assign w51915 = ~w51695 & ~w51696;
assign w51916 = ~w51697 & ~w51698;
assign w51917 = ~w51699 & ~w51700;
assign w51918 = ~w51701 & ~w51702;
assign w51919 = ~w51703 & ~w51704;
assign w51920 = ~w51705 & ~w51706;
assign w51921 = ~w51707 & ~w51708;
assign w51922 = ~w51709 & ~w51710;
assign w51923 = ~w51711 & ~w51712;
assign w51924 = ~w51713 & ~w51714;
assign w51925 = ~w51715 & ~w51716;
assign w51926 = ~w51717 & ~w51718;
assign w51927 = ~w51719 & ~w51720;
assign w51928 = ~w51721 & ~w51722;
assign w51929 = ~w51723 & ~w51724;
assign w51930 = ~w51725 & ~w51726;
assign w51931 = ~w51727 & ~w51728;
assign w51932 = ~w51729 & ~w51730;
assign w51933 = ~w51731 & ~w51732;
assign w51934 = ~w51733 & ~w51734;
assign w51935 = ~w51735 & ~w51736;
assign w51936 = ~w51737 & ~w51738;
assign w51937 = ~w51739 & ~w51740;
assign w51938 = ~w51741 & ~w51742;
assign w51939 = ~w51743 & ~w51744;
assign w51940 = ~w51745 & ~w51746;
assign w51941 = ~w51747 & ~w51748;
assign w51942 = ~w51749 & ~w51750;
assign w51943 = ~w51751 & ~w51752;
assign w51944 = ~w51753 & ~w51754;
assign w51945 = ~w51755 & ~w51756;
assign w51946 = ~w51757 & ~w51758;
assign w51947 = ~w51759 & ~w51760;
assign w51948 = ~w51761 & ~w51762;
assign w51949 = ~w51763 & ~w51764;
assign w51950 = ~w51765 & ~w51766;
assign w51951 = ~w51767 & ~w51768;
assign w51952 = ~w51769 & ~w51770;
assign w51953 = ~w51771 & ~w51772;
assign w51954 = ~w51773 & ~w51774;
assign w51955 = ~w51775 & ~w51776;
assign w51956 = ~w51777 & ~w51778;
assign w51957 = ~w51779 & ~w51780;
assign w51958 = ~w51781 & ~w51782;
assign w51959 = ~w51783 & ~w51784;
assign w51960 = ~w51785 & ~w51786;
assign w51961 = ~w51787 & ~w51788;
assign w51962 = ~w51789 & ~w51790;
assign w51963 = ~w51791 & ~w51792;
assign w51964 = ~w51793 & ~w51794;
assign w51965 = ~w51795 & ~w51796;
assign w51966 = ~w51797 & ~w51798;
assign w51967 = ~w51799 & ~w51800;
assign w51968 = ~w51801 & ~w51802;
assign w51969 = ~w51803 & ~w51804;
assign w51970 = ~w51805 & ~w51806;
assign w51971 = ~w51807 & ~w51808;
assign w51972 = ~w51809 & ~w51810;
assign w51973 = ~w51811 & ~w51812;
assign w51974 = ~w51813 & ~w51814;
assign w51975 = ~w51815 & ~w51816;
assign w51976 = ~w51817 & ~w51818;
assign w51977 = ~w51819 & ~w51820;
assign w51978 = ~w51821 & ~w51822;
assign w51979 = ~w51823 & ~w51824;
assign w51980 = ~w51825 & ~w51826;
assign w51981 = ~w51827 & ~w51828;
assign w51982 = ~w51829 & ~w51830;
assign w51983 = ~w51831 & ~w51832;
assign w51984 = ~w51833 & ~w51834;
assign w51985 = ~w51835 & ~w51836;
assign w51986 = ~w51837 & ~w51838;
assign w51987 = ~w51839 & ~w51840;
assign w51988 = ~w51841 & ~w51842;
assign w51989 = ~w51843 & ~w51844;
assign w51990 = ~w51845 & ~w51846;
assign w51991 = ~w51847 & ~w51848;
assign w51992 = ~w51849 & ~w51850;
assign w51993 = ~w51851 & ~w51852;
assign w51994 = ~w51853 & ~w51854;
assign w51995 = ~w51855 & ~w51856;
assign w51996 = ~w51857 & ~w51858;
assign w51997 = ~w51859 & ~w51860;
assign w51998 = ~w51861 & ~w51862;
assign w51999 = ~w51863 & ~w51864;
assign w52000 = ~w51865 & ~w51866;
assign w52001 = ~w51867 & ~w51868;
assign w52002 = ~w51869 & ~w51870;
assign w52003 = ~w51871 & ~w51872;
assign w52004 = ~w51873 & ~w51874;
assign w52005 = ~w51875 & ~w51876;
assign w52006 = ~w51877 & ~w51878;
assign w52007 = w52005 & w52006;
assign w52008 = w52003 & w52004;
assign w52009 = w52001 & w52002;
assign w52010 = w51999 & w52000;
assign w52011 = w51997 & w51998;
assign w52012 = w51995 & w51996;
assign w52013 = w51993 & w51994;
assign w52014 = w51991 & w51992;
assign w52015 = w51989 & w51990;
assign w52016 = w51987 & w51988;
assign w52017 = w51985 & w51986;
assign w52018 = w51983 & w51984;
assign w52019 = w51981 & w51982;
assign w52020 = w51979 & w51980;
assign w52021 = w51977 & w51978;
assign w52022 = w51975 & w51976;
assign w52023 = w51973 & w51974;
assign w52024 = w51971 & w51972;
assign w52025 = w51969 & w51970;
assign w52026 = w51967 & w51968;
assign w52027 = w51965 & w51966;
assign w52028 = w51963 & w51964;
assign w52029 = w51961 & w51962;
assign w52030 = w51959 & w51960;
assign w52031 = w51957 & w51958;
assign w52032 = w51955 & w51956;
assign w52033 = w51953 & w51954;
assign w52034 = w51951 & w51952;
assign w52035 = w51949 & w51950;
assign w52036 = w51947 & w51948;
assign w52037 = w51945 & w51946;
assign w52038 = w51943 & w51944;
assign w52039 = w51941 & w51942;
assign w52040 = w51939 & w51940;
assign w52041 = w51937 & w51938;
assign w52042 = w51935 & w51936;
assign w52043 = w51933 & w51934;
assign w52044 = w51931 & w51932;
assign w52045 = w51929 & w51930;
assign w52046 = w51927 & w51928;
assign w52047 = w51925 & w51926;
assign w52048 = w51923 & w51924;
assign w52049 = w51921 & w51922;
assign w52050 = w51919 & w51920;
assign w52051 = w51917 & w51918;
assign w52052 = w51915 & w51916;
assign w52053 = w51913 & w51914;
assign w52054 = w51911 & w51912;
assign w52055 = w51909 & w51910;
assign w52056 = w51907 & w51908;
assign w52057 = w51905 & w51906;
assign w52058 = w51903 & w51904;
assign w52059 = w51901 & w51902;
assign w52060 = w51899 & w51900;
assign w52061 = w51897 & w51898;
assign w52062 = w51895 & w51896;
assign w52063 = w51893 & w51894;
assign w52064 = w51891 & w51892;
assign w52065 = w51889 & w51890;
assign w52066 = w51887 & w51888;
assign w52067 = w51885 & w51886;
assign w52068 = w51883 & w51884;
assign w52069 = w51881 & w51882;
assign w52070 = w51879 & w51880;
assign w52071 = w52069 & w52070;
assign w52072 = w52067 & w52068;
assign w52073 = w52065 & w52066;
assign w52074 = w52063 & w52064;
assign w52075 = w52061 & w52062;
assign w52076 = w52059 & w52060;
assign w52077 = w52057 & w52058;
assign w52078 = w52055 & w52056;
assign w52079 = w52053 & w52054;
assign w52080 = w52051 & w52052;
assign w52081 = w52049 & w52050;
assign w52082 = w52047 & w52048;
assign w52083 = w52045 & w52046;
assign w52084 = w52043 & w52044;
assign w52085 = w52041 & w52042;
assign w52086 = w52039 & w52040;
assign w52087 = w52037 & w52038;
assign w52088 = w52035 & w52036;
assign w52089 = w52033 & w52034;
assign w52090 = w52031 & w52032;
assign w52091 = w52029 & w52030;
assign w52092 = w52027 & w52028;
assign w52093 = w52025 & w52026;
assign w52094 = w52023 & w52024;
assign w52095 = w52021 & w52022;
assign w52096 = w52019 & w52020;
assign w52097 = w52017 & w52018;
assign w52098 = w52015 & w52016;
assign w52099 = w52013 & w52014;
assign w52100 = w52011 & w52012;
assign w52101 = w52009 & w52010;
assign w52102 = w52007 & w52008;
assign w52103 = w52101 & w52102;
assign w52104 = w52099 & w52100;
assign w52105 = w52097 & w52098;
assign w52106 = w52095 & w52096;
assign w52107 = w52093 & w52094;
assign w52108 = w52091 & w52092;
assign w52109 = w52089 & w52090;
assign w52110 = w52087 & w52088;
assign w52111 = w52085 & w52086;
assign w52112 = w52083 & w52084;
assign w52113 = w52081 & w52082;
assign w52114 = w52079 & w52080;
assign w52115 = w52077 & w52078;
assign w52116 = w52075 & w52076;
assign w52117 = w52073 & w52074;
assign w52118 = w52071 & w52072;
assign w52119 = w52117 & w52118;
assign w52120 = w52115 & w52116;
assign w52121 = w52113 & w52114;
assign w52122 = w52111 & w52112;
assign w52123 = w52109 & w52110;
assign w52124 = w52107 & w52108;
assign w52125 = w52105 & w52106;
assign w52126 = w52103 & w52104;
assign w52127 = w52125 & w52126;
assign w52128 = w52123 & w52124;
assign w52129 = w52121 & w52122;
assign w52130 = w52119 & w52120;
assign w52131 = w52129 & w52130;
assign w52132 = w52127 & w52128;
assign w52133 = w52131 & w52132;
assign w52134 = ~pi10577 & ~w52133;
assign w52135 = pi09268 & w3584;
assign w52136 = pi08935 & w3620;
assign w52137 = pi09072 & w3458;
assign w52138 = pi09333 & w3096;
assign w52139 = pi04828 & w3574;
assign w52140 = pi08915 & w3225;
assign w52141 = pi08660 & w3203;
assign w52142 = pi04881 & w3326;
assign w52143 = pi08544 & w3550;
assign w52144 = pi04972 & w3562;
assign w52145 = pi08577 & w3378;
assign w52146 = pi09183 & w3532;
assign w52147 = pi09228 & w3440;
assign w52148 = pi08621 & w3538;
assign w52149 = pi04553 & w3336;
assign w52150 = pi01531 & w3436;
assign w52151 = pi09275 & w3106;
assign w52152 = pi09066 & w3476;
assign w52153 = pi05075 & w3242;
assign w52154 = pi08792 & w3506;
assign w52155 = pi08771 & w3442;
assign w52156 = pi08765 & w3518;
assign w52157 = pi01488 & w3394;
assign w52158 = pi01962 & w3103;
assign w52159 = pi04814 & w3071;
assign w52160 = pi09513 & w3510;
assign w52161 = pi04630 & w3534;
assign w52162 = pi04978 & w3169;
assign w52163 = pi04604 & w3330;
assign w52164 = pi08779 & w3384;
assign w52165 = pi04920 & w3328;
assign w52166 = pi08870 & w3410;
assign w52167 = pi08692 & w3304;
assign w52168 = pi09241 & w3366;
assign w52169 = pi08818 & w3466;
assign w52170 = pi08752 & w3078;
assign w52171 = pi09046 & w3590;
assign w52172 = pi09098 & w3464;
assign w52173 = pi08928 & w3221;
assign w52174 = pi09215 & w3446;
assign w52175 = pi02498 & w3524;
assign w52176 = pi09367 & w3229;
assign w52177 = pi09288 & w3320;
assign w52178 = pi02212 & w3438;
assign w52179 = pi08595 & w3586;
assign w52180 = pi09137 & w3596;
assign w52181 = pi02566 & w3568;
assign w52182 = pi09092 & w3390;
assign w52183 = pi09111 & w3270;
assign w52184 = pi01668 & w3498;
assign w52185 = pi08640 & w3298;
assign w52186 = pi08961 & w3448;
assign w52187 = pi08837 & w3406;
assign w52188 = pi01981 & w3520;
assign w52189 = pi09393 & w3294;
assign w52190 = pi05031 & w3388;
assign w52191 = pi08627 & w3450;
assign w52192 = pi09085 & w3360;
assign w52193 = pi08824 & w3127;
assign w52194 = pi09150 & w3093;
assign w52195 = pi08896 & w3156;
assign w52196 = pi01938 & w3296;
assign w52197 = pi09373 & w3560;
assign w52198 = pi04894 & w3214;
assign w52199 = pi05004 & w3162;
assign w52200 = pi09399 & w3316;
assign w52201 = pi05025 & w3556;
assign w52202 = pi08889 & w3364;
assign w52203 = pi09059 & w3171;
assign w52204 = pi04526 & w3380;
assign w52205 = pi04800 & w3132;
assign w52206 = pi08883 & w3135;
assign w52207 = pi04571 & w3268;
assign w52208 = pi09118 & w3386;
assign w52209 = pi04985 & w3302;
assign w52210 = pi09189 & w3616;
assign w52211 = pi08528 & w3554;
assign w52212 = pi08785 & w3432;
assign w52213 = pi04841 & w3428;
assign w52214 = pi08850 & w3340;
assign w52215 = pi04558 & w3544;
assign w52216 = pi01978 & w3404;
assign w52217 = pi08941 & w3272;
assign w52218 = pi04867 & w3454;
assign w52219 = pi08653 & w3392;
assign w52220 = pi08719 & w3082;
assign w52221 = pi04643 & w3322;
assign w52222 = pi01588 & w3248;
assign w52223 = pi09163 & w3426;
assign w52224 = pi01927 & w3262;
assign w52225 = pi04734 & w3490;
assign w52226 = pi04907 & w3115;
assign w52227 = pi04998 & w3122;
assign w52228 = pi09327 & w3280;
assign w52229 = pi09026 & w3374;
assign w52230 = pi08831 & w3139;
assign w52231 = pi09195 & w3175;
assign w52232 = pi02082 & w3306;
assign w52233 = pi04952 & w3618;
assign w52234 = pi09006 & w3165;
assign w52235 = pi08902 & w3205;
assign w52236 = pi09040 & w3194;
assign w52237 = pi09013 & w3201;
assign w52238 = pi05018 & w3184;
assign w52239 = pi02430 & w3414;
assign w52240 = pi04695 & w3292;
assign w52241 = pi01823 & w3548;
assign w52242 = pi08666 & w3129;
assign w52243 = pi09314 & w3546;
assign w52244 = pi09105 & w3207;
assign w52245 = pi08634 & w3236;
assign w52246 = pi01828 & w3260;
assign w52247 = pi04774 & w3348;
assign w52248 = pi08699 & w3462;
assign w52249 = pi09749 & w3522;
assign w52250 = pi08673 & w3199;
assign w52251 = pi09255 & w3468;
assign w52252 = pi05064 & w3582;
assign w52253 = pi08811 & w3234;
assign w52254 = pi04939 & w3564;
assign w52255 = pi05011 & w3504;
assign w52256 = pi09019 & w3372;
assign w52257 = pi09131 & w3352;
assign w52258 = pi08459 & w3143;
assign w52259 = pi08732 & w3514;
assign w52260 = pi08745 & w3284;
assign w52261 = pi09301 & w3282;
assign w52262 = pi01494 & w3368;
assign w52263 = pi05051 & w3396;
assign w52264 = pi08491 & w3492;
assign w52265 = pi09407 & w3324;
assign w52266 = pi09176 & w3474;
assign w52267 = pi09495 & w3314;
assign w52268 = pi04854 & w3181;
assign w52269 = pi04682 & w3137;
assign w52270 = pi08922 & w3472;
assign w52271 = pi03019 & w3362;
assign w52272 = pi09307 & w3264;
assign w52273 = pi08465 & w3308;
assign w52274 = pi09506 & w3408;
assign w52275 = pi04991 & w3258;
assign w52276 = pi09053 & w3430;
assign w52277 = pi05038 & w3177;
assign w52278 = pi08987 & w3508;
assign w52279 = pi09170 & w3516;
assign w52280 = pi08510 & w3612;
assign w52281 = pi09209 & w3606;
assign w52282 = pi04565 & w3500;
assign w52283 = pi09522 & w3160;
assign w52284 = pi08647 & w3354;
assign w52285 = pi08440 & w3232;
assign w52286 = pi02064 & w3346;
assign w52287 = pi08446 & w3240;
assign w52288 = pi04874 & w3290;
assign w52289 = pi04959 & w3512;
assign w52290 = pi09722 & w3502;
assign w52291 = pi01842 & w3310;
assign w52292 = pi08606 & w3540;
assign w52293 = pi09202 & w3223;
assign w52294 = pi04900 & w3086;
assign w52295 = pi04747 & w3350;
assign w52296 = pi09235 & w3608;
assign w52297 = pi01994 & w3530;
assign w52298 = pi04913 & w3190;
assign w52299 = pi08679 & w3422;
assign w52300 = pi09000 & w3312;
assign w52301 = pi08954 & w3358;
assign w52302 = pi09249 & w3594;
assign w52303 = pi09486 & w3110;
assign w52304 = pi02552 & w3179;
assign w52305 = pi09479 & w3246;
assign w52306 = pi08559 & w3480;
assign w52307 = pi08712 & w3153;
assign w52308 = pi08993 & w3167;
assign w52309 = pi08433 & w3486;
assign w52310 = pi04177 & w3252;
assign w52311 = pi08686 & w3227;
assign w52312 = pi09262 & w3173;
assign w52313 = pi09157 & w3238;
assign w52314 = pi09079 & w3192;
assign w52315 = pi01950 & w3536;
assign w52316 = pi09354 & w3402;
assign w52317 = pi08453 & w3266;
assign w52318 = pi08844 & w3572;
assign w52319 = pi01750 & w3456;
assign w52320 = pi01602 & w3578;
assign w52321 = pi04669 & w3424;
assign w52322 = pi09340 & w3318;
assign w52323 = pi09380 & w3342;
assign w52324 = pi09320 & w3542;
assign w52325 = pi01567 & w3598;
assign w52326 = pi08532 & w3452;
assign w52327 = pi04585 & w3470;
assign w52328 = pi08568 & w3217;
assign w52329 = pi03114 & w3482;
assign w52330 = pi02568 & w3158;
assign w52331 = pi02418 & w3602;
assign w52332 = pi09360 & w3580;
assign w52333 = pi08726 & w3278;
assign w52334 = pi08980 & w3434;
assign w52335 = pi05044 & w3588;
assign w52336 = pi04577 & w3416;
assign w52337 = pi05070 & w3488;
assign w52338 = pi04965 & w3412;
assign w52339 = pi04787 & w3592;
assign w52340 = pi04926 & w3484;
assign w52341 = pi08538 & w3528;
assign w52342 = pi09500 & w3558;
assign w52343 = pi04887 & w3334;
assign w52344 = pi04513 & w3614;
assign w52345 = pi09144 & w3125;
assign w52346 = pi08863 & w3552;
assign w52347 = pi08589 & w3460;
assign w52348 = pi09294 & w3478;
assign w52349 = pi09386 & w3148;
assign w52350 = pi01960 & w3064;
assign w52351 = pi04617 & w3250;
assign w52352 = pi08948 & w3376;
assign w52353 = pi04946 & w3370;
assign w52354 = pi08584 & w3356;
assign w52355 = pi01969 & w3400;
assign w52356 = pi08909 & w3254;
assign w52357 = pi04933 & w3146;
assign w52358 = pi09796 & w3494;
assign w52359 = pi08758 & w3256;
assign w52360 = pi08974 & w3276;
assign w52361 = pi05057 & w3211;
assign w52362 = pi09222 & w3570;
assign w52363 = pi04708 & w3610;
assign w52364 = pi09473 & w3418;
assign w52365 = pi08541 & w3219;
assign w52366 = pi09281 & w3444;
assign w52367 = pi08492 & w3604;
assign w52368 = pi08705 & w3496;
assign w52369 = pi09032 & w3600;
assign w52370 = pi08555 & w3288;
assign w52371 = pi02045 & w3197;
assign w52372 = pi09492 & w3150;
assign w52373 = pi08876 & w3420;
assign w52374 = pi08573 & w3112;
assign w52375 = pi01766 & w3338;
assign w52376 = pi01803 & w3526;
assign w52377 = pi08739 & w3186;
assign w52378 = pi09124 & w3382;
assign w52379 = pi04760 & w3209;
assign w52380 = pi08798 & w3300;
assign w52381 = pi08857 & w3286;
assign w52382 = pi09346 & w3188;
assign w52383 = pi01758 & w3576;
assign w52384 = pi04721 & w3244;
assign w52385 = pi04656 & w3274;
assign w52386 = pi08967 & w3566;
assign w52387 = pi01513 & w3118;
assign w52388 = pi08805 & w3398;
assign w52389 = pi09413 & w3332;
assign w52390 = pi08498 & w3344;
assign w52391 = ~w52135 & ~w52136;
assign w52392 = ~w52137 & ~w52138;
assign w52393 = ~w52139 & ~w52140;
assign w52394 = ~w52141 & ~w52142;
assign w52395 = ~w52143 & ~w52144;
assign w52396 = ~w52145 & ~w52146;
assign w52397 = ~w52147 & ~w52148;
assign w52398 = ~w52149 & ~w52150;
assign w52399 = ~w52151 & ~w52152;
assign w52400 = ~w52153 & ~w52154;
assign w52401 = ~w52155 & ~w52156;
assign w52402 = ~w52157 & ~w52158;
assign w52403 = ~w52159 & ~w52160;
assign w52404 = ~w52161 & ~w52162;
assign w52405 = ~w52163 & ~w52164;
assign w52406 = ~w52165 & ~w52166;
assign w52407 = ~w52167 & ~w52168;
assign w52408 = ~w52169 & ~w52170;
assign w52409 = ~w52171 & ~w52172;
assign w52410 = ~w52173 & ~w52174;
assign w52411 = ~w52175 & ~w52176;
assign w52412 = ~w52177 & ~w52178;
assign w52413 = ~w52179 & ~w52180;
assign w52414 = ~w52181 & ~w52182;
assign w52415 = ~w52183 & ~w52184;
assign w52416 = ~w52185 & ~w52186;
assign w52417 = ~w52187 & ~w52188;
assign w52418 = ~w52189 & ~w52190;
assign w52419 = ~w52191 & ~w52192;
assign w52420 = ~w52193 & ~w52194;
assign w52421 = ~w52195 & ~w52196;
assign w52422 = ~w52197 & ~w52198;
assign w52423 = ~w52199 & ~w52200;
assign w52424 = ~w52201 & ~w52202;
assign w52425 = ~w52203 & ~w52204;
assign w52426 = ~w52205 & ~w52206;
assign w52427 = ~w52207 & ~w52208;
assign w52428 = ~w52209 & ~w52210;
assign w52429 = ~w52211 & ~w52212;
assign w52430 = ~w52213 & ~w52214;
assign w52431 = ~w52215 & ~w52216;
assign w52432 = ~w52217 & ~w52218;
assign w52433 = ~w52219 & ~w52220;
assign w52434 = ~w52221 & ~w52222;
assign w52435 = ~w52223 & ~w52224;
assign w52436 = ~w52225 & ~w52226;
assign w52437 = ~w52227 & ~w52228;
assign w52438 = ~w52229 & ~w52230;
assign w52439 = ~w52231 & ~w52232;
assign w52440 = ~w52233 & ~w52234;
assign w52441 = ~w52235 & ~w52236;
assign w52442 = ~w52237 & ~w52238;
assign w52443 = ~w52239 & ~w52240;
assign w52444 = ~w52241 & ~w52242;
assign w52445 = ~w52243 & ~w52244;
assign w52446 = ~w52245 & ~w52246;
assign w52447 = ~w52247 & ~w52248;
assign w52448 = ~w52249 & ~w52250;
assign w52449 = ~w52251 & ~w52252;
assign w52450 = ~w52253 & ~w52254;
assign w52451 = ~w52255 & ~w52256;
assign w52452 = ~w52257 & ~w52258;
assign w52453 = ~w52259 & ~w52260;
assign w52454 = ~w52261 & ~w52262;
assign w52455 = ~w52263 & ~w52264;
assign w52456 = ~w52265 & ~w52266;
assign w52457 = ~w52267 & ~w52268;
assign w52458 = ~w52269 & ~w52270;
assign w52459 = ~w52271 & ~w52272;
assign w52460 = ~w52273 & ~w52274;
assign w52461 = ~w52275 & ~w52276;
assign w52462 = ~w52277 & ~w52278;
assign w52463 = ~w52279 & ~w52280;
assign w52464 = ~w52281 & ~w52282;
assign w52465 = ~w52283 & ~w52284;
assign w52466 = ~w52285 & ~w52286;
assign w52467 = ~w52287 & ~w52288;
assign w52468 = ~w52289 & ~w52290;
assign w52469 = ~w52291 & ~w52292;
assign w52470 = ~w52293 & ~w52294;
assign w52471 = ~w52295 & ~w52296;
assign w52472 = ~w52297 & ~w52298;
assign w52473 = ~w52299 & ~w52300;
assign w52474 = ~w52301 & ~w52302;
assign w52475 = ~w52303 & ~w52304;
assign w52476 = ~w52305 & ~w52306;
assign w52477 = ~w52307 & ~w52308;
assign w52478 = ~w52309 & ~w52310;
assign w52479 = ~w52311 & ~w52312;
assign w52480 = ~w52313 & ~w52314;
assign w52481 = ~w52315 & ~w52316;
assign w52482 = ~w52317 & ~w52318;
assign w52483 = ~w52319 & ~w52320;
assign w52484 = ~w52321 & ~w52322;
assign w52485 = ~w52323 & ~w52324;
assign w52486 = ~w52325 & ~w52326;
assign w52487 = ~w52327 & ~w52328;
assign w52488 = ~w52329 & ~w52330;
assign w52489 = ~w52331 & ~w52332;
assign w52490 = ~w52333 & ~w52334;
assign w52491 = ~w52335 & ~w52336;
assign w52492 = ~w52337 & ~w52338;
assign w52493 = ~w52339 & ~w52340;
assign w52494 = ~w52341 & ~w52342;
assign w52495 = ~w52343 & ~w52344;
assign w52496 = ~w52345 & ~w52346;
assign w52497 = ~w52347 & ~w52348;
assign w52498 = ~w52349 & ~w52350;
assign w52499 = ~w52351 & ~w52352;
assign w52500 = ~w52353 & ~w52354;
assign w52501 = ~w52355 & ~w52356;
assign w52502 = ~w52357 & ~w52358;
assign w52503 = ~w52359 & ~w52360;
assign w52504 = ~w52361 & ~w52362;
assign w52505 = ~w52363 & ~w52364;
assign w52506 = ~w52365 & ~w52366;
assign w52507 = ~w52367 & ~w52368;
assign w52508 = ~w52369 & ~w52370;
assign w52509 = ~w52371 & ~w52372;
assign w52510 = ~w52373 & ~w52374;
assign w52511 = ~w52375 & ~w52376;
assign w52512 = ~w52377 & ~w52378;
assign w52513 = ~w52379 & ~w52380;
assign w52514 = ~w52381 & ~w52382;
assign w52515 = ~w52383 & ~w52384;
assign w52516 = ~w52385 & ~w52386;
assign w52517 = ~w52387 & ~w52388;
assign w52518 = ~w52389 & ~w52390;
assign w52519 = w52517 & w52518;
assign w52520 = w52515 & w52516;
assign w52521 = w52513 & w52514;
assign w52522 = w52511 & w52512;
assign w52523 = w52509 & w52510;
assign w52524 = w52507 & w52508;
assign w52525 = w52505 & w52506;
assign w52526 = w52503 & w52504;
assign w52527 = w52501 & w52502;
assign w52528 = w52499 & w52500;
assign w52529 = w52497 & w52498;
assign w52530 = w52495 & w52496;
assign w52531 = w52493 & w52494;
assign w52532 = w52491 & w52492;
assign w52533 = w52489 & w52490;
assign w52534 = w52487 & w52488;
assign w52535 = w52485 & w52486;
assign w52536 = w52483 & w52484;
assign w52537 = w52481 & w52482;
assign w52538 = w52479 & w52480;
assign w52539 = w52477 & w52478;
assign w52540 = w52475 & w52476;
assign w52541 = w52473 & w52474;
assign w52542 = w52471 & w52472;
assign w52543 = w52469 & w52470;
assign w52544 = w52467 & w52468;
assign w52545 = w52465 & w52466;
assign w52546 = w52463 & w52464;
assign w52547 = w52461 & w52462;
assign w52548 = w52459 & w52460;
assign w52549 = w52457 & w52458;
assign w52550 = w52455 & w52456;
assign w52551 = w52453 & w52454;
assign w52552 = w52451 & w52452;
assign w52553 = w52449 & w52450;
assign w52554 = w52447 & w52448;
assign w52555 = w52445 & w52446;
assign w52556 = w52443 & w52444;
assign w52557 = w52441 & w52442;
assign w52558 = w52439 & w52440;
assign w52559 = w52437 & w52438;
assign w52560 = w52435 & w52436;
assign w52561 = w52433 & w52434;
assign w52562 = w52431 & w52432;
assign w52563 = w52429 & w52430;
assign w52564 = w52427 & w52428;
assign w52565 = w52425 & w52426;
assign w52566 = w52423 & w52424;
assign w52567 = w52421 & w52422;
assign w52568 = w52419 & w52420;
assign w52569 = w52417 & w52418;
assign w52570 = w52415 & w52416;
assign w52571 = w52413 & w52414;
assign w52572 = w52411 & w52412;
assign w52573 = w52409 & w52410;
assign w52574 = w52407 & w52408;
assign w52575 = w52405 & w52406;
assign w52576 = w52403 & w52404;
assign w52577 = w52401 & w52402;
assign w52578 = w52399 & w52400;
assign w52579 = w52397 & w52398;
assign w52580 = w52395 & w52396;
assign w52581 = w52393 & w52394;
assign w52582 = w52391 & w52392;
assign w52583 = w52581 & w52582;
assign w52584 = w52579 & w52580;
assign w52585 = w52577 & w52578;
assign w52586 = w52575 & w52576;
assign w52587 = w52573 & w52574;
assign w52588 = w52571 & w52572;
assign w52589 = w52569 & w52570;
assign w52590 = w52567 & w52568;
assign w52591 = w52565 & w52566;
assign w52592 = w52563 & w52564;
assign w52593 = w52561 & w52562;
assign w52594 = w52559 & w52560;
assign w52595 = w52557 & w52558;
assign w52596 = w52555 & w52556;
assign w52597 = w52553 & w52554;
assign w52598 = w52551 & w52552;
assign w52599 = w52549 & w52550;
assign w52600 = w52547 & w52548;
assign w52601 = w52545 & w52546;
assign w52602 = w52543 & w52544;
assign w52603 = w52541 & w52542;
assign w52604 = w52539 & w52540;
assign w52605 = w52537 & w52538;
assign w52606 = w52535 & w52536;
assign w52607 = w52533 & w52534;
assign w52608 = w52531 & w52532;
assign w52609 = w52529 & w52530;
assign w52610 = w52527 & w52528;
assign w52611 = w52525 & w52526;
assign w52612 = w52523 & w52524;
assign w52613 = w52521 & w52522;
assign w52614 = w52519 & w52520;
assign w52615 = w52613 & w52614;
assign w52616 = w52611 & w52612;
assign w52617 = w52609 & w52610;
assign w52618 = w52607 & w52608;
assign w52619 = w52605 & w52606;
assign w52620 = w52603 & w52604;
assign w52621 = w52601 & w52602;
assign w52622 = w52599 & w52600;
assign w52623 = w52597 & w52598;
assign w52624 = w52595 & w52596;
assign w52625 = w52593 & w52594;
assign w52626 = w52591 & w52592;
assign w52627 = w52589 & w52590;
assign w52628 = w52587 & w52588;
assign w52629 = w52585 & w52586;
assign w52630 = w52583 & w52584;
assign w52631 = w52629 & w52630;
assign w52632 = w52627 & w52628;
assign w52633 = w52625 & w52626;
assign w52634 = w52623 & w52624;
assign w52635 = w52621 & w52622;
assign w52636 = w52619 & w52620;
assign w52637 = w52617 & w52618;
assign w52638 = w52615 & w52616;
assign w52639 = w52637 & w52638;
assign w52640 = w52635 & w52636;
assign w52641 = w52633 & w52634;
assign w52642 = w52631 & w52632;
assign w52643 = w52641 & w52642;
assign w52644 = w52639 & w52640;
assign w52645 = w52643 & w52644;
assign w52646 = ~pi10577 & ~w52645;
assign w52647 = pi01985 & w3554;
assign w52648 = pi04374 & w3468;
assign w52649 = pi08269 & w3580;
assign w52650 = pi03627 & w3262;
assign w52651 = pi03744 & w3490;
assign w52652 = pi08123 & w3570;
assign w52653 = pi03178 & w3380;
assign w52654 = pi03258 & w3500;
assign w52655 = pi03191 & w3520;
assign w52656 = pi04360 & w3484;
assign w52657 = pi04428 & w3258;
assign w52658 = pi03490 & w3064;
assign w52659 = pi09746 & w3356;
assign w52660 = pi03704 & w3244;
assign w52661 = pi03265 & w3268;
assign w52662 = pi04381 & w3370;
assign w52663 = pi08060 & w3175;
assign w52664 = pi01850 & w3568;
assign w52665 = pi07004 & w3572;
assign w52666 = pi08393 & w3110;
assign w52667 = pi08328 & w3158;
assign w52668 = pi08256 & w3188;
assign w52669 = pi03908 & w3348;
assign w52670 = pi03986 & w3132;
assign w52671 = pi04395 & w3512;
assign w52672 = pi07121 & w3420;
assign w52673 = pi06325 & w3538;
assign w52674 = pi04354 & w3328;
assign w52675 = pi02322 & w3227;
assign w52676 = pi09765 & w3598;
assign w52677 = pi08367 & w3160;
assign w52678 = pi06895 & w3506;
assign w52679 = pi03881 & w3338;
assign w52680 = pi04235 & w3290;
assign w52681 = pi06676 & w3082;
assign w52682 = pi04441 & w3162;
assign w52683 = pi04071 & w3428;
assign w52684 = pi06251 & w3414;
assign w52685 = pi04401 & w3412;
assign w52686 = pi07108 & w3410;
assign w52687 = pi08380 & w3418;
assign w52688 = pi07966 & w3238;
assign w52689 = pi08000 & w3474;
assign w52690 = pi06077 & w3550;
assign w52691 = pi05921 & w3344;
assign w52692 = pi03665 & w3610;
assign w52693 = pi06500 & w3422;
assign w52694 = pi03542 & w3322;
assign w52695 = pi07330 & w3272;
assign w52696 = pi08236 & w3280;
assign w52697 = pi07677 & w3590;
assign w52698 = pi04415 & w3169;
assign w52699 = pi03159 & w3306;
assign w52700 = pi06854 & w3442;
assign w52701 = pi03920 & w3456;
assign w52702 = pi05112 & w3492;
assign w52703 = pi04091 & w3522;
assign w52704 = pi02526 & w3444;
assign w52705 = pi09537 & w3432;
assign w52706 = pi08275 & w3229;
assign w52707 = pi06316 & w3156;
assign w52708 = pi03563 & w3103;
assign w52709 = pi03143 & w3614;
assign w52710 = pi01774 & w3078;
assign w52711 = pi04373 & w3564;
assign w52712 = pi07821 & w3207;
assign w52713 = pi06272 & w3540;
assign w52714 = pi08027 & w3532;
assign w52715 = pi07838 & w3270;
assign w52716 = pi02374 & w3458;
assign w52717 = pi07637 & w3600;
assign w52718 = pi04461 & w3556;
assign w52719 = pi07048 & w3286;
assign w52720 = pi07286 & w3221;
assign w52721 = pi03219 & w3173;
assign w52722 = pi03868 & w3576;
assign w52723 = pi08072 & w3223;
assign w52724 = pi04467 & w3388;
assign w52725 = pi07687 & w3430;
assign w52726 = pi03217 & w3336;
assign w52727 = pi08230 & w3542;
assign w52728 = pi04388 & w3618;
assign w52729 = pi08387 & w3246;
assign w52730 = pi08321 & w3332;
assign w52731 = pi08354 & w3438;
assign w52732 = pi07707 & w3171;
assign w52733 = pi08427 & w3242;
assign w52734 = pi02664 & w3167;
assign w52735 = pi04150 & w3502;
assign w52736 = pi09612 & w3586;
assign w52737 = pi02426 & w3264;
assign w52738 = pi03472 & w3250;
assign w52739 = pi04435 & w3122;
assign w52740 = pi01989 & w3266;
assign w52741 = pi08301 & w3294;
assign w52742 = pi08406 & w3558;
assign w52743 = pi06730 & w3514;
assign w52744 = pi02462 & w3320;
assign w52745 = pi08143 & w3608;
assign w52746 = pi07233 & w3225;
assign w52747 = pi09695 & w3364;
assign w52748 = pi02101 & w3186;
assign w52749 = pi08340 & w3578;
assign w52750 = pi07440 & w3434;
assign w52751 = pi06935 & w3234;
assign w52752 = pi06291 & w3482;
assign w52753 = pi02634 & w3106;
assign w52754 = pi05668 & w3486;
assign w52755 = pi03521 & w3400;
assign w52756 = pi03446 & w3530;
assign w52757 = pi06921 & w3398;
assign w52758 = pi09674 & w3129;
assign w52759 = pi03503 & w3534;
assign w52760 = pi06533 & w3304;
assign w52761 = pi03621 & w3137;
assign w52762 = pi01796 & w3406;
assign w52763 = pi05691 & w3232;
assign w52764 = pi05876 & w3604;
assign w52765 = pi08249 & w3318;
assign w52766 = pi03211 & w3197;
assign w52767 = pi03614 & w3296;
assign w52768 = pi01770 & w3450;
assign w52769 = pi08243 & w3096;
assign w52770 = pi07795 & w3390;
assign w52771 = pi04487 & w3396;
assign w52772 = pi07590 & w3372;
assign w52773 = pi05772 & w3143;
assign w52774 = pi07772 & w3192;
assign w52775 = pi08362 & w3368;
assign w52776 = pi07912 & w3596;
assign w52777 = pi06420 & w3203;
assign w52778 = pi06467 & w3199;
assign w52779 = pi07991 & w3516;
assign w52780 = pi03582 & w3274;
assign w52781 = pi07320 & w3620;
assign w52782 = pi02098 & w3127;
assign w52783 = pi04448 & w3504;
assign w52784 = pi06587 & w3153;
assign w52785 = pi04506 & w3488;
assign w52786 = pi01626 & w3112;
assign w52787 = pi01609 & w3148;
assign w52788 = pi05834 & w3248;
assign w52789 = pi03940 & w3592;
assign w52790 = pi04058 & w3574;
assign w52791 = pi01920 & w3350;
assign w52792 = pi07220 & w3254;
assign w52793 = pi07257 & w3472;
assign w52794 = pi08282 & w3560;
assign w52795 = pi05969 & w3252;
assign w52796 = pi08314 & w3324;
assign w52797 = pi08400 & w3150;
assign w52798 = pi02645 & w3584;
assign w52799 = pi08334 & w3602;
assign w52800 = pi06828 & w3518;
assign w52801 = pi03185 & w3346;
assign w52802 = pi02168 & w3184;
assign w52803 = pi05814 & w3436;
assign w52804 = pi06043 & w3452;
assign w52805 = pi04157 & w3454;
assign w52806 = pi03966 & w3498;
assign w52807 = pi02519 & w3612;
assign w52808 = pi01639 & w3276;
assign w52809 = pi01826 & w3496;
assign w52810 = pi09658 & w3460;
assign w52811 = pi06908 & w3300;
assign w52812 = pi01676 & w3354;
assign w52813 = pi06408 & w3392;
assign w52814 = pi03390 & w3404;
assign w52815 = pi07786 & w3360;
assign w52816 = pi03596 & w3536;
assign w52817 = pi01814 & w3288;
assign w52818 = pi04018 & w3071;
assign w52819 = pi09400 & w3594;
assign w52820 = pi04493 & w3211;
assign w52821 = pi04065 & w3494;
assign w52822 = pi01684 & w3298;
assign w52823 = pi06064 & w3528;
assign w52824 = pi04276 & w3334;
assign w52825 = pi07852 & w3386;
assign w52826 = pi04480 & w3588;
assign w52827 = pi07578 & w3201;
assign w52828 = pi04500 & w3582;
assign w52829 = pi08086 & w3606;
assign w52830 = pi05988 & w3219;
assign w52831 = pi04031 & w3118;
assign w52832 = pi02128 & w3362;
assign w52833 = pi06774 & w3284;
assign w52834 = pi04110 & w3181;
assign w52835 = pi05719 & w3240;
assign w52836 = pi02436 & w3476;
assign w52837 = pi07932 & w3125;
assign w52838 = pi03874 & w3209;
assign w52839 = pi06658 & w3194;
assign w52840 = pi07979 & w3426;
assign w52841 = pi08137 & w3440;
assign w52842 = pi07093 & w3552;
assign w52843 = pi07342 & w3376;
assign w52844 = pi07207 & w3205;
assign w52845 = pi02432 & w3165;
assign w52846 = pi08308 & w3316;
assign w52847 = pi02464 & w3278;
assign w52848 = pi05794 & w3308;
assign w52849 = pi06311 & w3314;
assign w52850 = pi07372 & w3358;
assign w52851 = pi08262 & w3402;
assign w52852 = pi04474 & w3177;
assign w52853 = pi04341 & w3115;
assign w52854 = pi08046 & w3616;
assign w52855 = pi06947 & w3466;
assign w52856 = pi04302 & w3214;
assign w52857 = pi09738 & w3384;
assign w52858 = pi03345 & w3416;
assign w52859 = pi08375 & w3524;
assign w52860 = pi04334 & w3086;
assign w52861 = pi07812 & w3464;
assign w52862 = pi08419 & w3510;
assign w52863 = pi01699 & w3236;
assign w52864 = pi07891 & w3352;
assign w52865 = pi06553 & w3462;
assign w52866 = pi03231 & w3544;
assign w52867 = pi07017 & w3340;
assign w52868 = pi07411 & w3566;
assign w52869 = pi03718 & w3548;
assign w52870 = pi06124 & w3480;
assign w52871 = pi03608 & w3424;
assign w52872 = pi01690 & w3217;
assign w52873 = pi07871 & w3382;
assign w52874 = pi03403 & w3330;
assign w52875 = pi02151 & w3546;
assign w52876 = pi08288 & w3342;
assign w52877 = pi04254 & w3326;
assign w52878 = pi04422 & w3302;
assign w52879 = pi03634 & w3292;
assign w52880 = pi04347 & w3190;
assign w52881 = pi08107 & w3446;
assign w52882 = pi08347 & w3179;
assign w52883 = pi06973 & w3139;
assign w52884 = pi07954 & w3093;
assign w52885 = pi04409 & w3562;
assign w52886 = pi04367 & w3146;
assign w52887 = pi03653 & w3260;
assign w52888 = pi03757 & w3526;
assign w52889 = pi02457 & w3478;
assign w52890 = pi08413 & w3408;
assign w52891 = pi01653 & w3256;
assign w52892 = pi01612 & w3374;
assign w52893 = pi09560 & w3366;
assign w52894 = pi02423 & w3508;
assign w52895 = pi03686 & w3310;
assign w52896 = pi07390 & w3448;
assign w52897 = pi09778 & w3378;
assign w52898 = pi01743 & w3135;
assign w52899 = pi03992 & w3394;
assign w52900 = pi07935 & w3312;
assign w52901 = pi03351 & w3470;
assign w52902 = pi02441 & w3282;
assign w52903 = ~w52647 & ~w52648;
assign w52904 = ~w52649 & ~w52650;
assign w52905 = ~w52651 & ~w52652;
assign w52906 = ~w52653 & ~w52654;
assign w52907 = ~w52655 & ~w52656;
assign w52908 = ~w52657 & ~w52658;
assign w52909 = ~w52659 & ~w52660;
assign w52910 = ~w52661 & ~w52662;
assign w52911 = ~w52663 & ~w52664;
assign w52912 = ~w52665 & ~w52666;
assign w52913 = ~w52667 & ~w52668;
assign w52914 = ~w52669 & ~w52670;
assign w52915 = ~w52671 & ~w52672;
assign w52916 = ~w52673 & ~w52674;
assign w52917 = ~w52675 & ~w52676;
assign w52918 = ~w52677 & ~w52678;
assign w52919 = ~w52679 & ~w52680;
assign w52920 = ~w52681 & ~w52682;
assign w52921 = ~w52683 & ~w52684;
assign w52922 = ~w52685 & ~w52686;
assign w52923 = ~w52687 & ~w52688;
assign w52924 = ~w52689 & ~w52690;
assign w52925 = ~w52691 & ~w52692;
assign w52926 = ~w52693 & ~w52694;
assign w52927 = ~w52695 & ~w52696;
assign w52928 = ~w52697 & ~w52698;
assign w52929 = ~w52699 & ~w52700;
assign w52930 = ~w52701 & ~w52702;
assign w52931 = ~w52703 & ~w52704;
assign w52932 = ~w52705 & ~w52706;
assign w52933 = ~w52707 & ~w52708;
assign w52934 = ~w52709 & ~w52710;
assign w52935 = ~w52711 & ~w52712;
assign w52936 = ~w52713 & ~w52714;
assign w52937 = ~w52715 & ~w52716;
assign w52938 = ~w52717 & ~w52718;
assign w52939 = ~w52719 & ~w52720;
assign w52940 = ~w52721 & ~w52722;
assign w52941 = ~w52723 & ~w52724;
assign w52942 = ~w52725 & ~w52726;
assign w52943 = ~w52727 & ~w52728;
assign w52944 = ~w52729 & ~w52730;
assign w52945 = ~w52731 & ~w52732;
assign w52946 = ~w52733 & ~w52734;
assign w52947 = ~w52735 & ~w52736;
assign w52948 = ~w52737 & ~w52738;
assign w52949 = ~w52739 & ~w52740;
assign w52950 = ~w52741 & ~w52742;
assign w52951 = ~w52743 & ~w52744;
assign w52952 = ~w52745 & ~w52746;
assign w52953 = ~w52747 & ~w52748;
assign w52954 = ~w52749 & ~w52750;
assign w52955 = ~w52751 & ~w52752;
assign w52956 = ~w52753 & ~w52754;
assign w52957 = ~w52755 & ~w52756;
assign w52958 = ~w52757 & ~w52758;
assign w52959 = ~w52759 & ~w52760;
assign w52960 = ~w52761 & ~w52762;
assign w52961 = ~w52763 & ~w52764;
assign w52962 = ~w52765 & ~w52766;
assign w52963 = ~w52767 & ~w52768;
assign w52964 = ~w52769 & ~w52770;
assign w52965 = ~w52771 & ~w52772;
assign w52966 = ~w52773 & ~w52774;
assign w52967 = ~w52775 & ~w52776;
assign w52968 = ~w52777 & ~w52778;
assign w52969 = ~w52779 & ~w52780;
assign w52970 = ~w52781 & ~w52782;
assign w52971 = ~w52783 & ~w52784;
assign w52972 = ~w52785 & ~w52786;
assign w52973 = ~w52787 & ~w52788;
assign w52974 = ~w52789 & ~w52790;
assign w52975 = ~w52791 & ~w52792;
assign w52976 = ~w52793 & ~w52794;
assign w52977 = ~w52795 & ~w52796;
assign w52978 = ~w52797 & ~w52798;
assign w52979 = ~w52799 & ~w52800;
assign w52980 = ~w52801 & ~w52802;
assign w52981 = ~w52803 & ~w52804;
assign w52982 = ~w52805 & ~w52806;
assign w52983 = ~w52807 & ~w52808;
assign w52984 = ~w52809 & ~w52810;
assign w52985 = ~w52811 & ~w52812;
assign w52986 = ~w52813 & ~w52814;
assign w52987 = ~w52815 & ~w52816;
assign w52988 = ~w52817 & ~w52818;
assign w52989 = ~w52819 & ~w52820;
assign w52990 = ~w52821 & ~w52822;
assign w52991 = ~w52823 & ~w52824;
assign w52992 = ~w52825 & ~w52826;
assign w52993 = ~w52827 & ~w52828;
assign w52994 = ~w52829 & ~w52830;
assign w52995 = ~w52831 & ~w52832;
assign w52996 = ~w52833 & ~w52834;
assign w52997 = ~w52835 & ~w52836;
assign w52998 = ~w52837 & ~w52838;
assign w52999 = ~w52839 & ~w52840;
assign w53000 = ~w52841 & ~w52842;
assign w53001 = ~w52843 & ~w52844;
assign w53002 = ~w52845 & ~w52846;
assign w53003 = ~w52847 & ~w52848;
assign w53004 = ~w52849 & ~w52850;
assign w53005 = ~w52851 & ~w52852;
assign w53006 = ~w52853 & ~w52854;
assign w53007 = ~w52855 & ~w52856;
assign w53008 = ~w52857 & ~w52858;
assign w53009 = ~w52859 & ~w52860;
assign w53010 = ~w52861 & ~w52862;
assign w53011 = ~w52863 & ~w52864;
assign w53012 = ~w52865 & ~w52866;
assign w53013 = ~w52867 & ~w52868;
assign w53014 = ~w52869 & ~w52870;
assign w53015 = ~w52871 & ~w52872;
assign w53016 = ~w52873 & ~w52874;
assign w53017 = ~w52875 & ~w52876;
assign w53018 = ~w52877 & ~w52878;
assign w53019 = ~w52879 & ~w52880;
assign w53020 = ~w52881 & ~w52882;
assign w53021 = ~w52883 & ~w52884;
assign w53022 = ~w52885 & ~w52886;
assign w53023 = ~w52887 & ~w52888;
assign w53024 = ~w52889 & ~w52890;
assign w53025 = ~w52891 & ~w52892;
assign w53026 = ~w52893 & ~w52894;
assign w53027 = ~w52895 & ~w52896;
assign w53028 = ~w52897 & ~w52898;
assign w53029 = ~w52899 & ~w52900;
assign w53030 = ~w52901 & ~w52902;
assign w53031 = w53029 & w53030;
assign w53032 = w53027 & w53028;
assign w53033 = w53025 & w53026;
assign w53034 = w53023 & w53024;
assign w53035 = w53021 & w53022;
assign w53036 = w53019 & w53020;
assign w53037 = w53017 & w53018;
assign w53038 = w53015 & w53016;
assign w53039 = w53013 & w53014;
assign w53040 = w53011 & w53012;
assign w53041 = w53009 & w53010;
assign w53042 = w53007 & w53008;
assign w53043 = w53005 & w53006;
assign w53044 = w53003 & w53004;
assign w53045 = w53001 & w53002;
assign w53046 = w52999 & w53000;
assign w53047 = w52997 & w52998;
assign w53048 = w52995 & w52996;
assign w53049 = w52993 & w52994;
assign w53050 = w52991 & w52992;
assign w53051 = w52989 & w52990;
assign w53052 = w52987 & w52988;
assign w53053 = w52985 & w52986;
assign w53054 = w52983 & w52984;
assign w53055 = w52981 & w52982;
assign w53056 = w52979 & w52980;
assign w53057 = w52977 & w52978;
assign w53058 = w52975 & w52976;
assign w53059 = w52973 & w52974;
assign w53060 = w52971 & w52972;
assign w53061 = w52969 & w52970;
assign w53062 = w52967 & w52968;
assign w53063 = w52965 & w52966;
assign w53064 = w52963 & w52964;
assign w53065 = w52961 & w52962;
assign w53066 = w52959 & w52960;
assign w53067 = w52957 & w52958;
assign w53068 = w52955 & w52956;
assign w53069 = w52953 & w52954;
assign w53070 = w52951 & w52952;
assign w53071 = w52949 & w52950;
assign w53072 = w52947 & w52948;
assign w53073 = w52945 & w52946;
assign w53074 = w52943 & w52944;
assign w53075 = w52941 & w52942;
assign w53076 = w52939 & w52940;
assign w53077 = w52937 & w52938;
assign w53078 = w52935 & w52936;
assign w53079 = w52933 & w52934;
assign w53080 = w52931 & w52932;
assign w53081 = w52929 & w52930;
assign w53082 = w52927 & w52928;
assign w53083 = w52925 & w52926;
assign w53084 = w52923 & w52924;
assign w53085 = w52921 & w52922;
assign w53086 = w52919 & w52920;
assign w53087 = w52917 & w52918;
assign w53088 = w52915 & w52916;
assign w53089 = w52913 & w52914;
assign w53090 = w52911 & w52912;
assign w53091 = w52909 & w52910;
assign w53092 = w52907 & w52908;
assign w53093 = w52905 & w52906;
assign w53094 = w52903 & w52904;
assign w53095 = w53093 & w53094;
assign w53096 = w53091 & w53092;
assign w53097 = w53089 & w53090;
assign w53098 = w53087 & w53088;
assign w53099 = w53085 & w53086;
assign w53100 = w53083 & w53084;
assign w53101 = w53081 & w53082;
assign w53102 = w53079 & w53080;
assign w53103 = w53077 & w53078;
assign w53104 = w53075 & w53076;
assign w53105 = w53073 & w53074;
assign w53106 = w53071 & w53072;
assign w53107 = w53069 & w53070;
assign w53108 = w53067 & w53068;
assign w53109 = w53065 & w53066;
assign w53110 = w53063 & w53064;
assign w53111 = w53061 & w53062;
assign w53112 = w53059 & w53060;
assign w53113 = w53057 & w53058;
assign w53114 = w53055 & w53056;
assign w53115 = w53053 & w53054;
assign w53116 = w53051 & w53052;
assign w53117 = w53049 & w53050;
assign w53118 = w53047 & w53048;
assign w53119 = w53045 & w53046;
assign w53120 = w53043 & w53044;
assign w53121 = w53041 & w53042;
assign w53122 = w53039 & w53040;
assign w53123 = w53037 & w53038;
assign w53124 = w53035 & w53036;
assign w53125 = w53033 & w53034;
assign w53126 = w53031 & w53032;
assign w53127 = w53125 & w53126;
assign w53128 = w53123 & w53124;
assign w53129 = w53121 & w53122;
assign w53130 = w53119 & w53120;
assign w53131 = w53117 & w53118;
assign w53132 = w53115 & w53116;
assign w53133 = w53113 & w53114;
assign w53134 = w53111 & w53112;
assign w53135 = w53109 & w53110;
assign w53136 = w53107 & w53108;
assign w53137 = w53105 & w53106;
assign w53138 = w53103 & w53104;
assign w53139 = w53101 & w53102;
assign w53140 = w53099 & w53100;
assign w53141 = w53097 & w53098;
assign w53142 = w53095 & w53096;
assign w53143 = w53141 & w53142;
assign w53144 = w53139 & w53140;
assign w53145 = w53137 & w53138;
assign w53146 = w53135 & w53136;
assign w53147 = w53133 & w53134;
assign w53148 = w53131 & w53132;
assign w53149 = w53129 & w53130;
assign w53150 = w53127 & w53128;
assign w53151 = w53149 & w53150;
assign w53152 = w53147 & w53148;
assign w53153 = w53145 & w53146;
assign w53154 = w53143 & w53144;
assign w53155 = w53153 & w53154;
assign w53156 = w53151 & w53152;
assign w53157 = w53155 & w53156;
assign w53158 = ~pi10577 & ~w53157;
assign w53159 = pi04973 & w3562;
assign w53160 = pi05065 & w3582;
assign w53161 = pi05012 & w3504;
assign w53162 = pi01534 & w3580;
assign w53163 = pi08783 & w3384;
assign w53164 = pi01543 & w3096;
assign w53165 = pi08687 & w3227;
assign w53166 = pi01548 & w3566;
assign w53167 = pi04715 & w3310;
assign w53168 = pi04788 & w3592;
assign w53169 = pi05045 & w3588;
assign w53170 = pi08466 & w3308;
assign w53171 = pi04722 & w3244;
assign w53172 = pi01650 & w3320;
assign w53173 = pi04842 & w3428;
assign w53174 = pi02500 & w3372;
assign w53175 = pi02490 & w3173;
assign w53176 = pi04618 & w3250;
assign w53177 = pi04794 & w3498;
assign w53178 = pi09421 & w3158;
assign w53179 = pi01528 & w3318;
assign w53180 = pi04683 & w3137;
assign w53181 = pi01916 & w3468;
assign w53182 = pi02483 & w3374;
assign w53183 = pi08615 & w3314;
assign w53184 = pi05032 & w3388;
assign w53185 = pi02487 & w3518;
assign w53186 = pi09775 & w3286;
assign w53187 = pi04921 & w3328;
assign w53188 = pi08545 & w3550;
assign w53189 = pi04808 & w3394;
assign w53190 = pi04835 & w3494;
assign w53191 = pi09777 & w3276;
assign w53192 = pi04689 & w3262;
assign w53193 = pi02600 & w3508;
assign w53194 = pi01592 & w3402;
assign w53195 = pi01564 & w3596;
assign w53196 = pi02593 & w3093;
assign w53197 = pi09196 & w3175;
assign w53198 = pi01503 & w3332;
assign w53199 = pi05005 & w3162;
assign w53200 = pi02550 & w3112;
assign w53201 = pi04801 & w3132;
assign w53202 = pi04702 & w3260;
assign w53203 = pi04527 & w3380;
assign w53204 = pi02563 & w3410;
assign w53205 = pi09434 & w3578;
assign w53206 = pi08484 & w3598;
assign w53207 = pi09487 & w3110;
assign w53208 = pi04735 & w3490;
assign w53209 = pi04534 & w3294;
assign w53210 = pi05431 & w3217;
assign w53211 = pi08661 & w3203;
assign w53212 = pi04624 & w3064;
assign w53213 = pi02573 & w3082;
assign w53214 = pi05076 & w3242;
assign w53215 = pi01596 & w3127;
assign w53216 = pi02584 & w3532;
assign w53217 = pi02585 & w3167;
assign w53218 = pi04709 & w3610;
assign w53219 = pi01485 & w3516;
assign w53220 = pi04947 & w3370;
assign w53221 = pi02583 & w3312;
assign w53222 = pi04548 & w3197;
assign w53223 = pi02619 & w3420;
assign w53224 = pi09770 & w3192;
assign w53225 = pi04940 & w3564;
assign w53226 = pi08607 & w3540;
assign w53227 = pi02427 & w3156;
assign w53228 = pi01557 & w3358;
assign w53229 = pi09787 & w3280;
assign w53230 = pi01886 & w3352;
assign w53231 = pi08622 & w3538;
assign w53232 = pi04631 & w3534;
assign w53233 = pi09440 & w3179;
assign w53234 = pi05058 & w3211;
assign w53235 = pi04676 & w3296;
assign w53236 = pi02767 & w3219;
assign w53237 = pi09501 & w3558;
assign w53238 = pi04979 & w3169;
assign w53239 = pi01586 & w3376;
assign w53240 = pi08505 & w3492;
assign w53241 = pi09466 & w3524;
assign w53242 = pi02467 & w3324;
assign w53243 = pi02549 & w3078;
assign w53244 = pi08641 & w3298;
assign w53245 = pi02570 & w3360;
assign w53246 = pi04754 & w3576;
assign w53247 = pi02493 & w3382;
assign w53248 = pi01579 & w3476;
assign w53249 = pi08471 & w3436;
assign w53250 = pi05026 & w3556;
assign w53251 = pi02589 & w3616;
assign w53252 = pi01738 & w3608;
assign w53253 = pi04741 & w3526;
assign w53254 = pi05427 & w3460;
assign w53255 = pi01563 & w3542;
assign w53256 = pi08713 & w3153;
assign w53257 = pi01498 & w3560;
assign w53258 = pi04670 & w3424;
assign w53259 = pi02623 & w3390;
assign w53260 = pi09447 & w3438;
assign w53261 = pi02330 & w3594;
assign w53262 = pi01632 & w3264;
assign w53263 = pi01562 & w3466;
assign w53264 = pi04868 & w3454;
assign w53265 = pi01749 & w3106;
assign w53266 = pi02621 & w3238;
assign w53267 = pi01945 & w3254;
assign w53268 = pi01899 & w3300;
assign w53269 = pi04848 & w3522;
assign w53270 = pi02452 & w3148;
assign w53271 = pi02567 & w3165;
assign w53272 = pi01845 & w3478;
assign w53273 = pi04696 & w3292;
assign w53274 = pi02480 & w3364;
assign w53275 = pi09242 & w3229;
assign w53276 = pi04637 & w3400;
assign w53277 = pi08434 & w3486;
assign w53278 = pi04815 & w3071;
assign w53279 = pi08600 & w3414;
assign w53280 = pi04953 & w3618;
assign w53281 = pi04592 & w3362;
assign w53282 = pi09514 & w3510;
assign w53283 = pi08493 & w3604;
assign w53284 = pi08717 & w3554;
assign w53285 = pi02554 & w3284;
assign w53286 = pi01846 & w3398;
assign w53287 = pi02596 & w3135;
assign w53288 = pi04781 & w3456;
assign w53289 = pi08693 & w3304;
assign w53290 = pi04535 & w3346;
assign w53291 = pi01844 & w3430;
assign w53292 = pi08611 & w3482;
assign w53293 = pi02806 & w3440;
assign w53294 = pi09792 & w3125;
assign w53295 = pi05052 & w3396;
assign w53296 = pi01870 & w3205;
assign w53297 = pi08648 & w3354;
assign w53298 = pi08441 & w3232;
assign w53299 = pi01928 & w3194;
assign w53300 = pi04855 & w3181;
assign w53301 = pi04579 & w3416;
assign w53302 = pi02528 & w3356;
assign w53303 = pi08578 & w3378;
assign w53304 = pi01915 & w3506;
assign w53305 = pi02611 & w3464;
assign w53306 = pi04927 & w3484;
assign w53307 = pi08549 & w3568;
assign w53308 = pi04861 & w3502;
assign w53309 = pi01594 & w3272;
assign w53310 = pi01966 & w3600;
assign w53311 = pi02421 & w3366;
assign w53312 = pi04992 & w3258;
assign w53313 = pi04966 & w3412;
assign w53314 = pi02604 & w3514;
assign w53315 = pi04821 & w3118;
assign w53316 = pi08635 & w3236;
assign w53317 = pi04586 & w3470;
assign w53318 = pi01857 & w3472;
assign w53319 = pi04520 & w3306;
assign w53320 = pi04960 & w3512;
assign w53321 = pi08700 & w3462;
assign w53322 = pi01923 & w3225;
assign w53323 = pi08447 & w3240;
assign w53324 = pi01840 & w3221;
assign w53325 = pi04402 & w3552;
assign w53326 = pi04542 & w3520;
assign w53327 = pi01607 & w3234;
assign w53328 = pi08706 & w3496;
assign w53329 = pi04895 & w3214;
assign w53330 = pi09534 & w3342;
assign w53331 = pi04875 & w3290;
assign w53332 = pi02576 & w3288;
assign w53333 = pi08628 & w3450;
assign w53334 = pi04598 & w3404;
assign w53335 = pi04611 & w3530;
assign w53336 = pi04888 & w3334;
assign w53337 = pi04514 & w3614;
assign w53338 = pi04657 & w3274;
assign w53339 = pi02607 & w3278;
assign w53340 = pi08680 & w3422;
assign w53341 = pi04901 & w3086;
assign w53342 = pi01582 & w3546;
assign w53343 = pi03324 & w3500;
assign w53344 = pi09554 & w3606;
assign w53345 = pi05039 & w3177;
assign w53346 = pi04882 & w3326;
assign w53347 = pi09453 & w3368;
assign w53348 = pi01773 & w3282;
assign w53349 = pi09493 & w3150;
assign w53350 = pi04559 & w3544;
assign w53351 = pi05292 & w3528;
assign w53352 = pi04748 & w3350;
assign w53353 = pi09460 & w3160;
assign w53354 = pi01527 & w3572;
assign w53355 = pi01581 & w3171;
assign w53356 = pi04663 & w3536;
assign w53357 = pi04572 & w3268;
assign w53358 = pi02592 & w3186;
assign w53359 = pi04914 & w3190;
assign w53360 = pi09427 & w3602;
assign w53361 = pi01919 & w3432;
assign w53362 = pi02551 & w3426;
assign w53363 = pi09474 & w3418;
assign w53364 = pi01566 & w3406;
assign w53365 = pi01532 & w3442;
assign w53366 = pi05817 & w3143;
assign w53367 = pi02502 & w3256;
assign w53368 = pi04908 & w3115;
assign w53369 = pi01584 & w3139;
assign w53370 = pi09524 & w3570;
assign w53371 = pi08499 & w3344;
assign w53372 = pi03483 & w3316;
assign w53373 = pi02608 & w3207;
assign w53374 = pi08454 & w3266;
assign w53375 = pi04999 & w3122;
assign w53376 = pi01708 & w3446;
assign w53377 = pi04934 & w3146;
assign w53378 = pi08560 & w3480;
assign w53379 = pi02590 & w3434;
assign w53380 = pi04728 & w3548;
assign w53381 = pi01544 & w3340;
assign w53382 = pi02571 & w3458;
assign w53383 = pi08596 & w3586;
assign w53384 = pi08674 & w3199;
assign w53385 = pi08517 & w3252;
assign w53386 = pi04650 & w3103;
assign w53387 = pi04829 & w3574;
assign w53388 = pi05071 & w3488;
assign w53389 = pi09507 & w3408;
assign w53390 = pi04761 & w3209;
assign w53391 = pi02558 & w3201;
assign w53392 = pi08654 & w3392;
assign w53393 = pi04554 & w3336;
assign w53394 = pi09480 & w3246;
assign w53395 = pi04605 & w3330;
assign w53396 = pi05019 & w3184;
assign w53397 = pi08533 & w3452;
assign w53398 = pi02555 & w3386;
assign w53399 = pi02603 & w3270;
assign w53400 = pi01868 & w3584;
assign w53401 = pi08511 & w3612;
assign w53402 = pi02306 & w3444;
assign w53403 = pi04775 & w3348;
assign w53404 = pi09650 & w3188;
assign w53405 = pi01709 & w3620;
assign w53406 = pi01912 & w3590;
assign w53407 = pi09181 & w3474;
assign w53408 = pi01546 & w3448;
assign w53409 = pi04644 & w3322;
assign w53410 = pi08667 & w3129;
assign w53411 = pi08479 & w3248;
assign w53412 = pi04986 & w3302;
assign w53413 = pi04767 & w3338;
assign w53414 = pi05373 & w3223;
assign w53415 = ~w53159 & ~w53160;
assign w53416 = ~w53161 & ~w53162;
assign w53417 = ~w53163 & ~w53164;
assign w53418 = ~w53165 & ~w53166;
assign w53419 = ~w53167 & ~w53168;
assign w53420 = ~w53169 & ~w53170;
assign w53421 = ~w53171 & ~w53172;
assign w53422 = ~w53173 & ~w53174;
assign w53423 = ~w53175 & ~w53176;
assign w53424 = ~w53177 & ~w53178;
assign w53425 = ~w53179 & ~w53180;
assign w53426 = ~w53181 & ~w53182;
assign w53427 = ~w53183 & ~w53184;
assign w53428 = ~w53185 & ~w53186;
assign w53429 = ~w53187 & ~w53188;
assign w53430 = ~w53189 & ~w53190;
assign w53431 = ~w53191 & ~w53192;
assign w53432 = ~w53193 & ~w53194;
assign w53433 = ~w53195 & ~w53196;
assign w53434 = ~w53197 & ~w53198;
assign w53435 = ~w53199 & ~w53200;
assign w53436 = ~w53201 & ~w53202;
assign w53437 = ~w53203 & ~w53204;
assign w53438 = ~w53205 & ~w53206;
assign w53439 = ~w53207 & ~w53208;
assign w53440 = ~w53209 & ~w53210;
assign w53441 = ~w53211 & ~w53212;
assign w53442 = ~w53213 & ~w53214;
assign w53443 = ~w53215 & ~w53216;
assign w53444 = ~w53217 & ~w53218;
assign w53445 = ~w53219 & ~w53220;
assign w53446 = ~w53221 & ~w53222;
assign w53447 = ~w53223 & ~w53224;
assign w53448 = ~w53225 & ~w53226;
assign w53449 = ~w53227 & ~w53228;
assign w53450 = ~w53229 & ~w53230;
assign w53451 = ~w53231 & ~w53232;
assign w53452 = ~w53233 & ~w53234;
assign w53453 = ~w53235 & ~w53236;
assign w53454 = ~w53237 & ~w53238;
assign w53455 = ~w53239 & ~w53240;
assign w53456 = ~w53241 & ~w53242;
assign w53457 = ~w53243 & ~w53244;
assign w53458 = ~w53245 & ~w53246;
assign w53459 = ~w53247 & ~w53248;
assign w53460 = ~w53249 & ~w53250;
assign w53461 = ~w53251 & ~w53252;
assign w53462 = ~w53253 & ~w53254;
assign w53463 = ~w53255 & ~w53256;
assign w53464 = ~w53257 & ~w53258;
assign w53465 = ~w53259 & ~w53260;
assign w53466 = ~w53261 & ~w53262;
assign w53467 = ~w53263 & ~w53264;
assign w53468 = ~w53265 & ~w53266;
assign w53469 = ~w53267 & ~w53268;
assign w53470 = ~w53269 & ~w53270;
assign w53471 = ~w53271 & ~w53272;
assign w53472 = ~w53273 & ~w53274;
assign w53473 = ~w53275 & ~w53276;
assign w53474 = ~w53277 & ~w53278;
assign w53475 = ~w53279 & ~w53280;
assign w53476 = ~w53281 & ~w53282;
assign w53477 = ~w53283 & ~w53284;
assign w53478 = ~w53285 & ~w53286;
assign w53479 = ~w53287 & ~w53288;
assign w53480 = ~w53289 & ~w53290;
assign w53481 = ~w53291 & ~w53292;
assign w53482 = ~w53293 & ~w53294;
assign w53483 = ~w53295 & ~w53296;
assign w53484 = ~w53297 & ~w53298;
assign w53485 = ~w53299 & ~w53300;
assign w53486 = ~w53301 & ~w53302;
assign w53487 = ~w53303 & ~w53304;
assign w53488 = ~w53305 & ~w53306;
assign w53489 = ~w53307 & ~w53308;
assign w53490 = ~w53309 & ~w53310;
assign w53491 = ~w53311 & ~w53312;
assign w53492 = ~w53313 & ~w53314;
assign w53493 = ~w53315 & ~w53316;
assign w53494 = ~w53317 & ~w53318;
assign w53495 = ~w53319 & ~w53320;
assign w53496 = ~w53321 & ~w53322;
assign w53497 = ~w53323 & ~w53324;
assign w53498 = ~w53325 & ~w53326;
assign w53499 = ~w53327 & ~w53328;
assign w53500 = ~w53329 & ~w53330;
assign w53501 = ~w53331 & ~w53332;
assign w53502 = ~w53333 & ~w53334;
assign w53503 = ~w53335 & ~w53336;
assign w53504 = ~w53337 & ~w53338;
assign w53505 = ~w53339 & ~w53340;
assign w53506 = ~w53341 & ~w53342;
assign w53507 = ~w53343 & ~w53344;
assign w53508 = ~w53345 & ~w53346;
assign w53509 = ~w53347 & ~w53348;
assign w53510 = ~w53349 & ~w53350;
assign w53511 = ~w53351 & ~w53352;
assign w53512 = ~w53353 & ~w53354;
assign w53513 = ~w53355 & ~w53356;
assign w53514 = ~w53357 & ~w53358;
assign w53515 = ~w53359 & ~w53360;
assign w53516 = ~w53361 & ~w53362;
assign w53517 = ~w53363 & ~w53364;
assign w53518 = ~w53365 & ~w53366;
assign w53519 = ~w53367 & ~w53368;
assign w53520 = ~w53369 & ~w53370;
assign w53521 = ~w53371 & ~w53372;
assign w53522 = ~w53373 & ~w53374;
assign w53523 = ~w53375 & ~w53376;
assign w53524 = ~w53377 & ~w53378;
assign w53525 = ~w53379 & ~w53380;
assign w53526 = ~w53381 & ~w53382;
assign w53527 = ~w53383 & ~w53384;
assign w53528 = ~w53385 & ~w53386;
assign w53529 = ~w53387 & ~w53388;
assign w53530 = ~w53389 & ~w53390;
assign w53531 = ~w53391 & ~w53392;
assign w53532 = ~w53393 & ~w53394;
assign w53533 = ~w53395 & ~w53396;
assign w53534 = ~w53397 & ~w53398;
assign w53535 = ~w53399 & ~w53400;
assign w53536 = ~w53401 & ~w53402;
assign w53537 = ~w53403 & ~w53404;
assign w53538 = ~w53405 & ~w53406;
assign w53539 = ~w53407 & ~w53408;
assign w53540 = ~w53409 & ~w53410;
assign w53541 = ~w53411 & ~w53412;
assign w53542 = ~w53413 & ~w53414;
assign w53543 = w53541 & w53542;
assign w53544 = w53539 & w53540;
assign w53545 = w53537 & w53538;
assign w53546 = w53535 & w53536;
assign w53547 = w53533 & w53534;
assign w53548 = w53531 & w53532;
assign w53549 = w53529 & w53530;
assign w53550 = w53527 & w53528;
assign w53551 = w53525 & w53526;
assign w53552 = w53523 & w53524;
assign w53553 = w53521 & w53522;
assign w53554 = w53519 & w53520;
assign w53555 = w53517 & w53518;
assign w53556 = w53515 & w53516;
assign w53557 = w53513 & w53514;
assign w53558 = w53511 & w53512;
assign w53559 = w53509 & w53510;
assign w53560 = w53507 & w53508;
assign w53561 = w53505 & w53506;
assign w53562 = w53503 & w53504;
assign w53563 = w53501 & w53502;
assign w53564 = w53499 & w53500;
assign w53565 = w53497 & w53498;
assign w53566 = w53495 & w53496;
assign w53567 = w53493 & w53494;
assign w53568 = w53491 & w53492;
assign w53569 = w53489 & w53490;
assign w53570 = w53487 & w53488;
assign w53571 = w53485 & w53486;
assign w53572 = w53483 & w53484;
assign w53573 = w53481 & w53482;
assign w53574 = w53479 & w53480;
assign w53575 = w53477 & w53478;
assign w53576 = w53475 & w53476;
assign w53577 = w53473 & w53474;
assign w53578 = w53471 & w53472;
assign w53579 = w53469 & w53470;
assign w53580 = w53467 & w53468;
assign w53581 = w53465 & w53466;
assign w53582 = w53463 & w53464;
assign w53583 = w53461 & w53462;
assign w53584 = w53459 & w53460;
assign w53585 = w53457 & w53458;
assign w53586 = w53455 & w53456;
assign w53587 = w53453 & w53454;
assign w53588 = w53451 & w53452;
assign w53589 = w53449 & w53450;
assign w53590 = w53447 & w53448;
assign w53591 = w53445 & w53446;
assign w53592 = w53443 & w53444;
assign w53593 = w53441 & w53442;
assign w53594 = w53439 & w53440;
assign w53595 = w53437 & w53438;
assign w53596 = w53435 & w53436;
assign w53597 = w53433 & w53434;
assign w53598 = w53431 & w53432;
assign w53599 = w53429 & w53430;
assign w53600 = w53427 & w53428;
assign w53601 = w53425 & w53426;
assign w53602 = w53423 & w53424;
assign w53603 = w53421 & w53422;
assign w53604 = w53419 & w53420;
assign w53605 = w53417 & w53418;
assign w53606 = w53415 & w53416;
assign w53607 = w53605 & w53606;
assign w53608 = w53603 & w53604;
assign w53609 = w53601 & w53602;
assign w53610 = w53599 & w53600;
assign w53611 = w53597 & w53598;
assign w53612 = w53595 & w53596;
assign w53613 = w53593 & w53594;
assign w53614 = w53591 & w53592;
assign w53615 = w53589 & w53590;
assign w53616 = w53587 & w53588;
assign w53617 = w53585 & w53586;
assign w53618 = w53583 & w53584;
assign w53619 = w53581 & w53582;
assign w53620 = w53579 & w53580;
assign w53621 = w53577 & w53578;
assign w53622 = w53575 & w53576;
assign w53623 = w53573 & w53574;
assign w53624 = w53571 & w53572;
assign w53625 = w53569 & w53570;
assign w53626 = w53567 & w53568;
assign w53627 = w53565 & w53566;
assign w53628 = w53563 & w53564;
assign w53629 = w53561 & w53562;
assign w53630 = w53559 & w53560;
assign w53631 = w53557 & w53558;
assign w53632 = w53555 & w53556;
assign w53633 = w53553 & w53554;
assign w53634 = w53551 & w53552;
assign w53635 = w53549 & w53550;
assign w53636 = w53547 & w53548;
assign w53637 = w53545 & w53546;
assign w53638 = w53543 & w53544;
assign w53639 = w53637 & w53638;
assign w53640 = w53635 & w53636;
assign w53641 = w53633 & w53634;
assign w53642 = w53631 & w53632;
assign w53643 = w53629 & w53630;
assign w53644 = w53627 & w53628;
assign w53645 = w53625 & w53626;
assign w53646 = w53623 & w53624;
assign w53647 = w53621 & w53622;
assign w53648 = w53619 & w53620;
assign w53649 = w53617 & w53618;
assign w53650 = w53615 & w53616;
assign w53651 = w53613 & w53614;
assign w53652 = w53611 & w53612;
assign w53653 = w53609 & w53610;
assign w53654 = w53607 & w53608;
assign w53655 = w53653 & w53654;
assign w53656 = w53651 & w53652;
assign w53657 = w53649 & w53650;
assign w53658 = w53647 & w53648;
assign w53659 = w53645 & w53646;
assign w53660 = w53643 & w53644;
assign w53661 = w53641 & w53642;
assign w53662 = w53639 & w53640;
assign w53663 = w53661 & w53662;
assign w53664 = w53659 & w53660;
assign w53665 = w53657 & w53658;
assign w53666 = w53655 & w53656;
assign w53667 = w53665 & w53666;
assign w53668 = w53663 & w53664;
assign w53669 = w53667 & w53668;
assign w53670 = ~pi10577 & ~w53669;
assign w53671 = pi08210 & w3282;
assign w53672 = pi06140 & w3217;
assign w53673 = pi08401 & w3150;
assign w53674 = pi03266 & w3268;
assign w53675 = pi01674 & w3354;
assign w53676 = pi08355 & w3438;
assign w53677 = pi08374 & w3524;
assign w53678 = pi09632 & w3464;
assign w53679 = pi07209 & w3205;
assign w53680 = pi07442 & w3434;
assign w53681 = pi01971 & w3548;
assign w53682 = pi02134 & w3588;
assign w53683 = pi09600 & w3574;
assign w53684 = pi08341 & w3578;
assign w53685 = pi02016 & w3292;
assign w53686 = pi08420 & w3510;
assign w53687 = pi07481 & w3167;
assign w53688 = pi05732 & w3266;
assign w53689 = pi06937 & w3234;
assign w53690 = pi05944 & w3492;
assign w53691 = pi06790 & w3078;
assign w53692 = pi02120 & w3396;
assign w53693 = pi05924 & w3344;
assign w53694 = pi07394 & w3448;
assign w53695 = pi07234 & w3225;
assign w53696 = pi08263 & w3402;
assign w53697 = pi08165 & w3468;
assign w53698 = pi06028 & w3554;
assign w53699 = pi07892 & w3352;
assign w53700 = pi07344 & w3376;
assign w53701 = pi03179 & w3380;
assign w53702 = pi08348 & w3179;
assign w53703 = pi07005 & w3572;
assign w53704 = pi06924 & w3398;
assign w53705 = pi02809 & w3516;
assign w53706 = pi05796 & w3308;
assign w53707 = pi01956 & w3490;
assign w53708 = pi07968 & w3238;
assign w53709 = pi07913 & w3596;
assign w53710 = pi02112 & w3211;
assign w53711 = pi08368 & w3160;
assign w53712 = pi02232 & w3512;
assign w53713 = pi08335 & w3602;
assign w53714 = pi02200 & w3258;
assign w53715 = pi02122 & w3223;
assign w53716 = pi02367 & w3232;
assign w53717 = pi08223 & w3546;
assign w53718 = pi07678 & w3590;
assign w53719 = pi02266 & w3146;
assign w53720 = pi08158 & w3594;
assign w53721 = pi06731 & w3514;
assign w53722 = pi02117 & w3582;
assign w53723 = pi09663 & w3394;
assign w53724 = pi02760 & w3290;
assign w53725 = pi06088 & w3568;
assign w53726 = pi02059 & w3400;
assign w53727 = pi03780 & w3350;
assign w53728 = pi07287 & w3221;
assign w53729 = pi02030 & w3536;
assign w53730 = pi01614 & w3606;
assign w53731 = pi07498 & w3312;
assign w53732 = pi06536 & w3304;
assign w53733 = pi02778 & w3454;
assign w53734 = pi09797 & w3620;
assign w53735 = pi06501 & w3422;
assign w53736 = pi07611 & w3374;
assign w53737 = pi04454 & w3184;
assign w53738 = pi02617 & w3334;
assign w53739 = pi03450 & w3530;
assign w53740 = pi01977 & w3310;
assign w53741 = pi03505 & w3534;
assign w53742 = pi03212 & w3197;
assign w53743 = pi02224 & w3412;
assign w53744 = pi02269 & w3484;
assign w53745 = pi08191 & w3444;
assign w53746 = pi09698 & w3498;
assign w53747 = pi07981 & w3426;
assign w53748 = pi01620 & w3338;
assign w53749 = pi07854 & w3386;
assign w53750 = pi08315 & w3324;
assign w53751 = pi02508 & w3214;
assign w53752 = pi06356 & w3450;
assign w53753 = pi08244 & w3096;
assign w53754 = pi06455 & w3129;
assign w53755 = pi08322 & w3332;
assign w53756 = pi05877 & w3604;
assign w53757 = pi02158 & w3504;
assign w53758 = pi02140 & w3177;
assign w53759 = pi09677 & w3132;
assign w53760 = pi06327 & w3538;
assign w53761 = pi01556 & w3440;
assign w53762 = pi02072 & w3064;
assign w53763 = pi02004 & w3260;
assign w53764 = pi06880 & w3384;
assign w53765 = pi02132 & w3416;
assign w53766 = pi03195 & w3520;
assign w53767 = pi02209 & w3562;
assign w53768 = pi07876 & w3382;
assign w53769 = pi08327 & w3158;
assign w53770 = pi02129 & w3470;
assign w53771 = pi07689 & w3430;
assign w53772 = pi08125 & w3570;
assign w53773 = pi02243 & w3564;
assign w53774 = pi08353 & w3194;
assign w53775 = pi06254 & w3414;
assign w53776 = pi08171 & w3173;
assign w53777 = pi02036 & w3274;
assign w53778 = pi07110 & w3410;
assign w53779 = pi09543 & w3181;
assign w53780 = pi08361 & w3368;
assign w53781 = pi08426 & w3242;
assign w53782 = pi02154 & w3388;
assign w53783 = pi07167 & w3364;
assign w53784 = pi08152 & w3366;
assign w53785 = pi09588 & w3428;
assign w53786 = pi07196 & w3156;
assign w53787 = pi09592 & w3494;
assign w53788 = pi07331 & w3272;
assign w53789 = pi01511 & w3348;
assign w53790 = pi07724 & w3476;
assign w53791 = pi03394 & w3404;
assign w53792 = pi06822 & w3256;
assign w53793 = pi03259 & w3500;
assign w53794 = pi02145 & w3556;
assign w53795 = pi07774 & w3192;
assign w53796 = pi02241 & w3328;
assign w53797 = pi02693 & w3270;
assign w53798 = pi06369 & w3236;
assign w53799 = pi02299 & w3190;
assign w53800 = pi08414 & w3408;
assign w53801 = pi02026 & w3296;
assign w53802 = pi01713 & w3276;
assign w53803 = pi08276 & w3229;
assign w53804 = pi01801 & w3288;
assign w53805 = pi08388 & w3246;
assign w53806 = pi07640 & w3600;
assign w53807 = pi03147 & w3614;
assign w53808 = pi08283 & w3560;
assign w53809 = pi01872 & w3314;
assign w53810 = pi06777 & w3284;
assign w53811 = pi09638 & w3071;
assign w53812 = pi07095 & w3552;
assign w53813 = pi07413 & w3566;
assign w53814 = pi08302 & w3294;
assign w53815 = pi01576 & w3392;
assign w53816 = pi02274 & w3175;
assign w53817 = pi07122 & w3420;
assign w53818 = pi06468 & w3199;
assign w53819 = pi03186 & w3346;
assign w53820 = pi07936 & w3125;
assign w53821 = pi07579 & w3201;
assign w53822 = pi07592 & w3372;
assign w53823 = pi06179 & w3356;
assign w53824 = pi06207 & w3586;
assign w53825 = pi06991 & w3406;
assign w53826 = pi04382 & w3370;
assign w53827 = pi09795 & w3508;
assign w53828 = pi02334 & w3616;
assign w53829 = pi07258 & w3472;
assign w53830 = pi07546 & w3165;
assign w53831 = pi08184 & w3106;
assign w53832 = pi05670 & w3486;
assign w53833 = pi06423 & w3203;
assign w53834 = pi06079 & w3550;
assign w53835 = pi06589 & w3153;
assign w53836 = pi03218 & w3336;
assign w53837 = pi06705 & w3278;
assign w53838 = pi08289 & w3342;
assign w53839 = pi06194 & w3460;
assign w53840 = pi02127 & w3362;
assign w53841 = pi09574 & w3522;
assign w53842 = pi02779 & w3502;
assign w53843 = pi02091 & w3488;
assign w53844 = pi01980 & w3610;
assign w53845 = pi06976 & w3139;
assign w53846 = pi02052 & w3322;
assign w53847 = pi01776 & w3436;
assign w53848 = pi08309 & w3316;
assign w53849 = pi08237 & w3280;
assign w53850 = pi05991 & w3219;
assign w53851 = pi09626 & w3118;
assign w53852 = pi06950 & w3466;
assign w53853 = pi08029 & w3532;
assign w53854 = pi02752 & w3326;
assign w53855 = pi01944 & w3244;
assign w53856 = pi01654 & w3248;
assign w53857 = pi06382 & w3298;
assign w53858 = pi02215 & w3169;
assign w53859 = pi08002 & w3474;
assign w53860 = pi06168 & w3378;
assign w53861 = pi01700 & w3576;
assign w53862 = pi07709 & w3171;
assign w53863 = pi02027 & w3424;
assign w53864 = pi08108 & w3446;
assign w53865 = pi02239 & w3240;
assign w53866 = pi06857 & w3442;
assign w53867 = pi02380 & w3086;
assign w53868 = pi08231 & w3542;
assign w53869 = pi08296 & w3148;
assign w53870 = pi06516 & w3227;
assign w53871 = pi05970 & w3252;
assign w53872 = pi08270 & w3580;
assign w53873 = pi09724 & w3592;
assign w53874 = pi03923 & w3456;
assign w53875 = pi08178 & w3584;
assign w53876 = pi07955 & w3093;
assign w53877 = pi06887 & w3432;
assign w53878 = pi08394 & w3110;
assign w53879 = pi07796 & w3390;
assign w53880 = pi06965 & w3127;
assign w53881 = pi07050 & w3286;
assign w53882 = pi04442 & w3162;
assign w53883 = pi02111 & w3330;
assign w53884 = pi09776 & w3598;
assign w53885 = pi07018 & w3340;
assign w53886 = pi07223 & w3254;
assign w53887 = pi02376 & w3115;
assign w53888 = pi06831 & w3518;
assign w53889 = pi08381 & w3418;
assign w53890 = pi08197 & w3320;
assign w53891 = pi06069 & w3528;
assign w53892 = pi07822 & w3207;
assign w53893 = pi02024 & w3137;
assign w53894 = pi06911 & w3300;
assign w53895 = pi06274 & w3540;
assign w53896 = pi07374 & w3358;
assign w53897 = pi08204 & w3478;
assign w53898 = pi02185 & w3122;
assign w53899 = pi08250 & w3318;
assign w53900 = pi03477 & w3250;
assign w53901 = pi06294 & w3482;
assign w53902 = pi01655 & w3209;
assign w53903 = pi02174 & w3302;
assign w53904 = pi07737 & w3458;
assign w53905 = pi06573 & w3496;
assign w53906 = pi01723 & w3143;
assign w53907 = pi03232 & w3544;
assign w53908 = pi03565 & w3103;
assign w53909 = pi06153 & w3112;
assign w53910 = pi01924 & w3526;
assign w53911 = pi01983 & w3262;
assign w53912 = pi08257 & w3188;
assign w53913 = pi05957 & w3612;
assign w53914 = pi02248 & w3618;
assign w53915 = pi08145 & w3608;
assign w53916 = pi08218 & w3264;
assign w53917 = pi06750 & w3186;
assign w53918 = pi06046 & w3452;
assign w53919 = pi06555 & w3462;
assign w53920 = pi07788 & w3360;
assign w53921 = pi03160 & w3306;
assign w53922 = pi01687 & w3135;
assign w53923 = pi06127 & w3480;
assign w53924 = pi06898 & w3506;
assign w53925 = pi08407 & w3558;
assign w53926 = pi06678 & w3082;
assign w53927 = ~w53671 & ~w53672;
assign w53928 = ~w53673 & ~w53674;
assign w53929 = ~w53675 & ~w53676;
assign w53930 = ~w53677 & ~w53678;
assign w53931 = ~w53679 & ~w53680;
assign w53932 = ~w53681 & ~w53682;
assign w53933 = ~w53683 & ~w53684;
assign w53934 = ~w53685 & ~w53686;
assign w53935 = ~w53687 & ~w53688;
assign w53936 = ~w53689 & ~w53690;
assign w53937 = ~w53691 & ~w53692;
assign w53938 = ~w53693 & ~w53694;
assign w53939 = ~w53695 & ~w53696;
assign w53940 = ~w53697 & ~w53698;
assign w53941 = ~w53699 & ~w53700;
assign w53942 = ~w53701 & ~w53702;
assign w53943 = ~w53703 & ~w53704;
assign w53944 = ~w53705 & ~w53706;
assign w53945 = ~w53707 & ~w53708;
assign w53946 = ~w53709 & ~w53710;
assign w53947 = ~w53711 & ~w53712;
assign w53948 = ~w53713 & ~w53714;
assign w53949 = ~w53715 & ~w53716;
assign w53950 = ~w53717 & ~w53718;
assign w53951 = ~w53719 & ~w53720;
assign w53952 = ~w53721 & ~w53722;
assign w53953 = ~w53723 & ~w53724;
assign w53954 = ~w53725 & ~w53726;
assign w53955 = ~w53727 & ~w53728;
assign w53956 = ~w53729 & ~w53730;
assign w53957 = ~w53731 & ~w53732;
assign w53958 = ~w53733 & ~w53734;
assign w53959 = ~w53735 & ~w53736;
assign w53960 = ~w53737 & ~w53738;
assign w53961 = ~w53739 & ~w53740;
assign w53962 = ~w53741 & ~w53742;
assign w53963 = ~w53743 & ~w53744;
assign w53964 = ~w53745 & ~w53746;
assign w53965 = ~w53747 & ~w53748;
assign w53966 = ~w53749 & ~w53750;
assign w53967 = ~w53751 & ~w53752;
assign w53968 = ~w53753 & ~w53754;
assign w53969 = ~w53755 & ~w53756;
assign w53970 = ~w53757 & ~w53758;
assign w53971 = ~w53759 & ~w53760;
assign w53972 = ~w53761 & ~w53762;
assign w53973 = ~w53763 & ~w53764;
assign w53974 = ~w53765 & ~w53766;
assign w53975 = ~w53767 & ~w53768;
assign w53976 = ~w53769 & ~w53770;
assign w53977 = ~w53771 & ~w53772;
assign w53978 = ~w53773 & ~w53774;
assign w53979 = ~w53775 & ~w53776;
assign w53980 = ~w53777 & ~w53778;
assign w53981 = ~w53779 & ~w53780;
assign w53982 = ~w53781 & ~w53782;
assign w53983 = ~w53783 & ~w53784;
assign w53984 = ~w53785 & ~w53786;
assign w53985 = ~w53787 & ~w53788;
assign w53986 = ~w53789 & ~w53790;
assign w53987 = ~w53791 & ~w53792;
assign w53988 = ~w53793 & ~w53794;
assign w53989 = ~w53795 & ~w53796;
assign w53990 = ~w53797 & ~w53798;
assign w53991 = ~w53799 & ~w53800;
assign w53992 = ~w53801 & ~w53802;
assign w53993 = ~w53803 & ~w53804;
assign w53994 = ~w53805 & ~w53806;
assign w53995 = ~w53807 & ~w53808;
assign w53996 = ~w53809 & ~w53810;
assign w53997 = ~w53811 & ~w53812;
assign w53998 = ~w53813 & ~w53814;
assign w53999 = ~w53815 & ~w53816;
assign w54000 = ~w53817 & ~w53818;
assign w54001 = ~w53819 & ~w53820;
assign w54002 = ~w53821 & ~w53822;
assign w54003 = ~w53823 & ~w53824;
assign w54004 = ~w53825 & ~w53826;
assign w54005 = ~w53827 & ~w53828;
assign w54006 = ~w53829 & ~w53830;
assign w54007 = ~w53831 & ~w53832;
assign w54008 = ~w53833 & ~w53834;
assign w54009 = ~w53835 & ~w53836;
assign w54010 = ~w53837 & ~w53838;
assign w54011 = ~w53839 & ~w53840;
assign w54012 = ~w53841 & ~w53842;
assign w54013 = ~w53843 & ~w53844;
assign w54014 = ~w53845 & ~w53846;
assign w54015 = ~w53847 & ~w53848;
assign w54016 = ~w53849 & ~w53850;
assign w54017 = ~w53851 & ~w53852;
assign w54018 = ~w53853 & ~w53854;
assign w54019 = ~w53855 & ~w53856;
assign w54020 = ~w53857 & ~w53858;
assign w54021 = ~w53859 & ~w53860;
assign w54022 = ~w53861 & ~w53862;
assign w54023 = ~w53863 & ~w53864;
assign w54024 = ~w53865 & ~w53866;
assign w54025 = ~w53867 & ~w53868;
assign w54026 = ~w53869 & ~w53870;
assign w54027 = ~w53871 & ~w53872;
assign w54028 = ~w53873 & ~w53874;
assign w54029 = ~w53875 & ~w53876;
assign w54030 = ~w53877 & ~w53878;
assign w54031 = ~w53879 & ~w53880;
assign w54032 = ~w53881 & ~w53882;
assign w54033 = ~w53883 & ~w53884;
assign w54034 = ~w53885 & ~w53886;
assign w54035 = ~w53887 & ~w53888;
assign w54036 = ~w53889 & ~w53890;
assign w54037 = ~w53891 & ~w53892;
assign w54038 = ~w53893 & ~w53894;
assign w54039 = ~w53895 & ~w53896;
assign w54040 = ~w53897 & ~w53898;
assign w54041 = ~w53899 & ~w53900;
assign w54042 = ~w53901 & ~w53902;
assign w54043 = ~w53903 & ~w53904;
assign w54044 = ~w53905 & ~w53906;
assign w54045 = ~w53907 & ~w53908;
assign w54046 = ~w53909 & ~w53910;
assign w54047 = ~w53911 & ~w53912;
assign w54048 = ~w53913 & ~w53914;
assign w54049 = ~w53915 & ~w53916;
assign w54050 = ~w53917 & ~w53918;
assign w54051 = ~w53919 & ~w53920;
assign w54052 = ~w53921 & ~w53922;
assign w54053 = ~w53923 & ~w53924;
assign w54054 = ~w53925 & ~w53926;
assign w54055 = w54053 & w54054;
assign w54056 = w54051 & w54052;
assign w54057 = w54049 & w54050;
assign w54058 = w54047 & w54048;
assign w54059 = w54045 & w54046;
assign w54060 = w54043 & w54044;
assign w54061 = w54041 & w54042;
assign w54062 = w54039 & w54040;
assign w54063 = w54037 & w54038;
assign w54064 = w54035 & w54036;
assign w54065 = w54033 & w54034;
assign w54066 = w54031 & w54032;
assign w54067 = w54029 & w54030;
assign w54068 = w54027 & w54028;
assign w54069 = w54025 & w54026;
assign w54070 = w54023 & w54024;
assign w54071 = w54021 & w54022;
assign w54072 = w54019 & w54020;
assign w54073 = w54017 & w54018;
assign w54074 = w54015 & w54016;
assign w54075 = w54013 & w54014;
assign w54076 = w54011 & w54012;
assign w54077 = w54009 & w54010;
assign w54078 = w54007 & w54008;
assign w54079 = w54005 & w54006;
assign w54080 = w54003 & w54004;
assign w54081 = w54001 & w54002;
assign w54082 = w53999 & w54000;
assign w54083 = w53997 & w53998;
assign w54084 = w53995 & w53996;
assign w54085 = w53993 & w53994;
assign w54086 = w53991 & w53992;
assign w54087 = w53989 & w53990;
assign w54088 = w53987 & w53988;
assign w54089 = w53985 & w53986;
assign w54090 = w53983 & w53984;
assign w54091 = w53981 & w53982;
assign w54092 = w53979 & w53980;
assign w54093 = w53977 & w53978;
assign w54094 = w53975 & w53976;
assign w54095 = w53973 & w53974;
assign w54096 = w53971 & w53972;
assign w54097 = w53969 & w53970;
assign w54098 = w53967 & w53968;
assign w54099 = w53965 & w53966;
assign w54100 = w53963 & w53964;
assign w54101 = w53961 & w53962;
assign w54102 = w53959 & w53960;
assign w54103 = w53957 & w53958;
assign w54104 = w53955 & w53956;
assign w54105 = w53953 & w53954;
assign w54106 = w53951 & w53952;
assign w54107 = w53949 & w53950;
assign w54108 = w53947 & w53948;
assign w54109 = w53945 & w53946;
assign w54110 = w53943 & w53944;
assign w54111 = w53941 & w53942;
assign w54112 = w53939 & w53940;
assign w54113 = w53937 & w53938;
assign w54114 = w53935 & w53936;
assign w54115 = w53933 & w53934;
assign w54116 = w53931 & w53932;
assign w54117 = w53929 & w53930;
assign w54118 = w53927 & w53928;
assign w54119 = w54117 & w54118;
assign w54120 = w54115 & w54116;
assign w54121 = w54113 & w54114;
assign w54122 = w54111 & w54112;
assign w54123 = w54109 & w54110;
assign w54124 = w54107 & w54108;
assign w54125 = w54105 & w54106;
assign w54126 = w54103 & w54104;
assign w54127 = w54101 & w54102;
assign w54128 = w54099 & w54100;
assign w54129 = w54097 & w54098;
assign w54130 = w54095 & w54096;
assign w54131 = w54093 & w54094;
assign w54132 = w54091 & w54092;
assign w54133 = w54089 & w54090;
assign w54134 = w54087 & w54088;
assign w54135 = w54085 & w54086;
assign w54136 = w54083 & w54084;
assign w54137 = w54081 & w54082;
assign w54138 = w54079 & w54080;
assign w54139 = w54077 & w54078;
assign w54140 = w54075 & w54076;
assign w54141 = w54073 & w54074;
assign w54142 = w54071 & w54072;
assign w54143 = w54069 & w54070;
assign w54144 = w54067 & w54068;
assign w54145 = w54065 & w54066;
assign w54146 = w54063 & w54064;
assign w54147 = w54061 & w54062;
assign w54148 = w54059 & w54060;
assign w54149 = w54057 & w54058;
assign w54150 = w54055 & w54056;
assign w54151 = w54149 & w54150;
assign w54152 = w54147 & w54148;
assign w54153 = w54145 & w54146;
assign w54154 = w54143 & w54144;
assign w54155 = w54141 & w54142;
assign w54156 = w54139 & w54140;
assign w54157 = w54137 & w54138;
assign w54158 = w54135 & w54136;
assign w54159 = w54133 & w54134;
assign w54160 = w54131 & w54132;
assign w54161 = w54129 & w54130;
assign w54162 = w54127 & w54128;
assign w54163 = w54125 & w54126;
assign w54164 = w54123 & w54124;
assign w54165 = w54121 & w54122;
assign w54166 = w54119 & w54120;
assign w54167 = w54165 & w54166;
assign w54168 = w54163 & w54164;
assign w54169 = w54161 & w54162;
assign w54170 = w54159 & w54160;
assign w54171 = w54157 & w54158;
assign w54172 = w54155 & w54156;
assign w54173 = w54153 & w54154;
assign w54174 = w54151 & w54152;
assign w54175 = w54173 & w54174;
assign w54176 = w54171 & w54172;
assign w54177 = w54169 & w54170;
assign w54178 = w54167 & w54168;
assign w54179 = w54177 & w54178;
assign w54180 = w54175 & w54176;
assign w54181 = w54179 & w54180;
assign w54182 = ~pi10577 & ~w54181;
assign w54183 = pi09353 & w3402;
assign w54184 = pi04733 & w3490;
assign w54185 = pi09446 & w3438;
assign w54186 = pi08678 & w3422;
assign w54187 = pi08921 & w3472;
assign w54188 = pi02546 & w3378;
assign w54189 = pi08784 & w3432;
assign w54190 = pi09188 & w3616;
assign w54191 = pi08817 & w3466;
assign w54192 = pi04847 & w3522;
assign w54193 = pi08778 & w3384;
assign w54194 = pi08639 & w3298;
assign w54195 = pi09208 & w3606;
assign w54196 = pi09692 & w3334;
assign w54197 = pi08862 & w3552;
assign w54198 = pi09287 & w3320;
assign w54199 = pi04584 & w3470;
assign w54200 = pi08704 & w3496;
assign w54201 = pi04642 & w3322;
assign w54202 = pi08698 & w3462;
assign w54203 = pi04519 & w3306;
assign w54204 = pi08999 & w3312;
assign w54205 = pi04893 & w3214;
assign w54206 = pi08483 & w3598;
assign w54207 = pi04578 & w3416;
assign w54208 = pi04866 & w3454;
assign w54209 = pi09018 & w3372;
assign w54210 = pi04597 & w3404;
assign w54211 = pi08554 & w3288;
assign w54212 = pi08895 & w3156;
assign w54213 = pi08610 & w3482;
assign w54214 = pi09319 & w3542;
assign w54215 = pi09406 & w3324;
assign w54216 = pi08543 & w3550;
assign w54217 = pi05050 & w3396;
assign w54218 = pi04552 & w3336;
assign w54219 = pi09499 & w3558;
assign w54220 = pi09031 & w3600;
assign w54221 = pi04629 & w3534;
assign w54222 = pi04688 & w3262;
assign w54223 = pi09012 & w3201;
assign w54224 = pi09248 & w3594;
assign w54225 = pi04860 & w3502;
assign w54226 = pi08914 & w3225;
assign w54227 = pi04759 & w3209;
assign w54228 = pi04655 & w3274;
assign w54229 = pi04694 & w3292;
assign w54230 = pi09162 & w3426;
assign w54231 = pi08804 & w3398;
assign w54232 = pi04786 & w3592;
assign w54233 = pi09392 & w3294;
assign w54234 = pi09198 & w3175;
assign w54235 = pi08504 & w3492;
assign w54236 = pi08823 & w3127;
assign w54237 = pi09426 & w3602;
assign w54238 = pi08770 & w3442;
assign w54239 = pi02618 & w3452;
assign w54240 = pi09555 & w3184;
assign w54241 = pi09339 & w3318;
assign w54242 = pi04840 & w3428;
assign w54243 = pi09117 & w3386;
assign w54244 = pi04753 & w3576;
assign w54245 = pi08751 & w3078;
assign w54246 = pi04623 & w3064;
assign w54247 = pi09214 & w3446;
assign w54248 = pi04727 & w3548;
assign w54249 = pi02005 & w3418;
assign w54250 = pi09570 & w3162;
assign w54251 = pi08869 & w3410;
assign w54252 = pi04740 & w3526;
assign w54253 = pi08659 & w3203;
assign w54254 = pi08588 & w3460;
assign w54255 = pi08725 & w3278;
assign w54256 = pi09779 & w3110;
assign w54257 = pi04793 & w3498;
assign w54258 = pi09530 & w3388;
assign w54259 = pi09583 & w3258;
assign w54260 = pi09039 & w3194;
assign w54261 = pi04675 & w3296;
assign w54262 = pi08973 & w3276;
assign w54263 = pi09398 & w3316;
assign w54264 = pi02749 & w3211;
assign w54265 = pi09666 & w3484;
assign w54266 = pi04880 & w3326;
assign w54267 = pi04906 & w3115;
assign w54268 = pi08960 & w3448;
assign w54269 = pi08497 & w3344;
assign w54270 = pi08882 & w3135;
assign w54271 = pi09385 & w3148;
assign w54272 = pi02071 & w3380;
assign w54273 = pi08432 & w3486;
assign w54274 = pi04616 & w3250;
assign w54275 = pi08953 & w3358;
assign w54276 = pi04932 & w3146;
assign w54277 = pi09169 & w3516;
assign w54278 = pi02744 & w3488;
assign w54279 = pi04746 & w3350;
assign w54280 = pi04827 & w3574;
assign w54281 = pi04714 & w3310;
assign w54282 = pi08452 & w3266;
assign w54283 = pi09518 & w3408;
assign w54284 = pi05037 & w3177;
assign w54285 = pi08626 & w3450;
assign w54286 = pi09359 & w3580;
assign w54287 = pi04820 & w3118;
assign w54288 = pi05063 & w3582;
assign w54289 = pi08849 & w3340;
assign w54290 = pi09512 & w3510;
assign w54291 = pi08490 & w3604;
assign w54292 = pi04799 & w3132;
assign w54293 = pi04662 & w3536;
assign w54294 = pi04766 & w3338;
assign w54295 = pi08791 & w3506;
assign w54296 = pi09439 & w3179;
assign w54297 = pi08614 & w3314;
assign w54298 = pi08477 & w3248;
assign w54299 = pi08458 & w3143;
assign w54300 = pi04564 & w3500;
assign w54301 = pi08599 & w3414;
assign w54302 = pi08875 & w3420;
assign w54303 = pi08986 & w3508;
assign w54304 = pi04707 & w3610;
assign w54305 = pi09345 & w3188;
assign w54306 = pi09433 & w3578;
assign w54307 = pi09679 & w3190;
assign w54308 = pi09412 & w3332;
assign w54309 = pi09143 & w3125;
assign w54310 = pi02553 & w3150;
assign w54311 = pi04532 & w3346;
assign w54312 = pi09419 & w3158;
assign w54313 = pi04591 & w3362;
assign w54314 = pi09465 & w3524;
assign w54315 = pi02018 & w3544;
assign w54316 = pi09372 & w3560;
assign w54317 = pi09639 & w3618;
assign w54318 = pi09332 & w3096;
assign w54319 = pi04813 & w3071;
assign w54320 = pi08934 & w3620;
assign w54321 = pi08583 & w3356;
assign w54322 = pi04547 & w3197;
assign w54323 = pi08908 & w3254;
assign w54324 = pi08522 & w3219;
assign w54325 = pi09459 & w3160;
assign w54326 = pi09110 & w3270;
assign w54327 = pi09452 & w3368;
assign w54328 = pi08439 & w3232;
assign w54329 = pi02753 & w3588;
assign w54330 = pi08527 & w3554;
assign w54331 = pi08738 & w3186;
assign w54332 = pi08685 & w3227;
assign w54333 = pi08633 & w3236;
assign w54334 = pi09234 & w3608;
assign w54335 = pi09274 & w3106;
assign w54336 = pi09366 & w3229;
assign w54337 = pi09005 & w3165;
assign w54338 = pi09306 & w3264;
assign w54339 = pi09221 & w3570;
assign w54340 = pi04773 & w3348;
assign w54341 = pi09653 & w3564;
assign w54342 = pi09617 & w3412;
assign w54343 = pi09104 & w3207;
assign w54344 = pi09240 & w3366;
assign w54345 = pi09097 & w3464;
assign w54346 = pi04945 & w3370;
assign w54347 = pi08691 & w3304;
assign w54348 = pi04541 & w3520;
assign w54349 = pi04971 & w3562;
assign w54350 = pi09547 & w3169;
assign w54351 = pi09201 & w3223;
assign w54352 = pi09058 & w3171;
assign w54353 = pi08731 & w3514;
assign w54354 = pi08810 & w3234;
assign w54355 = pi01518 & w3246;
assign w54356 = pi02074 & w3614;
assign w54357 = pi04610 & w3530;
assign w54358 = pi09420 & w3568;
assign w54359 = pi09130 & w3352;
assign w54360 = pi09175 & w3474;
assign w54361 = pi08992 & w3167;
assign w54362 = pi05073 & w3242;
assign w54363 = pi09313 & w3546;
assign w54364 = pi03536 & w3612;
assign w54365 = pi09182 & w3532;
assign w54366 = pi04636 & w3400;
assign w54367 = pi08797 & w3300;
assign w54368 = pi05024 & w3556;
assign w54369 = pi04780 & w3456;
assign w54370 = pi08672 & w3199;
assign w54371 = pi08718 & w3082;
assign w54372 = pi09025 & w3374;
assign w54373 = pi08764 & w3518;
assign w54374 = pi08711 & w3153;
assign w54375 = pi09149 & w3093;
assign w54376 = pi09254 & w3468;
assign w54377 = pi04919 & w3328;
assign w54378 = pi09227 & w3440;
assign w54379 = pi04681 & w3137;
assign w54380 = pi04807 & w3394;
assign w54381 = pi09091 & w3390;
assign w54382 = pi08470 & w3436;
assign w54383 = pi08445 & w3240;
assign w54384 = pi08652 & w3392;
assign w54385 = pi09078 & w3192;
assign w54386 = pi05010 & w3504;
assign w54387 = pi08940 & w3272;
assign w54388 = pi04958 & w3512;
assign w54389 = pi08620 & w3538;
assign w54390 = pi04834 & w3494;
assign w54391 = pi09136 & w3596;
assign w54392 = pi09293 & w3478;
assign w54393 = pi08836 & w3406;
assign w54394 = pi05449 & w3480;
assign w54395 = pi08901 & w3205;
assign w54396 = pi09267 & w3584;
assign w54397 = pi08947 & w3376;
assign w54398 = pi09280 & w3444;
assign w54399 = pi09084 & w3360;
assign w54400 = pi09714 & w3290;
assign w54401 = pi09300 & w3282;
assign w54402 = pi04853 & w3181;
assign w54403 = pi09045 & w3590;
assign w54404 = pi08537 & w3528;
assign w54405 = pi08605 & w3540;
assign w54406 = pi04649 & w3103;
assign w54407 = pi09065 & w3476;
assign w54408 = pi08927 & w3221;
assign w54409 = pi09156 & w3238;
assign w54410 = pi09326 & w3280;
assign w54411 = pi08888 & w3364;
assign w54412 = pi08594 & w3586;
assign w54413 = pi08646 & w3354;
assign w54414 = pi09379 & w3342;
assign w54415 = pi09071 & w3458;
assign w54416 = pi08757 & w3256;
assign w54417 = pi08979 & w3434;
assign w54418 = pi08516 & w3252;
assign w54419 = pi04997 & w3122;
assign w54420 = pi08966 & w3566;
assign w54421 = pi08830 & w3139;
assign w54422 = pi08571 & w3112;
assign w54423 = pi08665 & w3129;
assign w54424 = pi02014 & w3268;
assign w54425 = pi08567 & w3217;
assign w54426 = pi04720 & w3244;
assign w54427 = pi04668 & w3424;
assign w54428 = pi04603 & w3330;
assign w54429 = pi08856 & w3286;
assign w54430 = pi09052 & w3430;
assign w54431 = pi04701 & w3260;
assign w54432 = pi01679 & w3308;
assign w54433 = pi09261 & w3173;
assign w54434 = pi08843 & w3572;
assign w54435 = pi09123 & w3382;
assign w54436 = pi09691 & w3086;
assign w54437 = pi04984 & w3302;
assign w54438 = pi08744 & w3284;
assign w54439 = ~w54183 & ~w54184;
assign w54440 = ~w54185 & ~w54186;
assign w54441 = ~w54187 & ~w54188;
assign w54442 = ~w54189 & ~w54190;
assign w54443 = ~w54191 & ~w54192;
assign w54444 = ~w54193 & ~w54194;
assign w54445 = ~w54195 & ~w54196;
assign w54446 = ~w54197 & ~w54198;
assign w54447 = ~w54199 & ~w54200;
assign w54448 = ~w54201 & ~w54202;
assign w54449 = ~w54203 & ~w54204;
assign w54450 = ~w54205 & ~w54206;
assign w54451 = ~w54207 & ~w54208;
assign w54452 = ~w54209 & ~w54210;
assign w54453 = ~w54211 & ~w54212;
assign w54454 = ~w54213 & ~w54214;
assign w54455 = ~w54215 & ~w54216;
assign w54456 = ~w54217 & ~w54218;
assign w54457 = ~w54219 & ~w54220;
assign w54458 = ~w54221 & ~w54222;
assign w54459 = ~w54223 & ~w54224;
assign w54460 = ~w54225 & ~w54226;
assign w54461 = ~w54227 & ~w54228;
assign w54462 = ~w54229 & ~w54230;
assign w54463 = ~w54231 & ~w54232;
assign w54464 = ~w54233 & ~w54234;
assign w54465 = ~w54235 & ~w54236;
assign w54466 = ~w54237 & ~w54238;
assign w54467 = ~w54239 & ~w54240;
assign w54468 = ~w54241 & ~w54242;
assign w54469 = ~w54243 & ~w54244;
assign w54470 = ~w54245 & ~w54246;
assign w54471 = ~w54247 & ~w54248;
assign w54472 = ~w54249 & ~w54250;
assign w54473 = ~w54251 & ~w54252;
assign w54474 = ~w54253 & ~w54254;
assign w54475 = ~w54255 & ~w54256;
assign w54476 = ~w54257 & ~w54258;
assign w54477 = ~w54259 & ~w54260;
assign w54478 = ~w54261 & ~w54262;
assign w54479 = ~w54263 & ~w54264;
assign w54480 = ~w54265 & ~w54266;
assign w54481 = ~w54267 & ~w54268;
assign w54482 = ~w54269 & ~w54270;
assign w54483 = ~w54271 & ~w54272;
assign w54484 = ~w54273 & ~w54274;
assign w54485 = ~w54275 & ~w54276;
assign w54486 = ~w54277 & ~w54278;
assign w54487 = ~w54279 & ~w54280;
assign w54488 = ~w54281 & ~w54282;
assign w54489 = ~w54283 & ~w54284;
assign w54490 = ~w54285 & ~w54286;
assign w54491 = ~w54287 & ~w54288;
assign w54492 = ~w54289 & ~w54290;
assign w54493 = ~w54291 & ~w54292;
assign w54494 = ~w54293 & ~w54294;
assign w54495 = ~w54295 & ~w54296;
assign w54496 = ~w54297 & ~w54298;
assign w54497 = ~w54299 & ~w54300;
assign w54498 = ~w54301 & ~w54302;
assign w54499 = ~w54303 & ~w54304;
assign w54500 = ~w54305 & ~w54306;
assign w54501 = ~w54307 & ~w54308;
assign w54502 = ~w54309 & ~w54310;
assign w54503 = ~w54311 & ~w54312;
assign w54504 = ~w54313 & ~w54314;
assign w54505 = ~w54315 & ~w54316;
assign w54506 = ~w54317 & ~w54318;
assign w54507 = ~w54319 & ~w54320;
assign w54508 = ~w54321 & ~w54322;
assign w54509 = ~w54323 & ~w54324;
assign w54510 = ~w54325 & ~w54326;
assign w54511 = ~w54327 & ~w54328;
assign w54512 = ~w54329 & ~w54330;
assign w54513 = ~w54331 & ~w54332;
assign w54514 = ~w54333 & ~w54334;
assign w54515 = ~w54335 & ~w54336;
assign w54516 = ~w54337 & ~w54338;
assign w54517 = ~w54339 & ~w54340;
assign w54518 = ~w54341 & ~w54342;
assign w54519 = ~w54343 & ~w54344;
assign w54520 = ~w54345 & ~w54346;
assign w54521 = ~w54347 & ~w54348;
assign w54522 = ~w54349 & ~w54350;
assign w54523 = ~w54351 & ~w54352;
assign w54524 = ~w54353 & ~w54354;
assign w54525 = ~w54355 & ~w54356;
assign w54526 = ~w54357 & ~w54358;
assign w54527 = ~w54359 & ~w54360;
assign w54528 = ~w54361 & ~w54362;
assign w54529 = ~w54363 & ~w54364;
assign w54530 = ~w54365 & ~w54366;
assign w54531 = ~w54367 & ~w54368;
assign w54532 = ~w54369 & ~w54370;
assign w54533 = ~w54371 & ~w54372;
assign w54534 = ~w54373 & ~w54374;
assign w54535 = ~w54375 & ~w54376;
assign w54536 = ~w54377 & ~w54378;
assign w54537 = ~w54379 & ~w54380;
assign w54538 = ~w54381 & ~w54382;
assign w54539 = ~w54383 & ~w54384;
assign w54540 = ~w54385 & ~w54386;
assign w54541 = ~w54387 & ~w54388;
assign w54542 = ~w54389 & ~w54390;
assign w54543 = ~w54391 & ~w54392;
assign w54544 = ~w54393 & ~w54394;
assign w54545 = ~w54395 & ~w54396;
assign w54546 = ~w54397 & ~w54398;
assign w54547 = ~w54399 & ~w54400;
assign w54548 = ~w54401 & ~w54402;
assign w54549 = ~w54403 & ~w54404;
assign w54550 = ~w54405 & ~w54406;
assign w54551 = ~w54407 & ~w54408;
assign w54552 = ~w54409 & ~w54410;
assign w54553 = ~w54411 & ~w54412;
assign w54554 = ~w54413 & ~w54414;
assign w54555 = ~w54415 & ~w54416;
assign w54556 = ~w54417 & ~w54418;
assign w54557 = ~w54419 & ~w54420;
assign w54558 = ~w54421 & ~w54422;
assign w54559 = ~w54423 & ~w54424;
assign w54560 = ~w54425 & ~w54426;
assign w54561 = ~w54427 & ~w54428;
assign w54562 = ~w54429 & ~w54430;
assign w54563 = ~w54431 & ~w54432;
assign w54564 = ~w54433 & ~w54434;
assign w54565 = ~w54435 & ~w54436;
assign w54566 = ~w54437 & ~w54438;
assign w54567 = w54565 & w54566;
assign w54568 = w54563 & w54564;
assign w54569 = w54561 & w54562;
assign w54570 = w54559 & w54560;
assign w54571 = w54557 & w54558;
assign w54572 = w54555 & w54556;
assign w54573 = w54553 & w54554;
assign w54574 = w54551 & w54552;
assign w54575 = w54549 & w54550;
assign w54576 = w54547 & w54548;
assign w54577 = w54545 & w54546;
assign w54578 = w54543 & w54544;
assign w54579 = w54541 & w54542;
assign w54580 = w54539 & w54540;
assign w54581 = w54537 & w54538;
assign w54582 = w54535 & w54536;
assign w54583 = w54533 & w54534;
assign w54584 = w54531 & w54532;
assign w54585 = w54529 & w54530;
assign w54586 = w54527 & w54528;
assign w54587 = w54525 & w54526;
assign w54588 = w54523 & w54524;
assign w54589 = w54521 & w54522;
assign w54590 = w54519 & w54520;
assign w54591 = w54517 & w54518;
assign w54592 = w54515 & w54516;
assign w54593 = w54513 & w54514;
assign w54594 = w54511 & w54512;
assign w54595 = w54509 & w54510;
assign w54596 = w54507 & w54508;
assign w54597 = w54505 & w54506;
assign w54598 = w54503 & w54504;
assign w54599 = w54501 & w54502;
assign w54600 = w54499 & w54500;
assign w54601 = w54497 & w54498;
assign w54602 = w54495 & w54496;
assign w54603 = w54493 & w54494;
assign w54604 = w54491 & w54492;
assign w54605 = w54489 & w54490;
assign w54606 = w54487 & w54488;
assign w54607 = w54485 & w54486;
assign w54608 = w54483 & w54484;
assign w54609 = w54481 & w54482;
assign w54610 = w54479 & w54480;
assign w54611 = w54477 & w54478;
assign w54612 = w54475 & w54476;
assign w54613 = w54473 & w54474;
assign w54614 = w54471 & w54472;
assign w54615 = w54469 & w54470;
assign w54616 = w54467 & w54468;
assign w54617 = w54465 & w54466;
assign w54618 = w54463 & w54464;
assign w54619 = w54461 & w54462;
assign w54620 = w54459 & w54460;
assign w54621 = w54457 & w54458;
assign w54622 = w54455 & w54456;
assign w54623 = w54453 & w54454;
assign w54624 = w54451 & w54452;
assign w54625 = w54449 & w54450;
assign w54626 = w54447 & w54448;
assign w54627 = w54445 & w54446;
assign w54628 = w54443 & w54444;
assign w54629 = w54441 & w54442;
assign w54630 = w54439 & w54440;
assign w54631 = w54629 & w54630;
assign w54632 = w54627 & w54628;
assign w54633 = w54625 & w54626;
assign w54634 = w54623 & w54624;
assign w54635 = w54621 & w54622;
assign w54636 = w54619 & w54620;
assign w54637 = w54617 & w54618;
assign w54638 = w54615 & w54616;
assign w54639 = w54613 & w54614;
assign w54640 = w54611 & w54612;
assign w54641 = w54609 & w54610;
assign w54642 = w54607 & w54608;
assign w54643 = w54605 & w54606;
assign w54644 = w54603 & w54604;
assign w54645 = w54601 & w54602;
assign w54646 = w54599 & w54600;
assign w54647 = w54597 & w54598;
assign w54648 = w54595 & w54596;
assign w54649 = w54593 & w54594;
assign w54650 = w54591 & w54592;
assign w54651 = w54589 & w54590;
assign w54652 = w54587 & w54588;
assign w54653 = w54585 & w54586;
assign w54654 = w54583 & w54584;
assign w54655 = w54581 & w54582;
assign w54656 = w54579 & w54580;
assign w54657 = w54577 & w54578;
assign w54658 = w54575 & w54576;
assign w54659 = w54573 & w54574;
assign w54660 = w54571 & w54572;
assign w54661 = w54569 & w54570;
assign w54662 = w54567 & w54568;
assign w54663 = w54661 & w54662;
assign w54664 = w54659 & w54660;
assign w54665 = w54657 & w54658;
assign w54666 = w54655 & w54656;
assign w54667 = w54653 & w54654;
assign w54668 = w54651 & w54652;
assign w54669 = w54649 & w54650;
assign w54670 = w54647 & w54648;
assign w54671 = w54645 & w54646;
assign w54672 = w54643 & w54644;
assign w54673 = w54641 & w54642;
assign w54674 = w54639 & w54640;
assign w54675 = w54637 & w54638;
assign w54676 = w54635 & w54636;
assign w54677 = w54633 & w54634;
assign w54678 = w54631 & w54632;
assign w54679 = w54677 & w54678;
assign w54680 = w54675 & w54676;
assign w54681 = w54673 & w54674;
assign w54682 = w54671 & w54672;
assign w54683 = w54669 & w54670;
assign w54684 = w54667 & w54668;
assign w54685 = w54665 & w54666;
assign w54686 = w54663 & w54664;
assign w54687 = w54685 & w54686;
assign w54688 = w54683 & w54684;
assign w54689 = w54681 & w54682;
assign w54690 = w54679 & w54680;
assign w54691 = w54689 & w54690;
assign w54692 = w54687 & w54688;
assign w54693 = w54691 & w54692;
assign w54694 = ~pi10577 & ~w54693;
assign w54695 = w168 & ~pi10236;
assign w54696 = pi00095 & pi00096;
assign w54697 = pi00098 & pi00099;
assign w54698 = pi00432 & pi00423;
assign w54699 = pi00424 & pi00425;
assign w54700 = ~pi10025 & ~pi00020;
assign w54701 = ~pi10234 & ~pi10235;
assign w54702 = pi10234 & pi10235;
assign w54703 = (~pi00016 & ~w185) | (~pi00016 & w54719) | (~w185 & w54719);
assign w54704 = ~w168 & pi10236;
assign w54705 = w222 & w54720;
assign w54706 = pi00119 & pi00120;
assign w54707 = pi00124 & pi00126;
assign w54708 = ~w1454 & ~w1430;
assign w54709 = ~w111 & ~pi09800;
assign w54710 = w111 & pi09800;
assign w54711 = ~w1528 & w1529;
assign w54712 = pi10377 & pi10391;
assign w54713 = pi10386 & pi10385;
assign w54714 = w1381 & pi00134;
assign w54715 = (~pi00146 & ~w1969) | (~pi00146 & w54743) | (~w1969 & w54743);
assign w54716 = ~w1980 & ~w2015;
assign w54717 = w2249 & w2383;
assign w54718 = w54699 & pi00426;
assign w54719 = ~pi00015 & ~pi00016;
assign w54720 = ~pi10025 & ~pi10239;
assign w54721 = w176 & ~pi00018;
assign w54722 = ~w54700 & pi00017;
assign w54723 = ~w54703 & ~w183;
assign w54724 = ~pi10025 & pi00020;
assign w54725 = w200 & ~w173;
assign w54726 = ~pi00017 & ~pi00018;
assign w54727 = ~pi10025 & ~pi10024;
assign w54728 = pi10025 & pi10024;
assign w54729 = ~w219 & ~w220;
assign w54730 = w54705 & ~pi10238;
assign w54731 = w229 & w54744;
assign w54732 = w242 & w54769;
assign w54733 = (~w221 & w54861) | (~w221 & w54862) | (w54861 & w54862);
assign w54734 = w54706 & w1354;
assign w54735 = w54707 & pi00181;
assign w54736 = pi00244 & pi00245;
assign w54737 = w1427 & w1456;
assign w54738 = ~w1523 & w1526;
assign w54739 = w54713 & pi10353;
assign w54740 = w1355 & pi00290;
assign w54741 = pi00427 & pi00428;
assign w54742 = w54741 & pi00429;
assign w54743 = ~pi00153 & ~pi00146;
assign w54744 = ~pi10021 & ~pi00010;
assign w54745 = ~pi09963 & ~pi09819;
assign w54746 = w186 & pi00016;
assign w54747 = ~w223 & pi10239;
assign w54748 = ~w54705 & pi10238;
assign w54749 = ~pi10021 & pi10234;
assign w54750 = ~pi10021 & ~pi10241;
assign w54751 = (~pi00030 & w522) | (~pi00030 & w54770) | (w522 & w54770);
assign w54752 = pi00127 & pi00136;
assign w54753 = w54736 & pi00246;
assign w54754 = (~pi00248 & ~w1410) | (~pi00248 & w54771) | (~w1410 & w54771);
assign w54755 = ~w54736 & ~pi00246;
assign w54756 = w1457 & ~w1456;
assign w54757 = w1457 & ~w54737;
assign w54758 = pi00247 & pi00248;
assign w54759 = pi00236 & pi00237;
assign w54760 = w1530 & ~w1529;
assign w54761 = w1530 & ~w54711;
assign w54762 = pi10361 & pi10347;
assign w54763 = w1582 & w54772;
assign w54764 = w2039 & w2030;
assign w54765 = pi00284 & pi00261;
assign w54766 = ~w2606 & w2597;
assign w54767 = w145 & pi00233;
assign w54768 = w54742 & pi00406;
assign w54769 = w245 & pi00022;
assign w54770 = w520 & ~pi00030;
assign w54771 = ~pi00247 & ~pi00248;
assign w54772 = w54762 & w1563;
assign w54773 = w54749 & w262;
assign w54774 = ~w295 & ~w287;
assign w54775 = (~w295 & w282) | (~w295 & w54774) | (w282 & w54774);
assign w54776 = w300 & w287;
assign w54777 = ~w282 & w54776;
assign w54778 = w536 & pi00025;
assign w54779 = w403 & w54830;
assign w54780 = ~w1482 & ~pi00234;
assign w54781 = w1482 & pi00234;
assign w54782 = ~w1459 & w1465;
assign w54783 = w1482 & w1468;
assign w54784 = (~w1500 & w1547) | (~w1500 & w54798) | (w1547 & w54798);
assign w54785 = w54752 & w54714;
assign w54786 = w1582 & w54799;
assign w54787 = ~w827 & w1789;
assign w54788 = w54765 & pi00285;
assign w54789 = w54788 & pi00286;
assign w54790 = pi00122 & w2396;
assign w54791 = ~pi00156 & ~pi00206;
assign w54792 = pi00190 & w2415;
assign w54793 = ~pi09969 & pi00249;
assign w54794 = w54767 & ~w2597;
assign w54795 = w54767 & ~w54766;
assign w54796 = w10846 & pi00413;
assign w54797 = pi00019 & pi00020;
assign w54798 = ~w1549 & ~w1500;
assign w54799 = w54772 & ~pi00150;
assign w54800 = w298 & ~w54774;
assign w54801 = w298 & ~w54775;
assign w54802 = w531 & ~w54776;
assign w54803 = w531 & ~w54777;
assign w54804 = w577 & ~w54776;
assign w54805 = w577 & ~w54777;
assign w54806 = w54779 & pi00021;
assign w54807 = w293 & w54774;
assign w54808 = w293 & w54775;
assign w54809 = w391 & ~w54776;
assign w54810 = w391 & ~w54777;
assign w54811 = w1471 & ~w1465;
assign w54812 = w1471 & ~w54782;
assign w54813 = w1553 & w54831;
assign w54814 = w1557 & w54784;
assign w54815 = w54786 & w1565;
assign w54816 = w54787 & pi00175;
assign w54817 = w54787 & ~pi00175;
assign w54818 = w2052 & ~w2042;
assign w54819 = w2053 & w2030;
assign w54820 = w139 & pi00250;
assign w54821 = w54789 & w2387;
assign w54822 = pi00135 & w54790;
assign w54823 = ~pi09949 & w1500;
assign w54824 = ~pi09949 & ~w54784;
assign w54825 = pi00240 & pi00241;
assign w54826 = pi00415 & pi00416;
assign w54827 = ~pi02648 & ~pi01206;
assign w54828 = pi00838 & pi00839;
assign w54829 = ~pi00868 & ~pi00852;
assign w54830 = w198 & w54797;
assign w54831 = w1556 & ~w1500;
assign w54832 = w223 & w262;
assign w54833 = ~w54750 & pi10240;
assign w54834 = w263 & ~pi10242;
assign w54835 = ~w263 & pi10242;
assign w54836 = w383 & ~w322;
assign w54837 = pi00015 & pi00016;
assign w54838 = ~w498 & w530;
assign w54839 = ~w498 & w576;
assign w54840 = ~w540 & w54806;
assign w54841 = pi00024 & ~w54800;
assign w54842 = pi00024 & ~w54801;
assign w54843 = w507 & w54805;
assign w54844 = w507 & w54804;
assign w54845 = pi00030 & w54805;
assign w54846 = pi00030 & w54804;
assign w54847 = pi00031 & ~w54807;
assign w54848 = pi00031 & ~w54808;
assign w54849 = w688 & w54809;
assign w54850 = w688 & w54810;
assign w54851 = w785 & ~w54809;
assign w54852 = w785 & ~w54810;
assign w54853 = pi00053 & w54809;
assign w54854 = pi00053 & w54810;
assign w54855 = w1469 & pi10021;
assign w54856 = ~w1478 & w1487;
assign w54857 = ~pi00238 & pi00239;
assign w54858 = pi00238 & ~pi00239;
assign w54859 = ~w1534 & w1541;
assign w54860 = ~pi00148 & w1564;
assign w54861 = ~w272 & w54732;
assign w54862 = ~w272 & w246;
assign w54863 = w507 & ~w54800;
assign w54864 = w507 & ~w54801;
assign w54865 = ~pi00241 & w26;
assign w54866 = pi00241 & w65;
assign w54867 = ~w54866 & w63;
assign w54868 = w54866 & w63;
assign w54869 = w73 & ~pi00188;
assign w54870 = ~w139 & w145;
assign w54871 = ~w78 & w152;
assign w54872 = ~w54871 & ~pi00023;
assign w54873 = w54871 & pi00023;
assign w54874 = w76 & pi00023;
assign w54875 = w76 & ~w54872;
assign w54876 = ~w78 & w161;
assign w54877 = ~w54876 & pi00027;
assign w54878 = w54876 & ~pi00027;
assign w54879 = w76 & ~pi00027;
assign w54880 = w76 & ~w54877;
assign w54881 = pi10025 & ~pi00020;
assign w54882 = w168 & ~w198;
assign w54883 = pi00019 & ~w212;
assign w54884 = pi00021 & ~w211;
assign w54885 = ~w54727 & pi10023;
assign w54886 = pi00008 & pi00022;
assign w54887 = ~w232 & w247;
assign w54888 = w248 & w220;
assign w54889 = w248 & ~w210;
assign w54890 = ~w232 & w250;
assign w54891 = ~w239 & pi00010;
assign w54892 = ~w255 & pi00010;
assign w54893 = ~w255 & ~w54731;
assign w54894 = pi10021 & pi10241;
assign w54895 = w263 & ~pi00012;
assign w54896 = w54773 & ~pi00012;
assign w54897 = ~w54896 & pi00011;
assign w54898 = ~w54773 & pi00012;
assign w54899 = ~pi10535 & w294;
assign w54900 = ~pi00031 & ~w297;
assign w54901 = pi00015 & ~pi00025;
assign w54902 = ~pi10263 & w302;
assign w54903 = pi10354 & ~pi10476;
assign w54904 = w54899 & w296;
assign w54905 = ~w397 & ~pi09952;
assign w54906 = w198 & pi00019;
assign w54907 = w441 & w406;
assign w54908 = w483 & ~w482;
assign w54909 = ~w488 & w489;
assign w54910 = ~w491 & w492;
assign w54911 = ~w401 & w391;
assign w54912 = pi10354 & pi10476;
assign w54913 = ~w505 & w288;
assign w54914 = ~pi00030 & ~w445;
assign w54915 = ~pi00030 & w523;
assign w54916 = ~w524 & w507;
assign w54917 = ~w540 & pi00006;
assign w54918 = w540 & ~pi00006;
assign w54919 = ~w561 & w562;
assign w54920 = w549 & ~w548;
assign w54921 = w547 & ~w546;
assign w54922 = w565 & w546;
assign w54923 = w565 & ~w54921;
assign w54924 = w567 & w450;
assign w54925 = ~w457 & w570;
assign w54926 = w520 & ~pi00007;
assign w54927 = ~w574 & ~pi00007;
assign w54928 = ~w574 & ~w44973;
assign w54929 = ~w540 & w405;
assign w54930 = ~w540 & w54779;
assign w54931 = ~pi00022 & ~pi00008;
assign w54932 = ~w54886 & ~pi00009;
assign w54933 = w54886 & pi00009;
assign w54934 = ~w54933 & ~pi00010;
assign w54935 = w54933 & pi00010;
assign w54936 = w54935 & pi00011;
assign w54937 = ~w54935 & ~pi00011;
assign w54938 = ~w54936 & ~pi00012;
assign w54939 = w54936 & pi00012;
assign w54940 = ~w54939 & ~pi00013;
assign w54941 = w54939 & pi00013;
assign w54942 = ~w540 & w188;
assign w54943 = ~w540 & w301;
assign w54944 = pi00016 & pi00017;
assign w54945 = ~pi00016 & ~pi00017;
assign w54946 = ~w540 & w404;
assign w54947 = pi00018 & ~w625;
assign w54948 = ~w78 & w648;
assign w54949 = pi00051 & w76;
assign w54950 = pi10263 & w302;
assign w54951 = ~w501 & pi00025;
assign w54952 = w54876 & ~w152;
assign w54953 = w54871 & ~w161;
assign w54954 = ~pi00054 & w76;
assign w54955 = ~w54914 & pi00032;
assign w54956 = pi00032 & ~w679;
assign w54957 = w401 & ~pi00033;
assign w54958 = ~w401 & pi00033;
assign w54959 = w520 & ~pi00929;
assign w54960 = ~pi00030 & w685;
assign w54961 = ~w319 & w687;
assign w54962 = w401 & w693;
assign w54963 = ~pi00035 & ~pi00036;
assign w54964 = ~w400 & pi00038;
assign w54965 = pi10418 & pi09920;
assign w54966 = ~pi10418 & pi00451;
assign w54967 = ~w708 & ~w713;
assign w54968 = pi10418 & pi00967;
assign w54969 = ~pi10418 & pi00452;
assign w54970 = ~w719 & ~w722;
assign w54971 = ~pi00024 & pi00055;
assign w54972 = pi00024 & ~pi00055;
assign w54973 = w671 & ~pi00055;
assign w54974 = w671 & ~w54971;
assign w54975 = pi10418 & pi09806;
assign w54976 = ~pi10418 & pi00453;
assign w54977 = ~w734 & ~w737;
assign w54978 = ~pi00024 & pi00057;
assign w54979 = pi00024 & ~pi00057;
assign w54980 = w671 & ~pi00057;
assign w54981 = w671 & ~w54978;
assign w54982 = ~w78 & w755;
assign w54983 = pi00060 & w76;
assign w54984 = ~w501 & ~w760;
assign w54985 = pi10418 & pi09922;
assign w54986 = ~pi10418 & pi00454;
assign w54987 = ~w765 & ~w768;
assign w54988 = ~pi00024 & pi00056;
assign w54989 = pi00024 & ~pi00056;
assign w54990 = w671 & ~pi00056;
assign w54991 = w671 & ~w54988;
assign w54992 = ~pi00024 & pi00059;
assign w54993 = pi00024 & ~pi00059;
assign w54994 = w671 & ~pi00059;
assign w54995 = w671 & ~w54992;
assign w54996 = ~w78 & w752;
assign w54997 = ~w54996 & pi00061;
assign w54998 = w54996 & ~pi00061;
assign w54999 = w76 & ~pi00061;
assign w55000 = w76 & ~w54997;
assign w55001 = w520 & pi00849;
assign w55002 = ~pi00024 & pi00065;
assign w55003 = pi00024 & ~pi00065;
assign w55004 = w671 & ~pi00065;
assign w55005 = w671 & ~w55002;
assign w55006 = ~pi00024 & pi00067;
assign w55007 = pi00024 & ~pi00067;
assign w55008 = w671 & ~pi00067;
assign w55009 = w671 & ~w55006;
assign w55010 = w803 & pi00066;
assign w55011 = ~w803 & ~pi00066;
assign w55012 = ~w78 & w645;
assign w55013 = ~w55012 & pi00069;
assign w55014 = w55012 & ~pi00069;
assign w55015 = w76 & ~pi00069;
assign w55016 = w76 & ~w55013;
assign w55017 = ~pi00024 & pi00068;
assign w55018 = pi00024 & ~pi00068;
assign w55019 = w671 & ~pi00068;
assign w55020 = w671 & ~w55017;
assign w55021 = ~w55012 & pi00070;
assign w55022 = w55012 & ~pi00070;
assign w55023 = w76 & ~pi00070;
assign w55024 = w76 & ~w55021;
assign w55025 = ~w54996 & pi00073;
assign w55026 = w54996 & ~pi00073;
assign w55027 = w76 & ~pi00073;
assign w55028 = w76 & ~w55025;
assign w55029 = ~pi09997 & ~pi00062;
assign w55030 = pi09997 & pi10563;
assign w55031 = ~w846 & w849;
assign w55032 = ~pi00310 & ~pi00296;
assign w55033 = pi00309 & ~pi10516;
assign w55034 = w860 & ~pi10511;
assign w55035 = w863 & w856;
assign w55036 = w898 & w896;
assign w55037 = w930 & w854;
assign w55038 = w935 & w896;
assign w55039 = ~w859 & ~pi00308;
assign w55040 = ~w857 & pi00308;
assign w55041 = ~w1004 & pi00309;
assign w55042 = w968 & w856;
assign w55043 = w898 & w1075;
assign w55044 = ~w78 & ~w1080;
assign w55045 = w54871 & w1080;
assign w55046 = w1083 & pi00141;
assign w55047 = ~w1083 & ~pi00141;
assign w55048 = ~pi00024 & pi00184;
assign w55049 = pi00024 & ~pi00184;
assign w55050 = ~pi00024 & pi00185;
assign w55051 = pi00024 & ~pi00185;
assign w55052 = w671 & ~pi00185;
assign w55053 = w671 & ~w55050;
assign w55054 = w54876 & ~w648;
assign w55055 = w1099 & ~pi00187;
assign w55056 = ~w1099 & pi00187;
assign w55057 = ~w54876 & pi00186;
assign w55058 = w54876 & ~pi00186;
assign w55059 = w897 & pi00308;
assign w55060 = w1113 & pi00309;
assign w55061 = ~w1114 & ~pi00071;
assign w55062 = w1113 & w1116;
assign w55063 = pi10345 & pi00105;
assign w55064 = ~pi00814 & pi01272;
assign w55065 = w1126 & w1125;
assign w55066 = pi00348 & pi00365;
assign w55067 = w54871 & ~w755;
assign w55068 = w1142 & pi00231;
assign w55069 = ~w1142 & ~pi00231;
assign w55070 = ~w1134 & ~pi10489;
assign w55071 = ~w1134 & ~pi10520;
assign w55072 = ~w1134 & ~pi10495;
assign w55073 = ~w1134 & ~pi10492;
assign w55074 = ~w1134 & ~pi10505;
assign w55075 = ~w1134 & pi10483;
assign w55076 = ~w1134 & pi10511;
assign w55077 = ~w1134 & pi10486;
assign w55078 = ~pi10471 & ~pi00089;
assign w55079 = pi10471 & ~pi10574;
assign w55080 = pi09928 & ~pi10563;
assign w55081 = ~pi09928 & pi00090;
assign w55082 = ~pi10663 & w1204;
assign w55083 = ~pi10662 & ~pi10578;
assign w55084 = ~w55083 & ~pi10575;
assign w55085 = ~pi10655 & ~pi10657;
assign w55086 = w1213 & w1216;
assign w55087 = ~pi10655 & pi10657;
assign w55088 = pi10654 & pi10656;
assign w55089 = pi10655 & pi10657;
assign w55090 = pi10655 & ~pi10657;
assign w55091 = w1213 & w1224;
assign w55092 = w1213 & w1239;
assign w55093 = w1248 & w1252;
assign w55094 = ~w55083 & ~pi10568;
assign w55095 = ~w55083 & ~pi10559;
assign w55096 = pi00131 & pi00115;
assign w55097 = w55096 & pi00094;
assign w55098 = ~w55096 & ~pi00094;
assign w55099 = ~w55097 & ~w1194;
assign w55100 = pi10471 & pi10575;
assign w55101 = pi10471 & pi10559;
assign w55102 = ~pi00095 & ~pi00096;
assign w55103 = pi10471 & pi10568;
assign w55104 = pi10432 & pi10575;
assign w55105 = w54752 & pi00130;
assign w55106 = ~w55105 & ~pi00097;
assign w55107 = w54752 & w1381;
assign w55108 = ~w55107 & ~w1371;
assign w55109 = pi10432 & pi10559;
assign w55110 = ~pi00098 & ~pi00099;
assign w55111 = pi10432 & pi10568;
assign w55112 = ~pi00024 & pi00297;
assign w55113 = pi00024 & ~pi00297;
assign w55114 = w671 & ~pi00297;
assign w55115 = w671 & ~w55112;
assign w55116 = ~pi00024 & pi00298;
assign w55117 = pi00024 & ~pi00298;
assign w55118 = w671 & ~pi00298;
assign w55119 = w671 & ~w55116;
assign w55120 = ~w1469 & ~pi10021;
assign w55121 = w1485 & pi10240;
assign w55122 = ~w1485 & ~pi10240;
assign w55123 = w1498 & ~w1487;
assign w55124 = w1498 & ~w54856;
assign w55125 = w1469 & pi09974;
assign w55126 = ~w1485 & ~pi09944;
assign w55127 = ~w1469 & ~pi09974;
assign w55128 = w1485 & pi09944;
assign w55129 = ~w1550 & w1556;
assign w55130 = ~w1499 & pi00333;
assign w55131 = w1584 & ~pi00147;
assign w55132 = w1499 & w1589;
assign w55133 = ~w1499 & ~pi00322;
assign w55134 = w54762 & ~pi00104;
assign w55135 = ~w54762 & pi00104;
assign w55136 = w1499 & w1596;
assign w55137 = ~pi10471 & ~pi00105;
assign w55138 = pi10471 & ~pi10572;
assign w55139 = ~w55083 & ~pi10571;
assign w55140 = w1616 & w1620;
assign w55141 = ~w55083 & ~pi10570;
assign w55142 = w1637 & w1641;
assign w55143 = ~w55083 & ~pi10564;
assign w55144 = w1660 & w1664;
assign w55145 = ~w55083 & ~pi10562;
assign w55146 = w1683 & w1687;
assign w55147 = ~w55083 & ~pi10567;
assign w55148 = ~w55083 & ~pi10573;
assign w55149 = w1740 & w1744;
assign w55150 = ~w55083 & ~pi10560;
assign w55151 = ~pi10432 & ~pi00113;
assign w55152 = pi10432 & pi10574;
assign w55153 = ~w1789 & ~pi00114;
assign w55154 = ~pi00131 & ~pi00115;
assign w55155 = ~w55096 & ~w1194;
assign w55156 = pi10471 & pi10570;
assign w55157 = ~w55083 & ~pi10566;
assign w55158 = w55097 & pi00128;
assign w55159 = ~pi00117 & ~w1194;
assign w55160 = pi10471 & pi10573;
assign w55161 = ~w55083 & ~pi10569;
assign w55162 = pi10471 & pi10560;
assign w55163 = ~pi00119 & ~pi00120;
assign w55164 = pi10471 & pi10567;
assign w55165 = pi10471 & pi10562;
assign w55166 = w54706 & pi00180;
assign w55167 = pi00123 & pi00135;
assign w55168 = w55167 & pi00122;
assign w55169 = ~w55167 & ~pi00122;
assign w55170 = ~w55168 & ~w1371;
assign w55171 = pi10432 & pi10566;
assign w55172 = ~pi00123 & ~w1371;
assign w55173 = pi10432 & pi10573;
assign w55174 = pi10432 & pi10560;
assign w55175 = w55096 & w1878;
assign w55176 = ~pi00125 & ~w1194;
assign w55177 = pi10471 & pi10566;
assign w55178 = ~pi00124 & ~pi00126;
assign w55179 = pi10432 & pi10567;
assign w55180 = ~pi00127 & ~w1371;
assign w55181 = pi10432 & pi10562;
assign w55182 = ~w55097 & ~pi00128;
assign w55183 = pi10471 & pi10571;
assign w55184 = pi10471 & pi10569;
assign w55185 = ~pi00117 & ~pi00129;
assign w55186 = ~w54752 & ~pi00130;
assign w55187 = ~w55105 & ~w1371;
assign w55188 = pi10432 & pi10570;
assign w55189 = ~pi00131 & ~w1194;
assign w55190 = pi10471 & pi10564;
assign w55191 = ~pi09928 & pi00132;
assign w55192 = pi09928 & ~pi10569;
assign w55193 = ~pi09928 & pi00133;
assign w55194 = pi09928 & ~pi10566;
assign w55195 = ~w55107 & ~pi00134;
assign w55196 = pi10432 & pi10571;
assign w55197 = ~pi00123 & ~pi00135;
assign w55198 = ~w55167 & ~w1371;
assign w55199 = pi10432 & pi10569;
assign w55200 = ~pi00127 & ~pi00136;
assign w55201 = pi10432 & pi10564;
assign w55202 = ~pi09997 & pi00137;
assign w55203 = pi09997 & pi10571;
assign w55204 = ~pi09997 & pi00138;
assign w55205 = pi09997 & pi10573;
assign w55206 = ~pi09997 & pi00139;
assign w55207 = pi09997 & ~pi10569;
assign w55208 = ~pi09997 & pi00140;
assign w55209 = pi09997 & ~pi10566;
assign w55210 = pi00343 & w76;
assign w55211 = ~w54860 & pi00142;
assign w55212 = w54860 & ~pi00142;
assign w55213 = w1499 & w1957;
assign w55214 = ~w1499 & pi00323;
assign w55215 = ~w55212 & pi00143;
assign w55216 = w55212 & ~pi00143;
assign w55217 = w1499 & w1963;
assign w55218 = ~w1499 & pi00324;
assign w55219 = w55216 & ~pi00152;
assign w55220 = ~w55219 & pi00144;
assign w55221 = w55219 & ~pi00144;
assign w55222 = w1499 & w1970;
assign w55223 = ~w1499 & pi00332;
assign w55224 = ~w1499 & pi00328;
assign w55225 = ~w55134 & pi00145;
assign w55226 = ~w1584 & ~w1975;
assign w55227 = w1499 & w1976;
assign w55228 = ~w1499 & ~pi00327;
assign w55229 = w1499 & w54715;
assign w55230 = ~w1584 & pi00147;
assign w55231 = w1499 & w1984;
assign w55232 = ~w1499 & pi00329;
assign w55233 = w1499 & w1989;
assign w55234 = ~w1499 & pi00335;
assign w55235 = ~w1499 & pi00336;
assign w55236 = ~pi00148 & ~pi00155;
assign w55237 = ~w55236 & pi00149;
assign w55238 = w1499 & w1996;
assign w55239 = ~w54763 & pi00150;
assign w55240 = w1499 & w2000;
assign w55241 = ~w1499 & pi00330;
assign w55242 = ~w54786 & pi00151;
assign w55243 = w54786 & ~pi00151;
assign w55244 = w1499 & w2006;
assign w55245 = ~w1499 & pi00331;
assign w55246 = ~w55216 & pi00152;
assign w55247 = w1499 & w2011;
assign w55248 = ~w1499 & pi00325;
assign w55249 = w1499 & w54716;
assign w55250 = ~w1499 & pi00326;
assign w55251 = ~w1499 & pi00334;
assign w55252 = w1499 & w2021;
assign w55253 = pi00148 & pi00155;
assign w55254 = w1499 & w2025;
assign w55255 = ~w1499 & pi00337;
assign w55256 = w827 & ~w2042;
assign w55257 = ~pi00114 & pi00292;
assign w55258 = pi00114 & ~w2048;
assign w55259 = ~w2046 & w2044;
assign w55260 = ~w2036 & w2057;
assign w55261 = pi09997 & pi00321;
assign w55262 = w2036 & ~pi00156;
assign w55263 = ~w2058 & ~w2057;
assign w55264 = ~w2058 & ~w55260;
assign w55265 = w1113 & pi10486;
assign w55266 = w1113 & ~pi00309;
assign w55267 = ~pi09997 & ~pi00174;
assign w55268 = ~w1789 & ~pi00175;
assign w55269 = ~w55083 & ~pi10565;
assign w55270 = ~pi10432 & ~pi00177;
assign w55271 = ~w55083 & ~pi10574;
assign w55272 = pi10654 & pi00842;
assign w55273 = w2169 & w1226;
assign w55274 = ~w55083 & ~pi10563;
assign w55275 = ~w54706 & ~pi00180;
assign w55276 = pi10471 & pi10565;
assign w55277 = ~w54707 & ~pi00181;
assign w55278 = pi10432 & pi10565;
assign w55279 = pi10471 & pi10563;
assign w55280 = ~pi00125 & ~pi00182;
assign w55281 = ~w55168 & ~pi00183;
assign w55282 = w55168 & pi00183;
assign w55283 = pi10432 & pi10563;
assign w55284 = ~pi00024 & pi00358;
assign w55285 = pi00024 & ~pi00358;
assign w55286 = w671 & ~pi00358;
assign w55287 = w671 & ~w55284;
assign w55288 = ~pi00024 & pi00359;
assign w55289 = pi00024 & ~pi00359;
assign w55290 = ~pi00361 & w76;
assign w55291 = w1142 & ~pi00360;
assign w55292 = ~w1142 & pi00360;
assign w55293 = ~w2275 & ~pi00271;
assign w55294 = w145 & w642;
assign w55295 = ~w2275 & pi00188;
assign w55296 = w145 & w2283;
assign w55297 = ~w2291 & ~pi09873;
assign w55298 = ~w2294 & ~w2290;
assign w55299 = ~w2296 & w145;
assign w55300 = ~w2289 & w2285;
assign w55301 = ~w2032 & w2301;
assign w55302 = pi09997 & pi00344;
assign w55303 = w2032 & ~pi00189;
assign w55304 = ~w2302 & ~w2301;
assign w55305 = ~w2302 & ~w55301;
assign w55306 = w55303 & ~pi00191;
assign w55307 = ~w827 & pi00190;
assign w55308 = ~w55306 & w2306;
assign w55309 = pi09997 & pi00346;
assign w55310 = w55306 & ~pi00190;
assign w55311 = ~w2307 & ~w2306;
assign w55312 = ~w2307 & ~w55308;
assign w55313 = ~w55303 & w2311;
assign w55314 = pi09997 & pi00345;
assign w55315 = ~w55306 & ~w2313;
assign w55316 = w1217 & pi09939;
assign w55317 = w1244 & pi10252;
assign w55318 = ~w55083 & pi00321;
assign w55319 = w1242 & pi10009;
assign w55320 = w1230 & pi10241;
assign w55321 = ~pi09997 & ~pi00193;
assign w55322 = ~pi09997 & ~pi00194;
assign w55323 = pi09997 & pi10558;
assign w55324 = ~pi09997 & ~pi00195;
assign w55325 = pi09997 & pi00347;
assign w55326 = ~pi09997 & ~pi00196;
assign w55327 = ~pi09997 & ~pi00197;
assign w55328 = ~w55083 & ~pi10572;
assign w55329 = w54821 & pi00220;
assign w55330 = pi00221 & pi00222;
assign w55331 = w55330 & pi00199;
assign w55332 = ~w55330 & ~pi00199;
assign w55333 = ~w55331 & ~w1194;
assign w55334 = pi10471 & pi00321;
assign w55335 = w54822 & w2399;
assign w55336 = w2403 & w2405;
assign w55337 = w55336 & pi00200;
assign w55338 = ~w55336 & ~pi00200;
assign w55339 = ~w55337 & ~w1371;
assign w55340 = pi10432 & pi00321;
assign w55341 = w2036 & w54791;
assign w55342 = w55341 & ~pi00208;
assign w55343 = ~w55342 & w2412;
assign w55344 = w54792 | w2415;
assign w55345 = (w2415 & w54792) | (w2415 & ~w55306) | (w54792 & ~w55306);
assign w55346 = pi00814 & ~pi00320;
assign w55347 = ~pi00230 & ~pi00203;
assign w55348 = w2423 & ~w2428;
assign w55349 = w144 & pi00249;
assign w55350 = ~pi00250 & ~w2431;
assign w55351 = pi00204 & ~w2431;
assign w55352 = pi00204 & w55350;
assign w55353 = ~pi00869 & ~w55351;
assign w55354 = ~pi00869 & ~w55352;
assign w55355 = ~w54996 & pi00366;
assign w55356 = w54996 & ~pi00366;
assign w55357 = ~w55262 & w2442;
assign w55358 = pi09997 & pi10561;
assign w55359 = ~w55341 & ~w2444;
assign w55360 = pi09997 & pi00363;
assign w55361 = ~w827 & pi00208;
assign w55362 = ~w55341 & w2456;
assign w55363 = pi09997 & pi00364;
assign w55364 = w54787 & pi00267;
assign w55365 = ~w2461 & w2044;
assign w55366 = w55365 & ~pi00268;
assign w55367 = w1217 & pi09988;
assign w55368 = w1244 & pi10253;
assign w55369 = ~w55083 & pi00347;
assign w55370 = w1242 & pi10008;
assign w55371 = w1230 & pi10022;
assign w55372 = w1217 & pi09941;
assign w55373 = w1242 & pi10260;
assign w55374 = ~w55083 & pi10558;
assign w55375 = w1244 & pi10251;
assign w55376 = w1230 & pi10021;
assign w55377 = w1217 & pi09981;
assign w55378 = w1244 & pi10249;
assign w55379 = ~w55083 & pi00344;
assign w55380 = w1242 & pi10011;
assign w55381 = w1230 & pi10023;
assign w55382 = w1217 & pi09982;
assign w55383 = w1244 & pi10013;
assign w55384 = ~w55083 & pi00346;
assign w55385 = w1242 & pi10010;
assign w55386 = w1230 & pi10238;
assign w55387 = w1217 & pi09942;
assign w55388 = w1242 & pi10259;
assign w55389 = ~w55083 & pi00345;
assign w55390 = w1244 & pi10250;
assign w55391 = w1230 & pi10239;
assign w55392 = ~pi09997 & ~pi00215;
assign w55393 = ~pi09997 & ~pi00216;
assign w55394 = ~pi09997 & ~pi00217;
assign w55395 = ~pi09997 & ~pi00218;
assign w55396 = pi09997 & pi00362;
assign w55397 = pi10471 & pi00344;
assign w55398 = w54789 & pi00262;
assign w55399 = ~w55398 & ~pi00219;
assign w55400 = ~w54821 & ~w1194;
assign w55401 = ~w54821 & ~pi00220;
assign w55402 = pi10471 & pi00345;
assign w55403 = ~pi00221 & ~w1194;
assign w55404 = pi10471 & pi00346;
assign w55405 = ~pi00221 & ~pi00222;
assign w55406 = pi10471 & pi10558;
assign w55407 = w55330 & w2542;
assign w55408 = w55407 & ~pi00251;
assign w55409 = ~w55408 & ~pi00223;
assign w55410 = w55408 & pi00223;
assign w55411 = pi10471 & pi00347;
assign w55412 = pi10432 & pi10558;
assign w55413 = w2403 & pi00225;
assign w55414 = ~w55413 & ~pi00224;
assign w55415 = ~w55336 & ~w1371;
assign w55416 = ~w2403 & ~pi00225;
assign w55417 = ~w55413 & ~w1371;
assign w55418 = pi10432 & pi00346;
assign w55419 = w55336 & w2560;
assign w55420 = pi00252 & ~pi00226;
assign w55421 = ~pi00252 & pi00226;
assign w55422 = pi10432 & pi00347;
assign w55423 = w2402 & pi00227;
assign w55424 = ~w2402 & ~pi00227;
assign w55425 = ~w55423 & ~w1371;
assign w55426 = pi10432 & pi00344;
assign w55427 = pi10432 & pi00345;
assign w55428 = ~w55423 & ~pi00228;
assign w55429 = ~pi00269 & ~pi00270;
assign w55430 = ~w55429 & w2579;
assign w55431 = ~w2032 & ~w2520;
assign w55432 = w1122 & ~w1123;
assign w55433 = w55012 & w1080;
assign w55434 = w2588 & ~pi00373;
assign w55435 = ~w2588 & pi00373;
assign w55436 = pi00232 & ~w2431;
assign w55437 = pi00232 & w55350;
assign w55438 = ~pi00869 & ~w55436;
assign w55439 = ~pi00869 & ~w55437;
assign w55440 = w145 & ~w2597;
assign w55441 = w145 & ~w54766;
assign w55442 = w2284 & w145;
assign w55443 = w54825 & w2598;
assign w55444 = w55443 & pi00244;
assign w55445 = w55444 & w1482;
assign w55446 = ~w55445 & ~pi00234;
assign w55447 = w55445 & pi00234;
assign w55448 = ~w55447 & ~pi00235;
assign w55449 = w55447 & pi00235;
assign w55450 = w55445 & w1481;
assign w55451 = w2616 & w1484;
assign w55452 = ~w55450 & ~pi00237;
assign w55453 = ~pi00238 & ~w2609;
assign w55454 = ~pi00240 & ~pi00241;
assign w55455 = ~w54825 & ~pi00242;
assign w55456 = w54825 & pi00242;
assign w55457 = ~w55456 & ~pi00243;
assign w55458 = ~w55443 & ~pi00244;
assign w55459 = ~w55444 & ~pi00245;
assign w55460 = w55444 & pi00245;
assign w55461 = ~w55460 & ~pi00246;
assign w55462 = w2616 & w1410;
assign w55463 = w2609 & pi00247;
assign w55464 = w2616 & w1411;
assign w55465 = pi00249 & ~pi00250;
assign w55466 = ~w55407 & pi00251;
assign w55467 = ~w55408 & ~w1194;
assign w55468 = pi10471 & pi00363;
assign w55469 = ~w55419 & pi00252;
assign w55470 = pi00252 & ~w1371;
assign w55471 = pi10432 & pi00363;
assign w55472 = w1217 & pi09985;
assign w55473 = w1242 & pi10261;
assign w55474 = ~w55083 & pi00363;
assign w55475 = w1244 & pi10015;
assign w55476 = w1230 & pi10242;
assign w55477 = w1217 & pi09903;
assign w55478 = w1242 & pi10258;
assign w55479 = ~w55083 & pi00362;
assign w55480 = w1244 & pi10248;
assign w55481 = w1230 & pi10024;
assign w55482 = w1217 & pi09900;
assign w55483 = w1242 & pi10257;
assign w55484 = ~w55083 & pi00364;
assign w55485 = w1244 & pi10246;
assign w55486 = w1230 & pi10237;
assign w55487 = w1217 & pi09984;
assign w55488 = w1244 & pi10017;
assign w55489 = ~w55083 & pi10561;
assign w55490 = w1242 & pi10007;
assign w55491 = w1230 & pi10240;
assign w55492 = ~pi09997 & ~pi00257;
assign w55493 = pi09997 & pi00369;
assign w55494 = ~pi09997 & ~pi00258;
assign w55495 = pi09997 & pi00370;
assign w55496 = ~pi09997 & ~pi00259;
assign w55497 = pi09997 & pi00368;
assign w55498 = ~pi09997 & ~pi00260;
assign w55499 = pi09997 & pi00367;
assign w55500 = ~pi00284 & ~pi00261;
assign w55501 = ~w54765 & ~w1194;
assign w55502 = pi10471 & pi00364;
assign w55503 = ~w54789 & ~pi00262;
assign w55504 = ~w55398 & ~w1194;
assign w55505 = pi10471 & pi00362;
assign w55506 = pi10471 & pi10561;
assign w55507 = ~w55331 & ~pi00263;
assign w55508 = pi10432 & pi00364;
assign w55509 = w54822 & pi00293;
assign w55510 = ~pi00287 & ~pi00264;
assign w55511 = ~w1371 & pi00264;
assign w55512 = ~w1371 & ~w55510;
assign w55513 = ~pi00288 & ~pi00265;
assign w55514 = ~w2402 & ~w1371;
assign w55515 = pi10432 & pi00362;
assign w55516 = pi10432 & pi10561;
assign w55517 = ~w55337 & ~pi00266;
assign w55518 = ~pi00267 & ~w2721;
assign w55519 = w2461 & pi00268;
assign w55520 = ~pi09997 & pi00269;
assign w55521 = w2046 & w2768;
assign w55522 = ~w827 & pi00270;
assign w55523 = ~w55429 & ~w2727;
assign w55524 = ~w2779 & pi00301;
assign w55525 = pi00272 & pi00277;
assign w55526 = w55525 & pi00275;
assign w55527 = ~w55526 & ~pi00273;
assign w55528 = w55526 & pi00273;
assign w55529 = ~w55525 & ~pi00275;
assign w55530 = w2296 & ~pi00276;
assign w55531 = ~pi00272 & ~pi00277;
assign w55532 = w1217 & pi09902;
assign w55533 = w1244 & pi10018;
assign w55534 = ~w55083 & pi00368;
assign w55535 = w1242 & pi10012;
assign w55536 = w1230 & pi10025;
assign w55537 = w1217 & pi09901;
assign w55538 = w1244 & pi10247;
assign w55539 = ~w55083 & pi00367;
assign w55540 = w1242 & pi10233;
assign w55541 = w1230 & pi10236;
assign w55542 = ~pi09997 & ~pi00280;
assign w55543 = pi09997 & pi00371;
assign w55544 = ~pi09997 & ~pi00281;
assign w55545 = pi09997 & pi00372;
assign w55546 = w1242 & pi10255;
assign w55547 = w1217 & pi09898;
assign w55548 = w1230 & pi10234;
assign w55549 = ~w55083 & pi00369;
assign w55550 = w1266 & pi09813;
assign w55551 = w1244 & pi10245;
assign w55552 = w1217 & pi09899;
assign w55553 = w1244 & pi10019;
assign w55554 = w1230 & pi10235;
assign w55555 = ~w55083 & pi00370;
assign w55556 = w1266 & pi09847;
assign w55557 = w1242 & pi10256;
assign w55558 = ~pi00284 & ~w1194;
assign w55559 = pi10471 & pi00370;
assign w55560 = ~w54765 & ~pi00285;
assign w55561 = pi10471 & pi00367;
assign w55562 = ~w54788 & ~pi00286;
assign w55563 = ~w54789 & ~w1194;
assign w55564 = pi10471 & pi00368;
assign w55565 = ~pi00287 & ~w1371;
assign w55566 = pi10432 & pi00370;
assign w55567 = ~pi00288 & ~w1371;
assign w55568 = pi10432 & pi00368;
assign w55569 = pi10432 & pi00367;
assign w55570 = ~w2397 & ~pi00289;
assign w55571 = ~w1355 & ~pi00290;
assign w55572 = pi10471 & pi00369;
assign w55573 = w2042 & pi00291;
assign w55574 = pi00291 & ~w2820;
assign w55575 = pi00114 & ~pi00292;
assign w55576 = ~w2887 & ~w2823;
assign w55577 = ~w54822 & ~pi00293;
assign w55578 = pi10432 & pi00369;
assign w55579 = ~w2900 & ~pi00320;
assign w55580 = w2902 & ~w2899;
assign w55581 = pi00308 & pi00309;
assign w55582 = ~w55581 & ~pi00295;
assign w55583 = w55581 & pi00295;
assign w55584 = pi00296 & ~pi00841;
assign w55585 = ~pi00024 & ~w793;
assign w55586 = ~pi00402 & w671;
assign w55587 = pi00024 & w742;
assign w55588 = pi00401 & w671;
assign w55589 = ~pi00241 & w2930;
assign w55590 = ~w55589 & ~w2928;
assign w55591 = ~pi00241 & pi00250;
assign w55592 = ~pi00241 & w2943;
assign w55593 = pi00241 & ~w78;
assign w55594 = w2954 & ~w2944;
assign w55595 = w2951 & w2950;
assign w55596 = ~w2958 & ~w2950;
assign w55597 = ~w2958 & ~w55595;
assign w55598 = w2779 & ~pi00301;
assign w55599 = ~w55083 & pi00371;
assign w55600 = w1242 & pi10014;
assign w55601 = w1217 & pi09897;
assign w55602 = w1266 & pi09846;
assign w55603 = ~pi00304 & ~w1194;
assign w55604 = pi10471 & pi00371;
assign w55605 = pi10471 & pi00372;
assign w55606 = ~pi00304 & ~pi00305;
assign w55607 = w55282 & pi00306;
assign w55608 = ~w55282 & ~pi00306;
assign w55609 = pi10432 & pi00371;
assign w55610 = pi10432 & pi00372;
assign w55611 = ~w54822 & ~w1371;
assign w55612 = w852 & w1116;
assign w55613 = ~pi00308 & ~pi00841;
assign w55614 = pi00296 & pi00310;
assign w55615 = ~pi00841 & pi00310;
assign w55616 = ~pi00841 & ~w55032;
assign w55617 = w852 & w856;
assign w55618 = pi01272 & ~pi00312;
assign w55619 = pi01272 & ~pi10520;
assign w55620 = pi01272 & ~pi00313;
assign w55621 = pi01272 & ~pi10495;
assign w55622 = pi01272 & ~pi00314;
assign w55623 = pi01272 & pi10486;
assign w55624 = pi01272 & ~pi00315;
assign w55625 = pi01272 & ~pi10492;
assign w55626 = pi01272 & ~pi00316;
assign w55627 = pi01272 & ~pi10505;
assign w55628 = pi01272 & ~pi00317;
assign w55629 = pi01272 & pi10483;
assign w55630 = pi01272 & ~pi00318;
assign w55631 = pi01272 & pi10511;
assign w55632 = pi01272 & ~pi00319;
assign w55633 = ~pi00342 & pi00320;
assign w55634 = pi00338 & ~pi00349;
assign w55635 = ~pi00338 & ~pi10516;
assign w55636 = ~pi00322 & ~pi10516;
assign w55637 = ~pi00322 & w55635;
assign w55638 = pi00338 & ~pi00312;
assign w55639 = ~pi00323 & ~pi10516;
assign w55640 = ~pi00323 & w55635;
assign w55641 = pi00338 & ~pi00314;
assign w55642 = ~pi00324 & ~pi10516;
assign w55643 = ~pi00324 & w55635;
assign w55644 = pi00338 & ~pi00313;
assign w55645 = ~pi00325 & ~pi10516;
assign w55646 = ~pi00325 & w55635;
assign w55647 = pi00338 & ~pi00316;
assign w55648 = ~pi00326 & ~pi10516;
assign w55649 = ~pi00326 & w55635;
assign w55650 = pi00338 & ~pi00317;
assign w55651 = ~pi00327 & ~pi10516;
assign w55652 = ~pi00327 & w55635;
assign w55653 = pi00338 & ~pi00355;
assign w55654 = ~pi00328 & ~pi10516;
assign w55655 = ~pi00328 & w55635;
assign w55656 = pi00338 & ~pi00352;
assign w55657 = ~pi00329 & ~pi10516;
assign w55658 = ~pi00329 & w55635;
assign w55659 = pi00338 & ~pi00350;
assign w55660 = ~pi00330 & ~pi10516;
assign w55661 = ~pi00330 & w55635;
assign w55662 = pi00338 & ~pi00351;
assign w55663 = ~pi00331 & ~pi10516;
assign w55664 = ~pi00331 & w55635;
assign w55665 = pi00338 & ~pi00315;
assign w55666 = ~pi00332 & ~pi10516;
assign w55667 = ~pi00332 & w55635;
assign w55668 = pi00338 & ~pi00354;
assign w55669 = ~pi00333 & ~pi10516;
assign w55670 = ~pi00333 & w55635;
assign w55671 = pi00338 & ~pi00353;
assign w55672 = ~pi00334 & ~pi10516;
assign w55673 = ~pi00334 & w55635;
assign w55674 = pi00338 & ~pi00356;
assign w55675 = ~pi00335 & ~pi10516;
assign w55676 = ~pi00335 & w55635;
assign w55677 = pi00338 & ~pi00319;
assign w55678 = ~pi00336 & ~pi10516;
assign w55679 = ~pi00336 & w55635;
assign w55680 = pi00338 & ~pi00318;
assign w55681 = w3933 & pi00063;
assign w55682 = ~w55681 & ~pi00338;
assign w55683 = w2900 & pi00340;
assign w55684 = ~pi00340 & ~pi00341;
assign w55685 = w1142 & ~pi00879;
assign w55686 = ~w1142 & pi00879;
assign w55687 = ~pi00365 & ~w1121;
assign w55688 = pi00365 & ~pi00348;
assign w55689 = w852 & w896;
assign w55690 = pi01272 & ~pi00349;
assign w55691 = pi01272 & ~pi00350;
assign w55692 = pi01272 & ~pi00351;
assign w55693 = pi01272 & ~pi00352;
assign w55694 = pi01272 & ~pi00353;
assign w55695 = pi01272 & ~pi00354;
assign w55696 = pi01272 & ~pi00355;
assign w55697 = pi01272 & ~pi10489;
assign w55698 = pi01272 & ~pi00356;
assign w55699 = ~w3933 & ~pi00357;
assign w55700 = ~pi00463 & w671;
assign w55701 = ~pi00024 & ~w743;
assign w55702 = ~pi00464 & w671;
assign w55703 = w2588 & ~pi01166;
assign w55704 = ~w2588 & pi01166;
assign w55705 = w2588 & ~pi00472;
assign w55706 = ~w2588 & pi00472;
assign w55707 = pi00465 & w76;
assign w55708 = w2286 & w78;
assign w55709 = ~pi01454 & ~pi01312;
assign w55710 = ~w10691 & w10685;
assign w55711 = pi01274 & ~pi00461;
assign w55712 = ~w10690 & ~pi00460;
assign w55713 = pi01274 & pi00474;
assign w55714 = ~w10683 & pi00474;
assign w55715 = ~w10683 & w55713;
assign w55716 = w10705 & w10717;
assign w55717 = ~pi00461 & ~pi00474;
assign w55718 = w10710 & pi00098;
assign w55719 = w10748 & pi00377;
assign w55720 = ~w10748 & ~pi10520;
assign w55721 = w10748 & pi00378;
assign w55722 = ~w10748 & pi10486;
assign w55723 = w10748 & pi00379;
assign w55724 = ~w10748 & ~pi10495;
assign w55725 = w10748 & pi00380;
assign w55726 = ~w10748 & ~pi10492;
assign w55727 = w10748 & pi00381;
assign w55728 = ~w10748 & ~pi10505;
assign w55729 = w10748 & pi00382;
assign w55730 = ~w10748 & pi10483;
assign w55731 = w10748 & pi00399;
assign w55732 = ~w10748 & pi10511;
assign w55733 = w10748 & pi00400;
assign w55734 = ~w10748 & ~pi10489;
assign w55735 = ~pi00024 & pi00537;
assign w55736 = pi00024 & ~pi00537;
assign w55737 = w671 & ~pi00537;
assign w55738 = w671 & ~w55735;
assign w55739 = ~pi00536 & w671;
assign w55740 = w54826 & w10851;
assign w55741 = w55740 & pi00405;
assign w55742 = w55741 & pi00419;
assign w55743 = w55742 & w10855;
assign w55744 = ~pi00403 & w10856;
assign w55745 = w10723 & pi00403;
assign w55746 = w10710 & ~pi00252;
assign w55747 = w10710 & pi00293;
assign w55748 = pi00407 & pi00431;
assign w55749 = w55748 & pi00408;
assign w55750 = w55749 & pi00409;
assign w55751 = w55750 & pi00410;
assign w55752 = w10723 & pi00404;
assign w55753 = ~w10873 & w10872;
assign w55754 = w10849 & pi00416;
assign w55755 = w10723 & pi00405;
assign w55756 = w10710 & pi00225;
assign w55757 = w10723 & pi00406;
assign w55758 = ~w10839 & w10838;
assign w55759 = w10710 & pi00123;
assign w55760 = w10723 & pi00407;
assign w55761 = w10710 & pi00135;
assign w55762 = ~pi00407 & w10839;
assign w55763 = ~pi00408 & w10869;
assign w55764 = w10723 & pi00408;
assign w55765 = w10710 & pi00183;
assign w55766 = w10723 & pi00409;
assign w55767 = ~w10871 & w10870;
assign w55768 = w10710 & pi00306;
assign w55769 = ~pi00410 & w10871;
assign w55770 = w10710 & pi00307;
assign w55771 = ~pi00411 & w10873;
assign w55772 = w10710 & pi00287;
assign w55773 = ~w10846 & pi00411;
assign w55774 = w55773 & w10873;
assign w55775 = w10939 & pi00412;
assign w55776 = w10710 & pi00264;
assign w55777 = w10939 & pi00413;
assign w55778 = ~pi00413 & w10847;
assign w55779 = w10723 & pi00414;
assign w55780 = w10710 & pi00288;
assign w55781 = ~w10849 & ~w10963;
assign w55782 = ~w10849 & ~pi00416;
assign w55783 = w10710 & pi00265;
assign w55784 = w10710 & pi00227;
assign w55785 = w10723 & pi00417;
assign w55786 = w54826 & pi00417;
assign w55787 = ~w10852 & w10985;
assign w55788 = w10723 & pi00418;
assign w55789 = w10710 & pi00228;
assign w55790 = w10710 & pi00224;
assign w55791 = w10723 & pi00419;
assign w55792 = ~w10854 & w10853;
assign w55793 = w10710 & pi00200;
assign w55794 = w10723 & pi00420;
assign w55795 = w10854 & ~pi00420;
assign w55796 = w10723 & pi00421;
assign w55797 = w10710 & pi00266;
assign w55798 = w10854 & w11011;
assign w55799 = w10857 & pi00422;
assign w55800 = w11019 & w10856;
assign w55801 = w10723 & pi00423;
assign w55802 = w10710 & pi00126;
assign w55803 = pi00432 & ~pi00423;
assign w55804 = w10710 & pi00181;
assign w55805 = w10723 & pi00424;
assign w55806 = ~w10833 & w10832;
assign w55807 = w10723 & pi00425;
assign w55808 = pi00424 & ~pi00425;
assign w55809 = w10710 & pi00136;
assign w55810 = w10723 & pi00426;
assign w55811 = ~w10835 & w10834;
assign w55812 = w10723 & pi00427;
assign w55813 = w10710 & pi00097;
assign w55814 = w10723 & pi00428;
assign w55815 = ~w10837 & w10836;
assign w55816 = w54741 & ~pi00429;
assign w55817 = w10723 & pi00429;
assign w55818 = w10710 & pi00122;
assign w55819 = w10723 & pi00431;
assign w55820 = w10710 & pi00124;
assign w55821 = w10723 & pi00432;
assign w55822 = ~pi01274 & ~w10694;
assign w55823 = w11106 & ~w11105;
assign w55824 = w54865 & w11115;
assign w55825 = ~w55824 & pi00250;
assign w55826 = ~pi10472 & ~pi00436;
assign w55827 = ~w831 & pi00438;
assign w55828 = ~w831 & ~pi00439;
assign w55829 = w2049 & w11132;
assign w55830 = pi00442 & pi00460;
assign w55831 = pi00461 & pi00474;
assign w55832 = pi00461 & w55713;
assign w55833 = ~w11104 & ~w11138;
assign w55834 = pi00457 & pi00458;
assign w55835 = ~pi00267 & ~pi00268;
assign w55836 = w11151 & w11152;
assign w55837 = w55589 & pi00812;
assign w55838 = ~w11176 & ~w11175;
assign w55839 = ~w11180 & pi00447;
assign w55840 = w11183 & pi01187;
assign w55841 = pi10000 & pi01270;
assign w55842 = ~w11184 & ~w11181;
assign w55843 = ~w11180 & pi00448;
assign w55844 = w11183 & pi01188;
assign w55845 = ~w11213 & ~w11212;
assign w55846 = ~w11180 & pi00449;
assign w55847 = w11183 & pi01189;
assign w55848 = ~w11230 & ~w11229;
assign w55849 = ~w11180 & pi00450;
assign w55850 = w11183 & pi01190;
assign w55851 = ~w11247 & ~w11246;
assign w55852 = w11183 & pi01191;
assign w55853 = ~w11180 & pi00451;
assign w55854 = w11183 & pi01195;
assign w55855 = ~w11180 & pi00452;
assign w55856 = w11183 & pi01194;
assign w55857 = ~w11180 & pi00453;
assign w55858 = w11183 & pi01192;
assign w55859 = ~w11180 & pi00454;
assign w55860 = ~pi01204 & ~pi01214;
assign w55861 = w55860 & ~pi00959;
assign w55862 = ~pi01205 & pi10231;
assign w55863 = ~w55862 & ~pi00455;
assign w55864 = w11347 & ~pi01307;
assign w55865 = ~pi01308 & ~pi01305;
assign w55866 = pi01309 & pi01307;
assign w55867 = w11347 & pi01307;
assign w55868 = pi09833 & ~w11362;
assign w55869 = ~w11365 & w11342;
assign w55870 = ~w55862 & pi00456;
assign w55871 = ~w11378 & w11368;
assign w55872 = ~w11105 & pi00458;
assign w55873 = ~w55834 & ~pi00459;
assign w55874 = w11140 & pi00460;
assign w55875 = w11140 & pi00461;
assign w55876 = ~pi00024 & pi00824;
assign w55877 = pi00024 & ~pi00824;
assign w55878 = ~pi00825 & w671;
assign w55879 = ~w55862 & ~pi00466;
assign w55880 = ~w11342 & ~w11410;
assign w55881 = ~w55862 & ~pi00467;
assign w55882 = ~w11342 & ~w11421;
assign w55883 = ~w55862 & ~pi00468;
assign w55884 = ~w11342 & ~w11432;
assign w55885 = ~w55862 & ~pi00469;
assign w55886 = ~w11342 & ~w11443;
assign w55887 = ~pi00089 & ~pi00105;
assign w55888 = ~pi01167 & w76;
assign w55889 = ~pi10472 & ~pi00473;
assign w55890 = ~pi00461 & pi01454;
assign w55891 = pi00540 & pi00488;
assign w55892 = ~pi10662 & pi10578;
assign w55893 = w55892 & pi10664;
assign w55894 = ~w11485 & pi00477;
assign w55895 = w11485 & pi10591;
assign w55896 = ~w11485 & pi00478;
assign w55897 = w11485 & pi10593;
assign w55898 = ~w11485 & pi00479;
assign w55899 = w11485 & pi10595;
assign w55900 = ~w11485 & pi00480;
assign w55901 = w11485 & pi10594;
assign w55902 = ~w11485 & pi00481;
assign w55903 = w11485 & pi10596;
assign w55904 = ~w11485 & pi00482;
assign w55905 = w11485 & pi10592;
assign w55906 = ~w11485 & pi00483;
assign w55907 = w11485 & pi10597;
assign w55908 = ~w11485 & pi00484;
assign w55909 = w11485 & pi10590;
assign w55910 = ~w55862 & ~pi00485;
assign w55911 = w11545 & w11342;
assign w55912 = ~w55862 & ~pi00486;
assign w55913 = w11553 & w11342;
assign w55914 = ~pi10254 & pi00876;
assign w55915 = ~w11568 & w11569;
assign w55916 = ~pi10243 & ~pi00876;
assign w55917 = ~w11574 & w11575;
assign w55918 = ~w11580 & pi00874;
assign w55919 = ~pi10252 & ~pi00876;
assign w55920 = ~w11602 & w11603;
assign w55921 = ~pi09917 & pi00876;
assign w55922 = ~w11608 & w11609;
assign w55923 = ~w11588 & ~pi00874;
assign w55924 = ~pi09915 & pi00876;
assign w55925 = ~w11635 & w11636;
assign w55926 = ~pi09906 & ~pi00876;
assign w55927 = ~w11641 & w11642;
assign w55928 = ~pi10018 & ~pi00876;
assign w55929 = ~w11667 & w11668;
assign w55930 = ~pi09994 & pi00876;
assign w55931 = ~w11673 & w11674;
assign w55932 = w11631 & w11560;
assign w55933 = ~pi01274 & w11707;
assign w55934 = ~pi00541 & w11710;
assign w55935 = ~w11705 & pi00489;
assign w55936 = w11705 & ~pi00074;
assign w55937 = ~w11705 & pi00490;
assign w55938 = w11705 & ~pi00080;
assign w55939 = ~w11705 & pi00491;
assign w55940 = w11705 & ~pi00168;
assign w55941 = ~w11705 & pi00492;
assign w55942 = w11705 & ~pi00160;
assign w55943 = ~w11705 & pi00493;
assign w55944 = w11705 & ~pi00164;
assign w55945 = ~w11705 & pi00494;
assign w55946 = w11705 & ~pi00082;
assign w55947 = ~w11705 & pi00495;
assign w55948 = w11705 & ~pi00085;
assign w55949 = ~w11733 & pi00496;
assign w55950 = w11733 & ~pi00075;
assign w55951 = ~w11733 & pi00497;
assign w55952 = w11733 & ~pi00080;
assign w55953 = ~w11733 & pi00498;
assign w55954 = w11733 & ~pi00078;
assign w55955 = ~w11733 & pi00499;
assign w55956 = w11733 & ~pi00165;
assign w55957 = ~w11733 & pi00500;
assign w55958 = w11733 & ~pi00166;
assign w55959 = ~w11733 & pi00501;
assign w55960 = w11733 & ~pi00167;
assign w55961 = ~w11733 & pi00502;
assign w55962 = w11733 & ~pi00170;
assign w55963 = ~w11733 & pi00503;
assign w55964 = w11733 & ~pi00157;
assign w55965 = ~w11733 & pi00504;
assign w55966 = w11733 & ~pi00085;
assign w55967 = pi00541 & w11761;
assign w55968 = ~w11705 & pi00505;
assign w55969 = ~w11705 & pi00506;
assign w55970 = ~w11705 & pi00507;
assign w55971 = w11705 & ~pi00167;
assign w55972 = ~w11705 & pi00508;
assign w55973 = w11705 & ~pi00157;
assign w55974 = ~w11705 & pi00509;
assign w55975 = w11705 & ~pi00161;
assign w55976 = ~w11705 & pi00510;
assign w55977 = w11705 & ~pi00162;
assign w55978 = ~w11705 & pi00511;
assign w55979 = w11705 & ~pi00163;
assign w55980 = ~w11705 & pi00512;
assign w55981 = ~w11705 & pi00513;
assign w55982 = w11705 & ~pi00072;
assign w55983 = ~w11733 & pi00514;
assign w55984 = w11733 & ~pi00076;
assign w55985 = ~w11733 & pi00515;
assign w55986 = ~w11733 & pi00516;
assign w55987 = w11733 & ~pi00088;
assign w55988 = ~pi00541 & w11761;
assign w55989 = ~w11799 & pi00517;
assign w55990 = w11799 & ~pi00075;
assign w55991 = ~w11799 & pi00518;
assign w55992 = w11799 & ~pi00079;
assign w55993 = ~w11799 & pi00519;
assign w55994 = w11799 & ~pi00169;
assign w55995 = ~w11799 & pi00520;
assign w55996 = w11799 & ~pi00170;
assign w55997 = ~w11799 & pi00521;
assign w55998 = w11799 & ~pi00171;
assign w55999 = ~w11799 & pi00522;
assign w56000 = w11799 & ~pi00157;
assign w56001 = ~w11799 & pi00523;
assign w56002 = w11799 & ~pi00158;
assign w56003 = ~w11799 & pi00524;
assign w56004 = w11799 & ~pi00083;
assign w56005 = w11826 & pi00810;
assign w56006 = ~w11825 & pi00525;
assign w56007 = w11825 & ~pi00087;
assign w56008 = ~w11825 & pi00526;
assign w56009 = w11825 & ~pi00167;
assign w56010 = ~w11825 & pi00527;
assign w56011 = w11825 & ~pi00168;
assign w56012 = ~w11825 & pi00528;
assign w56013 = w11825 & ~pi00170;
assign w56014 = ~w11825 & pi00529;
assign w56015 = w11825 & ~pi00171;
assign w56016 = ~w11825 & pi00530;
assign w56017 = w11825 & ~pi00158;
assign w56018 = ~w11825 & pi00531;
assign w56019 = w11825 & ~pi00081;
assign w56020 = ~w11825 & pi00532;
assign w56021 = w11825 & ~pi00083;
assign w56022 = ~w11825 & pi00533;
assign w56023 = w11825 & ~pi00085;
assign w56024 = ~w11825 & pi00534;
assign w56025 = w11825 & ~pi00072;
assign w56026 = ~pi09821 & w671;
assign w56027 = ~pi01276 & w671;
assign w56028 = ~pi00006 & ~pi09964;
assign w56029 = w11874 & w406;
assign w56030 = w54828 & pi00828;
assign w56031 = w56030 & pi00826;
assign w56032 = w56031 & pi00829;
assign w56033 = w56032 & pi00830;
assign w56034 = w56033 & pi00840;
assign w56035 = ~w400 & w11895;
assign w56036 = ~pi00539 & ~w789;
assign w56037 = ~w11107 & pi00540;
assign w56038 = ~w11705 & pi00542;
assign w56039 = w11705 & ~pi00165;
assign w56040 = ~w11705 & pi00543;
assign w56041 = w11705 & ~pi00077;
assign w56042 = ~w11705 & pi00544;
assign w56043 = w11705 & ~pi00079;
assign w56044 = ~w11705 & pi00545;
assign w56045 = ~w11705 & pi00546;
assign w56046 = ~w11705 & pi00547;
assign w56047 = w11705 & ~pi00083;
assign w56048 = ~w11705 & pi00548;
assign w56049 = ~w11733 & pi00549;
assign w56050 = w11733 & ~pi00077;
assign w56051 = ~w11733 & pi00550;
assign w56052 = w11733 & ~pi00169;
assign w56053 = ~w11733 & pi00551;
assign w56054 = w11733 & ~pi00171;
assign w56055 = ~w11733 & pi00552;
assign w56056 = w11733 & ~pi00160;
assign w56057 = ~w11733 & pi00553;
assign w56058 = w11733 & ~pi00164;
assign w56059 = ~w11733 & pi00554;
assign w56060 = w11733 & ~pi00161;
assign w56061 = ~w11733 & pi00555;
assign w56062 = w11733 & ~pi00082;
assign w56063 = ~w11705 & pi00556;
assign w56064 = w11705 & ~pi00076;
assign w56065 = ~w11705 & pi00557;
assign w56066 = ~w11705 & pi00558;
assign w56067 = w11705 & ~pi00172;
assign w56068 = ~w11705 & pi00559;
assign w56069 = w11705 & ~pi00159;
assign w56070 = ~w11705 & pi00560;
assign w56071 = w11705 & ~pi00081;
assign w56072 = ~w11705 & pi00561;
assign w56073 = ~w11705 & pi00562;
assign w56074 = ~w11705 & pi00563;
assign w56075 = w11705 & ~pi00086;
assign w56076 = ~w11733 & pi00564;
assign w56077 = w11733 & ~pi00074;
assign w56078 = ~w11733 & pi00565;
assign w56079 = ~w11733 & pi00566;
assign w56080 = ~w11733 & pi00567;
assign w56081 = w11733 & ~pi00079;
assign w56082 = ~w11733 & pi00568;
assign w56083 = w11733 & ~pi00168;
assign w56084 = ~w11733 & pi00569;
assign w56085 = ~w11733 & pi00570;
assign w56086 = ~w11733 & pi00571;
assign w56087 = ~w11733 & pi00572;
assign w56088 = ~w11733 & pi00573;
assign w56089 = ~w11733 & pi00574;
assign w56090 = w11733 & ~pi00159;
assign w56091 = ~w11733 & pi00575;
assign w56092 = w11733 & ~pi00084;
assign w56093 = ~w11799 & pi00576;
assign w56094 = w11799 & ~pi00087;
assign w56095 = ~w11799 & pi00577;
assign w56096 = w11799 & ~pi00074;
assign w56097 = ~w11799 & pi00578;
assign w56098 = w11799 & ~pi00077;
assign w56099 = ~w11799 & pi00579;
assign w56100 = w11799 & ~pi00078;
assign w56101 = ~w11799 & pi00580;
assign w56102 = w11799 & ~pi00165;
assign w56103 = ~w11799 & pi00581;
assign w56104 = w11799 & ~pi00172;
assign w56105 = ~w11733 & pi00582;
assign w56106 = w11733 & ~pi00086;
assign w56107 = ~w11799 & pi00583;
assign w56108 = w11799 & ~pi00167;
assign w56109 = ~w11799 & pi00584;
assign w56110 = w11799 & ~pi00159;
assign w56111 = ~w11799 & pi00585;
assign w56112 = w11799 & ~pi00160;
assign w56113 = ~w11799 & pi00586;
assign w56114 = w11799 & ~pi00081;
assign w56115 = ~w11799 & pi00587;
assign w56116 = w11799 & ~pi00164;
assign w56117 = ~w11799 & pi00588;
assign w56118 = w11799 & ~pi00161;
assign w56119 = ~w11799 & pi00589;
assign w56120 = w11799 & ~pi00084;
assign w56121 = ~w11799 & pi00590;
assign w56122 = w11799 & ~pi00085;
assign w56123 = ~w11799 & pi00591;
assign w56124 = w11799 & ~pi00072;
assign w56125 = ~w11825 & pi00592;
assign w56126 = w11825 & ~pi00074;
assign w56127 = ~w11825 & pi00593;
assign w56128 = w11825 & ~pi00075;
assign w56129 = ~w11825 & pi00594;
assign w56130 = w11825 & ~pi00076;
assign w56131 = ~w11825 & pi00595;
assign w56132 = w11825 & ~pi00166;
assign w56133 = ~w11825 & pi00596;
assign w56134 = w11825 & ~pi00165;
assign w56135 = ~w11825 & pi00597;
assign w56136 = w11825 & ~pi00172;
assign w56137 = ~w11825 & pi00598;
assign w56138 = w11825 & ~pi00169;
assign w56139 = ~w11825 & pi00599;
assign w56140 = w11825 & ~pi00157;
assign w56141 = ~w11825 & pi00600;
assign w56142 = w11825 & ~pi00079;
assign w56143 = ~w11825 & pi00601;
assign w56144 = w11825 & ~pi00159;
assign w56145 = ~w11825 & pi00602;
assign w56146 = w11825 & ~pi00160;
assign w56147 = ~w11825 & pi00603;
assign w56148 = w11825 & ~pi00162;
assign w56149 = ~w11825 & pi00604;
assign w56150 = w11825 & ~pi00163;
assign w56151 = ~w11825 & pi00605;
assign w56152 = w11825 & ~pi00082;
assign w56153 = ~w11733 & pi00606;
assign w56154 = w11733 & ~pi00083;
assign w56155 = ~w11733 & pi00607;
assign w56156 = ~w11799 & pi00608;
assign w56157 = ~pi00036 & pi01480;
assign w56158 = ~w54871 & ~pi00064;
assign w56159 = w54871 & pi00064;
assign w56160 = w11194 & pi01171;
assign w56161 = ~w11194 & pi00611;
assign w56162 = w11194 & pi01172;
assign w56163 = ~w11194 & pi00612;
assign w56164 = w11194 & pi01173;
assign w56165 = ~w11194 & pi00613;
assign w56166 = w11194 & pi01174;
assign w56167 = ~w11194 & pi00614;
assign w56168 = w11194 & pi01175;
assign w56169 = ~w11194 & pi00615;
assign w56170 = w11194 & pi01176;
assign w56171 = ~w11194 & pi00616;
assign w56172 = w11194 & pi01177;
assign w56173 = ~w11194 & pi00617;
assign w56174 = w11194 & pi01178;
assign w56175 = ~w11194 & pi00618;
assign w56176 = w11194 & pi01179;
assign w56177 = ~w11194 & pi00619;
assign w56178 = w11194 & pi01180;
assign w56179 = ~w11194 & pi00620;
assign w56180 = w11194 & pi01181;
assign w56181 = ~w11194 & pi00621;
assign w56182 = w11194 & pi01182;
assign w56183 = ~w11194 & pi00622;
assign w56184 = w11194 & pi01183;
assign w56185 = ~w11194 & pi00623;
assign w56186 = w11194 & pi01184;
assign w56187 = ~w11194 & pi00624;
assign w56188 = w11194 & pi01185;
assign w56189 = ~w11194 & pi00625;
assign w56190 = w11194 & pi01186;
assign w56191 = ~w11194 & pi00626;
assign w56192 = w11194 & pi01187;
assign w56193 = ~w11194 & pi00627;
assign w56194 = w11194 & pi01188;
assign w56195 = ~w11194 & pi00628;
assign w56196 = w11194 & pi01189;
assign w56197 = ~w11194 & pi00629;
assign w56198 = w11194 & pi01190;
assign w56199 = ~w11194 & pi00630;
assign w56200 = w11194 & pi01191;
assign w56201 = ~w11194 & pi00631;
assign w56202 = w11194 & pi01192;
assign w56203 = ~w11194 & pi00632;
assign w56204 = w11194 & pi01193;
assign w56205 = ~w11194 & pi00633;
assign w56206 = w11194 & pi01194;
assign w56207 = ~w11194 & pi00634;
assign w56208 = w11194 & pi01195;
assign w56209 = ~w11194 & pi00635;
assign w56210 = w11194 & pi01197;
assign w56211 = ~w11194 & pi00636;
assign w56212 = w11194 & pi01199;
assign w56213 = ~w11194 & pi00637;
assign w56214 = w11194 & pi01198;
assign w56215 = ~w11194 & pi00638;
assign w56216 = w11194 & pi01201;
assign w56217 = ~w11194 & pi00639;
assign w56218 = w11194 & pi01200;
assign w56219 = ~w11194 & pi00640;
assign w56220 = w11194 & pi01202;
assign w56221 = ~w11194 & pi00641;
assign w56222 = w11194 & pi01196;
assign w56223 = ~w11194 & pi00642;
assign w56224 = ~w55891 & ~pi00643;
assign w56225 = w12219 & pi00087;
assign w56226 = ~w12219 & ~pi00644;
assign w56227 = w12219 & pi00074;
assign w56228 = ~w12219 & ~pi00645;
assign w56229 = w12219 & pi00075;
assign w56230 = ~w12219 & ~pi00646;
assign w56231 = w12219 & pi00080;
assign w56232 = ~w12219 & ~pi00647;
assign w56233 = w12219 & pi00076;
assign w56234 = ~w12219 & ~pi00648;
assign w56235 = w12219 & pi00077;
assign w56236 = ~w12219 & ~pi00649;
assign w56237 = w12219 & pi00078;
assign w56238 = ~w12219 & ~pi00650;
assign w56239 = w12219 & pi00165;
assign w56240 = ~w12219 & ~pi00651;
assign w56241 = w12219 & pi00166;
assign w56242 = ~w12219 & ~pi00652;
assign w56243 = w12219 & pi00172;
assign w56244 = ~w12219 & ~pi00653;
assign w56245 = w12219 & pi00167;
assign w56246 = ~w12219 & ~pi00654;
assign w56247 = w12219 & pi00079;
assign w56248 = ~w12219 & ~pi00655;
assign w56249 = w12219 & pi00168;
assign w56250 = ~w12219 & ~pi00656;
assign w56251 = w12219 & pi00169;
assign w56252 = ~w12219 & ~pi00657;
assign w56253 = w12219 & pi00170;
assign w56254 = ~w12219 & ~pi00658;
assign w56255 = w12219 & pi00171;
assign w56256 = ~w12219 & ~pi00659;
assign w56257 = w12219 & pi00157;
assign w56258 = ~w12219 & ~pi00660;
assign w56259 = w12219 & pi00158;
assign w56260 = ~w12219 & ~pi00661;
assign w56261 = w12219 & pi00159;
assign w56262 = ~w12219 & ~pi00662;
assign w56263 = w12219 & pi00160;
assign w56264 = ~w12219 & ~pi00663;
assign w56265 = w12219 & pi00161;
assign w56266 = ~w12219 & ~pi00664;
assign w56267 = w12219 & pi00162;
assign w56268 = ~w12219 & ~pi00665;
assign w56269 = w12219 & pi00081;
assign w56270 = ~w12219 & ~pi00666;
assign w56271 = w12219 & pi00163;
assign w56272 = ~w12219 & ~pi00667;
assign w56273 = w12219 & pi00164;
assign w56274 = ~w12219 & ~pi00668;
assign w56275 = w12219 & pi00088;
assign w56276 = ~w12219 & ~pi00669;
assign w56277 = w12219 & pi00082;
assign w56278 = ~w12219 & ~pi00670;
assign w56279 = w12219 & pi00083;
assign w56280 = ~w12219 & ~pi00671;
assign w56281 = w12219 & pi00084;
assign w56282 = ~w12219 & ~pi00672;
assign w56283 = w12219 & pi00085;
assign w56284 = ~w12219 & ~pi00673;
assign w56285 = w12219 & pi00086;
assign w56286 = ~w12219 & ~pi00674;
assign w56287 = w12219 & pi00072;
assign w56288 = ~w12219 & ~pi00675;
assign w56289 = ~w11705 & pi00676;
assign w56290 = w11705 & ~pi00087;
assign w56291 = ~w11705 & pi00677;
assign w56292 = w11705 & ~pi00075;
assign w56293 = ~w11705 & pi00678;
assign w56294 = ~w11705 & pi00679;
assign w56295 = w11705 & ~pi00078;
assign w56296 = ~w11705 & pi00680;
assign w56297 = ~w11705 & pi00681;
assign w56298 = ~w11705 & pi00682;
assign w56299 = ~w11705 & pi00683;
assign w56300 = w11705 & ~pi00170;
assign w56301 = ~w11705 & pi00684;
assign w56302 = w11705 & ~pi00158;
assign w56303 = ~w11705 & pi00685;
assign w56304 = ~w11705 & pi00686;
assign w56305 = ~w11705 & pi00687;
assign w56306 = ~w11705 & pi00688;
assign w56307 = ~w11705 & pi00689;
assign w56308 = ~w11705 & pi00690;
assign w56309 = ~w11733 & pi00691;
assign w56310 = w11733 & ~pi00087;
assign w56311 = ~w11733 & pi00692;
assign w56312 = ~w11733 & pi00693;
assign w56313 = ~w11733 & pi00694;
assign w56314 = ~w11733 & pi00695;
assign w56315 = ~w11733 & pi00696;
assign w56316 = w11733 & ~pi00172;
assign w56317 = ~w11733 & pi00697;
assign w56318 = ~w11733 & pi00698;
assign w56319 = ~w11733 & pi00699;
assign w56320 = ~w11733 & pi00700;
assign w56321 = ~w11733 & pi00701;
assign w56322 = ~w11733 & pi00702;
assign w56323 = w11733 & ~pi00072;
assign w56324 = ~w11799 & pi00703;
assign w56325 = ~w11799 & pi00704;
assign w56326 = w11799 & ~pi00168;
assign w56327 = ~w11799 & pi00705;
assign w56328 = ~w11799 & pi00706;
assign w56329 = ~w11799 & pi00707;
assign w56330 = ~w11799 & pi00708;
assign w56331 = ~w11799 & pi00709;
assign w56332 = ~w11799 & pi00710;
assign w56333 = w11799 & ~pi00162;
assign w56334 = ~w11799 & pi00711;
assign w56335 = w11799 & ~pi00082;
assign w56336 = ~w11799 & pi00712;
assign w56337 = ~w11799 & pi00713;
assign w56338 = ~w11799 & pi00714;
assign w56339 = ~w11799 & pi00715;
assign w56340 = ~w11799 & pi00716;
assign w56341 = w11799 & ~pi00076;
assign w56342 = ~w11799 & pi00717;
assign w56343 = ~w11799 & pi00718;
assign w56344 = ~w11799 & pi00719;
assign w56345 = ~w11799 & pi00720;
assign w56346 = ~w11799 & pi00721;
assign w56347 = ~w11799 & pi00722;
assign w56348 = ~w11825 & pi00723;
assign w56349 = ~w11825 & pi00724;
assign w56350 = ~w11825 & pi00725;
assign w56351 = w11825 & ~pi00077;
assign w56352 = ~w11825 & pi00726;
assign w56353 = ~w11825 & pi00727;
assign w56354 = ~w11825 & pi00728;
assign w56355 = ~w11825 & pi00729;
assign w56356 = ~w11825 & pi00730;
assign w56357 = ~w11825 & pi00731;
assign w56358 = ~w11825 & pi00732;
assign w56359 = ~w11825 & pi00733;
assign w56360 = ~w11825 & pi00734;
assign w56361 = ~w11825 & pi00735;
assign w56362 = w11825 & ~pi00086;
assign w56363 = ~w11705 & pi00736;
assign w56364 = ~w11705 & pi00737;
assign w56365 = ~w11825 & pi00738;
assign w56366 = ~w11705 & pi00739;
assign w56367 = ~w11705 & pi00740;
assign w56368 = ~w11705 & pi00741;
assign w56369 = w11705 & ~pi00169;
assign w56370 = ~w11705 & pi00742;
assign w56371 = ~w11705 & pi00743;
assign w56372 = ~w11705 & pi00744;
assign w56373 = ~w11733 & pi00745;
assign w56374 = ~w11705 & pi00746;
assign w56375 = w11705 & ~pi00166;
assign w56376 = ~w11733 & pi00747;
assign w56377 = ~w11733 & pi00748;
assign w56378 = ~w11733 & pi00749;
assign w56379 = ~w11733 & pi00750;
assign w56380 = ~w11733 & pi00751;
assign w56381 = ~w11733 & pi00752;
assign w56382 = ~w11733 & pi00753;
assign w56383 = ~w11733 & pi00754;
assign w56384 = ~w11733 & pi00755;
assign w56385 = w11733 & ~pi00158;
assign w56386 = ~w11733 & pi00756;
assign w56387 = ~w11733 & pi00757;
assign w56388 = ~w11733 & pi00758;
assign w56389 = w11733 & ~pi00162;
assign w56390 = ~w11733 & pi00759;
assign w56391 = w11733 & ~pi00081;
assign w56392 = ~w11733 & pi00760;
assign w56393 = w11733 & ~pi00163;
assign w56394 = ~w11733 & pi00761;
assign w56395 = ~w11733 & pi00762;
assign w56396 = ~w11733 & pi00763;
assign w56397 = ~w11733 & pi00764;
assign w56398 = ~w11733 & pi00765;
assign w56399 = ~w11733 & pi00766;
assign w56400 = ~w11733 & pi00767;
assign w56401 = ~w11799 & pi00768;
assign w56402 = ~w11799 & pi00769;
assign w56403 = ~w11799 & pi00770;
assign w56404 = ~w11799 & pi00771;
assign w56405 = ~w11799 & pi00772;
assign w56406 = w11799 & ~pi00166;
assign w56407 = ~w11799 & pi00773;
assign w56408 = ~w11799 & pi00774;
assign w56409 = ~w11799 & pi00775;
assign w56410 = ~w11799 & pi00776;
assign w56411 = ~w11799 & pi00777;
assign w56412 = ~w11799 & pi00778;
assign w56413 = ~w11799 & pi00779;
assign w56414 = ~w11799 & pi00780;
assign w56415 = ~w11799 & pi00781;
assign w56416 = ~w11799 & pi00782;
assign w56417 = ~w11799 & pi00783;
assign w56418 = w11799 & ~pi00163;
assign w56419 = ~w11799 & pi00784;
assign w56420 = w11799 & ~pi00088;
assign w56421 = ~w11799 & pi00785;
assign w56422 = ~w11799 & pi00786;
assign w56423 = ~w11799 & pi00787;
assign w56424 = ~w11799 & pi00788;
assign w56425 = ~w11825 & pi00789;
assign w56426 = ~w11825 & pi00790;
assign w56427 = ~w11825 & pi00791;
assign w56428 = w11825 & ~pi00080;
assign w56429 = ~w11825 & pi00792;
assign w56430 = ~w11825 & pi00793;
assign w56431 = ~w11825 & pi00794;
assign w56432 = ~w11825 & pi00795;
assign w56433 = ~w11825 & pi00796;
assign w56434 = ~w11825 & pi00797;
assign w56435 = ~w11825 & pi00798;
assign w56436 = ~w11825 & pi00799;
assign w56437 = ~w11799 & pi00800;
assign w56438 = ~w11825 & pi00801;
assign w56439 = ~w11825 & pi00802;
assign w56440 = ~w11825 & pi00803;
assign w56441 = w11825 & ~pi00164;
assign w56442 = ~w11825 & pi00804;
assign w56443 = w11825 & ~pi00088;
assign w56444 = ~w11825 & pi00805;
assign w56445 = w11825 & ~pi00084;
assign w56446 = ~w11825 & pi00806;
assign w56447 = ~w11825 & pi00807;
assign w56448 = pi00541 & pi00808;
assign w56449 = ~pi00541 & ~pi00808;
assign w56450 = ~w56448 & ~pi00809;
assign w56451 = w56448 & pi00809;
assign w56452 = ~w56451 & ~w11706;
assign w56453 = ~w12723 & ~pi00811;
assign w56454 = ~pi00036 & pi09932;
assign w56455 = ~pi10472 & ~pi00818;
assign w56456 = ~pi10472 & ~pi00819;
assign w56457 = ~pi10472 & ~pi00820;
assign w56458 = ~pi10472 & ~pi00821;
assign w56459 = ~pi10472 & ~pi00822;
assign w56460 = ~pi10472 & ~pi00823;
assign w56461 = ~w56030 & ~pi00826;
assign w56462 = ~w406 & ~pi00827;
assign w56463 = w406 & pi00827;
assign w56464 = ~w54828 & ~pi00828;
assign w56465 = ~w56031 & ~pi00829;
assign w56466 = ~w56032 & ~pi00830;
assign w56467 = ~pi00831 & ~pi00832;
assign w56468 = pi00831 & pi00832;
assign w56469 = ~w56468 & ~pi00833;
assign w56470 = w56468 & pi00833;
assign w56471 = ~w56470 & ~pi00834;
assign w56472 = w56468 & w11868;
assign w56473 = ~w56472 & ~pi00835;
assign w56474 = w56472 & pi00835;
assign w56475 = ~w56474 & ~pi00836;
assign w56476 = w56474 & pi00836;
assign w56477 = ~w56476 & ~pi00837;
assign w56478 = ~pi00838 & ~pi00839;
assign w56479 = ~w56033 & ~pi00840;
assign w56480 = ~pi00241 & ~w2599;
assign w56481 = ~w1320 & ~pi00842;
assign w56482 = w1320 & ~pi10591;
assign w56483 = ~w1320 & ~pi00843;
assign w56484 = w1320 & ~pi10592;
assign w56485 = pi10381 & ~pi10577;
assign w56486 = ~pi02665 & ~pi00857;
assign w56487 = pi00858 & pi00867;
assign w56488 = ~w56487 & pi02665;
assign w56489 = ~pi09969 & pi10418;
assign w56490 = w12846 & w12856;
assign w56491 = ~w12848 & pi00867;
assign w56492 = ~w56491 & ~pi00844;
assign w56493 = w56491 & pi00844;
assign w56494 = ~w12867 & pi00848;
assign w56495 = w12867 & pi00469;
assign w56496 = pi10527 & pi00132;
assign w56497 = ~w12876 & pi00481;
assign w56498 = pi09519 & pi10364;
assign w56499 = pi01207 & pi01311;
assign w56500 = w56499 & pi01215;
assign w56501 = w56500 & ~pi00850;
assign w56502 = w12876 & pi00850;
assign w56503 = w12894 & ~pi00867;
assign w56504 = pi00858 & ~pi00867;
assign w56505 = w56504 & pi09947;
assign w56506 = w56487 & pi09884;
assign w56507 = w12894 & pi00867;
assign w56508 = w12903 & pi00852;
assign w56509 = ~pi00867 & ~pi00858;
assign w56510 = ~pi09896 & ~pi00857;
assign w56511 = ~w12911 & ~w12913;
assign w56512 = pi00852 & w12845;
assign w56513 = w1259 & pi10596;
assign w56514 = w1259 & pi10593;
assign w56515 = w1259 & pi10595;
assign w56516 = w1259 & pi10594;
assign w56517 = w12847 & ~pi00857;
assign w56518 = ~w12847 & pi00857;
assign w56519 = pi00852 & pi00868;
assign w56520 = ~w56519 & ~pi00858;
assign w56521 = w56519 & pi00858;
assign w56522 = w12845 & pi00858;
assign w56523 = w12845 & ~w56520;
assign w56524 = ~w12867 & pi00859;
assign w56525 = w12867 & pi00455;
assign w56526 = ~w12867 & pi00860;
assign w56527 = w12867 & pi00468;
assign w56528 = ~w12867 & pi00861;
assign w56529 = w12867 & pi00466;
assign w56530 = ~w12867 & pi00862;
assign w56531 = w12867 & pi00467;
assign w56532 = ~w12867 & pi00863;
assign w56533 = w12867 & pi00456;
assign w56534 = ~w12867 & pi00864;
assign w56535 = w12867 & pi00485;
assign w56536 = ~w12867 & pi00865;
assign w56537 = w12867 & ~pi10589;
assign w56538 = w1485 & pi00869;
assign w56539 = w12848 & ~pi00867;
assign w56540 = ~w56519 & w12845;
assign w56541 = pi01209 & w12984;
assign w56542 = ~w1320 & pi00872;
assign w56543 = w1320 & ~pi10590;
assign w56544 = w1469 & pi00869;
assign w56545 = ~pi02810 & pi02812;
assign w56546 = w13029 & ~pi00686;
assign w56547 = w13032 & ~pi01094;
assign w56548 = pi02810 & pi02812;
assign w56549 = w13035 & ~pi01042;
assign w56550 = pi02810 & ~pi02812;
assign w56551 = w13038 & ~pi00897;
assign w56552 = w13038 & ~pi00560;
assign w56553 = w11706 & ~pi00666;
assign w56554 = w13038 & ~pi01073;
assign w56555 = w13035 & ~pi00983;
assign w56556 = w13035 & ~pi00802;
assign w56557 = w13029 & ~pi00721;
assign w56558 = w13029 & ~pi00531;
assign w56559 = w13035 & ~pi00922;
assign w56560 = w13029 & ~pi01024;
assign w56561 = w13038 & ~pi01144;
assign w56562 = w13032 & ~pi00759;
assign w56563 = w13032 & ~pi00586;
assign w56564 = w13029 & ~pi01014;
assign w56565 = w13029 & ~pi00717;
assign w56566 = w13032 & ~pi01112;
assign w56567 = w13035 & ~pi00549;
assign w56568 = w13029 & ~pi00989;
assign w56569 = w11706 & ~pi00649;
assign w56570 = w13029 & ~pi00888;
assign w56571 = w13035 & ~pi00918;
assign w56572 = w13035 & ~pi00793;
assign w56573 = w13035 & ~pi00543;
assign w56574 = w13038 & ~pi00725;
assign w56575 = w13038 & ~pi01121;
assign w56576 = w13038 & ~pi00557;
assign w56577 = w13032 & ~pi00578;
assign w56578 = w13032 & ~pi01084;
assign w56579 = w13038 & ~pi00770;
assign w56580 = w13029 & ~pi00987;
assign w56581 = w13038 & ~pi00892;
assign w56582 = w13035 & ~pi00489;
assign w56583 = w13029 & ~pi00715;
assign w56584 = w13038 & ~pi00564;
assign w56585 = w11706 & ~pi00645;
assign w56586 = w13038 & ~pi00738;
assign w56587 = w13032 & ~pi01081;
assign w56588 = w13029 & ~pi00592;
assign w56589 = w13032 & ~pi01111;
assign w56590 = w13035 & ~pi00790;
assign w56591 = w13035 & ~pi01001;
assign w56592 = w13035 & ~pi00703;
assign w56593 = w13029 & ~pi00692;
assign w56594 = w13038 & ~pi00505;
assign w56595 = w13032 & ~pi00577;
assign w56596 = w13035 & ~pi01003;
assign w56597 = w13038 & ~pi00773;
assign w56598 = w13032 & ~pi00749;
assign w56599 = w13035 & ~pi00976;
assign w56600 = w13029 & ~pi00681;
assign w56601 = w11706 & ~pi00653;
assign w56602 = w13029 & ~pi00597;
assign w56603 = w13032 & ~pi00739;
assign w56604 = w13035 & ~pi01149;
assign w56605 = w13029 & ~pi01051;
assign w56606 = w13038 & ~pi01069;
assign w56607 = w13035 & ~pi01037;
assign w56608 = w13038 & ~pi00558;
assign w56609 = w13032 & ~pi00581;
assign w56610 = w13029 & ~pi00696;
assign w56611 = w13038 & ~pi01123;
assign w56612 = ~w11825 & pi00887;
assign w56613 = w11825 & ~pi00161;
assign w56614 = ~w11825 & pi00888;
assign w56615 = ~w11825 & pi00889;
assign w56616 = ~w11825 & pi00890;
assign w56617 = ~w11825 & pi00891;
assign w56618 = ~w11799 & pi00892;
assign w56619 = ~w11799 & pi00893;
assign w56620 = ~w11799 & pi00894;
assign w56621 = ~w11705 & pi00895;
assign w56622 = ~w11733 & pi00896;
assign w56623 = ~w11733 & pi00897;
assign w56624 = ~w11733 & pi00898;
assign w56625 = ~w11705 & pi00899;
assign w56626 = w11705 & ~pi00084;
assign w56627 = ~w11733 & pi00900;
assign w56628 = ~w11705 & pi00901;
assign w56629 = ~w11705 & pi00902;
assign w56630 = ~w11705 & pi00903;
assign w56631 = ~w11705 & pi00904;
assign w56632 = ~w11705 & pi00905;
assign w56633 = w11705 & ~pi00171;
assign w56634 = ~w11705 & pi00906;
assign w56635 = ~w11825 & pi00907;
assign w56636 = ~w11825 & pi00908;
assign w56637 = ~w11825 & pi00909;
assign w56638 = ~w11799 & pi00910;
assign w56639 = ~w11799 & pi00911;
assign w56640 = ~w11799 & pi00912;
assign w56641 = ~w11799 & pi00913;
assign w56642 = ~w11799 & pi00914;
assign w56643 = ~w11799 & pi00915;
assign w56644 = w11799 & ~pi00086;
assign w56645 = ~w11733 & pi00916;
assign w56646 = ~w11799 & pi00917;
assign w56647 = ~w11799 & pi00918;
assign w56648 = ~w11733 & pi00919;
assign w56649 = ~w11733 & pi00920;
assign w56650 = ~w11733 & pi00921;
assign w56651 = ~w11733 & pi00922;
assign w56652 = ~w11733 & pi00923;
assign w56653 = ~w11705 & pi00924;
assign w56654 = ~w11705 & pi00925;
assign w56655 = ~w11705 & pi00926;
assign w56656 = ~w11705 & pi00927;
assign w56657 = ~w11705 & pi00928;
assign w56658 = pi00030 & ~pi00929;
assign w56659 = w13029 & ~pi00687;
assign w56660 = w13038 & ~pi01127;
assign w56661 = w13035 & ~pi00553;
assign w56662 = w13038 & ~pi01145;
assign w56663 = w13029 & ~pi01060;
assign w56664 = w11706 & ~pi00668;
assign w56665 = w13035 & ~pi00803;
assign w56666 = w13038 & ~pi00512;
assign w56667 = w13029 & ~pi01161;
assign w56668 = w13032 & ~pi00761;
assign w56669 = w13038 & ~pi00907;
assign w56670 = w13035 & ~pi01044;
assign w56671 = w13032 & ~pi00587;
assign w56672 = w13035 & ~pi00493;
assign w56673 = w13029 & ~pi00700;
assign w56674 = w13032 & ~pi01095;
assign w56675 = w13032 & ~pi01136;
assign w56676 = w13035 & ~pi00927;
assign w56677 = w13032 & ~pi00760;
assign w56678 = w13035 & ~pi00911;
assign w56679 = w13038 & ~pi00783;
assign w56680 = w11706 & ~pi00667;
assign w56681 = w13029 & ~pi00604;
assign w56682 = w13032 & ~pi00904;
assign w56683 = w13038 & ~pi01074;
assign w56684 = w13029 & ~pi01025;
assign w56685 = w13035 & ~pi01153;
assign w56686 = w13038 & ~pi01126;
assign w56687 = w13029 & ~pi00996;
assign w56688 = w13038 & ~pi00511;
assign w56689 = w13035 & ~pi01008;
assign w56690 = w13029 & ~pi01059;
assign w56691 = w13035 & ~pi00710;
assign w56692 = w13038 & ~pi01125;
assign w56693 = w13029 & ~pi01023;
assign w56694 = w13035 & ~pi01007;
assign w56695 = w13035 & ~pi00546;
assign w56696 = w11706 & ~pi00665;
assign w56697 = w13035 & ~pi00801;
assign w56698 = w13029 & ~pi00925;
assign w56699 = w13029 & ~pi00603;
assign w56700 = w13029 & ~pi00912;
assign w56701 = w13038 & ~pi01072;
assign w56702 = w13038 & ~pi00782;
assign w56703 = w13032 & ~pi01135;
assign w56704 = w13038 & ~pi00510;
assign w56705 = w13032 & ~pi01093;
assign w56706 = w13032 & ~pi00758;
assign w56707 = w13035 & ~pi00545;
assign w56708 = w13032 & ~pi00588;
assign w56709 = w13038 & ~pi00509;
assign w56710 = w13035 & ~pi00709;
assign w56711 = w13029 & ~pi01058;
assign w56712 = w11706 & ~pi00664;
assign w56713 = w13038 & ~pi00908;
assign w56714 = w13029 & ~pi01022;
assign w56715 = w13035 & ~pi00887;
assign w56716 = w13038 & ~pi00781;
assign w56717 = w13029 & ~pi01160;
assign w56718 = w13029 & ~pi00995;
assign w56719 = w13035 & ~pi00554;
assign w56720 = w13032 & ~pi01092;
assign w56721 = w13038 & ~pi00573;
assign w56722 = w13032 & ~pi00757;
assign w56723 = w13032 & ~pi01091;
assign w56724 = w13029 & ~pi00994;
assign w56725 = w13029 & ~pi00919;
assign w56726 = w13029 & ~pi01057;
assign w56727 = w13035 & ~pi00552;
assign w56728 = w11706 & ~pi00663;
assign w56729 = w13038 & ~pi00734;
assign w56730 = w13038 & ~pi01108;
assign w56731 = w13029 & ~pi00602;
assign w56732 = w13038 & ~pi00780;
assign w56733 = w13035 & ~pi01152;
assign w56734 = w13035 & ~pi00708;
assign w56735 = w13032 & ~pi01116;
assign w56736 = w13032 & ~pi00585;
assign w56737 = w13035 & ~pi00492;
assign w56738 = w13038 & ~pi01124;
assign w56739 = w13038 & ~pi00574;
assign w56740 = w13029 & ~pi00720;
assign w56741 = w13038 & ~pi00779;
assign w56742 = w13035 & ~pi01006;
assign w56743 = w13035 & ~pi00707;
assign w56744 = w11706 & ~pi00662;
assign w56745 = w13035 & ~pi00807;
assign w56746 = w13032 & ~pi01090;
assign w56747 = w13038 & ~pi00733;
assign w56748 = w13032 & ~pi00584;
assign w56749 = w13029 & ~pi00601;
assign w56750 = w13038 & ~pi00559;
assign w56751 = w13032 & ~pi00756;
assign w56752 = w13035 & ~pi00982;
assign w56753 = w13029 & ~pi00685;
assign w56754 = w13029 & ~pi01021;
assign w56755 = w13035 & ~pi00921;
assign w56756 = w13032 & ~pi00523;
assign w56757 = w13029 & ~pi01056;
assign w56758 = w13032 & ~pi00755;
assign w56759 = w13032 & ~pi01089;
assign w56760 = w11706 & ~pi00661;
assign w56761 = w13038 & ~pi00732;
assign w56762 = w13038 & ~pi00898;
assign w56763 = w13035 & ~pi00799;
assign w56764 = w13035 & ~pi00706;
assign w56765 = w13029 & ~pi00530;
assign w56766 = w13038 & ~pi00901;
assign w56767 = w13038 & ~pi00778;
assign w56768 = w13029 & ~pi00684;
assign w56769 = w13035 & ~pi00981;
assign w56770 = w13029 & ~pi01020;
assign w56771 = w13035 & ~pi00928;
assign w56772 = w13032 & ~pi00753;
assign w56773 = w13038 & ~pi01143;
assign w56774 = w13029 & ~pi00916;
assign w56775 = w13035 & ~pi00551;
assign w56776 = w11706 & ~pi00659;
assign w56777 = w13029 & ~pi00529;
assign w56778 = w13032 & ~pi00905;
assign w56779 = w13035 & ~pi01151;
assign w56780 = w13029 & ~pi01055;
assign w56781 = w13038 & ~pi00730;
assign w56782 = w13035 & ~pi01040;
assign w56783 = w13032 & ~pi00521;
assign w56784 = w13029 & ~pi00924;
assign w56785 = w13038 & ~pi01106;
assign w56786 = w13038 & ~pi00570;
assign w56787 = w13029 & ~pi00913;
assign w56788 = w13029 & ~pi00993;
assign w56789 = w13029 & ~pi01019;
assign w56790 = w13035 & ~pi00980;
assign w56791 = w13038 & ~pi00508;
assign w56792 = w11706 & ~pi00660;
assign w56793 = w13029 & ~pi00599;
assign w56794 = w13035 & ~pi00503;
assign w56795 = w13035 & ~pi00798;
assign w56796 = w13032 & ~pi01088;
assign w56797 = w13038 & ~pi00731;
assign w56798 = w13038 & ~pi00571;
assign w56799 = w13032 & ~pi00522;
assign w56800 = w13035 & ~pi01041;
assign w56801 = w13032 & ~pi00754;
assign w56802 = w13038 & ~pi00777;
assign w56803 = w13032 & ~pi01115;
assign w56804 = w13038 & ~pi01105;
assign w56805 = w13038 & ~pi00569;
assign w56806 = w13029 & ~pi01018;
assign w56807 = w13029 & ~pi00719;
assign w56808 = w11706 & ~pi00658;
assign w56809 = w13029 & ~pi00528;
assign w56810 = w13035 & ~pi01039;
assign w56811 = w13035 & ~pi01150;
assign w56812 = w13032 & ~pi00520;
assign w56813 = w13038 & ~pi00729;
assign w56814 = w13029 & ~pi00683;
assign w56815 = w13038 & ~pi00776;
assign w56816 = w13035 & ~pi00502;
assign w56817 = w13032 & ~pi01087;
assign w56818 = w13035 & ~pi00979;
assign w56819 = w13032 & ~pi00519;
assign w56820 = w13035 & ~pi00550;
assign w56821 = w13029 & ~pi00991;
assign w56822 = w13035 & ~pi00705;
assign w56823 = w13032 & ~pi00741;
assign w56824 = w11706 & ~pi00657;
assign w56825 = w13038 & ~pi00728;
assign w56826 = w13029 & ~pi01017;
assign w56827 = w13035 & ~pi00797;
assign w56828 = w13035 & ~pi00978;
assign w56829 = w13029 & ~pi00598;
assign w56830 = w13032 & ~pi00752;
assign w56831 = w13029 & ~pi01054;
assign w56832 = w13038 & ~pi01104;
assign w56833 = w13038 & ~pi00775;
assign w56834 = w13038 & ~pi00572;
assign w56835 = w13035 & ~pi00704;
assign w56836 = w13032 & ~pi01134;
assign w56837 = w13038 & ~pi00568;
assign w56838 = w13029 & ~pi00698;
assign w56839 = w13038 & ~pi01142;
assign w56840 = w11706 & ~pi00656;
assign w56841 = w13038 & ~pi00727;
assign w56842 = w13032 & ~pi01114;
assign w56843 = w13029 & ~pi00527;
assign w56844 = w13035 & ~pi00491;
assign w56845 = w13035 & ~pi00890;
assign w56846 = w13038 & ~pi01103;
assign w56847 = w13029 & ~pi00992;
assign w56848 = w13029 & ~pi00718;
assign w56849 = w13035 & ~pi01005;
assign w56850 = w13032 & ~pi00740;
assign w56851 = w13029 & ~pi01052;
assign w56852 = w13038 & ~pi00566;
assign w56853 = w13032 & ~pi01085;
assign w56854 = w13038 & ~pi01141;
assign w56855 = w13032 & ~pi00583;
assign w56856 = w11706 & ~pi00654;
assign w56857 = w13038 & ~pi01071;
assign w56858 = w13035 & ~pi00977;
assign w56859 = w13029 & ~pi00526;
assign w56860 = w13032 & ~pi00750;
assign w56861 = w13035 & ~pi00795;
assign w56862 = w13029 & ~pi00682;
assign w56863 = w13038 & ~pi00507;
assign w56864 = w13035 & ~pi01036;
assign w56865 = w13035 & ~pi00501;
assign w56866 = w13029 & ~pi01016;
assign w56867 = w13035 & ~pi01035;
assign w56868 = w13032 & ~pi00893;
assign w56869 = w13029 & ~pi00926;
assign w56870 = w13029 & ~pi00695;
assign w56871 = w13038 & ~pi00772;
assign w56872 = w11706 & ~pi00652;
assign w56873 = w13038 & ~pi01070;
assign w56874 = w13035 & ~pi00975;
assign w56875 = w13035 & ~pi01148;
assign w56876 = w13032 & ~pi00746;
assign w56877 = w13029 & ~pi00595;
assign w56878 = w13038 & ~pi01101;
assign w56879 = w13032 & ~pi00900;
assign w56880 = w13035 & ~pi00500;
assign w56881 = w13038 & ~pi00515;
assign w56882 = w13029 & ~pi01050;
assign w56883 = w13038 & ~pi00608;
assign w56884 = w13038 & ~pi01122;
assign w56885 = w13035 & ~pi01034;
assign w56886 = w13029 & ~pi01049;
assign w56887 = w13032 & ~pi00895;
assign w56888 = w11706 & ~pi00651;
assign w56889 = w13035 & ~pi00794;
assign w56890 = w13029 & ~pi00680;
assign w56891 = w13029 & ~pi00596;
assign w56892 = w13032 & ~pi00580;
assign w56893 = w13038 & ~pi00909;
assign w56894 = w13038 & ~pi01102;
assign w56895 = w13035 & ~pi00499;
assign w56896 = w13029 & ~pi00920;
assign w56897 = w13035 & ~pi00542;
assign w56898 = w13032 & ~pi00748;
assign w56899 = w13038 & ~pi00771;
assign w56900 = w13035 & ~pi00974;
assign w56901 = w13035 & ~pi01033;
assign w56902 = w13038 & ~pi00565;
assign w56903 = w13035 & ~pi00498;
assign w56904 = w11706 & ~pi00650;
assign w56905 = w13029 & ~pi01159;
assign w56906 = w13029 & ~pi00914;
assign w56907 = w13038 & ~pi01068;
assign w56908 = w13029 & ~pi01015;
assign w56909 = w13035 & ~pi01147;
assign w56910 = w13038 & ~pi00902;
assign w56911 = w13032 & ~pi00579;
assign w56912 = w13032 & ~pi01113;
assign w56913 = w13032 & ~pi00737;
assign w56914 = w13029 & ~pi00679;
assign w56915 = w13032 & ~pi01133;
assign w56916 = w13029 & ~pi00694;
assign w56917 = w13035 & ~pi00923;
assign w56918 = w13029 & ~pi00716;
assign w56919 = w13029 & ~pi00678;
assign w56920 = w11706 & ~pi00648;
assign w56921 = w13038 & ~pi00724;
assign w56922 = w13038 & ~pi00769;
assign w56923 = w13035 & ~pi00792;
assign w56924 = w13032 & ~pi01083;
assign w56925 = w13029 & ~pi00594;
assign w56926 = w13035 & ~pi00973;
assign w56927 = w13032 & ~pi00747;
assign w56928 = w13038 & ~pi00514;
assign w56929 = w13038 & ~pi00556;
assign w56930 = w13035 & ~pi00917;
assign w56931 = w13035 & ~pi00490;
assign w56932 = w13029 & ~pi00988;
assign w56933 = w13032 & ~pi00607;
assign w56934 = w13035 & ~pi00497;
assign w56935 = w13038 & ~pi01140;
assign w56936 = w11706 & ~pi00647;
assign w56937 = w13029 & ~pi01158;
assign w56938 = w13038 & ~pi00506;
assign w56939 = w13038 & ~pi01067;
assign w56940 = w13038 & ~pi00896;
assign w56941 = w13035 & ~pi00791;
assign w56942 = w13029 & ~pi00693;
assign w56943 = w13035 & ~pi01032;
assign w56944 = w13032 & ~pi01132;
assign w56945 = w13029 & ~pi01048;
assign w56946 = w13032 & ~pi01082;
assign w56947 = w13038 & ~pi00768;
assign w56948 = w13032 & ~pi00906;
assign w56949 = w13029 & ~pi00699;
assign w56950 = w13038 & ~pi01100;
assign w56951 = w13032 & ~pi00767;
assign w56952 = w11706 & ~pi00646;
assign w56953 = w13038 & ~pi00723;
assign w56954 = w13032 & ~pi00517;
assign w56955 = w13035 & ~pi00891;
assign w56956 = w13029 & ~pi01047;
assign w56957 = w13029 & ~pi00593;
assign w56958 = w13029 & ~pi00677;
assign w56959 = w13035 & ~pi01031;
assign w56960 = w13035 & ~pi00496;
assign w56961 = w13035 & ~pi00972;
assign w56962 = w13038 & ~pi01120;
assign w56963 = w13038 & ~pi01146;
assign w56964 = w13029 & ~pi00701;
assign w56965 = w13035 & ~pi00986;
assign w56966 = w13029 & ~pi01064;
assign w56967 = w13032 & ~pi00742;
assign w56968 = w11706 & ~pi00674;
assign w56969 = w13029 & ~pi01163;
assign w56970 = w13032 & ~pi01118;
assign w56971 = w13035 & ~pi00806;
assign w56972 = w13038 & ~pi00563;
assign w56973 = w13038 & ~pi00735;
assign w56974 = w13032 & ~pi01138;
assign w56975 = w13035 & ~pi01012;
assign w56976 = w13038 & ~pi00582;
assign w56977 = w13029 & ~pi00999;
assign w56978 = w13035 & ~pi00915;
assign w56979 = w13038 & ~pi00562;
assign w56980 = w13029 & ~pi01063;
assign w56981 = w13032 & ~pi00590;
assign w56982 = w13029 & ~pi00690;
assign w56983 = w13038 & ~pi00787;
assign w56984 = w11706 & ~pi00673;
assign w56985 = w13029 & ~pi00533;
assign w56986 = w13029 & ~pi01029;
assign w56987 = w13035 & ~pi01156;
assign w56988 = w13038 & ~pi01128;
assign w56989 = w13038 & ~pi01079;
assign w56990 = w13032 & ~pi00744;
assign w56991 = w13035 & ~pi00713;
assign w56992 = w13035 & ~pi00495;
assign w56993 = w13032 & ~pi00766;
assign w56994 = w13035 & ~pi00504;
assign w56995 = w13038 & ~pi00575;
assign w56996 = w13035 & ~pi00712;
assign w56997 = w13035 & ~pi00985;
assign w56998 = w13038 & ~pi00786;
assign w56999 = w13032 & ~pi01117;
assign w57000 = w11706 & ~pi00672;
assign w57001 = w13038 & ~pi01078;
assign w57002 = w13035 & ~pi01011;
assign w57003 = w13029 & ~pi00889;
assign w57004 = w13029 & ~pi00998;
assign w57005 = w13035 & ~pi00805;
assign w57006 = w13032 & ~pi01098;
assign w57007 = w13038 & ~pi00899;
assign w57008 = w13029 & ~pi01028;
assign w57009 = w13029 & ~pi00722;
assign w57010 = w13032 & ~pi00589;
assign w57011 = w13032 & ~pi00903;
assign w57012 = w13029 & ~pi00606;
assign w57013 = w13029 & ~pi00689;
assign w57014 = w13029 & ~pi01062;
assign w57015 = w13038 & ~pi00785;
assign w57016 = w11706 & ~pi00671;
assign w57017 = w13035 & ~pi01154;
assign w57018 = w13038 & ~pi01131;
assign w57019 = w13038 & ~pi01077;
assign w57020 = w13035 & ~pi01010;
assign w57021 = w13029 & ~pi00532;
assign w57022 = w13038 & ~pi01110;
assign w57023 = w13032 & ~pi00764;
assign w57024 = w13035 & ~pi01045;
assign w57025 = w13035 & ~pi00547;
assign w57026 = w13032 & ~pi00524;
assign w57027 = w13029 & ~pi00997;
assign w57028 = w13035 & ~pi00984;
assign w57029 = w13032 & ~pi00762;
assign w57030 = w13038 & ~pi00516;
assign w57031 = w13038 & ~pi00784;
assign w57032 = w11706 & ~pi00669;
assign w57033 = w13029 & ~pi01162;
assign w57034 = w13032 & ~pi01096;
assign w57035 = w13038 & ~pi01075;
assign w57036 = w13029 & ~pi01027;
assign w57037 = w13035 & ~pi00804;
assign w57038 = w13035 & ~pi01009;
assign w57039 = w13035 & ~pi01043;
assign w57040 = w13032 & ~pi00894;
assign w57041 = w13038 & ~pi01109;
assign w57042 = w13029 & ~pi01061;
assign w57043 = w13032 & ~pi01097;
assign w57044 = w13035 & ~pi00555;
assign w57045 = w13032 & ~pi01137;
assign w57046 = w13038 & ~pi01130;
assign w57047 = w13038 & ~pi00800;
assign w57048 = w11706 & ~pi00670;
assign w57049 = w13038 & ~pi01076;
assign w57050 = w13029 & ~pi01026;
assign w57051 = w13035 & ~pi01155;
assign w57052 = w13035 & ~pi00494;
assign w57053 = w13029 & ~pi00605;
assign w57054 = w13029 & ~pi00688;
assign w57055 = w13038 & ~pi00561;
assign w57056 = w13035 & ~pi00711;
assign w57057 = w13032 & ~pi00763;
assign w57058 = w13029 & ~pi00910;
assign w57059 = w13029 & ~pi00697;
assign w57060 = w13032 & ~pi01086;
assign w57061 = w13032 & ~pi00518;
assign w57062 = w13035 & ~pi01038;
assign w57063 = w13038 & ~pi01107;
assign w57064 = w11706 & ~pi00655;
assign w57065 = w13035 & ~pi00796;
assign w57066 = w13032 & ~pi00751;
assign w57067 = w13029 & ~pi00600;
assign w57068 = w13038 & ~pi00567;
assign w57069 = w13038 & ~pi00726;
assign w57070 = w13029 & ~pi00990;
assign w57071 = w13029 & ~pi01053;
assign w57072 = w13035 & ~pi01004;
assign w57073 = w13038 & ~pi00774;
assign w57074 = w13035 & ~pi00544;
assign w57075 = w13038 & ~pi01139;
assign w57076 = w13029 & ~pi01046;
assign w57077 = w13035 & ~pi00971;
assign w57078 = w13038 & ~pi01099;
assign w57079 = w13035 & ~pi01002;
assign w57080 = w11706 & ~pi00644;
assign w57081 = w13035 & ~pi00789;
assign w57082 = w13029 & ~pi00691;
assign w57083 = w13038 & ~pi01066;
assign w57084 = w13029 & ~pi00676;
assign w57085 = w13029 & ~pi00525;
assign w57086 = w13035 & ~pi01030;
assign w57087 = w13038 & ~pi01119;
assign w57088 = w13032 & ~pi00576;
assign w57089 = w13032 & ~pi00736;
assign w57090 = w13032 & ~pi00745;
assign w57091 = ~pi01205 & ~pi10231;
assign w57092 = w57091 & ~pi00962;
assign w57093 = w57092 & w14135;
assign w57094 = w14148 & pi01309;
assign w57095 = w14144 & pi00957;
assign w57096 = w13038 & ~pi01129;
assign w57097 = w13038 & ~pi00788;
assign w57098 = w13029 & ~pi00702;
assign w57099 = w11706 & ~pi00675;
assign w57100 = w13032 & ~pi00591;
assign w57101 = w13035 & ~pi00714;
assign w57102 = w13038 & ~pi00513;
assign w57103 = w13035 & ~pi01013;
assign w57104 = w13029 & ~pi01065;
assign w57105 = ~w14187 & ~pi09809;
assign w57106 = ~pi09860 & ~pi09805;
assign w57107 = w57106 & ~pi09861;
assign w57108 = w57107 & ~pi09862;
assign w57109 = pi09808 & pi09864;
assign w57110 = ~pi01205 & ~pi09864;
assign w57111 = ~pi01205 & ~w57109;
assign w57112 = ~w55860 & pi00959;
assign w57113 = ~pi00024 & ~pi00043;
assign w57114 = w14144 & ~pi00962;
assign w57115 = w445 & ~pi00963;
assign w57116 = w1259 & pi10592;
assign w57117 = w1259 & pi10590;
assign w57118 = w1259 & pi10591;
assign w57119 = w56487 & pi09893;
assign w57120 = pi00858 & pi09977;
assign w57121 = ~w14227 & ~w14238;
assign w57122 = pi02123 & pi00455;
assign w57123 = ~pi02123 & pi00968;
assign w57124 = pi02123 & pi00469;
assign w57125 = ~pi02123 & pi00969;
assign w57126 = w55593 & w2599;
assign w57127 = ~w57126 & ~pi00970;
assign w57128 = w57126 & w14259;
assign w57129 = ~w11705 & pi00971;
assign w57130 = ~w11705 & pi00972;
assign w57131 = ~w11705 & pi00973;
assign w57132 = ~w11705 & pi00974;
assign w57133 = ~w11705 & pi00975;
assign w57134 = ~w11705 & pi00976;
assign w57135 = ~w11705 & pi00977;
assign w57136 = ~w11705 & pi00978;
assign w57137 = ~w11705 & pi00979;
assign w57138 = ~w11705 & pi00980;
assign w57139 = ~w11705 & pi00981;
assign w57140 = ~w11705 & pi00982;
assign w57141 = ~w11705 & pi00983;
assign w57142 = ~w11705 & pi00984;
assign w57143 = w11705 & ~pi00088;
assign w57144 = ~w11705 & pi00985;
assign w57145 = ~w11705 & pi00986;
assign w57146 = ~w11705 & pi00987;
assign w57147 = ~w11705 & pi00988;
assign w57148 = ~w11705 & pi00989;
assign w57149 = ~w11705 & pi00990;
assign w57150 = ~w11705 & pi00991;
assign w57151 = ~w11705 & pi00992;
assign w57152 = ~w11705 & pi00993;
assign w57153 = ~w11705 & pi00994;
assign w57154 = ~w11705 & pi00995;
assign w57155 = ~w11705 & pi00996;
assign w57156 = ~w11705 & pi00997;
assign w57157 = ~w11705 & pi00998;
assign w57158 = ~w11705 & pi00999;
assign w57159 = ~w11705 & pi01000;
assign w57160 = ~w11733 & pi01001;
assign w57161 = ~w11733 & pi01002;
assign w57162 = ~w11733 & pi01003;
assign w57163 = ~w11733 & pi01004;
assign w57164 = ~w11733 & pi01005;
assign w57165 = ~w11733 & pi01006;
assign w57166 = ~w11733 & pi01007;
assign w57167 = ~w11733 & pi01008;
assign w57168 = ~w11733 & pi01009;
assign w57169 = ~w11733 & pi01010;
assign w57170 = ~w11733 & pi01011;
assign w57171 = ~w11733 & pi01012;
assign w57172 = ~w11733 & pi01013;
assign w57173 = ~w11733 & pi01014;
assign w57174 = ~w11733 & pi01015;
assign w57175 = ~w11733 & pi01016;
assign w57176 = ~w11733 & pi01017;
assign w57177 = ~w11733 & pi01018;
assign w57178 = ~w11733 & pi01019;
assign w57179 = ~w11733 & pi01020;
assign w57180 = ~w11733 & pi01021;
assign w57181 = ~w11733 & pi01022;
assign w57182 = ~w11733 & pi01023;
assign w57183 = ~w11733 & pi01024;
assign w57184 = ~w11733 & pi01025;
assign w57185 = ~w11733 & pi01026;
assign w57186 = ~w11733 & pi01027;
assign w57187 = ~w11733 & pi01028;
assign w57188 = ~w11733 & pi01029;
assign w57189 = ~w11799 & pi01030;
assign w57190 = ~w11799 & pi01031;
assign w57191 = ~w11799 & pi01032;
assign w57192 = w11799 & ~pi00080;
assign w57193 = ~w11799 & pi01033;
assign w57194 = ~w11799 & pi01034;
assign w57195 = ~w11799 & pi01035;
assign w57196 = ~w11799 & pi01036;
assign w57197 = ~w11799 & pi01037;
assign w57198 = ~w11799 & pi01038;
assign w57199 = ~w11799 & pi01039;
assign w57200 = ~w11799 & pi01040;
assign w57201 = ~w11799 & pi01041;
assign w57202 = ~w11799 & pi01042;
assign w57203 = ~w11799 & pi01043;
assign w57204 = ~w11799 & pi01044;
assign w57205 = ~w11799 & pi01045;
assign w57206 = ~w11799 & pi01046;
assign w57207 = ~w11799 & pi01047;
assign w57208 = ~w11799 & pi01048;
assign w57209 = ~w11799 & pi01049;
assign w57210 = ~w11799 & pi01050;
assign w57211 = ~w11799 & pi01051;
assign w57212 = ~w11799 & pi01052;
assign w57213 = ~w11799 & pi01053;
assign w57214 = ~w11799 & pi01054;
assign w57215 = ~w11799 & pi01055;
assign w57216 = ~w11799 & pi01056;
assign w57217 = ~w11799 & pi01057;
assign w57218 = ~w11799 & pi01058;
assign w57219 = ~w11799 & pi01059;
assign w57220 = ~w11799 & pi01060;
assign w57221 = ~w11799 & pi01061;
assign w57222 = ~w11799 & pi01062;
assign w57223 = ~w11799 & pi01063;
assign w57224 = ~w11799 & pi01064;
assign w57225 = ~w11799 & pi01065;
assign w57226 = ~w11825 & pi01066;
assign w57227 = ~w11825 & pi01067;
assign w57228 = ~w11825 & pi01068;
assign w57229 = w11825 & ~pi00078;
assign w57230 = ~w11825 & pi01069;
assign w57231 = ~w11825 & pi01070;
assign w57232 = ~w11825 & pi01071;
assign w57233 = ~w11825 & pi01072;
assign w57234 = ~w11825 & pi01073;
assign w57235 = ~w11825 & pi01074;
assign w57236 = ~w11825 & pi01075;
assign w57237 = ~w11825 & pi01076;
assign w57238 = ~w11825 & pi01077;
assign w57239 = ~w11825 & pi01078;
assign w57240 = ~w11825 & pi01079;
assign w57241 = ~w11825 & pi01080;
assign w57242 = ~w11705 & pi01081;
assign w57243 = ~w11705 & pi01082;
assign w57244 = ~w11705 & pi01083;
assign w57245 = ~w11705 & pi01084;
assign w57246 = ~w11705 & pi01085;
assign w57247 = ~w11705 & pi01086;
assign w57248 = ~w11705 & pi01087;
assign w57249 = ~w11705 & pi01088;
assign w57250 = ~w11705 & pi01089;
assign w57251 = ~w11705 & pi01090;
assign w57252 = ~w11705 & pi01091;
assign w57253 = ~w11705 & pi01092;
assign w57254 = ~w11705 & pi01093;
assign w57255 = ~w11705 & pi01094;
assign w57256 = ~w11705 & pi01095;
assign w57257 = ~w11705 & pi01096;
assign w57258 = ~w11705 & pi01097;
assign w57259 = ~w11705 & pi01098;
assign w57260 = ~w11705 & pi01099;
assign w57261 = ~w11705 & pi01100;
assign w57262 = ~w11705 & pi01101;
assign w57263 = ~w11705 & pi01102;
assign w57264 = ~w11705 & pi01103;
assign w57265 = ~w11705 & pi01104;
assign w57266 = ~w11705 & pi01105;
assign w57267 = ~w11705 & pi01106;
assign w57268 = ~w11705 & pi01107;
assign w57269 = ~w11705 & pi01108;
assign w57270 = ~w11705 & pi01109;
assign w57271 = ~w11705 & pi01110;
assign w57272 = ~w11733 & pi01111;
assign w57273 = ~w11733 & pi01112;
assign w57274 = ~w11733 & pi01113;
assign w57275 = ~w11733 & pi01114;
assign w57276 = ~w11733 & pi01115;
assign w57277 = ~w11733 & pi01116;
assign w57278 = ~w11733 & pi01117;
assign w57279 = ~w11733 & pi01118;
assign w57280 = ~w11733 & pi01119;
assign w57281 = ~w11733 & pi01120;
assign w57282 = ~w11733 & pi01121;
assign w57283 = ~w11733 & pi01122;
assign w57284 = ~w11733 & pi01123;
assign w57285 = ~w11733 & pi01124;
assign w57286 = ~w11733 & pi01125;
assign w57287 = ~w11733 & pi01126;
assign w57288 = ~w11733 & pi01127;
assign w57289 = ~w11733 & pi01128;
assign w57290 = ~w11733 & pi01129;
assign w57291 = ~w11733 & pi01130;
assign w57292 = ~w11733 & pi01131;
assign w57293 = ~w11799 & pi01132;
assign w57294 = ~w11799 & pi01133;
assign w57295 = ~w11799 & pi01134;
assign w57296 = ~w11799 & pi01135;
assign w57297 = ~w11799 & pi01136;
assign w57298 = ~w11799 & pi01137;
assign w57299 = ~w11799 & pi01138;
assign w57300 = ~w11799 & pi01139;
assign w57301 = ~w11799 & pi01140;
assign w57302 = ~w11799 & pi01141;
assign w57303 = ~w11799 & pi01142;
assign w57304 = ~w11799 & pi01143;
assign w57305 = ~w11799 & pi01144;
assign w57306 = ~w11799 & pi01145;
assign w57307 = ~w11799 & pi01146;
assign w57308 = ~w11825 & pi01147;
assign w57309 = ~w11825 & pi01148;
assign w57310 = ~w11825 & pi01149;
assign w57311 = ~w11825 & pi01150;
assign w57312 = ~w11825 & pi01151;
assign w57313 = ~w11825 & pi01152;
assign w57314 = ~w11825 & pi01153;
assign w57315 = ~w11825 & pi01154;
assign w57316 = ~w11825 & pi01155;
assign w57317 = ~w11825 & pi01156;
assign w57318 = ~w11825 & pi01157;
assign w57319 = ~w11825 & pi01158;
assign w57320 = ~w11825 & pi01159;
assign w57321 = ~w11825 & pi01160;
assign w57322 = ~w11825 & pi01161;
assign w57323 = ~w11825 & pi01162;
assign w57324 = ~w11825 & pi01163;
assign w57325 = pi01274 & w1192;
assign w57326 = ~pi01209 & w1789;
assign w57327 = ~pi01451 & w14862;
assign w57328 = ~w14861 & pi01169;
assign w57329 = w14861 & ~pi10647;
assign w57330 = ~w506 & pi01170;
assign w57331 = ~w12993 & ~pi02670;
assign w57332 = w14877 & ~pi01427;
assign w57333 = ~w12993 & ~pi02668;
assign w57334 = w14877 & ~pi10049;
assign w57335 = ~w12993 & ~pi01336;
assign w57336 = w14877 & ~pi01281;
assign w57337 = ~w12993 & ~pi02669;
assign w57338 = w14877 & ~pi01429;
assign w57339 = ~w12993 & ~pi01337;
assign w57340 = w14877 & ~pi01428;
assign w57341 = ~w12993 & ~pi01338;
assign w57342 = w14877 & ~pi10194;
assign w57343 = ~w12993 & ~pi02671;
assign w57344 = w14877 & ~pi01430;
assign w57345 = ~w12993 & ~pi01339;
assign w57346 = w14877 & ~pi10195;
assign w57347 = ~w12993 & ~pi01340;
assign w57348 = w14877 & ~pi01431;
assign w57349 = ~w12993 & ~pi02256;
assign w57350 = w14877 & ~pi01432;
assign w57351 = ~w12993 & ~pi02673;
assign w57352 = w14877 & ~pi01434;
assign w57353 = ~w12993 & ~pi02672;
assign w57354 = w14877 & ~pi01433;
assign w57355 = ~w12993 & ~pi02253;
assign w57356 = w14877 & ~pi10196;
assign w57357 = ~w12993 & ~pi01341;
assign w57358 = w14877 & ~pi10153;
assign w57359 = ~w12993 & ~pi01342;
assign w57360 = w14877 & ~pi10197;
assign w57361 = ~w12993 & ~pi02674;
assign w57362 = w14877 & ~pi10198;
assign w57363 = ~w12993 & ~pi01343;
assign w57364 = w14877 & ~pi10199;
assign w57365 = ~w12993 & ~pi02675;
assign w57366 = w14877 & ~pi02193;
assign w57367 = ~w12993 & ~pi01344;
assign w57368 = w14877 & ~pi10051;
assign w57369 = ~w12993 & ~pi01345;
assign w57370 = w14877 & ~pi10200;
assign w57371 = ~w12993 & ~pi02676;
assign w57372 = w14877 & ~pi10201;
assign w57373 = ~w12993 & ~pi02250;
assign w57374 = w14877 & ~pi10202;
assign w57375 = ~w12993 & ~pi02677;
assign w57376 = w14877 & ~pi01435;
assign w57377 = ~w12993 & ~pi02678;
assign w57378 = w14877 & ~pi01436;
assign w57379 = ~w12993 & ~pi02246;
assign w57380 = w14877 & ~pi01437;
assign w57381 = ~w12993 & ~pi01346;
assign w57382 = w14877 & ~pi02191;
assign w57383 = ~w12993 & ~pi02680;
assign w57384 = w14877 & ~pi02692;
assign w57385 = ~w12993 & ~pi02679;
assign w57386 = w14877 & ~pi01438;
assign w57387 = ~w12993 & ~pi01347;
assign w57388 = w14877 & ~pi02189;
assign w57389 = ~w12993 & ~pi02238;
assign w57390 = w14877 & ~pi10052;
assign w57391 = ~w12993 & ~pi02682;
assign w57392 = w14877 & ~pi01439;
assign w57393 = ~w12993 & ~pi02681;
assign w57394 = ~w57107 & pi09862;
assign w57395 = pi02648 & pi01206;
assign w57396 = ~w57106 & pi09861;
assign w57397 = ~w12876 & pi00478;
assign w57398 = w1789 & w15945;
assign w57399 = ~w12984 & pi01209;
assign w57400 = pi01209 & w12993;
assign w57401 = ~w57091 & ~pi01210;
assign w57402 = w14148 & w11345;
assign w57403 = ~w57091 & ~pi01211;
assign w57404 = w57091 & pi00962;
assign w57405 = w57404 & w15959;
assign w57406 = pi01308 & w15964;
assign w57407 = ~w57404 & ~pi01213;
assign w57408 = w57091 & pi01213;
assign w57409 = pi01204 & pi01214;
assign w57410 = ~w12876 & pi00479;
assign w57411 = w12876 & pi01215;
assign w57412 = w1789 & w15944;
assign w57413 = ~w1789 & w12985;
assign w57414 = pi01262 & ~w12984;
assign w57415 = ~w15949 & ~pi01217;
assign w57416 = ~pi01451 & w16004;
assign w57417 = ~w16003 & pi01218;
assign w57418 = w16003 & ~pi10649;
assign w57419 = ~w16003 & pi01219;
assign w57420 = w16003 & ~pi10651;
assign w57421 = ~w16013 & pi01220;
assign w57422 = w16013 & ~pi10634;
assign w57423 = ~w16013 & pi01221;
assign w57424 = w16013 & ~pi10636;
assign w57425 = ~w16013 & pi01222;
assign w57426 = w16013 & ~pi10640;
assign w57427 = ~w16013 & pi01223;
assign w57428 = w16013 & ~pi10647;
assign w57429 = ~w16013 & pi01224;
assign w57430 = w16013 & ~pi10625;
assign w57431 = pi01451 & w14862;
assign w57432 = ~w16003 & pi01225;
assign w57433 = w16003 & ~pi10633;
assign w57434 = ~w16003 & pi01226;
assign w57435 = w16003 & ~pi10632;
assign w57436 = ~w16003 & pi01227;
assign w57437 = w16003 & ~pi10635;
assign w57438 = ~w16003 & pi01228;
assign w57439 = w16003 & ~pi10640;
assign w57440 = ~w16003 & pi01229;
assign w57441 = w16003 & ~pi10653;
assign w57442 = ~w16003 & pi01230;
assign w57443 = w16003 & ~pi10627;
assign w57444 = ~w16003 & pi01231;
assign w57445 = w16003 & ~pi10630;
assign w57446 = ~w16013 & pi01232;
assign w57447 = w16013 & ~pi10641;
assign w57448 = ~w16013 & pi01233;
assign w57449 = w16013 & ~pi10646;
assign w57450 = ~w16013 & pi01234;
assign w57451 = w16013 & ~pi10648;
assign w57452 = ~w16013 & pi01235;
assign w57453 = w16013 & ~pi10630;
assign w57454 = ~w14861 & pi01236;
assign w57455 = w14861 & ~pi10634;
assign w57456 = ~w14861 & pi01237;
assign w57457 = w14861 & ~pi10636;
assign w57458 = ~w14861 & pi01238;
assign w57459 = w14861 & ~pi10638;
assign w57460 = ~w14861 & pi01239;
assign w57461 = w14861 & ~pi10623;
assign w57462 = ~w14861 & pi01240;
assign w57463 = w14861 & ~pi10642;
assign w57464 = ~w14861 & pi01241;
assign w57465 = w14861 & ~pi10645;
assign w57466 = ~w14861 & pi01242;
assign w57467 = w14861 & ~pi10649;
assign w57468 = ~w14861 & pi01243;
assign w57469 = w14861 & ~pi10650;
assign w57470 = ~w14861 & pi01244;
assign w57471 = w14861 & ~pi10652;
assign w57472 = ~w14861 & pi01245;
assign w57473 = w14861 & ~pi10627;
assign w57474 = ~w14861 & pi01246;
assign w57475 = w14861 & ~pi10628;
assign w57476 = ~w14861 & pi01247;
assign w57477 = w14861 & ~pi10625;
assign w57478 = ~w14861 & pi01248;
assign w57479 = w14861 & ~pi10630;
assign w57480 = ~w55862 & ~pi01249;
assign w57481 = ~w1313 & pi01251;
assign w57482 = w1313 & pi10590;
assign w57483 = ~w1313 & pi01252;
assign w57484 = w1313 & pi10591;
assign w57485 = ~w1313 & pi01253;
assign w57486 = w1313 & pi10592;
assign w57487 = ~w1281 & pi01254;
assign w57488 = w1281 & pi10591;
assign w57489 = ~w1281 & pi01255;
assign w57490 = w1281 & pi10592;
assign w57491 = ~w1281 & pi01256;
assign w57492 = w1281 & pi10593;
assign w57493 = ~w1281 & pi01257;
assign w57494 = w1281 & pi10594;
assign w57495 = ~w1281 & pi01258;
assign w57496 = w1281 & pi10595;
assign w57497 = ~w1281 & pi01259;
assign w57498 = w1281 & pi10596;
assign w57499 = ~w1281 & pi01260;
assign w57500 = w1281 & pi10590;
assign w57501 = w55892 & pi10666;
assign w57502 = ~w1232 & ~pi01261;
assign w57503 = w1232 & ~pi10606;
assign w57504 = ~pi01262 & w12993;
assign w57505 = ~w1279 & pi01263;
assign w57506 = w1279 & pi10590;
assign w57507 = ~w1279 & pi01264;
assign w57508 = w1279 & pi10591;
assign w57509 = ~w1279 & pi01265;
assign w57510 = w1279 & pi10592;
assign w57511 = ~w1279 & pi01266;
assign w57512 = w1279 & pi10593;
assign w57513 = ~w1279 & pi01267;
assign w57514 = w1279 & pi10594;
assign w57515 = ~w1279 & pi01268;
assign w57516 = w1279 & pi10595;
assign w57517 = ~w1279 & pi01269;
assign w57518 = w1279 & pi10596;
assign w57519 = pi00845 & pi00177;
assign w57520 = ~pi00845 & pi01270;
assign w57521 = ~pi00845 & pi01271;
assign w57522 = ~pi01271 & w16172;
assign w57523 = ~w1192 & ~w16192;
assign w57524 = w1192 & ~w10686;
assign w57525 = ~pi01454 & ~w15985;
assign w57526 = w16198 & ~pi01274;
assign w57527 = ~w16198 & pi01274;
assign w57528 = ~w57091 & pi01275;
assign w57529 = w57404 & w16204;
assign w57530 = ~w139 & w12833;
assign w57531 = ~w1268 & pi01278;
assign w57532 = w1268 & pi10595;
assign w57533 = pi01451 & w16004;
assign w57534 = ~w16003 & pi01279;
assign w57535 = ~w16218 & pi01280;
assign w57536 = w16218 & ~pi10623;
assign w57537 = pi01451 & pi09825;
assign w57538 = w57537 & pi09856;
assign w57539 = w57538 & w14862;
assign w57540 = ~w16013 & pi01282;
assign w57541 = w16013 & ~pi10642;
assign w57542 = ~w16003 & pi01283;
assign w57543 = w16003 & ~pi10644;
assign w57544 = ~w16218 & pi01284;
assign w57545 = w16218 & ~pi10630;
assign w57546 = ~w16218 & pi01285;
assign w57547 = w16218 & ~pi10639;
assign w57548 = ~w14861 & pi01286;
assign w57549 = ~w14861 & pi01287;
assign w57550 = w14861 & ~pi10624;
assign w57551 = ~w14861 & pi01288;
assign w57552 = ~w14861 & pi01289;
assign w57553 = w14861 & ~pi10622;
assign w57554 = ~w14861 & pi01290;
assign w57555 = w14861 & ~pi10648;
assign w57556 = ~w16013 & pi01291;
assign w57557 = w16013 & ~pi10624;
assign w57558 = ~w16013 & pi01292;
assign w57559 = w16013 & ~pi10643;
assign w57560 = ~w16003 & pi01293;
assign w57561 = w16003 & ~pi10625;
assign w57562 = ~w16218 & pi01294;
assign w57563 = w16218 & ~pi10652;
assign w57564 = ~w16218 & pi01295;
assign w57565 = w16218 & ~pi10635;
assign w57566 = ~w14861 & pi01296;
assign w57567 = w14861 & ~pi10640;
assign w57568 = ~w14861 & pi01297;
assign w57569 = w14861 & ~pi10629;
assign w57570 = ~w14861 & pi01298;
assign w57571 = w14861 & ~pi10633;
assign w57572 = ~w16003 & pi01299;
assign w57573 = ~w16013 & pi01300;
assign w57574 = w16013 & ~pi10623;
assign w57575 = ~w16003 & pi01301;
assign w57576 = w16003 & ~pi10647;
assign w57577 = ~w16013 & pi01302;
assign w57578 = w16013 & ~pi10652;
assign w57579 = w16299 & pi01303;
assign w57580 = ~w16299 & w16301;
assign w57581 = ~w12876 & pi00482;
assign w57582 = ~pi10374 & ~pi01304;
assign w57583 = w14137 & pi01307;
assign w57584 = ~pi00962 & ~pi01305;
assign w57585 = ~w57092 & pi01306;
assign w57586 = ~pi01308 & ~pi01307;
assign w57587 = w11356 & pi09863;
assign w57588 = w14137 & pi01309;
assign w57589 = ~w57091 & pi01310;
assign w57590 = ~w12876 & pi00480;
assign w57591 = w12876 & pi01311;
assign w57592 = w16333 & ~pi01312;
assign w57593 = ~w16333 & pi01312;
assign w57594 = ~w16003 & pi01313;
assign w57595 = w16003 & ~pi10636;
assign w57596 = ~w16003 & pi01314;
assign w57597 = ~w16003 & pi01315;
assign w57598 = ~w16013 & pi01316;
assign w57599 = w16013 & ~pi10644;
assign w57600 = ~w16013 & pi01317;
assign w57601 = w16013 & ~pi10649;
assign w57602 = ~w16013 & pi01318;
assign w57603 = w16013 & ~pi10650;
assign w57604 = ~w16013 & pi01319;
assign w57605 = w16013 & ~pi10628;
assign w57606 = ~w16003 & pi01320;
assign w57607 = w16003 & ~pi10641;
assign w57608 = ~w16003 & pi01321;
assign w57609 = w16003 & ~pi10626;
assign w57610 = ~w16013 & pi01322;
assign w57611 = ~w16013 & pi01323;
assign w57612 = w16013 & ~pi10633;
assign w57613 = ~w16013 & pi01324;
assign w57614 = ~w16013 & pi01325;
assign w57615 = w16013 & ~pi10645;
assign w57616 = ~w16013 & pi01326;
assign w57617 = ~w16013 & pi01327;
assign w57618 = ~w14861 & pi01328;
assign w57619 = w14861 & ~pi10626;
assign w57620 = ~w16218 & pi01329;
assign w57621 = w16218 & ~pi10634;
assign w57622 = ~w16218 & pi01330;
assign w57623 = w16218 & ~pi10636;
assign w57624 = ~w16218 & pi01331;
assign w57625 = w16218 & ~pi10642;
assign w57626 = ~w16218 & pi01332;
assign w57627 = w16218 & ~pi10648;
assign w57628 = ~w16218 & pi01333;
assign w57629 = w16218 & ~pi10647;
assign w57630 = ~w16218 & pi01334;
assign w57631 = w16218 & ~pi10627;
assign w57632 = ~w16218 & pi01335;
assign w57633 = ~w16218 & ~w16407;
assign w57634 = ~pi01336 & ~w16407;
assign w57635 = ~pi01336 & w57633;
assign w57636 = pi10635 & w16407;
assign w57637 = pi10635 & ~w57633;
assign w57638 = ~pi01337 & ~w16407;
assign w57639 = ~pi01337 & w57633;
assign w57640 = pi10636 & w16407;
assign w57641 = pi10636 & ~w57633;
assign w57642 = ~pi01338 & ~w16407;
assign w57643 = ~pi01338 & w57633;
assign w57644 = pi10638 & w16407;
assign w57645 = pi10638 & ~w57633;
assign w57646 = ~pi01339 & ~w16407;
assign w57647 = ~pi01339 & w57633;
assign w57648 = pi10639 & w16407;
assign w57649 = pi10639 & ~w57633;
assign w57650 = ~pi01340 & ~w16407;
assign w57651 = ~pi01340 & w57633;
assign w57652 = pi10643 & w16407;
assign w57653 = pi10643 & ~w57633;
assign w57654 = ~pi01341 & ~w16407;
assign w57655 = ~pi01341 & w57633;
assign w57656 = pi10644 & w16407;
assign w57657 = pi10644 & ~w57633;
assign w57658 = ~pi01342 & ~w16407;
assign w57659 = ~pi01342 & w57633;
assign w57660 = pi10646 & w16407;
assign w57661 = pi10646 & ~w57633;
assign w57662 = ~pi01343 & ~w16407;
assign w57663 = ~pi01343 & w57633;
assign w57664 = pi10648 & w16407;
assign w57665 = pi10648 & ~w57633;
assign w57666 = ~pi01344 & ~w16407;
assign w57667 = ~pi01344 & w57633;
assign w57668 = pi10649 & w16407;
assign w57669 = pi10649 & ~w57633;
assign w57670 = ~pi01345 & ~w16407;
assign w57671 = ~pi01345 & w57633;
assign w57672 = pi10625 & w16407;
assign w57673 = pi10625 & ~w57633;
assign w57674 = ~pi01346 & ~w16407;
assign w57675 = ~pi01346 & w57633;
assign w57676 = pi10628 & w16407;
assign w57677 = pi10628 & ~w57633;
assign w57678 = ~pi01347 & ~w16407;
assign w57679 = ~pi01347 & w57633;
assign w57680 = ~w16003 & pi01348;
assign w57681 = ~w16003 & pi01349;
assign w57682 = ~w16003 & pi01350;
assign w57683 = w16003 & ~pi10637;
assign w57684 = ~w16003 & pi01351;
assign w57685 = w16003 & ~pi10638;
assign w57686 = ~w16003 & pi01352;
assign w57687 = w16003 & ~pi10639;
assign w57688 = ~w16003 & pi01353;
assign w57689 = ~w16003 & pi01354;
assign w57690 = w16003 & ~pi10645;
assign w57691 = ~w16003 & pi01355;
assign w57692 = w16003 & ~pi10624;
assign w57693 = ~w16003 & pi01356;
assign w57694 = ~w16003 & pi01357;
assign w57695 = w16003 & ~pi10629;
assign w57696 = ~w16003 & pi01358;
assign w57697 = w16003 & ~pi10631;
assign w57698 = ~w16013 & pi01359;
assign w57699 = w16013 & ~pi10622;
assign w57700 = ~w16013 & pi01360;
assign w57701 = ~w16013 & pi01361;
assign w57702 = ~w16013 & pi01362;
assign w57703 = w16013 & ~pi10637;
assign w57704 = ~w16013 & pi01363;
assign w57705 = ~w16013 & pi01364;
assign w57706 = ~w16013 & pi01365;
assign w57707 = ~w16013 & pi01366;
assign w57708 = w16013 & ~pi10651;
assign w57709 = ~w16013 & pi01367;
assign w57710 = ~w16013 & pi01368;
assign w57711 = w16013 & ~pi10626;
assign w57712 = ~w16013 & pi01369;
assign w57713 = ~w14861 & pi01370;
assign w57714 = w14861 & ~pi10632;
assign w57715 = ~w14861 & pi01371;
assign w57716 = ~w14861 & pi01372;
assign w57717 = ~w14861 & pi01373;
assign w57718 = w14861 & ~pi10635;
assign w57719 = ~w14861 & pi01374;
assign w57720 = w14861 & ~pi10637;
assign w57721 = ~w14861 & pi01375;
assign w57722 = ~w14861 & pi01376;
assign w57723 = w14861 & ~pi10643;
assign w57724 = ~w14861 & pi01377;
assign w57725 = ~w14861 & pi01378;
assign w57726 = ~w14861 & pi01379;
assign w57727 = ~w14861 & pi01380;
assign w57728 = w14861 & ~pi10651;
assign w57729 = ~w14861 & pi01381;
assign w57730 = ~w14861 & pi01382;
assign w57731 = w14861 & ~pi10653;
assign w57732 = ~w14861 & pi01383;
assign w57733 = ~w14861 & pi01384;
assign w57734 = ~w14861 & pi01385;
assign w57735 = ~w14861 & pi01386;
assign w57736 = ~w14861 & pi01387;
assign w57737 = ~w14861 & pi01388;
assign w57738 = ~w14861 & pi01389;
assign w57739 = ~w14861 & pi01390;
assign w57740 = w14861 & ~pi10639;
assign w57741 = ~w14861 & pi01391;
assign w57742 = w14861 & ~pi10641;
assign w57743 = ~w14861 & pi01392;
assign w57744 = ~w14861 & pi01393;
assign w57745 = ~w14861 & pi01394;
assign w57746 = ~w14861 & pi01395;
assign w57747 = ~w14861 & pi01396;
assign w57748 = ~w14861 & pi01397;
assign w57749 = ~w14861 & pi01398;
assign w57750 = ~w14861 & pi01399;
assign w57751 = ~w14861 & pi01400;
assign w57752 = w14861 & ~pi10631;
assign w57753 = ~w16218 & pi01401;
assign w57754 = w16218 & ~pi10622;
assign w57755 = ~w16218 & pi01402;
assign w57756 = ~w16218 & pi01403;
assign w57757 = ~w16218 & pi01404;
assign w57758 = ~w16218 & pi01405;
assign w57759 = w16218 & ~pi10650;
assign w57760 = ~w16218 & pi01406;
assign w57761 = w16218 & ~pi10625;
assign w57762 = ~w16218 & pi01407;
assign w57763 = w16218 & ~pi10626;
assign w57764 = ~w16218 & pi01408;
assign w57765 = ~w16218 & pi01409;
assign w57766 = w16218 & ~pi10629;
assign w57767 = ~w16003 & pi01410;
assign w57768 = ~w16003 & pi01411;
assign w57769 = ~w16003 & pi01412;
assign w57770 = ~w16003 & pi01413;
assign w57771 = ~w16003 & pi01414;
assign w57772 = ~w16013 & pi01415;
assign w57773 = ~w16013 & pi01416;
assign w57774 = w16013 & ~pi10632;
assign w57775 = ~w16013 & pi01417;
assign w57776 = ~w16013 & pi01418;
assign w57777 = w16013 & ~pi10638;
assign w57778 = ~w16013 & pi01419;
assign w57779 = w16013 & ~pi10639;
assign w57780 = ~w16013 & pi01420;
assign w57781 = ~w16013 & pi01421;
assign w57782 = ~w16013 & pi01422;
assign w57783 = ~w16013 & pi01423;
assign w57784 = ~w16013 & pi01424;
assign w57785 = ~w16013 & pi01425;
assign w57786 = ~w16013 & pi01426;
assign w57787 = ~w16218 & pi01440;
assign w57788 = ~w16218 & pi01441;
assign w57789 = ~w16218 & pi01442;
assign w57790 = w16218 & ~pi10638;
assign w57791 = ~w16218 & pi01443;
assign w57792 = ~w16218 & pi01444;
assign w57793 = w16218 & ~pi10641;
assign w57794 = ~w16218 & pi01445;
assign w57795 = ~w16218 & pi01446;
assign w57796 = w16218 & ~pi10631;
assign w57797 = ~w16218 & pi01447;
assign w57798 = w16218 & ~pi10646;
assign w57799 = ~w16218 & pi01448;
assign w57800 = w16218 & ~pi10633;
assign w57801 = w56504 & pi09973;
assign w57802 = w56487 & pi09887;
assign w57803 = ~w12894 & ~w16752;
assign w57804 = ~w16750 & ~w16751;
assign w57805 = ~w16748 & ~w16756;
assign w57806 = w1192 & ~w16764;
assign w57807 = ~w1192 & w16764;
assign w57808 = ~pi01451 & w12993;
assign w57809 = pi09804 & ~pi10438;
assign w57810 = ~w57809 & pi00139;
assign w57811 = w16789 & w16791;
assign w57812 = ~pi09866 & ~pi01452;
assign w57813 = ~w16792 & pi01453;
assign w57814 = ~pi01454 & ~w11706;
assign w57815 = pi02796 & w16788;
assign w57816 = ~w57815 & ~pi01455;
assign w57817 = ~w1268 & pi01456;
assign w57818 = w1268 & pi10590;
assign w57819 = ~w1268 & pi01457;
assign w57820 = w1268 & pi10591;
assign w57821 = ~w1268 & pi01458;
assign w57822 = w1268 & pi10592;
assign w57823 = ~w1268 & pi01459;
assign w57824 = w1268 & pi10593;
assign w57825 = ~w1268 & pi01460;
assign w57826 = w1268 & pi10594;
assign w57827 = ~w1268 & pi01461;
assign w57828 = w1268 & pi10596;
assign w57829 = ~w1264 & pi01462;
assign w57830 = w1264 & pi10591;
assign w57831 = ~w1789 & ~w16833;
assign w57832 = w1789 & w16833;
assign w57833 = ~w1264 & pi01464;
assign w57834 = w1264 & pi10592;
assign w57835 = ~w1264 & pi01465;
assign w57836 = w1264 & pi10593;
assign w57837 = ~w1264 & pi01466;
assign w57838 = w1264 & pi10594;
assign w57839 = ~w1264 & pi01467;
assign w57840 = w1264 & pi10596;
assign w57841 = ~w1264 & pi01468;
assign w57842 = w1264 & pi10595;
assign w57843 = ~w1240 & pi01469;
assign w57844 = w1240 & pi10591;
assign w57845 = ~w1240 & pi01470;
assign w57846 = w1240 & pi10592;
assign w57847 = ~w1240 & pi01471;
assign w57848 = w1240 & pi10593;
assign w57849 = ~w1240 & pi01472;
assign w57850 = w1240 & pi10594;
assign w57851 = ~w1240 & pi01473;
assign w57852 = w1240 & pi10596;
assign w57853 = ~w1240 & pi01474;
assign w57854 = w1240 & pi10597;
assign w57855 = ~w1240 & pi01475;
assign w57856 = w1240 & pi10590;
assign w57857 = ~w1240 & pi01476;
assign w57858 = w1240 & pi10595;
assign w57859 = pi01164 & pi02812;
assign w57860 = ~w57859 & ~w11706;
assign w57861 = ~w13027 & w11706;
assign w57862 = ~w13027 & ~w57860;
assign w57863 = ~w1264 & pi01478;
assign w57864 = w1264 & pi10590;
assign w57865 = pi01168 & ~w12877;
assign w57866 = w16891 & w16899;
assign w57867 = w16904 & w16912;
assign w57868 = w16891 & w16922;
assign w57869 = w16927 & w16931;
assign w57870 = w16904 & w16941;
assign w57871 = w16891 & w16948;
assign w57872 = w16927 & w16954;
assign w57873 = w16891 & w16961;
assign w57874 = w16904 & w16970;
assign w57875 = w16904 & ~pi02717;
assign w57876 = w16970 & ~pi02717;
assign w57877 = w16970 & w57875;
assign w57878 = w16904 & w16978;
assign w57879 = w16904 & w16986;
assign w57880 = w16991 & w16994;
assign w57881 = w16927 & w16999;
assign w57882 = w16904 & w17006;
assign w57883 = w16991 & w17011;
assign w57884 = w16904 & w17017;
assign w57885 = w16904 & ~pi02712;
assign w57886 = w17017 & ~pi02712;
assign w57887 = w17017 & w57885;
assign w57888 = w16927 & w17023;
assign w57889 = w16904 & w17028;
assign w57890 = w16891 & w17039;
assign w57891 = w16927 & w17047;
assign w57892 = w16904 & w17053;
assign w57893 = w16891 & w17060;
assign w57894 = w55589 & ~pi09969;
assign w57895 = w16904 & w16994;
assign w57896 = w16927 & w17078;
assign w57897 = w16927 & w17084;
assign w57898 = w16891 & w17098;
assign w57899 = w16927 & w17103;
assign w57900 = w16991 & w17108;
assign w57901 = w16991 & w17114;
assign w57902 = w16927 & w17119;
assign w57903 = w16927 & w17125;
assign w57904 = w16927 & ~pi02720;
assign w57905 = w17125 & ~pi02720;
assign w57906 = w17125 & w57904;
assign w57907 = w16891 & w17131;
assign w57908 = w16904 & w17137;
assign w57909 = w16927 & w17148;
assign w57910 = w16927 & w17153;
assign w57911 = w16927 & w16912;
assign w57912 = w16927 & w17162;
assign w57913 = w16927 & w17167;
assign w57914 = w16927 & w17172;
assign w57915 = w16927 & w17177;
assign w57916 = w16927 & w17183;
assign w57917 = w16927 & ~pi09848;
assign w57918 = w17183 & ~pi09848;
assign w57919 = w17183 & w57917;
assign w57920 = w16927 & w17190;
assign w57921 = w16927 & ~pi09812;
assign w57922 = w17190 & ~pi09812;
assign w57923 = w17190 & w57921;
assign w57924 = w16991 & w17047;
assign w57925 = w16927 & w17200;
assign w57926 = w17200 & ~pi09812;
assign w57927 = w17200 & w57921;
assign w57928 = w16991 & w17205;
assign w57929 = w16927 & w17210;
assign w57930 = w16891 & w17218;
assign w57931 = w16927 & w17226;
assign w57932 = w16927 & w17231;
assign w57933 = w16927 & w17239;
assign w57934 = w16927 & w17244;
assign w57935 = w17244 & ~pi09812;
assign w57936 = w17244 & w57921;
assign w57937 = w16991 & w17249;
assign w57938 = w16927 & w17254;
assign w57939 = w16927 & w17259;
assign w57940 = w16927 & w17264;
assign w57941 = w17264 & ~pi09812;
assign w57942 = w17264 & w57921;
assign w57943 = w16904 & w17205;
assign w57944 = w17254 & ~pi02720;
assign w57945 = w17254 & w57904;
assign w57946 = w16927 & w17279;
assign w57947 = w16927 & w17284;
assign w57948 = w16904 & w17289;
assign w57949 = w16927 & w17300;
assign w57950 = w16927 & w17305;
assign w57951 = w16927 & ~pi02704;
assign w57952 = w16912 & ~pi02704;
assign w57953 = w16912 & w57951;
assign w57954 = w16904 & w17314;
assign w57955 = w16904 & ~pi02716;
assign w57956 = w17314 & ~pi02716;
assign w57957 = w17314 & w57955;
assign w57958 = w16927 & w17320;
assign one = 1;
assign po00000 = pi00198;// level 0
assign po00001 = pi00178;// level 0
assign po00002 = pi00093;// level 0
assign po00003 = pi00092;// level 0
assign po00004 = pi00112;// level 0
assign po00005 = pi00110;// level 0
assign po00006 = pi00176;// level 0
assign po00007 = pi00109;// level 0
assign po00008 = pi00108;// level 0
assign po00009 = pi00107;// level 0
assign po00010 = pi00091;// level 0
assign po00011 = pi00106;// level 0
assign po00012 = pi00111;// level 0
assign po00013 = pi00118;// level 0
assign po00014 = pi00116;// level 0
assign po00015 = pi00179;// level 0
assign po00016 = pi00302;// level 0
assign po00017 = pi00303;// level 0
assign po00018 = pi00282;// level 0
assign po00019 = pi00283;// level 0
assign po00020 = pi00255;// level 0
assign po00021 = pi00279;// level 0
assign po00022 = pi00278;// level 0
assign po00023 = pi00254;// level 0
assign po00024 = pi00212;// level 0
assign po00025 = pi00214;// level 0
assign po00026 = pi00213;// level 0
assign po00027 = pi00211;// level 0
assign po00028 = pi00192;// level 0
assign po00029 = pi00256;// level 0
assign po00030 = pi00253;// level 0
assign po00031 = pi00210;// level 0
assign po00032 = pi00375;// level 0
assign po00033 = pi00414;// level 0
assign po00034 = pi00432;// level 0
assign po00035 = pi00423;// level 0
assign po00036 = pi00424;// level 0
assign po00037 = pi00425;// level 0
assign po00038 = pi00426;// level 0
assign po00039 = pi00427;// level 0
assign po00040 = pi00428;// level 0
assign po00041 = pi00429;// level 0
assign po00042 = pi00406;// level 0
assign po00043 = pi00407;// level 0
assign po00044 = pi00431;// level 0
assign po00045 = pi00408;// level 0
assign po00046 = pi00409;// level 0
assign po00047 = pi00410;// level 0
assign po00048 = pi00404;// level 0
assign po00049 = pi00411;// level 0
assign po00050 = pi00412;// level 0
assign po00051 = pi00413;// level 0
assign po00052 = pi00415;// level 0
assign po00053 = pi00416;// level 0
assign po00054 = pi00417;// level 0
assign po00055 = pi00418;// level 0
assign po00056 = pi00405;// level 0
assign po00057 = pi00419;// level 0
assign po00058 = pi00420;// level 0
assign po00059 = pi00421;// level 0
assign po00060 = pi00403;// level 0
assign po00061 = pi00422;// level 0
assign po00062 = pi00956;// level 0
assign po00063 = pi00955;// level 0
assign po00064 = pi00882;// level 0
assign po00065 = pi00953;// level 0
assign po00066 = pi00954;// level 0
assign po00067 = pi00952;// level 0
assign po00068 = pi00951;// level 0
assign po00069 = pi00950;// level 0
assign po00070 = pi00949;// level 0
assign po00071 = pi00958;// level 0
assign po00072 = pi00884;// level 0
assign po00073 = pi00948;// level 0
assign po00074 = pi00947;// level 0
assign po00075 = pi00946;// level 0
assign po00076 = pi00883;// level 0
assign po00077 = pi00945;// level 0
assign po00078 = pi00944;// level 0
assign po00079 = pi00943;// level 0
assign po00080 = pi00885;// level 0
assign po00081 = pi00942;// level 0
assign po00082 = pi00941;// level 0
assign po00083 = pi00940;// level 0
assign po00084 = pi00939;// level 0
assign po00085 = pi00937;// level 0
assign po00086 = pi00938;// level 0
assign po00087 = pi00936;// level 0
assign po00088 = pi00935;// level 0
assign po00089 = pi00934;// level 0
assign po00090 = pi00933;// level 0
assign po00091 = pi00932;// level 0
assign po00092 = pi00931;// level 0
assign po00093 = pi00930;// level 0
assign po00094 = pi10016;// level 0
assign po00095 = pi10473;// level 0
assign po00096 = pi00430;// level 0
assign po00097 = pi00440;// level 0
assign po00098 = pi00440;// level 0
assign po00099 = pi10447;// level 0
assign po00100 = pi01606;// level 0
assign po00101 = pi10231;// level 0
assign po00102 = pi09956;// level 0
assign po00103 = pi09957;// level 0
assign po00104 = ~w12;// level 4
assign po00105 = pi00433;// level 0
assign po00106 = pi00462;// level 0
assign po00107 = pi00470;// level 0
assign po00108 = pi00471;// level 0
assign po00109 = pi09933;// level 0
assign po00110 = pi10372;// level 0
assign po00111 = pi10370;// level 0
assign po00112 = pi00961;// level 0
assign po00113 = ~pi10577;// level 0
assign po00114 = one;// level 0
assign po00115 = pi10584;// level 0
assign po00116 = w62;// level 8
assign po00117 = ~w71;// level 7
assign po00118 = ~w77;// level 5
assign po00119 = ~w155;// level 9
assign po00120 = ~w164;// level 9
assign po00121 = ~w167;// level 7
assign po00122 = pi10583;// level 0
assign po00123 = w544;// level 15
assign po00124 = w580;// level 14
assign po00125 = w588;// level 15
assign po00126 = w592;// level 15
assign po00127 = w596;// level 15
assign po00128 = w600;// level 15
assign po00129 = w604;// level 15
assign po00130 = w608;// level 15
assign po00131 = w612;// level 15
assign po00132 = w616;// level 15
assign po00133 = w620;// level 15
assign po00134 = w624;// level 15
assign po00135 = w627;// level 15
assign po00136 = w630;// level 15
assign po00137 = w633;// level 15
assign po00138 = w636;// level 15
assign po00139 = w639;// level 15
assign po00140 = ~w652;// level 10
assign po00141 = w655;// level 15
assign po00142 = w660;// level 14
assign po00143 = ~w661;// level 5
assign po00144 = ~w667;// level 11
assign po00145 = ~w672;// level 4
assign po00146 = ~w673;// level 4
assign po00147 = w675;// level 15
assign po00148 = w678;// level 15
assign po00149 = w681;// level 14
assign po00150 = w691;// level 15
assign po00151 = w696;// level 15
assign po00152 = w700;// level 15
assign po00153 = w704;// level 15
assign po00154 = pi00042;// level 0
assign po00155 = w706;// level 14
assign po00156 = ~w733;// level 10
assign po00157 = ~w746;// level 8
assign po00158 = ~w759;// level 10
assign po00159 = ~w764;// level 14
assign po00160 = ~w776;// level 8
assign po00161 = ~w779;// level 8
assign po00162 = pi00045;// level 0
assign po00163 = ~w764;// level 14
assign po00164 = w780;// level 7
assign po00165 = pi00046;// level 0
assign po00166 = w781;// level 5
assign po00167 = pi00047;// level 0
assign po00168 = ~pi00033;// level 0
assign po00169 = pi00048;// level 0
assign po00170 = ~pi00034;// level 0
assign po00171 = pi00049;// level 0
assign po00172 = ~pi00035;// level 0
assign po00173 = pi00050;// level 0
assign po00174 = ~pi00036;// level 0
assign po00175 = ~w784;// level 9
assign po00176 = ~w788;// level 15
assign po00177 = w791;// level 15
assign po00178 = ~w792;// level 5
assign po00179 = ~w796;// level 8
assign po00180 = ~w802;// level 10
assign po00181 = ~w809;// level 11
assign po00182 = ~w813;// level 9
assign po00183 = ~w819;// level 10
assign po00184 = ~w822;// level 9
assign po00185 = ~w825;// level 9
assign po00186 = pi10576;// level 0
assign po00187 = ~w851;// level 6
assign po00188 = ~w1077;// level 11
assign po00189 = ~w1088;// level 12
assign po00190 = ~w1092;// level 9
assign po00191 = ~w1095;// level 8
assign po00192 = ~w1096;// level 4
assign po00193 = ~w1097;// level 4
assign po00194 = ~w1104;// level 12
assign po00195 = ~w1108;// level 10
assign po00196 = w1120;// level 7
assign po00197 = ~w1140;// level 8
assign po00198 = ~w1146;// level 12
assign po00199 = ~w1149;// level 8
assign po00200 = ~w1152;// level 8
assign po00201 = ~w1155;// level 8
assign po00202 = ~w1158;// level 8
assign po00203 = ~w1161;// level 8
assign po00204 = ~w1164;// level 6
assign po00205 = ~w1167;// level 8
assign po00206 = ~w1170;// level 6
assign po00207 = ~w1173;// level 6
assign po00208 = ~w1176;// level 6
assign po00209 = ~w1179;// level 6
assign po00210 = ~w1182;// level 6
assign po00211 = ~w1185;// level 8
assign po00212 = ~w1188;// level 6
assign po00213 = ~w1191;// level 6
assign po00214 = w1198;// level 4
assign po00215 = w1203;// level 4
assign po00216 = w1255;// level 9
assign po00217 = w1302;// level 10
assign po00218 = w1349;// level 10
assign po00219 = ~w1360;// level 6
assign po00220 = ~w1365;// level 5
assign po00221 = ~w1370;// level 5
assign po00222 = ~w1384;// level 6
assign po00223 = ~w1389;// level 5
assign po00224 = ~w1394;// level 5
assign po00225 = ~w1397;// level 8
assign po00226 = ~w1400;// level 8
assign po00227 = ~w1560;// level 14
assign po00228 = w1591;// level 14
assign po00229 = ~w1598;// level 14
assign po00230 = w1602;// level 4
assign po00231 = w1623;// level 9
assign po00232 = w1644;// level 9
assign po00233 = w1667;// level 9
assign po00234 = w1690;// level 9
assign po00235 = w1726;// level 10
assign po00236 = w1747;// level 9
assign po00237 = w1785;// level 10
assign po00238 = ~w1788;// level 3
assign po00239 = ~w1791;// level 4
assign po00240 = ~w1796;// level 6
assign po00241 = w1816;// level 9
assign po00242 = ~w1822;// level 7
assign po00243 = w1842;// level 9
assign po00244 = ~w1847;// level 6
assign po00245 = ~w1852;// level 6
assign po00246 = ~w1858;// level 6
assign po00247 = ~w1865;// level 7
assign po00248 = ~w1870;// level 7
assign po00249 = ~w1875;// level 6
assign po00250 = ~w1884;// level 7
assign po00251 = ~w1889;// level 6
assign po00252 = ~w1894;// level 6
assign po00253 = ~w1899;// level 7
assign po00254 = ~w1904;// level 7
assign po00255 = ~w1909;// level 6
assign po00256 = ~w1914;// level 6
assign po00257 = w1917;// level 3
assign po00258 = w1920;// level 3
assign po00259 = ~w1925;// level 7
assign po00260 = ~w1930;// level 7
assign po00261 = ~w1935;// level 7
assign po00262 = ~w1938;// level 3
assign po00263 = ~w1941;// level 3
assign po00264 = w1944;// level 3
assign po00265 = w1947;// level 3
assign po00266 = ~w1950;// level 11
assign po00267 = w1960;// level 14
assign po00268 = w1966;// level 14
assign po00269 = w1973;// level 14
assign po00270 = w1978;// level 14
assign po00271 = ~w1982;// level 14
assign po00272 = w1987;// level 14
assign po00273 = w1992;// level 14
assign po00274 = w1998;// level 14
assign po00275 = w2003;// level 14
assign po00276 = w2009;// level 14
assign po00277 = w2014;// level 14
assign po00278 = w2018;// level 14
assign po00279 = w2023;// level 14
assign po00280 = w2028;// level 14
assign po00281 = ~w2061;// level 10
assign po00282 = ~w2064;// level 6
assign po00283 = ~w2067;// level 6
assign po00284 = ~w2070;// level 6
assign po00285 = ~w2073;// level 6
assign po00286 = ~w2076;// level 6
assign po00287 = ~w2079;// level 6
assign po00288 = ~w2082;// level 6
assign po00289 = ~w2085;// level 6
assign po00290 = ~w2089;// level 8
assign po00291 = ~w2092;// level 8
assign po00292 = ~w2095;// level 8
assign po00293 = ~w2098;// level 8
assign po00294 = ~w2101;// level 8
assign po00295 = ~w2104;// level 8
assign po00296 = ~w2107;// level 8
assign po00297 = ~w2110;// level 8
assign po00298 = ~w2121;// level 6
assign po00299 = ~w2123;// level 3
assign po00300 = ~w2126;// level 4
assign po00301 = w2160;// level 10
assign po00302 = ~w2162;// level 4
assign po00303 = w2213;// level 10
assign po00304 = w2233;// level 9
assign po00305 = ~w2238;// level 6
assign po00306 = ~w2243;// level 6
assign po00307 = ~w2253;// level 7
assign po00308 = ~w2259;// level 8
assign po00309 = ~w2262;// level 10
assign po00310 = ~w2266;// level 9
assign po00311 = ~w2269;// level 10
assign po00312 = ~w2273;// level 12
assign po00313 = w2300;// level 10
assign po00314 = ~w2305;// level 10
assign po00315 = ~w2310;// level 10
assign po00316 = ~w2315;// level 10
assign po00317 = ~w2326;// level 8
assign po00318 = ~w2328;// level 3
assign po00319 = ~w2331;// level 3
assign po00320 = ~w2334;// level 3
assign po00321 = ~w2336;// level 3
assign po00322 = ~w2338;// level 3
assign po00323 = w2382;// level 10
assign po00324 = ~w2394;// level 9
assign po00325 = ~w2410;// level 9
assign po00326 = ~w2414;// level 10
assign po00327 = ~w2418;// level 11
assign po00328 = w2430;// level 6
assign po00329 = w2437;// level 13
assign po00330 = ~w2441;// level 10
assign po00331 = ~w2446;// level 10
assign po00332 = ~w2454;// level 4
assign po00333 = ~w2459;// level 11
assign po00334 = ~w2467;// level 10
assign po00335 = ~w2476;// level 8
assign po00336 = ~w2485;// level 8
assign po00337 = ~w2494;// level 8
assign po00338 = ~w2503;// level 8
assign po00339 = ~w2512;// level 8
assign po00340 = ~w2514;// level 3
assign po00341 = ~w2516;// level 3
assign po00342 = ~w2518;// level 3
assign po00343 = ~w2521;// level 3
assign po00344 = ~w2526;// level 8
assign po00345 = ~w2531;// level 9
assign po00346 = ~w2536;// level 9
assign po00347 = ~w2541;// level 10
assign po00348 = ~w2549;// level 10
assign po00349 = ~w2554;// level 9
assign po00350 = ~w2559;// level 9
assign po00351 = ~w2567;// level 11
assign po00352 = ~w2572;// level 9
assign po00353 = ~w2577;// level 10
assign po00354 = ~w2582;// level 10
assign po00355 = w2586;// level 6
assign po00356 = ~w2592;// level 12
assign po00357 = w2596;// level 14
assign po00358 = w2612;// level 9
assign po00359 = w2621;// level 10
assign po00360 = w2625;// level 10
assign po00361 = w2629;// level 10
assign po00362 = w2633;// level 11
assign po00363 = w2636;// level 11
assign po00364 = w2639;// level 12
assign po00365 = w2642;// level 10
assign po00366 = w2645;// level 10
assign po00367 = w2649;// level 10
assign po00368 = w2652;// level 10
assign po00369 = w2655;// level 10
assign po00370 = w2659;// level 10
assign po00371 = w2663;// level 11
assign po00372 = w2666;// level 11
assign po00373 = w2670;// level 11
assign po00374 = w2671;// level 10
assign po00375 = w2673;// level 10
assign po00376 = ~w2678;// level 9
assign po00377 = ~w2683;// level 10
assign po00378 = ~w2692;// level 8
assign po00379 = ~w2701;// level 8
assign po00380 = ~w2710;// level 8
assign po00381 = ~w2719;// level 8
assign po00382 = ~w2722;// level 3
assign po00383 = ~w2725;// level 3
assign po00384 = ~w2728;// level 3
assign po00385 = ~w2731;// level 3
assign po00386 = ~w2736;// level 8
assign po00387 = ~w2741;// level 8
assign po00388 = ~w2746;// level 10
assign po00389 = ~w2752;// level 9
assign po00390 = ~w2757;// level 9
assign po00391 = ~w2762;// level 10
assign po00392 = ~w2764;// level 9
assign po00393 = ~w2767;// level 10
assign po00394 = ~w2771;// level 10
assign po00395 = ~w2775;// level 11
assign po00396 = w2777;// level 10
assign po00397 = w2784;// level 8
assign po00398 = w2790;// level 8
assign po00399 = w2792;// level 4
assign po00400 = w2795;// level 8
assign po00401 = w2797;// level 9
assign po00402 = w2800;// level 8
assign po00403 = ~w2809;// level 8
assign po00404 = ~w2818;// level 8
assign po00405 = ~w2821;// level 3
assign po00406 = ~w2824;// level 3
assign po00407 = ~w2835;// level 8
assign po00408 = ~w2846;// level 8
assign po00409 = ~w2851;// level 8
assign po00410 = ~w2856;// level 9
assign po00411 = ~w2861;// level 8
assign po00412 = ~w2866;// level 9
assign po00413 = ~w2871;// level 9
assign po00414 = ~w2876;// level 9
assign po00415 = ~w2881;// level 8
assign po00416 = ~w2885;// level 7
assign po00417 = ~w2892;// level 9
assign po00418 = ~w2897;// level 9
assign po00419 = w2904;// level 6
assign po00420 = w2911;// level 5
assign po00421 = w2914;// level 5
assign po00422 = ~w2920;// level 12
assign po00423 = ~w2926;// level 12
assign po00424 = w2942;// level 6
assign po00425 = ~w2961;// level 11
assign po00426 = w2964;// level 7
assign po00427 = ~w2980;// level 9
assign po00428 = ~w2991;// level 9
assign po00429 = ~w2996;// level 7
assign po00430 = ~w3001;// level 8
assign po00431 = ~w3007;// level 8
assign po00432 = ~w3012;// level 8
assign po00433 = w3017;// level 5
assign po00434 = w3020;// level 5
assign po00435 = w3023;// level 5
assign po00436 = w3026;// level 6
assign po00437 = ~w3031;// level 5
assign po00438 = ~w3034;// level 5
assign po00439 = ~w3037;// level 5
assign po00440 = ~w3040;// level 5
assign po00441 = ~w3043;// level 5
assign po00442 = ~w3046;// level 5
assign po00443 = ~w3049;// level 5
assign po00444 = ~w3052;// level 6
assign po00445 = w3057;// level 5
assign po00446 = w3877;// level 13
assign po00447 = ~w3883;// level 5
assign po00448 = ~w3887;// level 5
assign po00449 = ~w3890;// level 5
assign po00450 = ~w3893;// level 5
assign po00451 = ~w3896;// level 5
assign po00452 = ~w3899;// level 5
assign po00453 = ~w3902;// level 5
assign po00454 = ~w3905;// level 5
assign po00455 = ~w3908;// level 5
assign po00456 = ~w3911;// level 5
assign po00457 = ~w3914;// level 5
assign po00458 = ~w3917;// level 5
assign po00459 = ~w3920;// level 5
assign po00460 = ~w3923;// level 5
assign po00461 = ~w3926;// level 5
assign po00462 = ~w3929;// level 5
assign po00463 = ~w3932;// level 6
assign po00464 = w3935;// level 5
assign po00465 = w3941;// level 4
assign po00466 = w3944;// level 4
assign po00467 = w3946;// level 4
assign po00468 = w3948;// level 5
assign po00469 = ~w3952;// level 12
assign po00470 = w4464;// level 13
assign po00471 = w4976;// level 13
assign po00472 = w5488;// level 13
assign po00473 = w6000;// level 13
assign po00474 = ~w6009;// level 5
assign po00475 = ~w6014;// level 5
assign po00476 = ~w6017;// level 5
assign po00477 = ~w6020;// level 5
assign po00478 = ~w6023;// level 5
assign po00479 = ~w6026;// level 5
assign po00480 = ~w6029;// level 5
assign po00481 = ~w6032;// level 5
assign po00482 = ~w6035;// level 6
assign po00483 = w6039;// level 5
assign po00484 = ~w6045;// level 12
assign po00485 = ~w6051;// level 12
assign po00486 = ~w6055;// level 12
assign po00487 = ~w6059;// level 12
assign po00488 = w6571;// level 13
assign po00489 = w7083;// level 13
assign po00490 = w7595;// level 13
assign po00491 = ~w7599;// level 5
assign po00492 = ~w7602;// level 10
assign po00493 = w8114;// level 13
assign po00494 = w8626;// level 13
assign po00495 = w9138;// level 13
assign po00496 = w9650;// level 13
assign po00497 = w10162;// level 13
assign po00498 = w10674;// level 13
assign po00499 = ~w10675;// level 11
assign po00500 = w10681;// level 5
assign po00501 = ~w10740;// level 10
assign po00502 = w10742;// level 4
assign po00503 = ~w10751;// level 6
assign po00504 = ~w10754;// level 6
assign po00505 = ~w10757;// level 6
assign po00506 = ~w10760;// level 6
assign po00507 = ~w10763;// level 6
assign po00508 = ~w10766;// level 6
assign po00509 = ~w10771;// level 8
assign po00510 = ~w10774;// level 8
assign po00511 = ~w10777;// level 8
assign po00512 = ~w10780;// level 8
assign po00513 = ~w10783;// level 8
assign po00514 = ~w10786;// level 8
assign po00515 = ~w10789;// level 8
assign po00516 = ~w10792;// level 8
assign po00517 = ~w10796;// level 8
assign po00518 = ~w10799;// level 8
assign po00519 = ~w10802;// level 8
assign po00520 = ~w10805;// level 8
assign po00521 = ~w10808;// level 8
assign po00522 = ~w10811;// level 8
assign po00523 = ~w10814;// level 8
assign po00524 = ~w10817;// level 8
assign po00525 = ~w10820;// level 6
assign po00526 = ~w10823;// level 6
assign po00527 = ~w10826;// level 10
assign po00528 = ~w10829;// level 12
assign po00529 = ~w10866;// level 11
assign po00530 = ~w10881;// level 11
assign po00531 = ~w10891;// level 11
assign po00532 = ~w10900;// level 11
assign po00533 = ~w10907;// level 11
assign po00534 = ~w10915;// level 11
assign po00535 = ~w10924;// level 11
assign po00536 = ~w10931;// level 11
assign po00537 = ~w10938;// level 11
assign po00538 = ~w10946;// level 12
assign po00539 = ~w10953;// level 11
assign po00540 = ~w10961;// level 11
assign po00541 = ~w10969;// level 11
assign po00542 = ~w10977;// level 11
assign po00543 = ~w10984;// level 11
assign po00544 = ~w10992;// level 11
assign po00545 = ~w11000;// level 11
assign po00546 = ~w11007;// level 11
assign po00547 = ~w11015;// level 11
assign po00548 = ~w11023;// level 11
assign po00549 = ~w11032;// level 11
assign po00550 = ~w11040;// level 11
assign po00551 = ~w11048;// level 11
assign po00552 = ~w11056;// level 11
assign po00553 = ~w11064;// level 11
assign po00554 = ~w11072;// level 11
assign po00555 = ~w11080;// level 11
assign po00556 = ~w11082;// level 8
assign po00557 = ~w11089;// level 11
assign po00558 = ~w11096;// level 11
assign po00559 = ~w11097;// level 8
assign po00560 = ~w11103;// level 6
assign po00561 = ~w11112;// level 8
assign po00562 = ~w11119;// level 7
assign po00563 = ~w11122;// level 3
assign po00564 = ~w11124;// level 4
assign po00565 = ~w11134;// level 6
assign po00566 = ~w11136;// level 8
assign po00567 = w11142;// level 7
assign po00568 = ~w11156;// level 9
assign po00569 = ~w11159;// level 6
assign po00570 = ~w11163;// level 3
assign po00571 = ~w11169;// level 6
assign po00572 = ~w11174;// level 6
assign po00573 = ~w11211;// level 7
assign po00574 = ~w11228;// level 7
assign po00575 = ~w11245;// level 7
assign po00576 = ~w11262;// level 7
assign po00577 = ~w11280;// level 8
assign po00578 = ~w11298;// level 8
assign po00579 = ~w11316;// level 8
assign po00580 = ~w11334;// level 8
assign po00581 = ~w11373;// level 9
assign po00582 = ~w11382;// level 9
assign po00583 = w11385;// level 8
assign po00584 = w11388;// level 8
assign po00585 = w11391;// level 9
assign po00586 = ~w11393;// level 8
assign po00587 = ~w11395;// level 8
assign po00588 = ~w11401;// level 10
assign po00589 = ~w11405;// level 11
assign po00590 = ~w11408;// level 12
assign po00591 = ~w11409;// level 5
assign po00592 = ~w11420;// level 9
assign po00593 = ~w11431;// level 9
assign po00594 = ~w11442;// level 9
assign po00595 = ~w11453;// level 9
assign po00596 = ~w11455;// level 9
assign po00597 = ~w11459;// level 9
assign po00598 = ~w11462;// level 11
assign po00599 = ~w11465;// level 7
assign po00600 = ~w11477;// level 9
assign po00601 = ~w11483;// level 4
assign po00602 = pi00535;// level 0
assign po00603 = ~w11520;// level 8
assign po00604 = ~w11523;// level 8
assign po00605 = ~w11526;// level 8
assign po00606 = ~w11529;// level 8
assign po00607 = ~w11532;// level 8
assign po00608 = ~w11535;// level 8
assign po00609 = ~w11538;// level 8
assign po00610 = ~w11541;// level 8
assign po00611 = ~w11550;// level 9
assign po00612 = ~w11559;// level 9
assign po00613 = w11702;// level 11
assign po00614 = w11704;// level 8
assign po00615 = w11714;// level 6
assign po00616 = w11717;// level 6
assign po00617 = w11720;// level 6
assign po00618 = w11723;// level 6
assign po00619 = w11726;// level 6
assign po00620 = w11729;// level 6
assign po00621 = w11732;// level 6
assign po00622 = w11736;// level 6
assign po00623 = w11739;// level 6
assign po00624 = w11742;// level 6
assign po00625 = w11745;// level 6
assign po00626 = w11748;// level 6
assign po00627 = w11751;// level 6
assign po00628 = w11754;// level 6
assign po00629 = w11757;// level 6
assign po00630 = w11760;// level 6
assign po00631 = w11765;// level 6
assign po00632 = w11768;// level 6
assign po00633 = w11771;// level 6
assign po00634 = w11774;// level 6
assign po00635 = w11777;// level 6
assign po00636 = w11780;// level 6
assign po00637 = w11783;// level 6
assign po00638 = w11786;// level 6
assign po00639 = w11789;// level 6
assign po00640 = w11792;// level 6
assign po00641 = w11795;// level 6
assign po00642 = w11798;// level 6
assign po00643 = w11803;// level 6
assign po00644 = w11806;// level 6
assign po00645 = w11809;// level 6
assign po00646 = w11812;// level 6
assign po00647 = w11815;// level 6
assign po00648 = w11818;// level 6
assign po00649 = w11821;// level 6
assign po00650 = w11824;// level 6
assign po00651 = w11831;// level 6
assign po00652 = w11834;// level 6
assign po00653 = w11837;// level 6
assign po00654 = w11840;// level 6
assign po00655 = w11843;// level 6
assign po00656 = w11846;// level 6
assign po00657 = w11849;// level 6
assign po00658 = w11852;// level 6
assign po00659 = w11855;// level 6
assign po00660 = w11858;// level 6
assign po00661 = w11861;// level 2
assign po00662 = ~w11864;// level 12
assign po00663 = ~w11867;// level 12
assign po00664 = w11898;// level 9
assign po00665 = ~w11900;// level 10
assign po00666 = w11903;// level 8
assign po00667 = w11905;// level 5
assign po00668 = w11908;// level 6
assign po00669 = w11911;// level 6
assign po00670 = w11914;// level 6
assign po00671 = w11917;// level 6
assign po00672 = w11920;// level 6
assign po00673 = w11923;// level 6
assign po00674 = w11926;// level 6
assign po00675 = w11929;// level 6
assign po00676 = w11932;// level 6
assign po00677 = w11935;// level 6
assign po00678 = w11938;// level 6
assign po00679 = w11941;// level 6
assign po00680 = w11944;// level 6
assign po00681 = w11947;// level 6
assign po00682 = w11950;// level 6
assign po00683 = w11953;// level 6
assign po00684 = w11956;// level 6
assign po00685 = w11959;// level 6
assign po00686 = w11962;// level 6
assign po00687 = w11965;// level 6
assign po00688 = w11968;// level 6
assign po00689 = w11971;// level 6
assign po00690 = w11974;// level 6
assign po00691 = w11977;// level 6
assign po00692 = w11980;// level 6
assign po00693 = w11983;// level 6
assign po00694 = w11986;// level 6
assign po00695 = w11989;// level 6
assign po00696 = w11992;// level 6
assign po00697 = w11995;// level 6
assign po00698 = w11998;// level 6
assign po00699 = w12001;// level 6
assign po00700 = w12004;// level 6
assign po00701 = w12007;// level 6
assign po00702 = w12010;// level 6
assign po00703 = w12013;// level 6
assign po00704 = w12016;// level 6
assign po00705 = w12019;// level 6
assign po00706 = w12022;// level 6
assign po00707 = w12025;// level 6
assign po00708 = w12028;// level 6
assign po00709 = w12031;// level 6
assign po00710 = w12034;// level 6
assign po00711 = w12037;// level 6
assign po00712 = w12040;// level 6
assign po00713 = w12043;// level 6
assign po00714 = w12046;// level 6
assign po00715 = w12049;// level 6
assign po00716 = w12052;// level 6
assign po00717 = w12055;// level 6
assign po00718 = w12058;// level 6
assign po00719 = w12061;// level 6
assign po00720 = w12064;// level 6
assign po00721 = w12067;// level 6
assign po00722 = w12070;// level 6
assign po00723 = w12073;// level 6
assign po00724 = w12076;// level 6
assign po00725 = w12079;// level 6
assign po00726 = w12082;// level 6
assign po00727 = w12085;// level 6
assign po00728 = w12088;// level 6
assign po00729 = w12091;// level 6
assign po00730 = w12094;// level 6
assign po00731 = w12097;// level 6
assign po00732 = w12100;// level 6
assign po00733 = w12103;// level 6
assign po00734 = w12107;// level 6
assign po00735 = ~w12112;// level 4
assign po00736 = ~w12116;// level 10
assign po00737 = ~w12122;// level 6
assign po00738 = ~w12125;// level 6
assign po00739 = ~w12128;// level 6
assign po00740 = ~w12131;// level 6
assign po00741 = ~w12134;// level 6
assign po00742 = ~w12137;// level 6
assign po00743 = ~w12140;// level 6
assign po00744 = ~w12143;// level 6
assign po00745 = ~w12146;// level 6
assign po00746 = ~w12149;// level 6
assign po00747 = ~w12152;// level 6
assign po00748 = ~w12155;// level 6
assign po00749 = ~w12158;// level 6
assign po00750 = ~w12161;// level 6
assign po00751 = ~w12164;// level 6
assign po00752 = ~w12167;// level 6
assign po00753 = ~w12170;// level 6
assign po00754 = ~w12173;// level 6
assign po00755 = ~w12176;// level 6
assign po00756 = ~w12179;// level 6
assign po00757 = ~w12182;// level 6
assign po00758 = ~w12185;// level 6
assign po00759 = ~w12188;// level 6
assign po00760 = ~w12191;// level 6
assign po00761 = ~w12194;// level 6
assign po00762 = ~w12197;// level 6
assign po00763 = ~w12200;// level 6
assign po00764 = ~w12203;// level 6
assign po00765 = ~w12206;// level 6
assign po00766 = ~w12209;// level 6
assign po00767 = ~w12212;// level 6
assign po00768 = ~w12215;// level 6
assign po00769 = w12218;// level 9
assign po00770 = ~w12223;// level 7
assign po00771 = ~w12226;// level 7
assign po00772 = ~w12229;// level 7
assign po00773 = ~w12232;// level 7
assign po00774 = ~w12235;// level 7
assign po00775 = ~w12238;// level 7
assign po00776 = ~w12241;// level 7
assign po00777 = ~w12244;// level 7
assign po00778 = ~w12247;// level 7
assign po00779 = ~w12250;// level 7
assign po00780 = ~w12253;// level 7
assign po00781 = ~w12256;// level 7
assign po00782 = ~w12259;// level 7
assign po00783 = ~w12262;// level 7
assign po00784 = ~w12265;// level 7
assign po00785 = ~w12268;// level 7
assign po00786 = ~w12271;// level 7
assign po00787 = ~w12274;// level 7
assign po00788 = ~w12277;// level 7
assign po00789 = ~w12280;// level 7
assign po00790 = ~w12283;// level 7
assign po00791 = ~w12286;// level 7
assign po00792 = ~w12289;// level 7
assign po00793 = ~w12292;// level 7
assign po00794 = ~w12295;// level 7
assign po00795 = ~w12298;// level 7
assign po00796 = ~w12301;// level 7
assign po00797 = ~w12304;// level 7
assign po00798 = ~w12307;// level 7
assign po00799 = ~w12310;// level 7
assign po00800 = ~w12313;// level 7
assign po00801 = ~w12316;// level 7
assign po00802 = w12319;// level 6
assign po00803 = w12322;// level 6
assign po00804 = w12325;// level 6
assign po00805 = w12328;// level 6
assign po00806 = w12331;// level 6
assign po00807 = w12334;// level 6
assign po00808 = w12337;// level 6
assign po00809 = w12340;// level 6
assign po00810 = w12343;// level 6
assign po00811 = w12346;// level 6
assign po00812 = w12349;// level 6
assign po00813 = w12352;// level 6
assign po00814 = w12355;// level 6
assign po00815 = w12358;// level 6
assign po00816 = w12361;// level 6
assign po00817 = w12364;// level 6
assign po00818 = w12367;// level 6
assign po00819 = w12370;// level 6
assign po00820 = w12373;// level 6
assign po00821 = w12376;// level 6
assign po00822 = w12379;// level 6
assign po00823 = w12382;// level 6
assign po00824 = w12385;// level 6
assign po00825 = w12388;// level 6
assign po00826 = w12391;// level 6
assign po00827 = w12394;// level 6
assign po00828 = w12397;// level 6
assign po00829 = w12400;// level 6
assign po00830 = w12403;// level 6
assign po00831 = w12406;// level 6
assign po00832 = w12409;// level 6
assign po00833 = w12412;// level 6
assign po00834 = w12415;// level 6
assign po00835 = w12418;// level 6
assign po00836 = w12421;// level 6
assign po00837 = w12424;// level 6
assign po00838 = w12427;// level 6
assign po00839 = w12430;// level 6
assign po00840 = w12433;// level 6
assign po00841 = w12436;// level 6
assign po00842 = w12439;// level 6
assign po00843 = w12442;// level 6
assign po00844 = w12445;// level 6
assign po00845 = w12448;// level 6
assign po00846 = w12451;// level 6
assign po00847 = w12454;// level 6
assign po00848 = w12457;// level 6
assign po00849 = w12460;// level 6
assign po00850 = w12463;// level 6
assign po00851 = w12466;// level 6
assign po00852 = w12469;// level 6
assign po00853 = w12472;// level 6
assign po00854 = w12475;// level 6
assign po00855 = w12478;// level 6
assign po00856 = w12481;// level 6
assign po00857 = w12484;// level 6
assign po00858 = w12487;// level 6
assign po00859 = w12490;// level 6
assign po00860 = w12493;// level 6
assign po00861 = w12496;// level 6
assign po00862 = w12499;// level 6
assign po00863 = w12502;// level 6
assign po00864 = w12505;// level 6
assign po00865 = w12508;// level 6
assign po00866 = w12511;// level 6
assign po00867 = w12514;// level 6
assign po00868 = w12517;// level 6
assign po00869 = w12520;// level 6
assign po00870 = w12523;// level 6
assign po00871 = w12526;// level 6
assign po00872 = w12529;// level 6
assign po00873 = w12532;// level 6
assign po00874 = w12535;// level 6
assign po00875 = w12538;// level 6
assign po00876 = w12541;// level 6
assign po00877 = w12544;// level 6
assign po00878 = w12547;// level 6
assign po00879 = w12550;// level 6
assign po00880 = w12553;// level 6
assign po00881 = w12556;// level 6
assign po00882 = w12559;// level 6
assign po00883 = w12562;// level 6
assign po00884 = w12565;// level 6
assign po00885 = w12568;// level 6
assign po00886 = w12571;// level 6
assign po00887 = w12574;// level 6
assign po00888 = w12577;// level 6
assign po00889 = w12580;// level 6
assign po00890 = w12583;// level 6
assign po00891 = w12586;// level 6
assign po00892 = w12589;// level 6
assign po00893 = w12592;// level 6
assign po00894 = w12595;// level 6
assign po00895 = w12598;// level 6
assign po00896 = w12601;// level 6
assign po00897 = w12604;// level 6
assign po00898 = w12607;// level 6
assign po00899 = w12610;// level 6
assign po00900 = w12613;// level 6
assign po00901 = w12616;// level 6
assign po00902 = w12619;// level 6
assign po00903 = w12622;// level 6
assign po00904 = w12625;// level 6
assign po00905 = w12628;// level 6
assign po00906 = w12631;// level 6
assign po00907 = w12634;// level 6
assign po00908 = w12637;// level 6
assign po00909 = w12640;// level 6
assign po00910 = w12643;// level 6
assign po00911 = w12646;// level 6
assign po00912 = w12649;// level 6
assign po00913 = w12652;// level 6
assign po00914 = w12655;// level 6
assign po00915 = w12658;// level 6
assign po00916 = w12661;// level 6
assign po00917 = w12664;// level 6
assign po00918 = w12667;// level 6
assign po00919 = w12670;// level 6
assign po00920 = w12673;// level 6
assign po00921 = w12676;// level 6
assign po00922 = w12679;// level 6
assign po00923 = w12682;// level 6
assign po00924 = w12685;// level 6
assign po00925 = w12688;// level 6
assign po00926 = w12691;// level 6
assign po00927 = w12694;// level 6
assign po00928 = w12697;// level 6
assign po00929 = w12700;// level 6
assign po00930 = w12703;// level 6
assign po00931 = w12706;// level 6
assign po00932 = w12709;// level 6
assign po00933 = w12712;// level 6
assign po00934 = w12716;// level 6
assign po00935 = w12719;// level 5
assign po00936 = ~w12721;// level 6
assign po00937 = w12727;// level 4
assign po00938 = pi00886;// level 0
assign po00939 = pi00847;// level 0
assign po00940 = pi00846;// level 0
assign po00941 = w12754;// level 9
assign po00942 = w12757;// level 2
assign po00943 = ~w12760;// level 3
assign po00944 = ~w12763;// level 7
assign po00945 = ~w12766;// level 7
assign po00946 = ~w12769;// level 7
assign po00947 = ~w12772;// level 7
assign po00948 = ~w12775;// level 7
assign po00949 = ~w12778;// level 7
assign po00950 = ~w12779;// level 11
assign po00951 = ~w12780;// level 11
assign po00952 = w12783;// level 9
assign po00953 = w12787;// level 8
assign po00954 = w12790;// level 9
assign po00955 = w12793;// level 9
assign po00956 = w12796;// level 9
assign po00957 = w12800;// level 9
assign po00958 = w12804;// level 9
assign po00959 = w12808;// level 9
assign po00960 = w12812;// level 9
assign po00961 = w12816;// level 9
assign po00962 = w12820;// level 9
assign po00963 = w12823;// level 8
assign po00964 = w12826;// level 9
assign po00965 = w12829;// level 9
assign po00966 = w12832;// level 9
assign po00967 = ~w12835;// level 7
assign po00968 = w12839;// level 7
assign po00969 = w12843;// level 7
assign po00970 = w12862;// level 7
assign po00971 = ~w12866;// level 3
assign po00972 = w11116;// level 5
assign po00973 = pi01203;// level 0
assign po00974 = w12870;// level 8
assign po00975 = w12873;// level 7
assign po00976 = ~w12892;// level 7
assign po00977 = w12930;// level 9
assign po00978 = w12933;// level 7
assign po00979 = ~w12936;// level 7
assign po00980 = ~w12939;// level 7
assign po00981 = ~w12942;// level 7
assign po00982 = ~w12946;// level 7
assign po00983 = w12950;// level 7
assign po00984 = w12953;// level 7
assign po00985 = w12956;// level 8
assign po00986 = w12959;// level 8
assign po00987 = w12962;// level 8
assign po00988 = w12965;// level 8
assign po00989 = w12968;// level 8
assign po00990 = w12971;// level 8
assign po00991 = w12974;// level 8
assign po00992 = w12977;// level 7
assign po00993 = w12980;// level 7
assign po00994 = w12983;// level 7
assign po00995 = ~w2433;// level 8
assign po00996 = ~w12997;// level 7
assign po00997 = w13000;// level 8
assign po00998 = w13003;// level 6
assign po00999 = w13006;// level 7
assign po01000 = ~w13009;// level 7
assign po01001 = ~w13012;// level 7
assign po01002 = ~w13015;// level 7
assign po01003 = ~w13018;// level 7
assign po01004 = ~w13025;// level 5
assign po01005 = ~w13026;// level 9
assign po01006 = w12724;// level 3
assign po01007 = pi01480;// level 0
assign po01008 = ~w13076;// level 7
assign po01009 = ~w13107;// level 7
assign po01010 = ~w13138;// level 7
assign po01011 = ~w13169;// level 7
assign po01012 = ~w749;// level 2
assign po01013 = w13172;// level 6
assign po01014 = w13175;// level 6
assign po01015 = w13178;// level 6
assign po01016 = w13181;// level 6
assign po01017 = w13184;// level 6
assign po01018 = w13187;// level 6
assign po01019 = w13190;// level 6
assign po01020 = w13193;// level 6
assign po01021 = w13196;// level 6
assign po01022 = w13199;// level 6
assign po01023 = w13202;// level 6
assign po01024 = w13205;// level 6
assign po01025 = w13208;// level 6
assign po01026 = w13211;// level 6
assign po01027 = w13214;// level 6
assign po01028 = w13217;// level 6
assign po01029 = w13220;// level 6
assign po01030 = w13223;// level 6
assign po01031 = w13226;// level 6
assign po01032 = w13229;// level 6
assign po01033 = w13232;// level 6
assign po01034 = w13235;// level 6
assign po01035 = w13238;// level 6
assign po01036 = w13241;// level 6
assign po01037 = w13244;// level 6
assign po01038 = w13247;// level 6
assign po01039 = w13250;// level 6
assign po01040 = w13253;// level 6
assign po01041 = w13256;// level 6
assign po01042 = w13259;// level 6
assign po01043 = w13262;// level 6
assign po01044 = w13265;// level 6
assign po01045 = w13268;// level 6
assign po01046 = w13271;// level 6
assign po01047 = w13274;// level 6
assign po01048 = w13277;// level 6
assign po01049 = w13280;// level 6
assign po01050 = w13283;// level 6
assign po01051 = w13286;// level 6
assign po01052 = w13289;// level 6
assign po01053 = w13292;// level 6
assign po01054 = w13295;// level 6
assign po01055 = w13297;// level 6
assign po01056 = ~w13328;// level 7
assign po01057 = ~w13359;// level 7
assign po01058 = ~w13390;// level 7
assign po01059 = ~w13421;// level 7
assign po01060 = ~w13452;// level 7
assign po01061 = ~w13483;// level 7
assign po01062 = ~w13514;// level 7
assign po01063 = ~w13545;// level 7
assign po01064 = ~w13576;// level 7
assign po01065 = ~w13607;// level 7
assign po01066 = ~w13638;// level 7
assign po01067 = ~w13669;// level 7
assign po01068 = ~w13700;// level 7
assign po01069 = ~w13731;// level 7
assign po01070 = ~w13762;// level 7
assign po01071 = ~w13793;// level 7
assign po01072 = ~w13824;// level 7
assign po01073 = ~w13855;// level 7
assign po01074 = ~w13886;// level 7
assign po01075 = ~w13917;// level 7
assign po01076 = ~w13948;// level 7
assign po01077 = ~w13979;// level 7
assign po01078 = ~w14010;// level 7
assign po01079 = ~w14041;// level 7
assign po01080 = ~w14072;// level 7
assign po01081 = ~w14103;// level 7
assign po01082 = ~w14134;// level 7
assign po01083 = ~w14155;// level 8
assign po01084 = ~w14186;// level 8
assign po01085 = ~w14200;// level 7
assign po01086 = w14203;// level 7
assign po01087 = ~w14209;// level 6
assign po01088 = w14211;// level 7
assign po01089 = w14217;// level 7
assign po01090 = ~w14220;// level 7
assign po01091 = ~w14223;// level 7
assign po01092 = ~w14226;// level 7
assign po01093 = ~w14249;// level 9
assign po01094 = w14253;// level 8
assign po01095 = w14256;// level 8
assign po01096 = ~w14264;// level 7
assign po01097 = w14267;// level 6
assign po01098 = w14270;// level 6
assign po01099 = w14273;// level 6
assign po01100 = w14276;// level 6
assign po01101 = w14279;// level 6
assign po01102 = w14282;// level 6
assign po01103 = w14285;// level 6
assign po01104 = w14288;// level 6
assign po01105 = w14291;// level 6
assign po01106 = w14294;// level 6
assign po01107 = w14297;// level 6
assign po01108 = w14300;// level 6
assign po01109 = w14303;// level 6
assign po01110 = w14306;// level 6
assign po01111 = w14309;// level 6
assign po01112 = w14312;// level 6
assign po01113 = w14315;// level 6
assign po01114 = w14318;// level 6
assign po01115 = w14321;// level 6
assign po01116 = w14324;// level 6
assign po01117 = w14327;// level 6
assign po01118 = w14330;// level 6
assign po01119 = w14333;// level 6
assign po01120 = w14336;// level 6
assign po01121 = w14339;// level 6
assign po01122 = w14342;// level 6
assign po01123 = w14345;// level 6
assign po01124 = w14348;// level 6
assign po01125 = w14351;// level 6
assign po01126 = w14354;// level 6
assign po01127 = w14357;// level 6
assign po01128 = w14360;// level 6
assign po01129 = w14363;// level 6
assign po01130 = w14366;// level 6
assign po01131 = w14369;// level 6
assign po01132 = w14372;// level 6
assign po01133 = w14375;// level 6
assign po01134 = w14378;// level 6
assign po01135 = w14381;// level 6
assign po01136 = w14384;// level 6
assign po01137 = w14387;// level 6
assign po01138 = w14390;// level 6
assign po01139 = w14393;// level 6
assign po01140 = w14396;// level 6
assign po01141 = w14399;// level 6
assign po01142 = w14402;// level 6
assign po01143 = w14405;// level 6
assign po01144 = w14408;// level 6
assign po01145 = w14411;// level 6
assign po01146 = w14414;// level 6
assign po01147 = w14417;// level 6
assign po01148 = w14420;// level 6
assign po01149 = w14423;// level 6
assign po01150 = w14426;// level 6
assign po01151 = w14429;// level 6
assign po01152 = w14432;// level 6
assign po01153 = w14435;// level 6
assign po01154 = w14438;// level 6
assign po01155 = w14441;// level 6
assign po01156 = w14444;// level 6
assign po01157 = w14447;// level 6
assign po01158 = w14450;// level 6
assign po01159 = w14453;// level 6
assign po01160 = w14456;// level 6
assign po01161 = w14459;// level 6
assign po01162 = w14462;// level 6
assign po01163 = w14465;// level 6
assign po01164 = w14468;// level 6
assign po01165 = w14471;// level 6
assign po01166 = w14474;// level 6
assign po01167 = w14477;// level 6
assign po01168 = w14480;// level 6
assign po01169 = w14483;// level 6
assign po01170 = w14486;// level 6
assign po01171 = w14489;// level 6
assign po01172 = w14492;// level 6
assign po01173 = w14495;// level 6
assign po01174 = w14498;// level 6
assign po01175 = w14501;// level 6
assign po01176 = w14504;// level 6
assign po01177 = w14507;// level 6
assign po01178 = w14510;// level 6
assign po01179 = w14513;// level 6
assign po01180 = w14516;// level 6
assign po01181 = w14519;// level 6
assign po01182 = w14522;// level 6
assign po01183 = w14525;// level 6
assign po01184 = w14528;// level 6
assign po01185 = w14531;// level 6
assign po01186 = w14534;// level 6
assign po01187 = w14537;// level 6
assign po01188 = w14540;// level 6
assign po01189 = w14543;// level 6
assign po01190 = w14546;// level 6
assign po01191 = w14549;// level 6
assign po01192 = w14552;// level 6
assign po01193 = w14555;// level 6
assign po01194 = w14558;// level 6
assign po01195 = w14561;// level 6
assign po01196 = w14564;// level 6
assign po01197 = w14567;// level 6
assign po01198 = w14570;// level 6
assign po01199 = w14573;// level 6
assign po01200 = w14576;// level 6
assign po01201 = w14579;// level 6
assign po01202 = w14582;// level 6
assign po01203 = w14585;// level 6
assign po01204 = w14588;// level 6
assign po01205 = w14591;// level 6
assign po01206 = w14594;// level 6
assign po01207 = w14597;// level 6
assign po01208 = w14600;// level 6
assign po01209 = w14603;// level 6
assign po01210 = w14606;// level 6
assign po01211 = w14609;// level 6
assign po01212 = w14612;// level 6
assign po01213 = w14615;// level 6
assign po01214 = w14618;// level 6
assign po01215 = w14621;// level 6
assign po01216 = w14624;// level 6
assign po01217 = w14627;// level 6
assign po01218 = w14630;// level 6
assign po01219 = w14633;// level 6
assign po01220 = w14636;// level 6
assign po01221 = w14639;// level 6
assign po01222 = w14642;// level 6
assign po01223 = w14645;// level 6
assign po01224 = w14648;// level 6
assign po01225 = w14651;// level 6
assign po01226 = w14654;// level 6
assign po01227 = w14657;// level 6
assign po01228 = w14660;// level 6
assign po01229 = w14663;// level 6
assign po01230 = w14666;// level 6
assign po01231 = w14669;// level 6
assign po01232 = w14672;// level 6
assign po01233 = w14675;// level 6
assign po01234 = w14678;// level 6
assign po01235 = w14681;// level 6
assign po01236 = w14684;// level 6
assign po01237 = w14687;// level 6
assign po01238 = w14690;// level 6
assign po01239 = w14693;// level 6
assign po01240 = w14696;// level 6
assign po01241 = w14699;// level 6
assign po01242 = w14702;// level 6
assign po01243 = w14705;// level 6
assign po01244 = w14708;// level 6
assign po01245 = w14711;// level 6
assign po01246 = w14714;// level 6
assign po01247 = w14717;// level 6
assign po01248 = w14720;// level 6
assign po01249 = w14723;// level 6
assign po01250 = w14726;// level 6
assign po01251 = w14729;// level 6
assign po01252 = w14732;// level 6
assign po01253 = w14735;// level 6
assign po01254 = w14738;// level 6
assign po01255 = w14741;// level 6
assign po01256 = w14744;// level 6
assign po01257 = w14747;// level 6
assign po01258 = w14750;// level 6
assign po01259 = w14753;// level 6
assign po01260 = w14756;// level 6
assign po01261 = w14759;// level 6
assign po01262 = w14762;// level 6
assign po01263 = w14765;// level 6
assign po01264 = w14768;// level 6
assign po01265 = w14771;// level 6
assign po01266 = w14774;// level 6
assign po01267 = w14777;// level 6
assign po01268 = w14780;// level 6
assign po01269 = w14783;// level 6
assign po01270 = w14786;// level 6
assign po01271 = w14789;// level 6
assign po01272 = w14792;// level 6
assign po01273 = w14795;// level 6
assign po01274 = w14798;// level 6
assign po01275 = w14801;// level 6
assign po01276 = w14804;// level 6
assign po01277 = w14807;// level 6
assign po01278 = w14810;// level 6
assign po01279 = w14813;// level 6
assign po01280 = w14816;// level 6
assign po01281 = w14819;// level 6
assign po01282 = w14822;// level 6
assign po01283 = w14825;// level 6
assign po01284 = w14828;// level 6
assign po01285 = w14831;// level 6
assign po01286 = w14834;// level 6
assign po01287 = w14837;// level 6
assign po01288 = w14840;// level 6
assign po01289 = w14843;// level 6
assign po01290 = ~w14850;// level 6
assign po01291 = w14853;// level 3
assign po01292 = ~w14854;// level 9
assign po01293 = ~w14855;// level 11
assign po01294 = w14860;// level 5
assign po01295 = w14869;// level 6
assign po01296 = w14871;// level 7
assign po01297 = ~w14928;// level 9
assign po01298 = ~w14960;// level 9
assign po01299 = ~w14992;// level 9
assign po01300 = ~w15024;// level 9
assign po01301 = ~w15056;// level 9
assign po01302 = ~w15088;// level 9
assign po01303 = ~w15120;// level 9
assign po01304 = ~w15152;// level 9
assign po01305 = ~w15184;// level 9
assign po01306 = ~w15216;// level 9
assign po01307 = ~w15248;// level 9
assign po01308 = ~w15280;// level 9
assign po01309 = ~w15312;// level 9
assign po01310 = ~w15344;// level 9
assign po01311 = ~w15376;// level 9
assign po01312 = ~w15408;// level 9
assign po01313 = ~w15440;// level 9
assign po01314 = ~w15472;// level 9
assign po01315 = ~w15504;// level 9
assign po01316 = ~w15536;// level 9
assign po01317 = ~w15568;// level 9
assign po01318 = ~w15600;// level 9
assign po01319 = ~w15632;// level 9
assign po01320 = ~w15664;// level 9
assign po01321 = ~w15696;// level 9
assign po01322 = ~w15728;// level 9
assign po01323 = ~w15760;// level 9
assign po01324 = ~w15792;// level 9
assign po01325 = ~w15824;// level 9
assign po01326 = ~w15856;// level 9
assign po01327 = ~w15888;// level 9
assign po01328 = ~w15920;// level 9
assign po01329 = ~w15921;// level 5
assign po01330 = w15927;// level 7
assign po01331 = w15928;// level 4
assign po01332 = w15934;// level 7
assign po01333 = ~w15940;// level 7
assign po01334 = w15943;// level 8
assign po01335 = w15952;// level 7
assign po01336 = ~w15956;// level 7
assign po01337 = ~w15966;// level 6
assign po01338 = w15969;// level 6
assign po01339 = w15972;// level 5
assign po01340 = w15978;// level 8
assign po01341 = ~w15983;// level 8
assign po01342 = ~w15990;// level 7
assign po01343 = w16002;// level 8
assign po01344 = w16009;// level 6
assign po01345 = w16012;// level 6
assign po01346 = w16017;// level 6
assign po01347 = w16020;// level 6
assign po01348 = w16023;// level 6
assign po01349 = w16026;// level 6
assign po01350 = w16029;// level 6
assign po01351 = w16035;// level 6
assign po01352 = w16038;// level 6
assign po01353 = w16041;// level 6
assign po01354 = w16044;// level 6
assign po01355 = w16047;// level 6
assign po01356 = w16050;// level 6
assign po01357 = w16053;// level 6
assign po01358 = w16057;// level 6
assign po01359 = w16060;// level 6
assign po01360 = w16063;// level 6
assign po01361 = w16066;// level 6
assign po01362 = w16069;// level 6
assign po01363 = w16072;// level 6
assign po01364 = w16075;// level 6
assign po01365 = w16078;// level 6
assign po01366 = w16081;// level 6
assign po01367 = w16084;// level 6
assign po01368 = w16087;// level 6
assign po01369 = w16090;// level 6
assign po01370 = w16093;// level 6
assign po01371 = w16096;// level 6
assign po01372 = w16099;// level 6
assign po01373 = w16102;// level 6
assign po01374 = w16105;// level 6
assign po01375 = ~w16109;// level 7
assign po01376 = w16112;// level 7
assign po01377 = ~w16115;// level 6
assign po01378 = ~w16118;// level 6
assign po01379 = ~w16121;// level 6
assign po01380 = ~w16124;// level 6
assign po01381 = ~w16127;// level 6
assign po01382 = ~w16130;// level 6
assign po01383 = ~w16133;// level 6
assign po01384 = ~w16136;// level 6
assign po01385 = ~w16139;// level 6
assign po01386 = ~w16142;// level 6
assign po01387 = w16147;// level 7
assign po01388 = w16150;// level 7
assign po01389 = ~w16153;// level 6
assign po01390 = ~w16156;// level 6
assign po01391 = ~w16159;// level 6
assign po01392 = ~w16162;// level 6
assign po01393 = ~w16165;// level 6
assign po01394 = ~w16168;// level 6
assign po01395 = ~w16171;// level 6
assign po01396 = w16179;// level 5
assign po01397 = w16186;// level 5
assign po01398 = pi01506;// level 0
assign po01399 = ~w16191;// level 4
assign po01400 = w16202;// level 9
assign po01401 = ~w16206;// level 5
assign po01402 = ~w16207;// level 10
assign po01403 = w16209;// level 9
assign po01404 = ~w16212;// level 6
assign po01405 = w16217;// level 6
assign po01406 = w16222;// level 6
assign po01407 = w16228;// level 6
assign po01408 = w16232;// level 6
assign po01409 = w16236;// level 6
assign po01410 = w16240;// level 6
assign po01411 = w16243;// level 6
assign po01412 = w16247;// level 6
assign po01413 = w16250;// level 6
assign po01414 = w16254;// level 6
assign po01415 = w16257;// level 6
assign po01416 = w16260;// level 6
assign po01417 = w16264;// level 6
assign po01418 = w16267;// level 6
assign po01419 = w16270;// level 6
assign po01420 = w16274;// level 6
assign po01421 = w16277;// level 6
assign po01422 = w16280;// level 6
assign po01423 = w16283;// level 6
assign po01424 = w16286;// level 6
assign po01425 = w16289;// level 6
assign po01426 = w16292;// level 6
assign po01427 = w16295;// level 6
assign po01428 = w16298;// level 6
assign po01429 = ~w16303;// level 5
assign po01430 = ~w16307;// level 7
assign po01431 = w16312;// level 8
assign po01432 = ~w16315;// level 7
assign po01433 = w16317;// level 7
assign po01434 = w16319;// level 7
assign po01435 = w16325;// level 7
assign po01436 = ~w16327;// level 5
assign po01437 = ~w16332;// level 8
assign po01438 = w16337;// level 9
assign po01439 = w16340;// level 6
assign po01440 = w16343;// level 6
assign po01441 = w16346;// level 6
assign po01442 = w16349;// level 6
assign po01443 = w16352;// level 6
assign po01444 = w16355;// level 6
assign po01445 = w16358;// level 6
assign po01446 = w16361;// level 6
assign po01447 = w16364;// level 6
assign po01448 = w16367;// level 6
assign po01449 = w16370;// level 6
assign po01450 = w16373;// level 6
assign po01451 = w16376;// level 6
assign po01452 = w16379;// level 6
assign po01453 = w16382;// level 6
assign po01454 = w16385;// level 6
assign po01455 = w16388;// level 6
assign po01456 = w16391;// level 6
assign po01457 = w16394;// level 6
assign po01458 = w16397;// level 6
assign po01459 = w16400;// level 6
assign po01460 = w16403;// level 6
assign po01461 = w16406;// level 6
assign po01462 = ~w16411;// level 7
assign po01463 = ~w16414;// level 6
assign po01464 = ~w16417;// level 6
assign po01465 = ~w16420;// level 6
assign po01466 = ~w16423;// level 6
assign po01467 = ~w16426;// level 6
assign po01468 = ~w16429;// level 6
assign po01469 = ~w16432;// level 6
assign po01470 = ~w16435;// level 6
assign po01471 = ~w16438;// level 6
assign po01472 = ~w16441;// level 6
assign po01473 = ~w16444;// level 6
assign po01474 = w16447;// level 6
assign po01475 = w16450;// level 6
assign po01476 = w16453;// level 6
assign po01477 = w16456;// level 6
assign po01478 = w16459;// level 6
assign po01479 = w16462;// level 6
assign po01480 = w16465;// level 6
assign po01481 = w16468;// level 6
assign po01482 = w16471;// level 6
assign po01483 = w16474;// level 6
assign po01484 = w16477;// level 6
assign po01485 = w16480;// level 6
assign po01486 = w16483;// level 6
assign po01487 = w16486;// level 6
assign po01488 = w16489;// level 6
assign po01489 = w16492;// level 6
assign po01490 = w16495;// level 6
assign po01491 = w16498;// level 6
assign po01492 = w16501;// level 6
assign po01493 = w16504;// level 6
assign po01494 = w16507;// level 6
assign po01495 = w16510;// level 6
assign po01496 = w16513;// level 6
assign po01497 = w16516;// level 6
assign po01498 = w16519;// level 6
assign po01499 = w16522;// level 6
assign po01500 = w16525;// level 6
assign po01501 = w16528;// level 6
assign po01502 = w16531;// level 6
assign po01503 = w16534;// level 6
assign po01504 = w16537;// level 6
assign po01505 = w16540;// level 6
assign po01506 = w16543;// level 6
assign po01507 = w16546;// level 6
assign po01508 = w16549;// level 6
assign po01509 = w16552;// level 6
assign po01510 = w16555;// level 6
assign po01511 = w16558;// level 6
assign po01512 = w16561;// level 6
assign po01513 = w16564;// level 6
assign po01514 = w16567;// level 6
assign po01515 = w16570;// level 6
assign po01516 = w16573;// level 6
assign po01517 = w16576;// level 6
assign po01518 = w16579;// level 6
assign po01519 = w16582;// level 6
assign po01520 = w16585;// level 6
assign po01521 = w16588;// level 6
assign po01522 = w16591;// level 6
assign po01523 = w16594;// level 6
assign po01524 = w16597;// level 6
assign po01525 = w16600;// level 6
assign po01526 = w16603;// level 6
assign po01527 = w16606;// level 6
assign po01528 = w16609;// level 6
assign po01529 = w16612;// level 6
assign po01530 = w16615;// level 6
assign po01531 = w16618;// level 6
assign po01532 = w16621;// level 6
assign po01533 = w16624;// level 6
assign po01534 = w16627;// level 6
assign po01535 = w16630;// level 6
assign po01536 = w16633;// level 6
assign po01537 = w16636;// level 6
assign po01538 = w16639;// level 6
assign po01539 = w16642;// level 6
assign po01540 = w16645;// level 6
assign po01541 = w16648;// level 6
assign po01542 = w16651;// level 6
assign po01543 = w16654;// level 6
assign po01544 = w16657;// level 6
assign po01545 = w16660;// level 6
assign po01546 = w16663;// level 6
assign po01547 = w16666;// level 6
assign po01548 = w16669;// level 6
assign po01549 = w16672;// level 6
assign po01550 = w16675;// level 6
assign po01551 = w16678;// level 6
assign po01552 = w16681;// level 6
assign po01553 = w16684;// level 6
assign po01554 = w16687;// level 6
assign po01555 = w16690;// level 6
assign po01556 = w16693;// level 6
assign po01557 = w16696;// level 6
assign po01558 = w16699;// level 6
assign po01559 = w16702;// level 6
assign po01560 = w16705;// level 6
assign po01561 = w16708;// level 6
assign po01562 = w16711;// level 6
assign po01563 = w16714;// level 6
assign po01564 = w16717;// level 6
assign po01565 = w16720;// level 6
assign po01566 = w16723;// level 6
assign po01567 = w16726;// level 6
assign po01568 = w16729;// level 6
assign po01569 = w16732;// level 6
assign po01570 = w16735;// level 6
assign po01571 = w16738;// level 6
assign po01572 = w16741;// level 6
assign po01573 = w16744;// level 6
assign po01574 = w16747;// level 6
assign po01575 = ~w16763;// level 8
assign po01576 = w16770;// level 8
assign po01577 = ~w16774;// level 6
assign po01578 = w16799;// level 8
assign po01579 = w16803;// level 8
assign po01580 = w16806;// level 7
assign po01581 = w16810;// level 7
assign po01582 = ~w16813;// level 6
assign po01583 = ~w16816;// level 6
assign po01584 = ~w16819;// level 6
assign po01585 = ~w16822;// level 6
assign po01586 = ~w16825;// level 6
assign po01587 = ~w16828;// level 6
assign po01588 = ~w16831;// level 6
assign po01589 = w16838;// level 8
assign po01590 = ~w16841;// level 6
assign po01591 = ~w16844;// level 6
assign po01592 = ~w16847;// level 6
assign po01593 = ~w16850;// level 6
assign po01594 = ~w16853;// level 6
assign po01595 = ~w16856;// level 6
assign po01596 = ~w16859;// level 6
assign po01597 = ~w16862;// level 6
assign po01598 = ~w16865;// level 6
assign po01599 = ~w16868;// level 6
assign po01600 = ~w16871;// level 6
assign po01601 = ~w16874;// level 6
assign po01602 = ~w16877;// level 6
assign po01603 = ~w16883;// level 6
assign po01604 = ~w16886;// level 6
assign po01605 = w16889;// level 7
assign po01606 = pi09932;// level 0
assign po01607 = pi10020;// level 0
assign po01608 = ~w16903;// level 7
assign po01609 = ~w16916;// level 7
assign po01610 = ~w16926;// level 7
assign po01611 = ~w16935;// level 7
assign po01612 = ~w16945;// level 7
assign po01613 = ~w16952;// level 7
assign po01614 = ~w16958;// level 7
assign po01615 = ~w16965;// level 7
assign po01616 = ~w16975;// level 7
assign po01617 = ~w16982;// level 7
assign po01618 = ~w16990;// level 7
assign po01619 = ~w16998;// level 7
assign po01620 = ~w17003;// level 7
assign po01621 = ~w17010;// level 7
assign po01622 = ~w17015;// level 7
assign po01623 = ~w17022;// level 7
assign po01624 = ~w17027;// level 7
assign po01625 = ~w17032;// level 7
assign po01626 = ~w17035;// level 7
assign po01627 = ~w17043;// level 7
assign po01628 = ~w17046;// level 7
assign po01629 = ~w17051;// level 7
assign po01630 = ~w17057;// level 7
assign po01631 = ~w17064;// level 7
assign po01632 = w17070;// level 7
assign po01633 = ~w17074;// level 7
assign po01634 = ~w17077;// level 7
assign po01635 = ~w17082;// level 7
assign po01636 = ~w17088;// level 7
assign po01637 = ~w17091;// level 7
assign po01638 = ~w17094;// level 7
assign po01639 = ~w17097;// level 7
assign po01640 = ~w17102;// level 7
assign po01641 = ~w17107;// level 7
assign po01642 = ~w17112;// level 7
assign po01643 = ~w17118;// level 7
assign po01644 = ~w17123;// level 7
assign po01645 = ~w17130;// level 7
assign po01646 = ~w17135;// level 7
assign po01647 = ~w17141;// level 7
assign po01648 = ~w17144;// level 7
assign po01649 = ~w17147;// level 7
assign po01650 = ~w17152;// level 7
assign po01651 = ~w17157;// level 7
assign po01652 = ~w17161;// level 7
assign po01653 = ~w17166;// level 7
assign po01654 = ~w17171;// level 7
assign po01655 = ~w17176;// level 7
assign po01656 = ~w17181;// level 7
assign po01657 = ~w17188;// level 7
assign po01658 = ~w17195;// level 7
assign po01659 = ~w17199;// level 7
assign po01660 = ~w17204;// level 7
assign po01661 = ~w17209;// level 7
assign po01662 = ~w17214;// level 7
assign po01663 = ~w17217;// level 7
assign po01664 = ~w17222;// level 7
assign po01665 = ~w17225;// level 7
assign po01666 = ~w17230;// level 7
assign po01667 = ~w17235;// level 7
assign po01668 = ~w17238;// level 7
assign po01669 = ~w17243;// level 7
assign po01670 = ~w17248;// level 7
assign po01671 = ~w17253;// level 7
assign po01672 = ~w17258;// level 7
assign po01673 = ~w17263;// level 7
assign po01674 = ~w17268;// level 7
assign po01675 = ~w17272;// level 7
assign po01676 = ~w17275;// level 7
assign po01677 = ~w17278;// level 7
assign po01678 = ~w17283;// level 7
assign po01679 = ~w17288;// level 7
assign po01680 = ~w17293;// level 7
assign po01681 = ~w17296;// level 7
assign po01682 = ~w17299;// level 7
assign po01683 = ~w17304;// level 7
assign po01684 = ~w17309;// level 7
assign po01685 = ~w17313;// level 7
assign po01686 = ~w17319;// level 7
assign po01687 = ~w17324;// level 7
assign po01688 = ~w17329;// level 8
assign po01689 = ~w17333;// level 8
assign po01690 = ~w17338;// level 8
assign po01691 = ~w17343;// level 8
assign po01692 = ~w17348;// level 8
assign po01693 = ~w17353;// level 8
assign po01694 = ~w17357;// level 8
assign po01695 = ~w17360;// level 7
assign po01696 = ~w17365;// level 8
assign po01697 = ~w17370;// level 8
assign po01698 = ~w17373;// level 7
assign po01699 = ~w17379;// level 8
assign po01700 = ~w17384;// level 8
assign po01701 = ~w17389;// level 8
assign po01702 = ~w17394;// level 8
assign po01703 = ~w17397;// level 7
assign po01704 = ~w17402;// level 8
assign po01705 = ~w17405;// level 7
assign po01706 = ~w17410;// level 8
assign po01707 = ~w17415;// level 8
assign po01708 = ~w17420;// level 8
assign po01709 = ~w17424;// level 8
assign po01710 = ~w17427;// level 7
assign po01711 = ~w17432;// level 8
assign po01712 = ~w17435;// level 8
assign po01713 = ~w17441;// level 8
assign po01714 = ~w17444;// level 8
assign po01715 = ~w17449;// level 8
assign po01716 = ~w17454;// level 8
assign po01717 = ~w17457;// level 8
assign po01718 = ~w17460;// level 8
assign po01719 = ~w17465;// level 8
assign po01720 = ~w17470;// level 8
assign po01721 = ~w17473;// level 8
assign po01722 = ~w17478;// level 8
assign po01723 = ~w17483;// level 8
assign po01724 = ~w17486;// level 8
assign po01725 = ~w17489;// level 8
assign po01726 = ~w17494;// level 8
assign po01727 = ~w17499;// level 8
assign po01728 = ~w17504;// level 8
assign po01729 = ~w17509;// level 8
assign po01730 = ~w17515;// level 8
assign po01731 = ~w17520;// level 8
assign po01732 = ~w761;// level 8
assign po01733 = ~w17525;// level 8
assign po01734 = ~w17530;// level 8
assign po01735 = ~w17534;// level 8
assign po01736 = ~w17539;// level 8
assign po01737 = ~w17544;// level 8
assign po01738 = ~w17547;// level 8
assign po01739 = ~w17551;// level 8
assign po01740 = ~w17555;// level 8
assign po01741 = ~w17560;// level 8
assign po01742 = ~w17564;// level 8
assign po01743 = ~w17569;// level 8
assign po01744 = ~w17572;// level 8
assign po01745 = ~w17577;// level 8
assign po01746 = ~w17581;// level 8
assign po01747 = ~w17588;// level 8
assign po01748 = ~w17591;// level 8
assign po01749 = ~w17596;// level 8
assign po01750 = ~w17599;// level 7
assign po01751 = ~w17605;// level 8
assign po01752 = ~w17608;// level 8
assign po01753 = ~w17613;// level 8
assign po01754 = ~w17618;// level 8
assign po01755 = ~w17622;// level 8
assign po01756 = ~w17625;// level 8
assign po01757 = ~w17630;// level 8
assign po01758 = ~w17635;// level 8
assign po01759 = ~w17640;// level 8
assign po01760 = ~w17645;// level 8
assign po01761 = ~w17649;// level 8
assign po01762 = ~w17654;// level 8
assign po01763 = ~w17657;// level 7
assign po01764 = ~w17662;// level 8
assign po01765 = ~w17667;// level 8
assign po01766 = ~w17673;// level 8
assign po01767 = ~w17677;// level 8
assign po01768 = ~w17680;// level 8
assign po01769 = ~w17685;// level 8
assign po01770 = ~w17690;// level 8
assign po01771 = ~w17693;// level 8
assign po01772 = ~w17698;// level 8
assign po01773 = ~w17701;// level 8
assign po01774 = ~w17705;// level 8
assign po01775 = ~w17709;// level 8
assign po01776 = ~w17714;// level 8
assign po01777 = ~w17717;// level 8
assign po01778 = ~w17722;// level 8
assign po01779 = ~w17725;// level 8
assign po01780 = ~w17729;// level 8
assign po01781 = ~w17733;// level 8
assign po01782 = ~w17738;// level 8
assign po01783 = ~w17744;// level 8
assign po01784 = ~w17748;// level 8
assign po01785 = ~w17753;// level 8
assign po01786 = ~w17758;// level 8
assign po01787 = ~w17761;// level 8
assign po01788 = ~w17766;// level 8
assign po01789 = ~w17771;// level 8
assign po01790 = ~w17774;// level 8
assign po01791 = ~w17779;// level 8
assign po01792 = ~w17783;// level 8
assign po01793 = ~w17786;// level 8
assign po01794 = ~w17789;// level 8
assign po01795 = ~w17793;// level 8
assign po01796 = ~w17797;// level 8
assign po01797 = ~w17801;// level 8
assign po01798 = ~w17804;// level 7
assign po01799 = ~w17807;// level 8
assign po01800 = ~w17813;// level 8
assign po01801 = ~w17818;// level 8
assign po01802 = ~w17821;// level 8
assign po01803 = ~w17826;// level 8
assign po01804 = ~w17830;// level 8
assign po01805 = ~w17833;// level 7
assign po01806 = ~w17836;// level 8
assign po01807 = ~w17841;// level 8
assign po01808 = ~w17844;// level 8
assign po01809 = ~w17847;// level 8
assign po01810 = ~w17851;// level 8
assign po01811 = ~w17854;// level 8
assign po01812 = ~w17859;// level 8
assign po01813 = ~w17862;// level 8
assign po01814 = ~w17865;// level 8
assign po01815 = ~w17869;// level 8
assign po01816 = ~w17872;// level 8
assign po01817 = ~w17876;// level 8
assign po01818 = ~w17879;// level 8
assign po01819 = ~w17882;// level 8
assign po01820 = ~w17885;// level 8
assign po01821 = ~w17888;// level 8
assign po01822 = ~w17892;// level 8
assign po01823 = ~w17895;// level 8
assign po01824 = ~w17899;// level 8
assign po01825 = ~w17903;// level 8
assign po01826 = ~w17906;// level 8
assign po01827 = ~w17911;// level 8
assign po01828 = ~w17916;// level 8
assign po01829 = ~w17921;// level 8
assign po01830 = ~w17927;// level 8
assign po01831 = ~w17931;// level 8
assign po01832 = ~w17934;// level 8
assign po01833 = ~w17937;// level 8
assign po01834 = ~w17942;// level 8
assign po01835 = ~w17945;// level 7
assign po01836 = ~w17949;// level 8
assign po01837 = ~w17953;// level 8
assign po01838 = ~w17957;// level 8
assign po01839 = ~w17960;// level 8
assign po01840 = ~w17964;// level 8
assign po01841 = ~w17969;// level 8
assign po01842 = ~w17972;// level 8
assign po01843 = ~w17976;// level 8
assign po01844 = ~w17981;// level 8
assign po01845 = ~w17984;// level 8
assign po01846 = ~w17987;// level 8
assign po01847 = ~w17991;// level 8
assign po01848 = ~w17995;// level 8
assign po01849 = ~w18000;// level 8
assign po01850 = ~w18005;// level 8
assign po01851 = ~w18008;// level 8
assign po01852 = ~w18013;// level 8
assign po01853 = ~w18017;// level 8
assign po01854 = ~w18021;// level 8
assign po01855 = ~w18026;// level 8
assign po01856 = ~w18031;// level 8
assign po01857 = ~w18036;// level 8
assign po01858 = ~w18039;// level 8
assign po01859 = ~w18044;// level 8
assign po01860 = ~w18047;// level 8
assign po01861 = ~w18050;// level 8
assign po01862 = ~w18055;// level 8
assign po01863 = ~w18061;// level 8
assign po01864 = ~w18065;// level 8
assign po01865 = ~w18069;// level 8
assign po01866 = ~w18074;// level 8
assign po01867 = ~w18078;// level 8
assign po01868 = ~w18082;// level 8
assign po01869 = ~w18085;// level 8
assign po01870 = ~w18089;// level 8
assign po01871 = ~w18094;// level 8
assign po01872 = ~w18097;// level 8
assign po01873 = ~w18100;// level 8
assign po01874 = ~w18104;// level 8
assign po01875 = ~w18108;// level 8
assign po01876 = ~w18111;// level 8
assign po01877 = ~w18115;// level 8
assign po01878 = ~w18120;// level 8
assign po01879 = ~w18123;// level 8
assign po01880 = ~w18126;// level 8
assign po01881 = ~w18130;// level 8
assign po01882 = ~w18133;// level 8
assign po01883 = ~w18137;// level 8
assign po01884 = ~w18141;// level 8
assign po01885 = ~w18145;// level 8
assign po01886 = ~w18150;// level 8
assign po01887 = ~w18154;// level 8
assign po01888 = ~w18159;// level 8
assign po01889 = ~w18163;// level 8
assign po01890 = ~w18167;// level 8
assign po01891 = ~w18170;// level 8
assign po01892 = ~w18173;// level 8
assign po01893 = ~w18176;// level 8
assign po01894 = ~w18181;// level 8
assign po01895 = ~w18185;// level 8
assign po01896 = ~w18190;// level 8
assign po01897 = ~w18193;// level 8
assign po01898 = ~w18197;// level 8
assign po01899 = ~w18200;// level 8
assign po01900 = ~w18203;// level 8
assign po01901 = ~w18206;// level 8
assign po01902 = ~w18209;// level 8
assign po01903 = ~w18213;// level 8
assign po01904 = ~w18216;// level 8
assign po01905 = ~w18221;// level 8
assign po01906 = ~w18225;// level 8
assign po01907 = ~w18228;// level 8
assign po01908 = ~w18232;// level 8
assign po01909 = ~w18236;// level 8
assign po01910 = ~w18239;// level 8
assign po01911 = ~w18242;// level 8
assign po01912 = ~w18246;// level 8
assign po01913 = ~w18251;// level 8
assign po01914 = ~w18255;// level 8
assign po01915 = ~w18259;// level 8
assign po01916 = ~w18262;// level 8
assign po01917 = ~w18267;// level 8
assign po01918 = ~w18270;// level 8
assign po01919 = ~w18274;// level 8
assign po01920 = ~w18277;// level 7
assign po01921 = ~w18282;// level 8
assign po01922 = ~w18286;// level 8
assign po01923 = ~w18290;// level 8
assign po01924 = ~w18295;// level 8
assign po01925 = ~w18299;// level 8
assign po01926 = ~w18304;// level 8
assign po01927 = ~w18307;// level 8
assign po01928 = ~w18312;// level 8
assign po01929 = ~w18315;// level 8
assign po01930 = ~w18318;// level 8
assign po01931 = ~w18322;// level 8
assign po01932 = ~w18325;// level 8
assign po01933 = ~w18329;// level 8
assign po01934 = ~w18333;// level 8
assign po01935 = ~w18336;// level 8
assign po01936 = ~w18340;// level 8
assign po01937 = ~w18343;// level 8
assign po01938 = ~w18347;// level 8
assign po01939 = ~w18352;// level 8
assign po01940 = ~w18355;// level 8
assign po01941 = ~w18358;// level 7
assign po01942 = ~w18361;// level 8
assign po01943 = ~w18366;// level 8
assign po01944 = ~w18369;// level 7
assign po01945 = ~w18374;// level 8
assign po01946 = ~w18377;// level 8
assign po01947 = ~w18381;// level 8
assign po01948 = ~w18385;// level 8
assign po01949 = ~w18388;// level 8
assign po01950 = ~w18392;// level 8
assign po01951 = ~w18396;// level 8
assign po01952 = ~w18399;// level 8
assign po01953 = ~w18403;// level 8
assign po01954 = ~w18407;// level 8
assign po01955 = ~w18410;// level 8
assign po01956 = ~w18414;// level 8
assign po01957 = ~w18417;// level 8
assign po01958 = ~w18421;// level 8
assign po01959 = ~w18426;// level 8
assign po01960 = ~w18430;// level 8
assign po01961 = ~w18435;// level 8
assign po01962 = ~w18438;// level 8
assign po01963 = ~w18442;// level 8
assign po01964 = ~w18445;// level 8
assign po01965 = ~w18448;// level 8
assign po01966 = ~w18453;// level 8
assign po01967 = ~w18458;// level 8
assign po01968 = ~w18461;// level 8
assign po01969 = ~w18464;// level 8
assign po01970 = ~w18467;// level 8
assign po01971 = ~w18472;// level 8
assign po01972 = ~w18475;// level 8
assign po01973 = ~w18478;// level 8
assign po01974 = ~w18481;// level 8
assign po01975 = ~w18485;// level 8
assign po01976 = ~w18488;// level 8
assign po01977 = ~w18491;// level 8
assign po01978 = ~w18495;// level 8
assign po01979 = ~w18499;// level 8
assign po01980 = ~w18502;// level 8
assign po01981 = ~w18506;// level 8
assign po01982 = ~w18510;// level 8
assign po01983 = ~w18513;// level 8
assign po01984 = ~w18517;// level 8
assign po01985 = ~w18521;// level 8
assign po01986 = ~w18525;// level 8
assign po01987 = ~w18530;// level 8
assign po01988 = ~w18534;// level 8
assign po01989 = ~w18538;// level 8
assign po01990 = ~w18541;// level 7
assign po01991 = ~w18546;// level 8
assign po01992 = ~w18550;// level 8
assign po01993 = ~w18553;// level 8
assign po01994 = ~w18558;// level 8
assign po01995 = ~w18562;// level 8
assign po01996 = ~w18567;// level 8
assign po01997 = ~w18571;// level 8
assign po01998 = ~w18576;// level 8
assign po01999 = ~w18580;// level 8
assign po02000 = ~w18584;// level 8
assign po02001 = ~w18589;// level 8
assign po02002 = ~w18593;// level 8
assign po02003 = ~w18596;// level 7
assign po02004 = ~w18600;// level 8
assign po02005 = ~w18604;// level 8
assign po02006 = ~w18608;// level 8
assign po02007 = ~w18611;// level 8
assign po02008 = ~w18616;// level 8
assign po02009 = ~w18621;// level 8
assign po02010 = ~w18626;// level 8
assign po02011 = ~w18630;// level 8
assign po02012 = ~w18635;// level 8
assign po02013 = ~w18640;// level 8
assign po02014 = ~w18644;// level 8
assign po02015 = ~w18649;// level 8
assign po02016 = ~w18652;// level 8
assign po02017 = ~w18655;// level 8
assign po02018 = ~w18658;// level 8
assign po02019 = ~w18661;// level 8
assign po02020 = ~w18666;// level 8
assign po02021 = ~w18670;// level 8
assign po02022 = ~w18674;// level 8
assign po02023 = ~w18678;// level 8
assign po02024 = ~w18682;// level 8
assign po02025 = ~w18687;// level 8
assign po02026 = ~w18691;// level 8
assign po02027 = ~w18695;// level 8
assign po02028 = ~w18699;// level 8
assign po02029 = ~w18702;// level 8
assign po02030 = ~w18706;// level 8
assign po02031 = ~w18709;// level 8
assign po02032 = ~w18713;// level 8
assign po02033 = ~w18717;// level 8
assign po02034 = ~w18721;// level 8
assign po02035 = ~w18725;// level 8
assign po02036 = ~w18730;// level 8
assign po02037 = ~w18735;// level 8
assign po02038 = ~w18739;// level 8
assign po02039 = ~w18744;// level 8
assign po02040 = ~w18749;// level 8
assign po02041 = ~w18752;// level 8
assign po02042 = ~w18756;// level 8
assign po02043 = ~w18760;// level 8
assign po02044 = ~w18764;// level 8
assign po02045 = ~w18768;// level 8
assign po02046 = ~w18771;// level 8
assign po02047 = ~w18776;// level 8
assign po02048 = ~w18780;// level 8
assign po02049 = ~w18785;// level 8
assign po02050 = ~w18789;// level 8
assign po02051 = ~w18793;// level 8
assign po02052 = ~w18797;// level 8
assign po02053 = ~w18800;// level 8
assign po02054 = ~w18803;// level 8
assign po02055 = ~w18807;// level 8
assign po02056 = ~w18812;// level 8
assign po02057 = ~w18817;// level 8
assign po02058 = ~w18821;// level 8
assign po02059 = ~w18826;// level 8
assign po02060 = ~w18830;// level 8
assign po02061 = ~w18835;// level 8
assign po02062 = ~w18838;// level 8
assign po02063 = ~w18841;// level 8
assign po02064 = ~w18844;// level 8
assign po02065 = ~w18847;// level 8
assign po02066 = ~w18851;// level 8
assign po02067 = ~w18855;// level 8
assign po02068 = ~w18859;// level 8
assign po02069 = ~w18863;// level 8
assign po02070 = ~w18867;// level 8
assign po02071 = ~w18870;// level 8
assign po02072 = ~w18875;// level 8
assign po02073 = ~w18878;// level 8
assign po02074 = ~w18882;// level 8
assign po02075 = ~w18885;// level 8
assign po02076 = ~w18888;// level 8
assign po02077 = ~w18892;// level 8
assign po02078 = ~w18896;// level 8
assign po02079 = ~w18901;// level 8
assign po02080 = ~w18904;// level 8
assign po02081 = ~w18908;// level 8
assign po02082 = ~w18912;// level 8
assign po02083 = ~w18917;// level 8
assign po02084 = ~w18921;// level 8
assign po02085 = ~w18924;// level 8
assign po02086 = ~w18929;// level 8
assign po02087 = ~w18932;// level 8
assign po02088 = ~w18935;// level 8
assign po02089 = ~w18939;// level 8
assign po02090 = ~w18943;// level 8
assign po02091 = ~w18948;// level 8
assign po02092 = ~w18953;// level 8
assign po02093 = ~w18957;// level 8
assign po02094 = ~w18960;// level 8
assign po02095 = ~w18963;// level 8
assign po02096 = ~w18966;// level 8
assign po02097 = ~w18970;// level 8
assign po02098 = ~w18974;// level 8
assign po02099 = ~w18977;// level 8
assign po02100 = ~w18981;// level 8
assign po02101 = ~w18985;// level 8
assign po02102 = ~w18990;// level 8
assign po02103 = ~w18994;// level 8
assign po02104 = ~w18999;// level 8
assign po02105 = ~w19003;// level 8
assign po02106 = ~w19007;// level 8
assign po02107 = ~w19011;// level 8
assign po02108 = ~w19016;// level 8
assign po02109 = ~w19020;// level 8
assign po02110 = ~w19023;// level 8
assign po02111 = ~w19026;// level 8
assign po02112 = ~w19030;// level 8
assign po02113 = ~w19033;// level 8
assign po02114 = ~w19038;// level 8
assign po02115 = ~w19042;// level 8
assign po02116 = ~w19046;// level 8
assign po02117 = ~w19049;// level 8
assign po02118 = ~w19052;// level 8
assign po02119 = ~w19057;// level 8
assign po02120 = ~w19060;// level 8
assign po02121 = ~w19064;// level 8
assign po02122 = ~w19068;// level 8
assign po02123 = ~w19071;// level 8
assign po02124 = ~w19074;// level 8
assign po02125 = ~w19079;// level 8
assign po02126 = ~w19083;// level 8
assign po02127 = ~w19086;// level 8
assign po02128 = ~w19091;// level 8
assign po02129 = ~w19095;// level 8
assign po02130 = ~w19099;// level 8
assign po02131 = ~w19102;// level 8
assign po02132 = ~w19105;// level 8
assign po02133 = ~w19110;// level 8
assign po02134 = ~w19114;// level 8
assign po02135 = ~w19119;// level 8
assign po02136 = ~w19123;// level 8
assign po02137 = ~w19126;// level 8
assign po02138 = ~w19129;// level 8
assign po02139 = ~w19134;// level 8
assign po02140 = ~w19137;// level 8
assign po02141 = ~w19141;// level 8
assign po02142 = ~w19144;// level 8
assign po02143 = ~w19148;// level 8
assign po02144 = ~w19153;// level 8
assign po02145 = ~w19157;// level 8
assign po02146 = ~w19161;// level 8
assign po02147 = ~w19165;// level 8
assign po02148 = ~w19170;// level 8
assign po02149 = ~w19174;// level 8
assign po02150 = ~w19177;// level 8
assign po02151 = ~w19180;// level 8
assign po02152 = ~w19184;// level 8
assign po02153 = ~w19187;// level 8
assign po02154 = ~w19191;// level 8
assign po02155 = ~w19195;// level 8
assign po02156 = ~w19198;// level 8
assign po02157 = ~w19201;// level 8
assign po02158 = ~w19205;// level 8
assign po02159 = ~w19209;// level 8
assign po02160 = ~w19213;// level 8
assign po02161 = ~w19216;// level 8
assign po02162 = ~w19220;// level 8
assign po02163 = ~w19223;// level 8
assign po02164 = ~w19227;// level 8
assign po02165 = ~w19231;// level 8
assign po02166 = ~w19234;// level 8
assign po02167 = ~w19237;// level 8
assign po02168 = ~w19241;// level 8
assign po02169 = ~w19245;// level 8
assign po02170 = ~w19248;// level 8
assign po02171 = ~w19252;// level 8
assign po02172 = ~w19256;// level 8
assign po02173 = ~w19259;// level 8
assign po02174 = ~w19262;// level 8
assign po02175 = ~w19265;// level 8
assign po02176 = ~w19270;// level 8
assign po02177 = ~w19275;// level 8
assign po02178 = ~w19278;// level 8
assign po02179 = ~w19281;// level 8
assign po02180 = ~w19286;// level 8
assign po02181 = ~w19290;// level 8
assign po02182 = ~w19294;// level 8
assign po02183 = ~w19297;// level 8
assign po02184 = ~w19301;// level 8
assign po02185 = ~w19305;// level 8
assign po02186 = ~w19310;// level 8
assign po02187 = ~w19314;// level 8
assign po02188 = ~w19318;// level 8
assign po02189 = ~w19322;// level 8
assign po02190 = ~w19326;// level 8
assign po02191 = ~w19331;// level 8
assign po02192 = ~w19334;// level 8
assign po02193 = ~w19338;// level 8
assign po02194 = ~w19342;// level 8
assign po02195 = ~w19347;// level 8
assign po02196 = ~w19352;// level 8
assign po02197 = ~w19355;// level 8
assign po02198 = ~w19358;// level 8
assign po02199 = ~w19362;// level 8
assign po02200 = ~w19367;// level 8
assign po02201 = ~w19370;// level 8
assign po02202 = ~w19373;// level 8
assign po02203 = ~w19378;// level 8
assign po02204 = ~w19383;// level 8
assign po02205 = ~w19387;// level 8
assign po02206 = ~w19391;// level 8
assign po02207 = ~w19394;// level 8
assign po02208 = ~w19398;// level 8
assign po02209 = ~w19401;// level 8
assign po02210 = ~w19405;// level 8
assign po02211 = ~w19409;// level 8
assign po02212 = ~w19412;// level 8
assign po02213 = ~w19415;// level 8
assign po02214 = ~w19419;// level 8
assign po02215 = ~w19424;// level 8
assign po02216 = ~w19427;// level 8
assign po02217 = ~w19431;// level 8
assign po02218 = ~w19434;// level 8
assign po02219 = ~w19439;// level 8
assign po02220 = ~w19443;// level 8
assign po02221 = ~w19448;// level 8
assign po02222 = ~w19451;// level 8
assign po02223 = ~w19454;// level 8
assign po02224 = ~w19458;// level 8
assign po02225 = ~w19463;// level 8
assign po02226 = ~w19466;// level 8
assign po02227 = ~w19469;// level 8
assign po02228 = ~w19472;// level 8
assign po02229 = ~w19475;// level 8
assign po02230 = ~w19479;// level 8
assign po02231 = ~w19484;// level 8
assign po02232 = ~w19488;// level 8
assign po02233 = ~w19491;// level 8
assign po02234 = ~w19496;// level 8
assign po02235 = ~w19500;// level 8
assign po02236 = ~w19504;// level 8
assign po02237 = ~w19507;// level 8
assign po02238 = ~w19511;// level 8
assign po02239 = ~w19514;// level 8
assign po02240 = ~w19517;// level 8
assign po02241 = ~w19522;// level 8
assign po02242 = ~w19526;// level 8
assign po02243 = ~w19529;// level 8
assign po02244 = ~w19534;// level 8
assign po02245 = ~w19537;// level 8
assign po02246 = ~w19540;// level 8
assign po02247 = ~w19544;// level 8
assign po02248 = ~w19548;// level 8
assign po02249 = ~w19551;// level 6
assign po02250 = ~w19556;// level 8
assign po02251 = ~w19560;// level 8
assign po02252 = ~w19565;// level 8
assign po02253 = ~w19568;// level 8
assign po02254 = ~w19571;// level 8
assign po02255 = ~w19575;// level 8
assign po02256 = ~w19580;// level 8
assign po02257 = ~w19583;// level 8
assign po02258 = ~w19587;// level 8
assign po02259 = ~w19590;// level 8
assign po02260 = ~w19595;// level 8
assign po02261 = ~w19600;// level 8
assign po02262 = ~w19605;// level 8
assign po02263 = ~w19610;// level 8
assign po02264 = ~w19614;// level 8
assign po02265 = ~w19617;// level 8
assign po02266 = ~w19620;// level 8
assign po02267 = ~w19623;// level 8
assign po02268 = ~w19628;// level 8
assign po02269 = ~w19633;// level 8
assign po02270 = ~w19637;// level 8
assign po02271 = ~w19641;// level 8
assign po02272 = ~w19644;// level 8
assign po02273 = ~w19649;// level 8
assign po02274 = ~w19654;// level 8
assign po02275 = ~w19659;// level 8
assign po02276 = ~w19664;// level 8
assign po02277 = ~w19668;// level 8
assign po02278 = ~w19671;// level 8
assign po02279 = ~w19674;// level 8
assign po02280 = ~w19678;// level 8
assign po02281 = ~w19683;// level 8
assign po02282 = ~w19686;// level 8
assign po02283 = w19689;// level 9
assign po02284 = ~w19693;// level 8
assign po02285 = ~w19697;// level 8
assign po02286 = ~w19719;// level 9
assign po02287 = ~w19722;// level 8
assign po02288 = ~w19727;// level 8
assign po02289 = ~w19732;// level 8
assign po02290 = ~w19739;// level 9
assign po02291 = ~w19744;// level 8
assign po02292 = ~w19747;// level 8
assign po02293 = ~w19754;// level 9
assign po02294 = ~w19758;// level 8
assign po02295 = ~w19765;// level 9
assign po02296 = ~w19772;// level 9
assign po02297 = ~w19776;// level 8
assign po02298 = ~w19779;// level 8
assign po02299 = ~w19782;// level 8
assign po02300 = ~w19786;// level 8
assign po02301 = ~w19790;// level 8
assign po02302 = ~w19794;// level 8
assign po02303 = ~w19799;// level 8
assign po02304 = ~w19806;// level 9
assign po02305 = ~w19810;// level 8
assign po02306 = ~w19817;// level 9
assign po02307 = ~w19822;// level 8
assign po02308 = ~w19825;// level 8
assign po02309 = ~w19830;// level 8
assign po02310 = ~w19834;// level 8
assign po02311 = ~w19837;// level 8
assign po02312 = ~w19842;// level 8
assign po02313 = ~w19845;// level 8
assign po02314 = ~w19848;// level 8
assign po02315 = w19851;// level 6
assign po02316 = ~w19856;// level 8
assign po02317 = w19859;// level 6
assign po02318 = ~w19863;// level 8
assign po02319 = w19866;// level 6
assign po02320 = w19869;// level 7
assign po02321 = ~w19872;// level 8
assign po02322 = ~w19875;// level 8
assign po02323 = ~w19879;// level 8
assign po02324 = ~w19883;// level 8
assign po02325 = ~w19887;// level 8
assign po02326 = ~w19891;// level 8
assign po02327 = w19894;// level 7
assign po02328 = ~w19898;// level 8
assign po02329 = ~w19902;// level 8
assign po02330 = ~w19905;// level 8
assign po02331 = ~w19908;// level 8
assign po02332 = ~w19913;// level 8
assign po02333 = ~w19917;// level 8
assign po02334 = ~w19921;// level 8
assign po02335 = ~w19925;// level 8
assign po02336 = ~w19929;// level 8
assign po02337 = ~w19934;// level 8
assign po02338 = ~w19937;// level 8
assign po02339 = ~w19940;// level 8
assign po02340 = ~w19945;// level 8
assign po02341 = ~w19949;// level 8
assign po02342 = w19952;// level 7
assign po02343 = w19955;// level 7
assign po02344 = ~w19958;// level 8
assign po02345 = ~w19962;// level 8
assign po02346 = ~w19966;// level 8
assign po02347 = ~w19970;// level 8
assign po02348 = ~w19973;// level 8
assign po02349 = ~w19977;// level 8
assign po02350 = ~w19981;// level 8
assign po02351 = ~w19984;// level 8
assign po02352 = w19987;// level 7
assign po02353 = ~w19992;// level 8
assign po02354 = w19995;// level 7
assign po02355 = ~w19999;// level 8
assign po02356 = ~w20003;// level 8
assign po02357 = ~w20006;// level 8
assign po02358 = ~w20010;// level 8
assign po02359 = ~w20013;// level 8
assign po02360 = ~w20018;// level 8
assign po02361 = w20021;// level 7
assign po02362 = ~w20024;// level 8
assign po02363 = ~w20027;// level 8
assign po02364 = ~w20030;// level 7
assign po02365 = ~w20033;// level 8
assign po02366 = ~w20037;// level 8
assign po02367 = ~w20041;// level 8
assign po02368 = ~w20044;// level 8
assign po02369 = ~w20048;// level 8
assign po02370 = ~w20051;// level 8
assign po02371 = ~w20055;// level 8
assign po02372 = ~w20058;// level 7
assign po02373 = ~w20063;// level 8
assign po02374 = ~w20067;// level 8
assign po02375 = ~w20071;// level 8
assign po02376 = ~w20074;// level 7
assign po02377 = ~w20079;// level 8
assign po02378 = ~w20083;// level 8
assign po02379 = ~w20086;// level 7
assign po02380 = ~w20089;// level 8
assign po02381 = ~w20093;// level 8
assign po02382 = ~w20096;// level 7
assign po02383 = ~w20100;// level 8
assign po02384 = ~w20103;// level 8
assign po02385 = ~w20107;// level 8
assign po02386 = ~w20110;// level 8
assign po02387 = ~w20114;// level 8
assign po02388 = ~w20118;// level 8
assign po02389 = ~w20123;// level 8
assign po02390 = ~w20126;// level 8
assign po02391 = ~w20129;// level 8
assign po02392 = ~w20132;// level 8
assign po02393 = ~w20135;// level 8
assign po02394 = ~w20139;// level 8
assign po02395 = ~w20143;// level 8
assign po02396 = ~w20146;// level 8
assign po02397 = ~w20150;// level 8
assign po02398 = ~w20154;// level 8
assign po02399 = ~w20158;// level 8
assign po02400 = ~w20161;// level 8
assign po02401 = ~w20165;// level 8
assign po02402 = ~w20169;// level 8
assign po02403 = ~w20174;// level 8
assign po02404 = ~w20177;// level 8
assign po02405 = ~w20180;// level 8
assign po02406 = ~w20184;// level 8
assign po02407 = ~w20188;// level 8
assign po02408 = ~w20192;// level 8
assign po02409 = ~w20196;// level 8
assign po02410 = ~w20199;// level 8
assign po02411 = ~w20203;// level 8
assign po02412 = ~w20207;// level 8
assign po02413 = ~w20211;// level 8
assign po02414 = ~w20214;// level 8
assign po02415 = ~w20218;// level 8
assign po02416 = ~w20221;// level 8
assign po02417 = ~w20225;// level 8
assign po02418 = ~w20229;// level 8
assign po02419 = ~w20233;// level 8
assign po02420 = ~w20236;// level 8
assign po02421 = ~w20240;// level 8
assign po02422 = ~w20243;// level 8
assign po02423 = ~w20248;// level 8
assign po02424 = ~w20252;// level 8
assign po02425 = ~w20256;// level 8
assign po02426 = ~w20260;// level 8
assign po02427 = ~w20264;// level 8
assign po02428 = ~w20268;// level 8
assign po02429 = ~w20272;// level 8
assign po02430 = ~w20276;// level 8
assign po02431 = ~w20280;// level 8
assign po02432 = ~w20284;// level 8
assign po02433 = ~w20288;// level 8
assign po02434 = ~w20291;// level 8
assign po02435 = ~w20295;// level 8
assign po02436 = ~w20298;// level 8
assign po02437 = ~w20302;// level 8
assign po02438 = ~w20305;// level 8
assign po02439 = ~w20309;// level 8
assign po02440 = ~w20313;// level 8
assign po02441 = ~w20317;// level 8
assign po02442 = ~w20321;// level 8
assign po02443 = ~w20325;// level 8
assign po02444 = ~w20329;// level 8
assign po02445 = ~w20333;// level 8
assign po02446 = ~w20336;// level 8
assign po02447 = ~w20340;// level 8
assign po02448 = ~w20343;// level 8
assign po02449 = ~w20346;// level 8
assign po02450 = ~w20349;// level 8
assign po02451 = ~w20352;// level 8
assign po02452 = ~w20356;// level 8
assign po02453 = ~w20359;// level 8
assign po02454 = ~w20362;// level 8
assign po02455 = ~w20365;// level 8
assign po02456 = ~w20369;// level 8
assign po02457 = ~w20373;// level 8
assign po02458 = ~w20376;// level 8
assign po02459 = ~w20379;// level 8
assign po02460 = ~w20382;// level 8
assign po02461 = ~w20385;// level 8
assign po02462 = ~w20389;// level 8
assign po02463 = ~w20393;// level 8
assign po02464 = ~w20397;// level 8
assign po02465 = ~w20400;// level 8
assign po02466 = ~w20403;// level 8
assign po02467 = ~w20406;// level 6
assign po02468 = ~w20410;// level 8
assign po02469 = ~w20414;// level 8
assign po02470 = ~w20418;// level 8
assign po02471 = ~w20421;// level 8
assign po02472 = ~w20424;// level 8
assign po02473 = ~w20428;// level 8
assign po02474 = ~w20438;// level 8
assign po02475 = ~w20441;// level 8
assign po02476 = ~w20445;// level 8
assign po02477 = ~w20449;// level 8
assign po02478 = ~w20453;// level 8
assign po02479 = ~w20456;// level 8
assign po02480 = ~w20460;// level 8
assign po02481 = ~w20464;// level 8
assign po02482 = ~w20469;// level 8
assign po02483 = ~w20474;// level 8
assign po02484 = ~w20477;// level 8
assign po02485 = ~w20481;// level 8
assign po02486 = ~w20484;// level 8
assign po02487 = ~w20488;// level 8
assign po02488 = ~w20492;// level 8
assign po02489 = ~w20496;// level 8
assign po02490 = ~w20500;// level 8
assign po02491 = ~w20504;// level 8
assign po02492 = ~w20508;// level 8
assign po02493 = ~w20511;// level 8
assign po02494 = ~w20515;// level 8
assign po02495 = ~w20518;// level 8
assign po02496 = ~w20522;// level 8
assign po02497 = ~w20526;// level 8
assign po02498 = ~w20530;// level 8
assign po02499 = ~w20534;// level 8
assign po02500 = ~w20537;// level 8
assign po02501 = ~w20541;// level 8
assign po02502 = ~w20544;// level 8
assign po02503 = ~w20548;// level 8
assign po02504 = ~w20552;// level 8
assign po02505 = ~w20556;// level 8
assign po02506 = ~w20560;// level 8
assign po02507 = ~w20565;// level 8
assign po02508 = ~w20570;// level 8
assign po02509 = ~w20573;// level 8
assign po02510 = ~w20577;// level 8
assign po02511 = ~w20580;// level 8
assign po02512 = ~w20584;// level 8
assign po02513 = ~w20587;// level 8
assign po02514 = ~w20591;// level 8
assign po02515 = ~w20595;// level 8
assign po02516 = ~w20599;// level 8
assign po02517 = ~w20603;// level 8
assign po02518 = ~w20607;// level 8
assign po02519 = ~w20610;// level 8
assign po02520 = ~w20613;// level 8
assign po02521 = ~w20616;// level 8
assign po02522 = ~w20620;// level 8
assign po02523 = ~w20624;// level 8
assign po02524 = ~w20628;// level 8
assign po02525 = ~w20632;// level 8
assign po02526 = ~w20636;// level 8
assign po02527 = ~w20640;// level 8
assign po02528 = ~w20643;// level 8
assign po02529 = ~w20646;// level 8
assign po02530 = ~w20650;// level 8
assign po02531 = ~w20653;// level 8
assign po02532 = ~w20656;// level 8
assign po02533 = ~w20659;// level 8
assign po02534 = ~w20663;// level 8
assign po02535 = ~w20667;// level 8
assign po02536 = ~w20670;// level 8
assign po02537 = ~w20673;// level 8
assign po02538 = ~w20676;// level 8
assign po02539 = ~w20679;// level 8
assign po02540 = ~w20683;// level 8
assign po02541 = ~w20687;// level 8
assign po02542 = ~w20690;// level 8
assign po02543 = ~w20693;// level 8
assign po02544 = ~w20697;// level 8
assign po02545 = ~w20701;// level 8
assign po02546 = ~w20705;// level 8
assign po02547 = ~w20709;// level 8
assign po02548 = ~w20712;// level 8
assign po02549 = ~w20716;// level 8
assign po02550 = ~w20719;// level 8
assign po02551 = ~w20724;// level 8
assign po02552 = ~w20727;// level 8
assign po02553 = ~w20730;// level 7
assign po02554 = ~w20734;// level 8
assign po02555 = ~w20738;// level 8
assign po02556 = ~w20742;// level 8
assign po02557 = ~w20746;// level 8
assign po02558 = ~w20750;// level 8
assign po02559 = ~w20754;// level 8
assign po02560 = ~w20757;// level 8
assign po02561 = ~w20761;// level 8
assign po02562 = ~w20764;// level 8
assign po02563 = ~w20767;// level 8
assign po02564 = ~w20770;// level 8
assign po02565 = ~w20774;// level 8
assign po02566 = ~w20779;// level 8
assign po02567 = ~w20783;// level 8
assign po02568 = ~w20786;// level 8
assign po02569 = ~w20790;// level 8
assign po02570 = ~w20794;// level 8
assign po02571 = ~w20798;// level 8
assign po02572 = ~w20802;// level 8
assign po02573 = ~w20805;// level 8
assign po02574 = ~w20809;// level 8
assign po02575 = ~w20813;// level 8
assign po02576 = ~w20816;// level 8
assign po02577 = ~w20820;// level 8
assign po02578 = ~w20824;// level 8
assign po02579 = ~w20828;// level 8
assign po02580 = ~w20831;// level 8
assign po02581 = ~w20834;// level 8
assign po02582 = ~w20838;// level 8
assign po02583 = ~w20842;// level 8
assign po02584 = ~w20846;// level 8
assign po02585 = ~w20849;// level 8
assign po02586 = ~w20852;// level 8
assign po02587 = ~w20855;// level 8
assign po02588 = ~w20859;// level 8
assign po02589 = ~w20863;// level 8
assign po02590 = ~w20866;// level 8
assign po02591 = ~w20870;// level 8
assign po02592 = ~w20874;// level 8
assign po02593 = ~w20878;// level 8
assign po02594 = ~w20882;// level 8
assign po02595 = ~w20886;// level 8
assign po02596 = ~w20890;// level 8
assign po02597 = ~w20894;// level 8
assign po02598 = ~w20898;// level 8
assign po02599 = ~w20901;// level 8
assign po02600 = ~w20905;// level 8
assign po02601 = ~w20909;// level 8
assign po02602 = ~w20912;// level 8
assign po02603 = ~w20915;// level 7
assign po02604 = ~w20918;// level 8
assign po02605 = ~w20922;// level 8
assign po02606 = ~w20927;// level 8
assign po02607 = ~w20931;// level 8
assign po02608 = ~w20935;// level 8
assign po02609 = ~w20938;// level 8
assign po02610 = ~w20942;// level 8
assign po02611 = ~w20945;// level 7
assign po02612 = ~w20949;// level 8
assign po02613 = ~w20952;// level 8
assign po02614 = ~w20956;// level 8
assign po02615 = ~w20959;// level 8
assign po02616 = ~w20962;// level 8
assign po02617 = ~w20965;// level 8
assign po02618 = ~w20969;// level 8
assign po02619 = ~w20973;// level 8
assign po02620 = ~w20977;// level 8
assign po02621 = ~w20980;// level 8
assign po02622 = ~w20984;// level 8
assign po02623 = ~w20987;// level 8
assign po02624 = ~w20991;// level 8
assign po02625 = ~w20995;// level 8
assign po02626 = ~w20999;// level 8
assign po02627 = ~w21003;// level 8
assign po02628 = ~w21007;// level 8
assign po02629 = ~w21010;// level 8
assign po02630 = ~w21014;// level 8
assign po02631 = ~w21017;// level 8
assign po02632 = ~w21021;// level 8
assign po02633 = ~w21025;// level 8
assign po02634 = ~w21029;// level 8
assign po02635 = ~w21033;// level 8
assign po02636 = ~w21036;// level 8
assign po02637 = ~w21040;// level 8
assign po02638 = ~w21044;// level 8
assign po02639 = ~w21048;// level 8
assign po02640 = ~w21051;// level 8
assign po02641 = ~w21055;// level 8
assign po02642 = ~w21059;// level 8
assign po02643 = ~w21063;// level 8
assign po02644 = ~w21066;// level 8
assign po02645 = ~w21069;// level 8
assign po02646 = ~w21073;// level 8
assign po02647 = ~w21076;// level 8
assign po02648 = ~w21079;// level 8
assign po02649 = ~w21083;// level 8
assign po02650 = ~w21087;// level 8
assign po02651 = ~w21091;// level 8
assign po02652 = ~w21094;// level 8
assign po02653 = ~w21098;// level 8
assign po02654 = ~w21101;// level 8
assign po02655 = ~w21104;// level 8
assign po02656 = ~w21108;// level 8
assign po02657 = ~w21111;// level 8
assign po02658 = ~w21114;// level 8
assign po02659 = ~w21118;// level 8
assign po02660 = ~w21121;// level 8
assign po02661 = ~w21125;// level 8
assign po02662 = ~w21128;// level 8
assign po02663 = ~w21131;// level 8
assign po02664 = ~w21134;// level 8
assign po02665 = ~w21138;// level 8
assign po02666 = ~w21141;// level 8
assign po02667 = ~w21145;// level 8
assign po02668 = ~w21149;// level 8
assign po02669 = ~w21153;// level 8
assign po02670 = ~w21158;// level 8
assign po02671 = ~w21161;// level 8
assign po02672 = ~w21165;// level 8
assign po02673 = ~w21169;// level 8
assign po02674 = ~w21173;// level 8
assign po02675 = ~w21176;// level 8
assign po02676 = ~w21180;// level 8
assign po02677 = ~w21184;// level 8
assign po02678 = ~w21188;// level 8
assign po02679 = ~w21191;// level 7
assign po02680 = ~w21195;// level 8
assign po02681 = ~w21198;// level 8
assign po02682 = ~w21201;// level 8
assign po02683 = ~w21205;// level 8
assign po02684 = ~w21208;// level 8
assign po02685 = ~w21212;// level 8
assign po02686 = ~w21215;// level 7
assign po02687 = ~w21219;// level 8
assign po02688 = ~w21223;// level 8
assign po02689 = ~w21227;// level 8
assign po02690 = ~w21231;// level 8
assign po02691 = ~w21235;// level 8
assign po02692 = ~w21238;// level 8
assign po02693 = ~w21242;// level 8
assign po02694 = ~w21245;// level 8
assign po02695 = ~w21249;// level 8
assign po02696 = ~w21253;// level 8
assign po02697 = ~w21257;// level 8
assign po02698 = ~w21261;// level 8
assign po02699 = ~w21265;// level 8
assign po02700 = ~w21269;// level 8
assign po02701 = ~w21273;// level 8
assign po02702 = ~w21276;// level 8
assign po02703 = ~w21280;// level 8
assign po02704 = ~w21284;// level 8
assign po02705 = ~w21288;// level 8
assign po02706 = ~w21292;// level 8
assign po02707 = ~w21296;// level 8
assign po02708 = ~w21299;// level 8
assign po02709 = ~w21302;// level 8
assign po02710 = ~w21306;// level 8
assign po02711 = ~w21310;// level 8
assign po02712 = ~w21314;// level 8
assign po02713 = ~w21317;// level 8
assign po02714 = ~w21321;// level 8
assign po02715 = ~w21325;// level 8
assign po02716 = ~w21329;// level 8
assign po02717 = ~w21333;// level 8
assign po02718 = ~w21336;// level 8
assign po02719 = ~w21340;// level 8
assign po02720 = ~w21344;// level 8
assign po02721 = ~w21348;// level 8
assign po02722 = ~w21351;// level 8
assign po02723 = ~w21355;// level 8
assign po02724 = ~w21359;// level 8
assign po02725 = ~w21363;// level 8
assign po02726 = ~w21366;// level 8
assign po02727 = ~w21370;// level 8
assign po02728 = ~w21373;// level 8
assign po02729 = ~w21377;// level 8
assign po02730 = ~w21381;// level 8
assign po02731 = ~w21384;// level 8
assign po02732 = ~w21388;// level 8
assign po02733 = ~w21391;// level 8
assign po02734 = ~w21395;// level 8
assign po02735 = ~w21398;// level 8
assign po02736 = ~w21402;// level 8
assign po02737 = ~w21406;// level 8
assign po02738 = ~w21410;// level 8
assign po02739 = ~w21414;// level 8
assign po02740 = ~w21417;// level 8
assign po02741 = ~w21421;// level 8
assign po02742 = ~w21424;// level 8
assign po02743 = ~w21428;// level 8
assign po02744 = ~w21431;// level 8
assign po02745 = ~w21435;// level 8
assign po02746 = ~w21439;// level 8
assign po02747 = ~w21442;// level 8
assign po02748 = ~w21446;// level 8
assign po02749 = ~w21449;// level 8
assign po02750 = ~w21452;// level 8
assign po02751 = ~w21455;// level 7
assign po02752 = ~w21459;// level 8
assign po02753 = ~w21463;// level 8
assign po02754 = ~w21466;// level 8
assign po02755 = ~w21470;// level 8
assign po02756 = ~w21473;// level 8
assign po02757 = ~w21476;// level 7
assign po02758 = ~w21480;// level 8
assign po02759 = ~w21483;// level 8
assign po02760 = ~w21487;// level 8
assign po02761 = ~w21491;// level 8
assign po02762 = ~w21495;// level 8
assign po02763 = ~w21499;// level 8
assign po02764 = ~w21503;// level 8
assign po02765 = ~w21506;// level 8
assign po02766 = ~w21509;// level 8
assign po02767 = ~w21513;// level 8
assign po02768 = ~w21516;// level 8
assign po02769 = ~w21520;// level 8
assign po02770 = ~w21523;// level 8
assign po02771 = ~w21526;// level 8
assign po02772 = ~w21530;// level 8
assign po02773 = ~w21533;// level 8
assign po02774 = w21539;// level 8
assign po02775 = ~w21543;// level 8
assign po02776 = ~w21547;// level 8
assign po02777 = ~w21551;// level 8
assign po02778 = ~w21554;// level 8
assign po02779 = ~w21558;// level 8
assign po02780 = ~w21562;// level 8
assign po02781 = ~w21566;// level 8
assign po02782 = w21578;// level 9
assign po02783 = ~w21581;// level 6
assign po02784 = ~w21584;// level 6
assign po02785 = ~w21587;// level 6
assign po02786 = ~w21590;// level 6
assign po02787 = ~w21593;// level 6
assign po02788 = ~w21596;// level 6
assign po02789 = ~w21599;// level 6
assign po02790 = ~w21603;// level 8
assign po02791 = ~w21605;// level 9
assign po02792 = w21609;// level 10
assign po02793 = ~w21613;// level 8
assign po02794 = ~w21616;// level 7
assign po02795 = ~w21619;// level 7
assign po02796 = ~w21622;// level 7
assign po02797 = ~w21625;// level 7
assign po02798 = ~w21628;// level 7
assign po02799 = ~w21631;// level 7
assign po02800 = ~w21634;// level 7
assign po02801 = ~w21637;// level 7
assign po02802 = ~w21640;// level 7
assign po02803 = ~w21643;// level 7
assign po02804 = ~w21646;// level 7
assign po02805 = ~w21649;// level 7
assign po02806 = ~w21652;// level 7
assign po02807 = ~w21655;// level 7
assign po02808 = ~w21658;// level 7
assign po02809 = w21661;// level 7
assign po02810 = w21664;// level 7
assign po02811 = w21667;// level 7
assign po02812 = w21670;// level 7
assign po02813 = w21673;// level 7
assign po02814 = w21676;// level 7
assign po02815 = w21679;// level 7
assign po02816 = w21682;// level 7
assign po02817 = w21685;// level 7
assign po02818 = w21688;// level 6
assign po02819 = ~w21692;// level 8
assign po02820 = w21695;// level 7
assign po02821 = w21698;// level 7
assign po02822 = ~w21705;// level 9
assign po02823 = ~w21712;// level 9
assign po02824 = ~w21719;// level 9
assign po02825 = ~w21726;// level 9
assign po02826 = ~w21733;// level 9
assign po02827 = ~w21740;// level 9
assign po02828 = ~w21747;// level 9
assign po02829 = ~w21754;// level 9
assign po02830 = ~w21761;// level 9
assign po02831 = ~w21768;// level 9
assign po02832 = ~w21775;// level 9
assign po02833 = ~w21782;// level 9
assign po02834 = ~w21789;// level 9
assign po02835 = ~w21796;// level 9
assign po02836 = ~w21803;// level 9
assign po02837 = ~w21810;// level 9
assign po02838 = ~w21817;// level 9
assign po02839 = ~w21824;// level 9
assign po02840 = ~w21831;// level 9
assign po02841 = ~w21838;// level 9
assign po02842 = ~w21845;// level 9
assign po02843 = ~w21852;// level 9
assign po02844 = ~w21859;// level 9
assign po02845 = ~w21866;// level 9
assign po02846 = ~w21873;// level 9
assign po02847 = ~w21880;// level 9
assign po02848 = ~w21887;// level 9
assign po02849 = ~w21894;// level 9
assign po02850 = w21902;// level 10
assign po02851 = w21905;// level 9
assign po02852 = w21908;// level 9
assign po02853 = w21911;// level 9
assign po02854 = w21914;// level 9
assign po02855 = w21917;// level 6
assign po02856 = w21920;// level 9
assign po02857 = ~w21924;// level 8
assign po02858 = ~w21928;// level 8
assign po02859 = ~w21932;// level 8
assign po02860 = ~w21936;// level 8
assign po02861 = ~w21940;// level 8
assign po02862 = ~w21943;// level 8
assign po02863 = ~w21947;// level 8
assign po02864 = ~w21951;// level 8
assign po02865 = ~w21954;// level 8
assign po02866 = ~w21957;// level 8
assign po02867 = ~w21961;// level 8
assign po02868 = ~w21965;// level 8
assign po02869 = ~w21968;// level 8
assign po02870 = ~w21971;// level 8
assign po02871 = ~w21975;// level 8
assign po02872 = ~w21979;// level 8
assign po02873 = ~w21982;// level 8
assign po02874 = ~w21986;// level 8
assign po02875 = ~w21989;// level 8
assign po02876 = ~w21993;// level 8
assign po02877 = ~w21997;// level 8
assign po02878 = ~w22001;// level 8
assign po02879 = ~w22005;// level 8
assign po02880 = ~w22008;// level 8
assign po02881 = ~w22012;// level 8
assign po02882 = ~w22016;// level 8
assign po02883 = ~w22019;// level 8
assign po02884 = ~w22023;// level 8
assign po02885 = ~w22027;// level 8
assign po02886 = ~w22030;// level 8
assign po02887 = ~w22034;// level 8
assign po02888 = ~w22038;// level 8
assign po02889 = ~w22041;// level 8
assign po02890 = ~w22045;// level 8
assign po02891 = ~w22049;// level 8
assign po02892 = ~w22052;// level 8
assign po02893 = ~w22056;// level 8
assign po02894 = ~w22059;// level 8
assign po02895 = ~w22063;// level 8
assign po02896 = ~w22067;// level 8
assign po02897 = ~w22070;// level 8
assign po02898 = ~w22074;// level 8
assign po02899 = ~w22077;// level 8
assign po02900 = ~w22081;// level 8
assign po02901 = ~w22084;// level 8
assign po02902 = ~w22088;// level 8
assign po02903 = ~w22092;// level 8
assign po02904 = ~w22095;// level 8
assign po02905 = ~w22099;// level 8
assign po02906 = ~w22103;// level 8
assign po02907 = ~w22106;// level 8
assign po02908 = ~w22110;// level 8
assign po02909 = ~w22114;// level 8
assign po02910 = ~w22117;// level 8
assign po02911 = w22120;// level 8
assign po02912 = ~w22124;// level 8
assign po02913 = ~w22127;// level 8
assign po02914 = ~w22130;// level 8
assign po02915 = ~w22133;// level 8
assign po02916 = ~w22136;// level 8
assign po02917 = ~w22139;// level 8
assign po02918 = ~w22142;// level 8
assign po02919 = ~w22145;// level 8
assign po02920 = ~w22149;// level 8
assign po02921 = w22152;// level 6
assign po02922 = w22156;// level 7
assign po02923 = ~w22160;// level 7
assign po02924 = ~w22163;// level 7
assign po02925 = ~w22166;// level 7
assign po02926 = ~w22169;// level 7
assign po02927 = ~w22172;// level 7
assign po02928 = ~w22175;// level 7
assign po02929 = ~w22178;// level 7
assign po02930 = ~w22181;// level 7
assign po02931 = ~w22184;// level 8
assign po02932 = ~w22188;// level 8
assign po02933 = ~w22192;// level 8
assign po02934 = ~w22196;// level 8
assign po02935 = ~w22199;// level 8
assign po02936 = w22201;// level 6
assign po02937 = w22203;// level 6
assign po02938 = w22205;// level 6
assign po02939 = ~w22208;// level 8
assign po02940 = ~w22211;// level 8
assign po02941 = ~w22214;// level 8
assign po02942 = ~w22217;// level 8
assign po02943 = ~w22220;// level 8
assign po02944 = ~w22223;// level 8
assign po02945 = ~w22226;// level 8
assign po02946 = ~w22229;// level 8
assign po02947 = ~w22232;// level 8
assign po02948 = ~w22235;// level 8
assign po02949 = ~w22238;// level 7
assign po02950 = ~w22241;// level 8
assign po02951 = ~w22244;// level 7
assign po02952 = ~w22247;// level 7
assign po02953 = ~w22250;// level 7
assign po02954 = ~w22253;// level 7
assign po02955 = ~w22256;// level 7
assign po02956 = ~w22259;// level 7
assign po02957 = ~w22262;// level 7
assign po02958 = ~w22265;// level 7
assign po02959 = ~w22268;// level 7
assign po02960 = ~w22271;// level 7
assign po02961 = ~w22274;// level 7
assign po02962 = ~w22277;// level 7
assign po02963 = ~w22280;// level 7
assign po02964 = ~w22283;// level 8
assign po02965 = ~w22286;// level 7
assign po02966 = ~w22289;// level 7
assign po02967 = ~w22292;// level 8
assign po02968 = ~w22295;// level 7
assign po02969 = ~w22298;// level 7
assign po02970 = ~w22301;// level 7
assign po02971 = ~w22304;// level 7
assign po02972 = ~w22307;// level 8
assign po02973 = ~w22310;// level 7
assign po02974 = ~w22313;// level 7
assign po02975 = ~w22316;// level 7
assign po02976 = ~w22319;// level 7
assign po02977 = ~w22322;// level 7
assign po02978 = ~w22325;// level 7
assign po02979 = ~w22328;// level 7
assign po02980 = ~w22331;// level 7
assign po02981 = ~w22335;// level 8
assign po02982 = ~w22338;// level 8
assign po02983 = ~w22341;// level 8
assign po02984 = ~w22344;// level 8
assign po02985 = ~w22347;// level 8
assign po02986 = ~w22350;// level 8
assign po02987 = ~w22353;// level 8
assign po02988 = ~w22357;// level 8
assign po02989 = ~w22360;// level 8
assign po02990 = ~w22363;// level 8
assign po02991 = ~w22366;// level 8
assign po02992 = ~w22369;// level 8
assign po02993 = ~w22372;// level 8
assign po02994 = ~w22376;// level 8
assign po02995 = ~w22379;// level 8
assign po02996 = ~w22382;// level 8
assign po02997 = ~w22385;// level 8
assign po02998 = ~w22388;// level 8
assign po02999 = ~w22391;// level 8
assign po03000 = ~w22394;// level 8
assign po03001 = ~w22398;// level 8
assign po03002 = ~w22401;// level 8
assign po03003 = ~w22404;// level 8
assign po03004 = ~w22407;// level 8
assign po03005 = ~w22410;// level 8
assign po03006 = ~w22413;// level 8
assign po03007 = ~w22417;// level 8
assign po03008 = ~w22420;// level 8
assign po03009 = ~w22423;// level 8
assign po03010 = ~w22426;// level 8
assign po03011 = ~w22429;// level 8
assign po03012 = ~w22432;// level 8
assign po03013 = ~w22435;// level 8
assign po03014 = ~w22439;// level 8
assign po03015 = ~w22442;// level 8
assign po03016 = ~w22445;// level 8
assign po03017 = ~w22448;// level 8
assign po03018 = ~w22451;// level 8
assign po03019 = ~w22454;// level 8
assign po03020 = ~w22458;// level 8
assign po03021 = ~w22461;// level 8
assign po03022 = ~w22464;// level 8
assign po03023 = ~w22467;// level 8
assign po03024 = ~w22470;// level 8
assign po03025 = ~w22473;// level 8
assign po03026 = ~w22476;// level 8
assign po03027 = ~w22480;// level 8
assign po03028 = ~w22483;// level 8
assign po03029 = ~w22486;// level 8
assign po03030 = ~w22489;// level 8
assign po03031 = ~w22492;// level 8
assign po03032 = ~w22495;// level 8
assign po03033 = ~w22499;// level 8
assign po03034 = ~w22502;// level 8
assign po03035 = ~w22505;// level 8
assign po03036 = ~w22508;// level 8
assign po03037 = ~w22511;// level 8
assign po03038 = ~w22514;// level 8
assign po03039 = ~w22517;// level 8
assign po03040 = ~w22520;// level 8
assign po03041 = ~w22524;// level 8
assign po03042 = ~w22527;// level 8
assign po03043 = ~w22530;// level 8
assign po03044 = ~w22533;// level 8
assign po03045 = ~w22536;// level 8
assign po03046 = ~w22539;// level 8
assign po03047 = ~w22543;// level 8
assign po03048 = ~w22546;// level 8
assign po03049 = ~w22549;// level 8
assign po03050 = ~w22552;// level 8
assign po03051 = ~w22555;// level 8
assign po03052 = ~w22558;// level 8
assign po03053 = ~w22561;// level 8
assign po03054 = ~w22565;// level 8
assign po03055 = ~w22568;// level 8
assign po03056 = ~w22571;// level 8
assign po03057 = ~w22574;// level 8
assign po03058 = ~w22577;// level 8
assign po03059 = ~w22580;// level 8
assign po03060 = ~w22584;// level 8
assign po03061 = ~w22587;// level 8
assign po03062 = ~w22590;// level 8
assign po03063 = ~w22593;// level 8
assign po03064 = ~w22596;// level 8
assign po03065 = ~w22599;// level 8
assign po03066 = ~w22602;// level 8
assign po03067 = ~w22606;// level 8
assign po03068 = ~w22609;// level 8
assign po03069 = ~w22612;// level 8
assign po03070 = ~w22615;// level 8
assign po03071 = ~w22618;// level 8
assign po03072 = ~w22621;// level 8
assign po03073 = ~w22625;// level 8
assign po03074 = ~w22628;// level 8
assign po03075 = ~w22631;// level 8
assign po03076 = ~w22634;// level 8
assign po03077 = ~w22637;// level 8
assign po03078 = ~w22640;// level 8
assign po03079 = ~w22643;// level 8
assign po03080 = ~w22647;// level 8
assign po03081 = ~w22650;// level 8
assign po03082 = ~w22653;// level 8
assign po03083 = ~w22656;// level 8
assign po03084 = ~w22659;// level 8
assign po03085 = ~w22662;// level 8
assign po03086 = ~w22666;// level 8
assign po03087 = ~w22669;// level 8
assign po03088 = ~w22672;// level 8
assign po03089 = ~w22675;// level 8
assign po03090 = ~w22678;// level 8
assign po03091 = ~w22681;// level 8
assign po03092 = ~w22684;// level 8
assign po03093 = ~w22688;// level 8
assign po03094 = ~w22691;// level 8
assign po03095 = ~w22694;// level 8
assign po03096 = ~w22697;// level 8
assign po03097 = ~w22700;// level 8
assign po03098 = ~w22703;// level 8
assign po03099 = ~w22706;// level 8
assign po03100 = ~w22710;// level 8
assign po03101 = ~w22713;// level 8
assign po03102 = ~w22716;// level 8
assign po03103 = ~w22719;// level 8
assign po03104 = ~w22722;// level 8
assign po03105 = ~w22725;// level 8
assign po03106 = ~w22729;// level 8
assign po03107 = ~w22732;// level 8
assign po03108 = ~w22735;// level 8
assign po03109 = ~w22738;// level 8
assign po03110 = ~w22741;// level 8
assign po03111 = ~w22744;// level 8
assign po03112 = ~w22747;// level 8
assign po03113 = ~w22751;// level 8
assign po03114 = ~w22754;// level 8
assign po03115 = ~w22757;// level 8
assign po03116 = ~w22760;// level 8
assign po03117 = ~w22763;// level 8
assign po03118 = ~w22766;// level 8
assign po03119 = ~w22770;// level 8
assign po03120 = ~w22773;// level 8
assign po03121 = ~w22776;// level 8
assign po03122 = ~w22779;// level 8
assign po03123 = ~w22782;// level 8
assign po03124 = ~w22785;// level 8
assign po03125 = ~w22788;// level 8
assign po03126 = ~w22791;// level 8
assign po03127 = ~w22794;// level 8
assign po03128 = ~w22797;// level 8
assign po03129 = ~w22800;// level 8
assign po03130 = ~w22803;// level 8
assign po03131 = ~w22806;// level 8
assign po03132 = ~w22810;// level 8
assign po03133 = ~w22813;// level 8
assign po03134 = ~w22816;// level 8
assign po03135 = ~w22819;// level 8
assign po03136 = ~w22822;// level 8
assign po03137 = ~w22825;// level 8
assign po03138 = ~w22828;// level 8
assign po03139 = ~w22831;// level 8
assign po03140 = ~w22834;// level 8
assign po03141 = ~w22837;// level 8
assign po03142 = ~w22840;// level 8
assign po03143 = ~w22843;// level 8
assign po03144 = ~w22846;// level 8
assign po03145 = ~w22849;// level 8
assign po03146 = ~w22852;// level 8
assign po03147 = ~w22855;// level 8
assign po03148 = ~w22858;// level 8
assign po03149 = ~w22861;// level 8
assign po03150 = ~w22864;// level 8
assign po03151 = ~w22867;// level 8
assign po03152 = ~w22870;// level 8
assign po03153 = ~w22873;// level 8
assign po03154 = ~w22876;// level 8
assign po03155 = ~w22879;// level 8
assign po03156 = ~w22882;// level 8
assign po03157 = ~w22885;// level 8
assign po03158 = ~w22888;// level 8
assign po03159 = ~w22891;// level 8
assign po03160 = ~w22894;// level 8
assign po03161 = ~w22897;// level 8
assign po03162 = ~w22900;// level 8
assign po03163 = ~w22903;// level 8
assign po03164 = ~w22906;// level 8
assign po03165 = ~w22909;// level 8
assign po03166 = ~w22912;// level 8
assign po03167 = ~w22915;// level 8
assign po03168 = ~w22918;// level 8
assign po03169 = ~w22921;// level 8
assign po03170 = ~w22924;// level 8
assign po03171 = ~w22927;// level 8
assign po03172 = ~w22930;// level 8
assign po03173 = ~w22933;// level 8
assign po03174 = ~w22936;// level 8
assign po03175 = ~w22939;// level 8
assign po03176 = ~w22942;// level 8
assign po03177 = ~w22945;// level 8
assign po03178 = ~w22948;// level 8
assign po03179 = ~w22951;// level 8
assign po03180 = ~w22954;// level 8
assign po03181 = ~w22957;// level 8
assign po03182 = ~w22960;// level 8
assign po03183 = ~w22963;// level 8
assign po03184 = ~w22966;// level 8
assign po03185 = ~w22969;// level 8
assign po03186 = ~w22972;// level 8
assign po03187 = ~w22975;// level 8
assign po03188 = ~w22978;// level 8
assign po03189 = ~w22981;// level 8
assign po03190 = ~w22984;// level 8
assign po03191 = ~w22987;// level 8
assign po03192 = ~w22990;// level 8
assign po03193 = ~w22993;// level 8
assign po03194 = ~w22996;// level 8
assign po03195 = ~w22999;// level 8
assign po03196 = ~w23002;// level 8
assign po03197 = ~w23005;// level 8
assign po03198 = ~w23008;// level 8
assign po03199 = ~w23011;// level 8
assign po03200 = ~w23014;// level 8
assign po03201 = ~w23017;// level 8
assign po03202 = ~w23020;// level 8
assign po03203 = ~w23023;// level 8
assign po03204 = ~w23026;// level 8
assign po03205 = ~w23029;// level 8
assign po03206 = ~w23032;// level 8
assign po03207 = ~w23035;// level 8
assign po03208 = ~w23038;// level 8
assign po03209 = ~w23041;// level 8
assign po03210 = ~w23044;// level 8
assign po03211 = ~w23047;// level 8
assign po03212 = ~w23050;// level 8
assign po03213 = ~w23053;// level 8
assign po03214 = ~w23056;// level 8
assign po03215 = ~w23059;// level 8
assign po03216 = ~w23062;// level 8
assign po03217 = ~w23065;// level 8
assign po03218 = ~w23068;// level 8
assign po03219 = ~w23071;// level 8
assign po03220 = ~w23074;// level 8
assign po03221 = ~w23077;// level 8
assign po03222 = ~w23080;// level 8
assign po03223 = ~w23083;// level 8
assign po03224 = ~w23086;// level 8
assign po03225 = ~w23089;// level 8
assign po03226 = ~w23092;// level 8
assign po03227 = ~w23095;// level 8
assign po03228 = ~w23098;// level 8
assign po03229 = ~w23101;// level 8
assign po03230 = ~w23104;// level 8
assign po03231 = ~w23107;// level 8
assign po03232 = ~w23110;// level 8
assign po03233 = ~w23113;// level 8
assign po03234 = ~w23116;// level 8
assign po03235 = ~w23119;// level 8
assign po03236 = ~w23122;// level 8
assign po03237 = ~w23125;// level 8
assign po03238 = ~w23128;// level 8
assign po03239 = ~w23131;// level 8
assign po03240 = ~w23134;// level 8
assign po03241 = ~w23137;// level 8
assign po03242 = ~w23140;// level 8
assign po03243 = ~w23143;// level 8
assign po03244 = ~w23146;// level 8
assign po03245 = ~w23149;// level 8
assign po03246 = ~w23152;// level 8
assign po03247 = ~w23155;// level 8
assign po03248 = ~w23158;// level 8
assign po03249 = ~w23161;// level 8
assign po03250 = ~w23164;// level 8
assign po03251 = ~w23167;// level 8
assign po03252 = ~w23170;// level 8
assign po03253 = ~w23173;// level 8
assign po03254 = ~w23176;// level 8
assign po03255 = ~w23179;// level 8
assign po03256 = ~w23182;// level 8
assign po03257 = ~w23185;// level 8
assign po03258 = ~w23188;// level 8
assign po03259 = ~w23191;// level 8
assign po03260 = ~w23194;// level 8
assign po03261 = ~w23197;// level 8
assign po03262 = ~w23200;// level 8
assign po03263 = ~w23203;// level 8
assign po03264 = ~w23206;// level 8
assign po03265 = ~w23209;// level 8
assign po03266 = ~w23212;// level 8
assign po03267 = ~w23215;// level 8
assign po03268 = ~w23218;// level 8
assign po03269 = ~w23221;// level 8
assign po03270 = ~w23224;// level 8
assign po03271 = ~w23227;// level 8
assign po03272 = ~w23230;// level 8
assign po03273 = ~w23233;// level 8
assign po03274 = ~w23236;// level 8
assign po03275 = ~w23239;// level 8
assign po03276 = ~w23242;// level 8
assign po03277 = ~w23245;// level 8
assign po03278 = ~w23248;// level 8
assign po03279 = ~w23251;// level 8
assign po03280 = ~w23254;// level 8
assign po03281 = ~w23257;// level 8
assign po03282 = ~w23260;// level 8
assign po03283 = ~w23263;// level 8
assign po03284 = ~w23266;// level 8
assign po03285 = ~w23269;// level 8
assign po03286 = ~w23272;// level 8
assign po03287 = ~w23275;// level 8
assign po03288 = ~w23278;// level 8
assign po03289 = ~w23281;// level 8
assign po03290 = ~w23284;// level 8
assign po03291 = ~w23287;// level 8
assign po03292 = ~w23290;// level 8
assign po03293 = ~w23293;// level 8
assign po03294 = ~w23296;// level 8
assign po03295 = ~w23299;// level 8
assign po03296 = ~w23302;// level 8
assign po03297 = ~w23305;// level 8
assign po03298 = ~w23308;// level 8
assign po03299 = ~w23311;// level 8
assign po03300 = ~w23314;// level 8
assign po03301 = ~w23317;// level 8
assign po03302 = ~w23320;// level 8
assign po03303 = ~w23323;// level 8
assign po03304 = ~w23326;// level 8
assign po03305 = ~w23329;// level 8
assign po03306 = ~w23332;// level 8
assign po03307 = ~w23335;// level 8
assign po03308 = ~w23338;// level 8
assign po03309 = ~w23341;// level 8
assign po03310 = ~w23344;// level 8
assign po03311 = ~w23347;// level 8
assign po03312 = ~w23350;// level 8
assign po03313 = ~w23353;// level 8
assign po03314 = ~w23356;// level 8
assign po03315 = ~w23359;// level 8
assign po03316 = ~w23362;// level 8
assign po03317 = ~w23365;// level 8
assign po03318 = ~w23368;// level 8
assign po03319 = ~w23371;// level 8
assign po03320 = ~w23374;// level 8
assign po03321 = ~w23377;// level 8
assign po03322 = ~w23380;// level 8
assign po03323 = ~w23383;// level 8
assign po03324 = ~w23386;// level 8
assign po03325 = ~w23389;// level 8
assign po03326 = ~w23392;// level 8
assign po03327 = ~w23395;// level 8
assign po03328 = ~w23398;// level 8
assign po03329 = ~w23401;// level 8
assign po03330 = ~w23404;// level 8
assign po03331 = ~w23407;// level 8
assign po03332 = ~w23410;// level 8
assign po03333 = ~w23413;// level 8
assign po03334 = ~w23416;// level 8
assign po03335 = ~w23419;// level 8
assign po03336 = ~w23422;// level 8
assign po03337 = ~w23425;// level 8
assign po03338 = ~w23428;// level 8
assign po03339 = ~w23431;// level 8
assign po03340 = ~w23434;// level 8
assign po03341 = ~w23437;// level 8
assign po03342 = ~w23440;// level 8
assign po03343 = ~w23443;// level 8
assign po03344 = ~w23446;// level 8
assign po03345 = ~w23450;// level 8
assign po03346 = ~w23453;// level 8
assign po03347 = ~w23456;// level 8
assign po03348 = ~w23459;// level 8
assign po03349 = ~w23462;// level 8
assign po03350 = ~w23465;// level 8
assign po03351 = ~w23468;// level 8
assign po03352 = ~w23471;// level 8
assign po03353 = ~w23474;// level 8
assign po03354 = ~w23477;// level 8
assign po03355 = ~w23480;// level 8
assign po03356 = ~w23483;// level 8
assign po03357 = ~w23486;// level 8
assign po03358 = ~w23489;// level 8
assign po03359 = ~w23492;// level 8
assign po03360 = ~w23495;// level 8
assign po03361 = ~w23498;// level 8
assign po03362 = ~w23501;// level 8
assign po03363 = ~w23504;// level 8
assign po03364 = ~w23507;// level 8
assign po03365 = ~w23510;// level 8
assign po03366 = ~w23513;// level 8
assign po03367 = ~w23516;// level 8
assign po03368 = ~w23519;// level 8
assign po03369 = ~w23522;// level 8
assign po03370 = ~w23525;// level 8
assign po03371 = ~w23528;// level 8
assign po03372 = ~w23532;// level 8
assign po03373 = ~w23535;// level 8
assign po03374 = ~w23538;// level 8
assign po03375 = ~w23541;// level 8
assign po03376 = ~w23544;// level 8
assign po03377 = ~w23547;// level 8
assign po03378 = ~w23550;// level 8
assign po03379 = ~w23553;// level 8
assign po03380 = ~w23556;// level 8
assign po03381 = ~w23559;// level 8
assign po03382 = ~w23562;// level 8
assign po03383 = ~w23565;// level 8
assign po03384 = ~w23568;// level 8
assign po03385 = ~w23571;// level 8
assign po03386 = ~w23574;// level 8
assign po03387 = ~w23577;// level 8
assign po03388 = ~w23580;// level 8
assign po03389 = ~w23583;// level 8
assign po03390 = ~w23586;// level 8
assign po03391 = ~w23589;// level 8
assign po03392 = ~w23592;// level 8
assign po03393 = ~w23595;// level 8
assign po03394 = ~w23598;// level 8
assign po03395 = ~w23601;// level 8
assign po03396 = ~w23604;// level 8
assign po03397 = ~w23607;// level 8
assign po03398 = ~w23610;// level 8
assign po03399 = ~w23613;// level 8
assign po03400 = ~w23616;// level 8
assign po03401 = ~w23619;// level 8
assign po03402 = ~w23622;// level 8
assign po03403 = ~w23625;// level 8
assign po03404 = ~w23628;// level 8
assign po03405 = ~w23631;// level 8
assign po03406 = ~w23634;// level 8
assign po03407 = ~w23637;// level 8
assign po03408 = ~w23640;// level 8
assign po03409 = ~w23643;// level 8
assign po03410 = ~w23646;// level 8
assign po03411 = ~w23649;// level 8
assign po03412 = ~w23652;// level 8
assign po03413 = ~w23655;// level 8
assign po03414 = ~w23658;// level 8
assign po03415 = ~w23661;// level 8
assign po03416 = ~w23664;// level 8
assign po03417 = ~w23667;// level 8
assign po03418 = ~w23670;// level 8
assign po03419 = ~w23673;// level 8
assign po03420 = ~w23676;// level 8
assign po03421 = ~w23679;// level 8
assign po03422 = ~w23682;// level 8
assign po03423 = ~w23685;// level 8
assign po03424 = ~w23688;// level 8
assign po03425 = ~w23691;// level 8
assign po03426 = ~w23694;// level 8
assign po03427 = ~w23697;// level 8
assign po03428 = ~w23700;// level 8
assign po03429 = ~w23703;// level 8
assign po03430 = ~w23706;// level 8
assign po03431 = ~w23709;// level 8
assign po03432 = ~w23712;// level 8
assign po03433 = ~w23715;// level 8
assign po03434 = ~w23718;// level 8
assign po03435 = ~w23721;// level 8
assign po03436 = ~w23724;// level 8
assign po03437 = ~w23727;// level 8
assign po03438 = ~w23730;// level 8
assign po03439 = ~w23733;// level 8
assign po03440 = ~w23736;// level 8
assign po03441 = ~w23739;// level 8
assign po03442 = ~w23742;// level 8
assign po03443 = ~w23745;// level 8
assign po03444 = ~w23748;// level 8
assign po03445 = ~w23751;// level 8
assign po03446 = ~w23754;// level 8
assign po03447 = ~w23757;// level 8
assign po03448 = ~w23760;// level 8
assign po03449 = ~w23763;// level 8
assign po03450 = ~w23766;// level 8
assign po03451 = ~w23769;// level 8
assign po03452 = ~w23772;// level 8
assign po03453 = ~w23775;// level 8
assign po03454 = ~w23778;// level 8
assign po03455 = ~w23781;// level 8
assign po03456 = ~w23784;// level 8
assign po03457 = ~w23787;// level 8
assign po03458 = ~w23790;// level 8
assign po03459 = ~w23793;// level 8
assign po03460 = ~w23796;// level 8
assign po03461 = ~w23799;// level 8
assign po03462 = ~w23802;// level 8
assign po03463 = ~w23805;// level 8
assign po03464 = ~w23808;// level 8
assign po03465 = ~w23811;// level 8
assign po03466 = ~w23814;// level 8
assign po03467 = ~w23817;// level 8
assign po03468 = ~w23820;// level 8
assign po03469 = ~w23823;// level 8
assign po03470 = ~w23826;// level 8
assign po03471 = ~w23829;// level 8
assign po03472 = ~w23832;// level 8
assign po03473 = ~w23835;// level 8
assign po03474 = ~w23838;// level 8
assign po03475 = ~w23841;// level 8
assign po03476 = ~w23844;// level 8
assign po03477 = ~w23847;// level 8
assign po03478 = ~w23850;// level 8
assign po03479 = ~w23853;// level 8
assign po03480 = ~w23856;// level 8
assign po03481 = ~w23859;// level 8
assign po03482 = ~w23862;// level 8
assign po03483 = ~w23865;// level 8
assign po03484 = ~w23868;// level 8
assign po03485 = ~w23871;// level 8
assign po03486 = ~w23874;// level 8
assign po03487 = ~w23877;// level 8
assign po03488 = ~w23880;// level 8
assign po03489 = ~w23883;// level 8
assign po03490 = ~w23886;// level 8
assign po03491 = ~w23889;// level 8
assign po03492 = ~w23892;// level 8
assign po03493 = ~w23895;// level 8
assign po03494 = ~w23898;// level 8
assign po03495 = ~w23901;// level 8
assign po03496 = ~w23904;// level 8
assign po03497 = ~w23907;// level 8
assign po03498 = ~w23910;// level 8
assign po03499 = ~w23913;// level 8
assign po03500 = ~w23916;// level 8
assign po03501 = ~w23919;// level 8
assign po03502 = ~w23922;// level 8
assign po03503 = ~w23925;// level 8
assign po03504 = ~w23928;// level 8
assign po03505 = ~w23931;// level 8
assign po03506 = ~w23934;// level 8
assign po03507 = ~w23937;// level 8
assign po03508 = ~w23940;// level 8
assign po03509 = ~w23943;// level 8
assign po03510 = ~w23946;// level 8
assign po03511 = ~w23949;// level 8
assign po03512 = ~w23952;// level 8
assign po03513 = ~w23955;// level 8
assign po03514 = ~w23958;// level 8
assign po03515 = ~w23961;// level 8
assign po03516 = ~w23964;// level 8
assign po03517 = ~w23967;// level 8
assign po03518 = ~w23970;// level 8
assign po03519 = ~w23973;// level 8
assign po03520 = ~w23976;// level 8
assign po03521 = ~w23979;// level 8
assign po03522 = ~w23982;// level 8
assign po03523 = ~w23985;// level 8
assign po03524 = ~w23988;// level 8
assign po03525 = ~w23991;// level 8
assign po03526 = ~w23994;// level 8
assign po03527 = ~w23997;// level 8
assign po03528 = ~w24000;// level 8
assign po03529 = ~w24003;// level 8
assign po03530 = ~w24007;// level 8
assign po03531 = ~w24010;// level 8
assign po03532 = ~w24013;// level 8
assign po03533 = ~w24016;// level 8
assign po03534 = ~w24019;// level 8
assign po03535 = ~w24022;// level 8
assign po03536 = ~w24025;// level 8
assign po03537 = ~w24028;// level 8
assign po03538 = ~w24031;// level 8
assign po03539 = ~w24034;// level 8
assign po03540 = ~w24037;// level 8
assign po03541 = ~w24040;// level 8
assign po03542 = ~w24043;// level 8
assign po03543 = ~w24046;// level 8
assign po03544 = ~w24049;// level 8
assign po03545 = ~w24052;// level 8
assign po03546 = ~w24055;// level 8
assign po03547 = ~w24058;// level 8
assign po03548 = ~w24061;// level 8
assign po03549 = ~w24064;// level 8
assign po03550 = ~w24067;// level 8
assign po03551 = ~w24070;// level 8
assign po03552 = ~w24073;// level 8
assign po03553 = ~w24076;// level 8
assign po03554 = ~w24079;// level 8
assign po03555 = ~w24082;// level 8
assign po03556 = ~w24085;// level 8
assign po03557 = ~w24088;// level 8
assign po03558 = ~w24091;// level 8
assign po03559 = ~w24094;// level 8
assign po03560 = ~w24097;// level 8
assign po03561 = ~w24100;// level 8
assign po03562 = ~w24103;// level 8
assign po03563 = ~w24106;// level 8
assign po03564 = ~w24109;// level 8
assign po03565 = ~w24112;// level 8
assign po03566 = ~w24115;// level 8
assign po03567 = ~w24118;// level 8
assign po03568 = ~w24121;// level 8
assign po03569 = ~w24124;// level 8
assign po03570 = ~w24127;// level 8
assign po03571 = ~w24130;// level 8
assign po03572 = ~w24133;// level 8
assign po03573 = ~w24136;// level 8
assign po03574 = ~w24139;// level 8
assign po03575 = ~w24142;// level 8
assign po03576 = ~w24145;// level 8
assign po03577 = ~w24148;// level 8
assign po03578 = ~w24151;// level 8
assign po03579 = ~w24154;// level 8
assign po03580 = ~w24158;// level 8
assign po03581 = ~w24161;// level 8
assign po03582 = ~w24164;// level 8
assign po03583 = ~w24167;// level 8
assign po03584 = ~w24170;// level 8
assign po03585 = ~w24173;// level 8
assign po03586 = ~w24176;// level 8
assign po03587 = ~w24179;// level 8
assign po03588 = ~w24182;// level 8
assign po03589 = ~w24185;// level 8
assign po03590 = ~w24188;// level 8
assign po03591 = ~w24191;// level 8
assign po03592 = ~w24194;// level 8
assign po03593 = ~w24197;// level 8
assign po03594 = ~w24200;// level 8
assign po03595 = ~w24203;// level 8
assign po03596 = ~w24206;// level 8
assign po03597 = ~w24209;// level 8
assign po03598 = ~w24212;// level 8
assign po03599 = ~w24215;// level 8
assign po03600 = ~w24218;// level 8
assign po03601 = ~w24221;// level 8
assign po03602 = ~w24224;// level 8
assign po03603 = ~w24227;// level 8
assign po03604 = ~w24230;// level 8
assign po03605 = ~w24233;// level 8
assign po03606 = ~w24236;// level 8
assign po03607 = ~w24239;// level 8
assign po03608 = ~w24242;// level 8
assign po03609 = ~w24246;// level 8
assign po03610 = ~w24249;// level 8
assign po03611 = ~w24252;// level 8
assign po03612 = ~w24255;// level 8
assign po03613 = ~w24258;// level 8
assign po03614 = ~w24261;// level 8
assign po03615 = ~w24264;// level 8
assign po03616 = ~w24267;// level 8
assign po03617 = ~w24270;// level 8
assign po03618 = ~w24273;// level 8
assign po03619 = ~w24276;// level 8
assign po03620 = ~w24279;// level 8
assign po03621 = ~w24282;// level 8
assign po03622 = ~w24285;// level 8
assign po03623 = ~w24288;// level 8
assign po03624 = ~w24291;// level 8
assign po03625 = ~w24294;// level 8
assign po03626 = ~w24297;// level 8
assign po03627 = ~w24300;// level 8
assign po03628 = ~w24303;// level 8
assign po03629 = ~w24306;// level 8
assign po03630 = ~w24309;// level 8
assign po03631 = ~w24312;// level 8
assign po03632 = ~w24315;// level 8
assign po03633 = ~w24318;// level 8
assign po03634 = ~w24321;// level 8
assign po03635 = ~w24324;// level 8
assign po03636 = ~w24327;// level 8
assign po03637 = ~w24330;// level 8
assign po03638 = ~w24333;// level 8
assign po03639 = ~w24336;// level 8
assign po03640 = ~w24339;// level 8
assign po03641 = ~w24342;// level 8
assign po03642 = ~w24345;// level 8
assign po03643 = ~w24348;// level 8
assign po03644 = ~w24351;// level 8
assign po03645 = ~w24354;// level 8
assign po03646 = ~w24357;// level 8
assign po03647 = ~w24360;// level 8
assign po03648 = ~w24363;// level 8
assign po03649 = ~w24366;// level 8
assign po03650 = ~w24369;// level 8
assign po03651 = ~w24372;// level 8
assign po03652 = ~w24375;// level 8
assign po03653 = ~w24378;// level 8
assign po03654 = ~w24381;// level 8
assign po03655 = ~w24384;// level 8
assign po03656 = ~w24387;// level 8
assign po03657 = ~w24390;// level 8
assign po03658 = ~w24393;// level 8
assign po03659 = ~w24396;// level 8
assign po03660 = ~w24399;// level 8
assign po03661 = ~w24402;// level 8
assign po03662 = ~w24406;// level 8
assign po03663 = ~w24409;// level 8
assign po03664 = ~w24412;// level 8
assign po03665 = ~w24415;// level 8
assign po03666 = ~w24418;// level 8
assign po03667 = ~w24421;// level 8
assign po03668 = ~w24424;// level 8
assign po03669 = ~w24427;// level 8
assign po03670 = ~w24430;// level 8
assign po03671 = ~w24433;// level 8
assign po03672 = ~w24436;// level 8
assign po03673 = ~w24439;// level 8
assign po03674 = ~w24442;// level 8
assign po03675 = ~w24445;// level 8
assign po03676 = ~w24448;// level 8
assign po03677 = ~w24451;// level 8
assign po03678 = ~w24454;// level 8
assign po03679 = ~w24457;// level 8
assign po03680 = ~w24460;// level 8
assign po03681 = ~w24463;// level 8
assign po03682 = ~w24466;// level 8
assign po03683 = ~w24469;// level 8
assign po03684 = ~w24472;// level 8
assign po03685 = ~w24475;// level 8
assign po03686 = ~w24478;// level 8
assign po03687 = ~w24481;// level 8
assign po03688 = ~w24484;// level 8
assign po03689 = ~w24487;// level 8
assign po03690 = ~w24490;// level 8
assign po03691 = ~w24493;// level 8
assign po03692 = ~w24496;// level 8
assign po03693 = ~w24499;// level 8
assign po03694 = ~w24502;// level 8
assign po03695 = ~w24505;// level 8
assign po03696 = ~w24508;// level 8
assign po03697 = ~w24511;// level 8
assign po03698 = ~w24514;// level 8
assign po03699 = ~w24517;// level 8
assign po03700 = ~w24520;// level 8
assign po03701 = ~w24523;// level 8
assign po03702 = ~w24526;// level 8
assign po03703 = ~w24529;// level 8
assign po03704 = ~w24532;// level 8
assign po03705 = ~w24535;// level 8
assign po03706 = ~w24538;// level 8
assign po03707 = ~w24541;// level 8
assign po03708 = ~w24544;// level 8
assign po03709 = ~w24547;// level 8
assign po03710 = ~w24550;// level 8
assign po03711 = ~w24553;// level 8
assign po03712 = ~w24556;// level 8
assign po03713 = ~w24559;// level 8
assign po03714 = ~w24562;// level 8
assign po03715 = ~w24565;// level 8
assign po03716 = ~w24568;// level 8
assign po03717 = ~w24571;// level 8
assign po03718 = ~w24574;// level 8
assign po03719 = ~w24577;// level 8
assign po03720 = ~w24580;// level 8
assign po03721 = ~w24583;// level 8
assign po03722 = ~w24586;// level 8
assign po03723 = ~w24589;// level 8
assign po03724 = ~w24592;// level 8
assign po03725 = ~w24595;// level 8
assign po03726 = ~w24598;// level 8
assign po03727 = ~w24601;// level 8
assign po03728 = ~w24604;// level 8
assign po03729 = ~w24607;// level 8
assign po03730 = ~w24610;// level 8
assign po03731 = ~w24613;// level 8
assign po03732 = ~w24616;// level 8
assign po03733 = ~w24619;// level 8
assign po03734 = ~w24622;// level 8
assign po03735 = ~w24625;// level 8
assign po03736 = ~w24628;// level 8
assign po03737 = ~w24631;// level 8
assign po03738 = ~w24634;// level 8
assign po03739 = ~w24637;// level 8
assign po03740 = ~w24640;// level 8
assign po03741 = ~w24643;// level 8
assign po03742 = ~w24646;// level 8
assign po03743 = ~w24649;// level 8
assign po03744 = ~w24652;// level 8
assign po03745 = ~w24655;// level 8
assign po03746 = ~w24658;// level 8
assign po03747 = ~w24661;// level 8
assign po03748 = ~w24664;// level 8
assign po03749 = ~w24667;// level 8
assign po03750 = ~w24670;// level 8
assign po03751 = ~w24673;// level 8
assign po03752 = ~w24676;// level 8
assign po03753 = ~w24679;// level 8
assign po03754 = ~w24682;// level 8
assign po03755 = ~w24685;// level 8
assign po03756 = ~w24688;// level 8
assign po03757 = ~w24691;// level 8
assign po03758 = ~w24694;// level 8
assign po03759 = ~w24697;// level 8
assign po03760 = ~w24700;// level 8
assign po03761 = ~w24703;// level 8
assign po03762 = ~w24706;// level 8
assign po03763 = ~w24709;// level 8
assign po03764 = ~w24713;// level 8
assign po03765 = ~w24716;// level 8
assign po03766 = ~w24719;// level 8
assign po03767 = ~w24722;// level 8
assign po03768 = ~w24725;// level 8
assign po03769 = ~w24728;// level 8
assign po03770 = ~w24731;// level 8
assign po03771 = ~w24734;// level 8
assign po03772 = ~w24737;// level 8
assign po03773 = ~w24740;// level 8
assign po03774 = ~w24743;// level 8
assign po03775 = ~w24746;// level 8
assign po03776 = ~w24749;// level 8
assign po03777 = ~w24752;// level 8
assign po03778 = ~w24755;// level 8
assign po03779 = ~w24758;// level 8
assign po03780 = ~w24761;// level 8
assign po03781 = ~w24764;// level 8
assign po03782 = ~w24767;// level 8
assign po03783 = ~w24770;// level 8
assign po03784 = ~w24773;// level 8
assign po03785 = ~w24776;// level 8
assign po03786 = ~w24779;// level 8
assign po03787 = ~w24782;// level 8
assign po03788 = ~w24785;// level 8
assign po03789 = ~w24788;// level 8
assign po03790 = ~w24791;// level 8
assign po03791 = ~w24794;// level 8
assign po03792 = ~w24797;// level 8
assign po03793 = ~w24800;// level 8
assign po03794 = ~w24803;// level 8
assign po03795 = ~w24806;// level 8
assign po03796 = ~w24809;// level 8
assign po03797 = ~w24812;// level 8
assign po03798 = ~w24815;// level 8
assign po03799 = ~w24818;// level 8
assign po03800 = ~w24821;// level 8
assign po03801 = ~w24824;// level 8
assign po03802 = ~w24827;// level 8
assign po03803 = ~w24830;// level 8
assign po03804 = ~w24833;// level 8
assign po03805 = ~w24836;// level 8
assign po03806 = ~w24839;// level 8
assign po03807 = ~w24842;// level 8
assign po03808 = ~w24845;// level 8
assign po03809 = ~w24848;// level 8
assign po03810 = ~w24851;// level 8
assign po03811 = ~w24854;// level 8
assign po03812 = ~w24857;// level 8
assign po03813 = ~w24860;// level 8
assign po03814 = ~w24863;// level 8
assign po03815 = ~w24866;// level 8
assign po03816 = ~w24869;// level 8
assign po03817 = ~w24872;// level 8
assign po03818 = ~w24875;// level 8
assign po03819 = ~w24878;// level 8
assign po03820 = ~w24881;// level 8
assign po03821 = ~w24884;// level 8
assign po03822 = ~w24887;// level 8
assign po03823 = ~w24890;// level 8
assign po03824 = ~w24893;// level 8
assign po03825 = ~w24896;// level 8
assign po03826 = ~w24899;// level 8
assign po03827 = ~w24902;// level 8
assign po03828 = ~w24905;// level 8
assign po03829 = ~w24908;// level 8
assign po03830 = ~w24911;// level 8
assign po03831 = ~w24914;// level 8
assign po03832 = ~w24917;// level 8
assign po03833 = ~w24920;// level 8
assign po03834 = ~w24923;// level 8
assign po03835 = ~w24926;// level 8
assign po03836 = ~w24929;// level 8
assign po03837 = ~w24932;// level 8
assign po03838 = ~w24935;// level 8
assign po03839 = ~w24938;// level 8
assign po03840 = ~w24941;// level 8
assign po03841 = ~w24944;// level 8
assign po03842 = ~w24947;// level 8
assign po03843 = ~w24950;// level 8
assign po03844 = ~w24953;// level 8
assign po03845 = ~w24956;// level 8
assign po03846 = ~w24959;// level 8
assign po03847 = ~w24962;// level 8
assign po03848 = ~w24965;// level 8
assign po03849 = ~w24968;// level 8
assign po03850 = ~w24971;// level 8
assign po03851 = ~w24974;// level 8
assign po03852 = ~w24977;// level 8
assign po03853 = ~w24980;// level 8
assign po03854 = ~w24983;// level 8
assign po03855 = ~w24986;// level 8
assign po03856 = ~w24989;// level 8
assign po03857 = ~w24992;// level 8
assign po03858 = ~w24995;// level 8
assign po03859 = ~w24998;// level 8
assign po03860 = ~w25001;// level 8
assign po03861 = ~w25004;// level 8
assign po03862 = ~w25007;// level 8
assign po03863 = ~w25010;// level 8
assign po03864 = ~w25013;// level 8
assign po03865 = ~w25016;// level 8
assign po03866 = ~w25019;// level 8
assign po03867 = ~w25022;// level 8
assign po03868 = ~w25025;// level 8
assign po03869 = ~w25028;// level 8
assign po03870 = ~w25031;// level 8
assign po03871 = ~w25034;// level 8
assign po03872 = ~w25037;// level 8
assign po03873 = ~w25040;// level 8
assign po03874 = ~w25043;// level 8
assign po03875 = ~w25046;// level 8
assign po03876 = ~w25049;// level 8
assign po03877 = ~w25052;// level 8
assign po03878 = ~w25055;// level 8
assign po03879 = ~w25058;// level 8
assign po03880 = ~w25061;// level 8
assign po03881 = ~w25064;// level 8
assign po03882 = ~w25067;// level 8
assign po03883 = ~w25070;// level 8
assign po03884 = ~w25073;// level 8
assign po03885 = ~w25076;// level 8
assign po03886 = ~w25079;// level 8
assign po03887 = ~w25082;// level 8
assign po03888 = ~w25085;// level 8
assign po03889 = ~w25088;// level 8
assign po03890 = ~w25091;// level 8
assign po03891 = ~w25094;// level 8
assign po03892 = ~w25097;// level 8
assign po03893 = ~w25100;// level 8
assign po03894 = ~w25103;// level 8
assign po03895 = ~w25106;// level 8
assign po03896 = ~w25109;// level 8
assign po03897 = ~w25112;// level 8
assign po03898 = ~w25115;// level 8
assign po03899 = ~w25118;// level 8
assign po03900 = ~w25121;// level 8
assign po03901 = ~w25124;// level 8
assign po03902 = ~w25127;// level 8
assign po03903 = ~w25130;// level 8
assign po03904 = ~w25133;// level 8
assign po03905 = ~w25136;// level 8
assign po03906 = ~w25139;// level 8
assign po03907 = ~w25142;// level 8
assign po03908 = ~w25145;// level 8
assign po03909 = ~w25148;// level 8
assign po03910 = ~w25151;// level 8
assign po03911 = ~w25154;// level 8
assign po03912 = ~w25157;// level 8
assign po03913 = ~w25160;// level 8
assign po03914 = ~w25163;// level 8
assign po03915 = ~w25166;// level 8
assign po03916 = ~w25169;// level 8
assign po03917 = ~w25172;// level 8
assign po03918 = ~w25175;// level 8
assign po03919 = ~w25178;// level 8
assign po03920 = ~w25181;// level 8
assign po03921 = ~w25184;// level 8
assign po03922 = ~w25187;// level 8
assign po03923 = ~w25190;// level 8
assign po03924 = ~w25193;// level 8
assign po03925 = ~w25196;// level 8
assign po03926 = ~w25199;// level 8
assign po03927 = ~w25202;// level 8
assign po03928 = ~w25205;// level 8
assign po03929 = ~w25208;// level 8
assign po03930 = ~w25211;// level 8
assign po03931 = ~w25214;// level 8
assign po03932 = ~w25217;// level 8
assign po03933 = ~w25220;// level 8
assign po03934 = ~w25223;// level 8
assign po03935 = ~w25226;// level 8
assign po03936 = ~w25229;// level 8
assign po03937 = ~w25232;// level 8
assign po03938 = ~w25235;// level 8
assign po03939 = ~w25238;// level 8
assign po03940 = ~w25241;// level 8
assign po03941 = ~w25244;// level 8
assign po03942 = ~w25247;// level 8
assign po03943 = ~w25250;// level 8
assign po03944 = ~w25253;// level 8
assign po03945 = ~w25256;// level 8
assign po03946 = ~w25259;// level 8
assign po03947 = ~w25262;// level 8
assign po03948 = ~w25265;// level 8
assign po03949 = ~w25268;// level 8
assign po03950 = ~w25271;// level 8
assign po03951 = ~w25274;// level 8
assign po03952 = ~w25277;// level 8
assign po03953 = ~w25280;// level 8
assign po03954 = ~w25283;// level 8
assign po03955 = ~w25286;// level 8
assign po03956 = ~w25289;// level 8
assign po03957 = ~w25292;// level 8
assign po03958 = ~w25295;// level 8
assign po03959 = ~w25298;// level 8
assign po03960 = ~w25301;// level 8
assign po03961 = ~w25304;// level 8
assign po03962 = ~w25307;// level 8
assign po03963 = ~w25310;// level 8
assign po03964 = ~w25313;// level 8
assign po03965 = ~w25316;// level 8
assign po03966 = ~w25319;// level 8
assign po03967 = ~w25322;// level 8
assign po03968 = ~w25325;// level 8
assign po03969 = ~w25328;// level 8
assign po03970 = ~w25331;// level 8
assign po03971 = ~w25334;// level 8
assign po03972 = ~w25337;// level 8
assign po03973 = ~w25340;// level 8
assign po03974 = ~w25343;// level 8
assign po03975 = ~w25346;// level 8
assign po03976 = ~w25349;// level 8
assign po03977 = ~w25352;// level 8
assign po03978 = ~w25355;// level 8
assign po03979 = ~w25358;// level 8
assign po03980 = ~w25361;// level 8
assign po03981 = ~w25364;// level 8
assign po03982 = ~w25367;// level 8
assign po03983 = ~w25370;// level 8
assign po03984 = ~w25373;// level 8
assign po03985 = ~w25376;// level 8
assign po03986 = ~w25379;// level 8
assign po03987 = ~w25382;// level 8
assign po03988 = ~w25385;// level 8
assign po03989 = ~w25388;// level 8
assign po03990 = ~w25391;// level 8
assign po03991 = ~w25394;// level 8
assign po03992 = ~w25397;// level 8
assign po03993 = ~w25400;// level 8
assign po03994 = ~w25403;// level 8
assign po03995 = ~w25406;// level 8
assign po03996 = ~w25409;// level 8
assign po03997 = ~w25412;// level 8
assign po03998 = ~w25415;// level 8
assign po03999 = ~w25418;// level 8
assign po04000 = ~w25421;// level 8
assign po04001 = ~w25424;// level 8
assign po04002 = ~w25427;// level 8
assign po04003 = ~w25430;// level 8
assign po04004 = ~w25433;// level 8
assign po04005 = ~w25436;// level 8
assign po04006 = ~w25439;// level 8
assign po04007 = ~w25442;// level 8
assign po04008 = ~w25445;// level 8
assign po04009 = ~w25448;// level 8
assign po04010 = ~w25451;// level 8
assign po04011 = ~w25454;// level 8
assign po04012 = ~w25457;// level 8
assign po04013 = ~w25460;// level 8
assign po04014 = ~w25463;// level 8
assign po04015 = ~w25466;// level 8
assign po04016 = ~w25469;// level 8
assign po04017 = ~w25472;// level 8
assign po04018 = ~w25475;// level 8
assign po04019 = ~w25478;// level 8
assign po04020 = ~w25481;// level 7
assign po04021 = ~w25484;// level 7
assign po04022 = ~w25487;// level 7
assign po04023 = ~w25490;// level 7
assign po04024 = ~w25493;// level 7
assign po04025 = ~w25496;// level 7
assign po04026 = ~w25499;// level 7
assign po04027 = ~w25503;// level 8
assign po04028 = ~w25506;// level 7
assign po04029 = ~w25509;// level 7
assign po04030 = ~w25512;// level 7
assign po04031 = ~w25515;// level 7
assign po04032 = ~w25518;// level 7
assign po04033 = ~w25521;// level 7
assign po04034 = ~w25524;// level 7
assign po04035 = ~w25527;// level 8
assign po04036 = ~w25530;// level 7
assign po04037 = ~w25533;// level 7
assign po04038 = ~w25536;// level 7
assign po04039 = ~w25539;// level 7
assign po04040 = ~w25542;// level 7
assign po04041 = ~w25545;// level 7
assign po04042 = ~w25548;// level 7
assign po04043 = ~w25551;// level 7
assign po04044 = ~w25554;// level 7
assign po04045 = ~w25557;// level 7
assign po04046 = ~w25561;// level 8
assign po04047 = ~w25564;// level 7
assign po04048 = ~w25568;// level 8
assign po04049 = ~w25571;// level 8
assign po04050 = ~w25574;// level 8
assign po04051 = ~w25577;// level 8
assign po04052 = ~w25580;// level 8
assign po04053 = ~w25583;// level 8
assign po04054 = ~w25586;// level 8
assign po04055 = ~w25589;// level 8
assign po04056 = ~w25592;// level 8
assign po04057 = ~w25595;// level 8
assign po04058 = ~w25598;// level 8
assign po04059 = ~w25601;// level 8
assign po04060 = ~w25605;// level 8
assign po04061 = ~w25608;// level 8
assign po04062 = ~w25611;// level 8
assign po04063 = ~w25614;// level 8
assign po04064 = ~w25617;// level 8
assign po04065 = ~w25620;// level 8
assign po04066 = ~w25624;// level 8
assign po04067 = ~w25627;// level 8
assign po04068 = ~w25630;// level 8
assign po04069 = ~w25633;// level 8
assign po04070 = ~w25636;// level 8
assign po04071 = ~w25639;// level 8
assign po04072 = ~w25642;// level 8
assign po04073 = ~w25646;// level 8
assign po04074 = ~w25649;// level 8
assign po04075 = ~w25652;// level 8
assign po04076 = ~w25655;// level 8
assign po04077 = ~w25658;// level 8
assign po04078 = ~w25661;// level 8
assign po04079 = ~w25665;// level 8
assign po04080 = ~w25668;// level 8
assign po04081 = ~w25671;// level 8
assign po04082 = ~w25674;// level 8
assign po04083 = ~w25677;// level 8
assign po04084 = ~w25680;// level 8
assign po04085 = ~w25683;// level 8
assign po04086 = ~w25687;// level 8
assign po04087 = ~w25690;// level 8
assign po04088 = ~w25693;// level 8
assign po04089 = ~w25696;// level 8
assign po04090 = ~w25699;// level 8
assign po04091 = ~w25702;// level 8
assign po04092 = ~w25706;// level 8
assign po04093 = ~w25709;// level 8
assign po04094 = ~w25713;// level 8
assign po04095 = ~w25716;// level 8
assign po04096 = ~w25719;// level 8
assign po04097 = ~w25722;// level 8
assign po04098 = ~w25725;// level 8
assign po04099 = ~w25728;// level 8
assign po04100 = ~w25731;// level 8
assign po04101 = ~w25734;// level 8
assign po04102 = ~w25737;// level 8
assign po04103 = ~w25740;// level 8
assign po04104 = ~w25743;// level 8
assign po04105 = ~w25747;// level 8
assign po04106 = ~w25750;// level 8
assign po04107 = ~w25753;// level 8
assign po04108 = ~w25756;// level 8
assign po04109 = ~w25759;// level 8
assign po04110 = ~w25762;// level 8
assign po04111 = ~w25765;// level 8
assign po04112 = ~w25769;// level 8
assign po04113 = ~w25772;// level 8
assign po04114 = ~w25775;// level 8
assign po04115 = ~w25778;// level 8
assign po04116 = ~w25781;// level 8
assign po04117 = ~w25784;// level 8
assign po04118 = ~w25788;// level 8
assign po04119 = ~w25791;// level 8
assign po04120 = ~w25794;// level 8
assign po04121 = ~w25797;// level 8
assign po04122 = ~w25800;// level 8
assign po04123 = ~w25803;// level 8
assign po04124 = ~w25806;// level 8
assign po04125 = ~w25810;// level 8
assign po04126 = ~w25813;// level 8
assign po04127 = ~w25816;// level 8
assign po04128 = ~w25819;// level 8
assign po04129 = ~w25822;// level 8
assign po04130 = ~w25825;// level 8
assign po04131 = ~w25829;// level 8
assign po04132 = ~w25832;// level 8
assign po04133 = ~w25835;// level 8
assign po04134 = ~w25838;// level 8
assign po04135 = ~w25841;// level 8
assign po04136 = ~w25844;// level 8
assign po04137 = ~w25847;// level 8
assign po04138 = ~w25851;// level 8
assign po04139 = ~w25854;// level 8
assign po04140 = ~w25857;// level 8
assign po04141 = ~w25860;// level 8
assign po04142 = ~w25863;// level 8
assign po04143 = ~w25866;// level 8
assign po04144 = ~w25870;// level 8
assign po04145 = ~w25874;// level 8
assign po04146 = ~w25877;// level 8
assign po04147 = ~w25880;// level 8
assign po04148 = ~w25883;// level 8
assign po04149 = ~w25886;// level 8
assign po04150 = ~w25889;// level 8
assign po04151 = ~w25892;// level 8
assign po04152 = ~w25895;// level 8
assign po04153 = ~w25898;// level 8
assign po04154 = ~w25901;// level 8
assign po04155 = ~w25904;// level 8
assign po04156 = ~w25907;// level 8
assign po04157 = ~w25911;// level 8
assign po04158 = ~w25915;// level 8
assign po04159 = ~w25918;// level 8
assign po04160 = ~w25922;// level 8
assign po04161 = ~w25925;// level 8
assign po04162 = ~w25928;// level 8
assign po04163 = ~w25931;// level 8
assign po04164 = ~w25934;// level 8
assign po04165 = ~w25937;// level 8
assign po04166 = ~w25940;// level 8
assign po04167 = ~w25943;// level 8
assign po04168 = ~w25946;// level 8
assign po04169 = ~w25949;// level 8
assign po04170 = ~w25952;// level 8
assign po04171 = ~w25956;// level 8
assign po04172 = ~w25959;// level 8
assign po04173 = ~w25962;// level 8
assign po04174 = ~w25965;// level 8
assign po04175 = ~w25968;// level 8
assign po04176 = ~w25971;// level 8
assign po04177 = ~w25974;// level 8
assign po04178 = ~w25978;// level 8
assign po04179 = ~w25981;// level 8
assign po04180 = ~w25984;// level 8
assign po04181 = ~w25987;// level 8
assign po04182 = ~w25990;// level 8
assign po04183 = ~w25993;// level 8
assign po04184 = ~w25997;// level 8
assign po04185 = ~w26000;// level 8
assign po04186 = ~w26003;// level 8
assign po04187 = ~w26006;// level 8
assign po04188 = ~w26009;// level 8
assign po04189 = ~w26012;// level 8
assign po04190 = ~w26015;// level 8
assign po04191 = ~w26019;// level 8
assign po04192 = ~w26022;// level 8
assign po04193 = ~w26025;// level 8
assign po04194 = ~w26028;// level 8
assign po04195 = ~w26031;// level 8
assign po04196 = ~w26034;// level 8
assign po04197 = ~w26038;// level 8
assign po04198 = ~w26041;// level 8
assign po04199 = ~w26044;// level 8
assign po04200 = ~w26047;// level 8
assign po04201 = ~w26050;// level 8
assign po04202 = ~w26053;// level 8
assign po04203 = ~w26056;// level 8
assign po04204 = ~w26060;// level 8
assign po04205 = ~w26063;// level 8
assign po04206 = ~w26066;// level 8
assign po04207 = ~w26069;// level 8
assign po04208 = ~w26072;// level 8
assign po04209 = ~w26075;// level 8
assign po04210 = ~w26079;// level 8
assign po04211 = ~w26082;// level 8
assign po04212 = ~w26085;// level 8
assign po04213 = ~w26088;// level 8
assign po04214 = ~w26091;// level 8
assign po04215 = ~w26094;// level 8
assign po04216 = ~w26097;// level 8
assign po04217 = ~w26101;// level 8
assign po04218 = ~w26105;// level 8
assign po04219 = ~w26108;// level 8
assign po04220 = ~w26111;// level 8
assign po04221 = ~w26114;// level 8
assign po04222 = ~w26117;// level 8
assign po04223 = ~w26120;// level 8
assign po04224 = ~w26123;// level 8
assign po04225 = ~w26126;// level 8
assign po04226 = ~w26129;// level 8
assign po04227 = ~w26132;// level 8
assign po04228 = ~w26135;// level 8
assign po04229 = ~w26138;// level 8
assign po04230 = ~w26142;// level 8
assign po04231 = ~w26145;// level 8
assign po04232 = ~w26148;// level 8
assign po04233 = ~w26151;// level 8
assign po04234 = ~w26154;// level 8
assign po04235 = ~w26157;// level 8
assign po04236 = ~w26161;// level 8
assign po04237 = ~w26165;// level 8
assign po04238 = ~w26168;// level 8
assign po04239 = ~w26171;// level 8
assign po04240 = ~w26174;// level 8
assign po04241 = ~w26177;// level 8
assign po04242 = ~w26180;// level 8
assign po04243 = ~w26183;// level 8
assign po04244 = ~w26187;// level 8
assign po04245 = ~w26190;// level 8
assign po04246 = ~w26193;// level 8
assign po04247 = ~w26196;// level 8
assign po04248 = ~w26199;// level 8
assign po04249 = ~w26202;// level 8
assign po04250 = ~w26205;// level 8
assign po04251 = ~w26208;// level 8
assign po04252 = ~w26211;// level 8
assign po04253 = ~w26214;// level 8
assign po04254 = ~w26217;// level 8
assign po04255 = ~w26220;// level 8
assign po04256 = ~w26223;// level 8
assign po04257 = ~w26226;// level 8
assign po04258 = ~w26229;// level 8
assign po04259 = ~w26232;// level 8
assign po04260 = ~w26235;// level 8
assign po04261 = ~w26238;// level 8
assign po04262 = ~w26241;// level 8
assign po04263 = ~w26244;// level 8
assign po04264 = ~w26247;// level 8
assign po04265 = ~w26250;// level 8
assign po04266 = ~w26253;// level 8
assign po04267 = ~w26256;// level 8
assign po04268 = ~w26259;// level 8
assign po04269 = ~w26262;// level 8
assign po04270 = ~w26265;// level 8
assign po04271 = ~w26268;// level 8
assign po04272 = ~w26271;// level 8
assign po04273 = ~w26274;// level 8
assign po04274 = ~w26277;// level 8
assign po04275 = ~w26280;// level 8
assign po04276 = ~w26283;// level 8
assign po04277 = ~w26286;// level 8
assign po04278 = ~w26289;// level 8
assign po04279 = ~w26292;// level 8
assign po04280 = ~w26295;// level 8
assign po04281 = ~w26298;// level 8
assign po04282 = ~w26301;// level 8
assign po04283 = ~w26304;// level 8
assign po04284 = ~w26307;// level 8
assign po04285 = ~w26310;// level 8
assign po04286 = ~w26313;// level 8
assign po04287 = ~w26316;// level 8
assign po04288 = ~w26319;// level 8
assign po04289 = ~w26322;// level 8
assign po04290 = ~w26325;// level 8
assign po04291 = ~w26328;// level 8
assign po04292 = ~w26331;// level 8
assign po04293 = ~w26334;// level 8
assign po04294 = ~w26337;// level 8
assign po04295 = ~w26340;// level 8
assign po04296 = ~w26343;// level 8
assign po04297 = ~w26346;// level 8
assign po04298 = ~w26349;// level 8
assign po04299 = ~w26352;// level 8
assign po04300 = ~w26355;// level 8
assign po04301 = ~w26358;// level 8
assign po04302 = ~w26361;// level 8
assign po04303 = ~w26364;// level 8
assign po04304 = ~w26367;// level 8
assign po04305 = ~w26370;// level 8
assign po04306 = ~w26373;// level 8
assign po04307 = ~w26376;// level 8
assign po04308 = ~w26379;// level 8
assign po04309 = ~w26382;// level 8
assign po04310 = ~w26385;// level 8
assign po04311 = ~w26388;// level 8
assign po04312 = ~w26391;// level 8
assign po04313 = ~w26394;// level 8
assign po04314 = ~w26397;// level 8
assign po04315 = ~w26400;// level 8
assign po04316 = ~w26403;// level 8
assign po04317 = ~w26406;// level 8
assign po04318 = ~w26409;// level 8
assign po04319 = ~w26412;// level 8
assign po04320 = ~w26415;// level 8
assign po04321 = ~w26418;// level 8
assign po04322 = ~w26421;// level 8
assign po04323 = ~w26424;// level 8
assign po04324 = ~w26427;// level 8
assign po04325 = ~w26430;// level 8
assign po04326 = ~w26433;// level 8
assign po04327 = ~w26436;// level 8
assign po04328 = ~w26439;// level 8
assign po04329 = ~w26442;// level 8
assign po04330 = ~w26445;// level 8
assign po04331 = ~w26448;// level 8
assign po04332 = ~w26451;// level 8
assign po04333 = ~w26454;// level 8
assign po04334 = ~w26457;// level 8
assign po04335 = ~w26460;// level 8
assign po04336 = ~w26463;// level 8
assign po04337 = ~w26466;// level 8
assign po04338 = ~w26469;// level 8
assign po04339 = ~w26472;// level 8
assign po04340 = ~w26475;// level 8
assign po04341 = ~w26478;// level 8
assign po04342 = ~w26481;// level 8
assign po04343 = ~w26484;// level 8
assign po04344 = ~w26487;// level 8
assign po04345 = ~w26490;// level 8
assign po04346 = ~w26493;// level 8
assign po04347 = ~w26496;// level 8
assign po04348 = ~w26499;// level 8
assign po04349 = ~w26502;// level 8
assign po04350 = ~w26505;// level 8
assign po04351 = ~w26508;// level 8
assign po04352 = ~w26511;// level 8
assign po04353 = ~w26514;// level 8
assign po04354 = ~w26517;// level 8
assign po04355 = ~w26520;// level 8
assign po04356 = ~w26523;// level 8
assign po04357 = ~w26526;// level 8
assign po04358 = ~w26529;// level 8
assign po04359 = ~w26532;// level 8
assign po04360 = ~w26535;// level 8
assign po04361 = ~w26538;// level 8
assign po04362 = ~w26541;// level 8
assign po04363 = ~w26544;// level 8
assign po04364 = ~w26547;// level 8
assign po04365 = ~w26550;// level 8
assign po04366 = ~w26553;// level 8
assign po04367 = ~w26556;// level 8
assign po04368 = ~w26559;// level 8
assign po04369 = ~w26562;// level 8
assign po04370 = ~w26565;// level 8
assign po04371 = ~w26568;// level 8
assign po04372 = ~w26571;// level 8
assign po04373 = ~w26574;// level 8
assign po04374 = ~w26577;// level 8
assign po04375 = ~w26580;// level 8
assign po04376 = ~w26583;// level 8
assign po04377 = ~w26586;// level 8
assign po04378 = ~w26589;// level 8
assign po04379 = ~w26592;// level 8
assign po04380 = ~w26595;// level 8
assign po04381 = ~w26598;// level 8
assign po04382 = ~w26601;// level 8
assign po04383 = ~w26604;// level 8
assign po04384 = ~w26607;// level 8
assign po04385 = ~w26610;// level 8
assign po04386 = ~w26613;// level 8
assign po04387 = ~w26616;// level 8
assign po04388 = ~w26619;// level 8
assign po04389 = ~w26622;// level 8
assign po04390 = ~w26625;// level 8
assign po04391 = ~w26628;// level 8
assign po04392 = ~w26631;// level 8
assign po04393 = ~w26634;// level 8
assign po04394 = ~w26638;// level 8
assign po04395 = ~w26641;// level 8
assign po04396 = ~w26644;// level 8
assign po04397 = ~w26647;// level 8
assign po04398 = ~w26650;// level 8
assign po04399 = ~w26653;// level 8
assign po04400 = ~w26656;// level 8
assign po04401 = ~w26659;// level 8
assign po04402 = ~w26662;// level 8
assign po04403 = ~w26665;// level 8
assign po04404 = ~w26668;// level 8
assign po04405 = ~w26671;// level 8
assign po04406 = ~w26674;// level 8
assign po04407 = ~w26677;// level 8
assign po04408 = ~w26680;// level 8
assign po04409 = ~w26683;// level 8
assign po04410 = ~w26686;// level 8
assign po04411 = ~w26689;// level 8
assign po04412 = ~w26692;// level 8
assign po04413 = ~w26695;// level 8
assign po04414 = ~w26698;// level 8
assign po04415 = ~w26701;// level 8
assign po04416 = ~w26704;// level 8
assign po04417 = ~w26707;// level 8
assign po04418 = ~w26710;// level 8
assign po04419 = ~w26713;// level 8
assign po04420 = ~w26716;// level 8
assign po04421 = ~w26719;// level 8
assign po04422 = ~w26722;// level 8
assign po04423 = ~w26725;// level 8
assign po04424 = ~w26728;// level 8
assign po04425 = ~w26731;// level 8
assign po04426 = ~w26734;// level 8
assign po04427 = ~w26737;// level 8
assign po04428 = ~w26740;// level 8
assign po04429 = ~w26743;// level 8
assign po04430 = ~w26746;// level 8
assign po04431 = ~w26749;// level 8
assign po04432 = ~w26752;// level 8
assign po04433 = ~w26755;// level 8
assign po04434 = ~w26758;// level 8
assign po04435 = ~w26761;// level 8
assign po04436 = ~w26764;// level 8
assign po04437 = ~w26767;// level 8
assign po04438 = ~w26770;// level 8
assign po04439 = ~w26773;// level 8
assign po04440 = ~w26776;// level 8
assign po04441 = ~w26779;// level 8
assign po04442 = ~w26782;// level 8
assign po04443 = ~w26785;// level 8
assign po04444 = ~w26788;// level 8
assign po04445 = ~w26791;// level 8
assign po04446 = ~w26794;// level 8
assign po04447 = ~w26797;// level 8
assign po04448 = ~w26800;// level 8
assign po04449 = ~w26803;// level 8
assign po04450 = ~w26806;// level 8
assign po04451 = ~w26809;// level 8
assign po04452 = ~w26812;// level 8
assign po04453 = ~w26815;// level 8
assign po04454 = ~w26818;// level 8
assign po04455 = ~w26821;// level 8
assign po04456 = ~w26824;// level 8
assign po04457 = ~w26827;// level 8
assign po04458 = ~w26830;// level 8
assign po04459 = ~w26833;// level 8
assign po04460 = ~w26836;// level 8
assign po04461 = ~w26839;// level 8
assign po04462 = ~w26842;// level 8
assign po04463 = ~w26845;// level 8
assign po04464 = ~w26848;// level 8
assign po04465 = ~w26851;// level 8
assign po04466 = ~w26854;// level 8
assign po04467 = ~w26857;// level 8
assign po04468 = ~w26860;// level 8
assign po04469 = ~w26863;// level 8
assign po04470 = ~w26866;// level 8
assign po04471 = ~w26869;// level 8
assign po04472 = ~w26872;// level 8
assign po04473 = ~w26875;// level 8
assign po04474 = ~w26878;// level 8
assign po04475 = ~w26881;// level 8
assign po04476 = ~w26884;// level 8
assign po04477 = ~w26887;// level 8
assign po04478 = ~w26890;// level 8
assign po04479 = ~w26893;// level 8
assign po04480 = ~w26896;// level 8
assign po04481 = ~w26899;// level 8
assign po04482 = ~w26902;// level 8
assign po04483 = ~w26905;// level 8
assign po04484 = ~w26908;// level 8
assign po04485 = ~w26911;// level 8
assign po04486 = ~w26914;// level 8
assign po04487 = ~w26917;// level 8
assign po04488 = ~w26920;// level 8
assign po04489 = ~w26923;// level 8
assign po04490 = ~w26926;// level 8
assign po04491 = ~w26929;// level 8
assign po04492 = ~w26932;// level 8
assign po04493 = ~w26935;// level 8
assign po04494 = ~w26938;// level 8
assign po04495 = ~w26941;// level 8
assign po04496 = ~w26944;// level 8
assign po04497 = ~w26947;// level 8
assign po04498 = ~w26950;// level 8
assign po04499 = ~w26953;// level 8
assign po04500 = ~w26956;// level 8
assign po04501 = ~w26959;// level 8
assign po04502 = ~w26962;// level 8
assign po04503 = ~w26965;// level 8
assign po04504 = ~w26968;// level 8
assign po04505 = ~w26971;// level 8
assign po04506 = ~w26974;// level 8
assign po04507 = ~w26977;// level 8
assign po04508 = ~w26980;// level 8
assign po04509 = ~w26983;// level 8
assign po04510 = ~w26986;// level 8
assign po04511 = ~w26989;// level 8
assign po04512 = ~w26992;// level 8
assign po04513 = ~w26995;// level 8
assign po04514 = ~w26998;// level 8
assign po04515 = ~w27001;// level 8
assign po04516 = ~w27004;// level 8
assign po04517 = ~w27007;// level 8
assign po04518 = ~w27010;// level 8
assign po04519 = ~w27013;// level 8
assign po04520 = ~w27016;// level 8
assign po04521 = ~w27019;// level 8
assign po04522 = ~w27022;// level 8
assign po04523 = ~w27025;// level 8
assign po04524 = ~w27028;// level 8
assign po04525 = ~w27031;// level 8
assign po04526 = ~w27034;// level 8
assign po04527 = ~w27037;// level 8
assign po04528 = ~w27041;// level 8
assign po04529 = ~w27044;// level 8
assign po04530 = ~w27047;// level 8
assign po04531 = ~w27050;// level 8
assign po04532 = ~w27053;// level 8
assign po04533 = ~w27056;// level 8
assign po04534 = ~w27059;// level 8
assign po04535 = ~w27062;// level 8
assign po04536 = ~w27065;// level 8
assign po04537 = ~w27068;// level 8
assign po04538 = ~w27071;// level 8
assign po04539 = ~w27074;// level 8
assign po04540 = ~w27077;// level 8
assign po04541 = ~w27080;// level 8
assign po04542 = ~w27083;// level 8
assign po04543 = ~w27086;// level 8
assign po04544 = ~w27089;// level 8
assign po04545 = ~w27092;// level 8
assign po04546 = ~w27095;// level 8
assign po04547 = ~w27098;// level 8
assign po04548 = ~w27101;// level 8
assign po04549 = ~w27104;// level 8
assign po04550 = ~w27107;// level 8
assign po04551 = ~w27110;// level 8
assign po04552 = ~w27113;// level 8
assign po04553 = ~w27116;// level 8
assign po04554 = ~w27119;// level 8
assign po04555 = ~w27122;// level 8
assign po04556 = ~w27125;// level 8
assign po04557 = ~w27128;// level 8
assign po04558 = ~w27131;// level 8
assign po04559 = ~w27134;// level 8
assign po04560 = ~w27137;// level 8
assign po04561 = ~w27140;// level 8
assign po04562 = ~w27143;// level 8
assign po04563 = ~w27146;// level 8
assign po04564 = ~w27149;// level 8
assign po04565 = ~w27152;// level 8
assign po04566 = ~w27155;// level 8
assign po04567 = ~w27158;// level 8
assign po04568 = ~w27161;// level 8
assign po04569 = ~w27164;// level 8
assign po04570 = ~w27167;// level 8
assign po04571 = ~w27170;// level 8
assign po04572 = ~w27173;// level 8
assign po04573 = ~w27176;// level 8
assign po04574 = ~w27179;// level 8
assign po04575 = ~w27182;// level 8
assign po04576 = ~w27185;// level 8
assign po04577 = ~w27188;// level 8
assign po04578 = ~w27191;// level 8
assign po04579 = ~w27194;// level 8
assign po04580 = ~w27197;// level 8
assign po04581 = ~w27200;// level 8
assign po04582 = ~w27203;// level 8
assign po04583 = ~w27206;// level 8
assign po04584 = ~w27209;// level 8
assign po04585 = ~w27212;// level 8
assign po04586 = ~w27215;// level 8
assign po04587 = ~w27218;// level 8
assign po04588 = ~w27221;// level 8
assign po04589 = ~w27224;// level 8
assign po04590 = ~w27227;// level 8
assign po04591 = ~w27230;// level 8
assign po04592 = ~w27233;// level 8
assign po04593 = ~w27236;// level 8
assign po04594 = ~w27239;// level 8
assign po04595 = ~w27242;// level 8
assign po04596 = ~w27245;// level 8
assign po04597 = ~w27248;// level 8
assign po04598 = ~w27251;// level 8
assign po04599 = ~w27254;// level 8
assign po04600 = ~w27257;// level 8
assign po04601 = ~w27260;// level 8
assign po04602 = ~w27263;// level 8
assign po04603 = ~w27266;// level 8
assign po04604 = ~w27269;// level 8
assign po04605 = ~w27272;// level 8
assign po04606 = ~w27275;// level 8
assign po04607 = ~w27278;// level 8
assign po04608 = ~w27281;// level 8
assign po04609 = ~w27284;// level 8
assign po04610 = ~w27287;// level 8
assign po04611 = ~w27290;// level 8
assign po04612 = ~w27293;// level 8
assign po04613 = ~w27296;// level 8
assign po04614 = ~w27299;// level 8
assign po04615 = ~w27302;// level 8
assign po04616 = ~w27305;// level 8
assign po04617 = ~w27308;// level 8
assign po04618 = ~w27311;// level 8
assign po04619 = ~w27314;// level 8
assign po04620 = ~w27317;// level 8
assign po04621 = ~w27320;// level 8
assign po04622 = ~w27323;// level 8
assign po04623 = ~w27326;// level 8
assign po04624 = ~w27329;// level 8
assign po04625 = ~w27332;// level 8
assign po04626 = ~w27335;// level 8
assign po04627 = ~w27338;// level 8
assign po04628 = ~w27341;// level 8
assign po04629 = ~w27344;// level 8
assign po04630 = ~w27347;// level 8
assign po04631 = ~w27350;// level 8
assign po04632 = ~w27353;// level 8
assign po04633 = ~w27356;// level 8
assign po04634 = ~w27359;// level 8
assign po04635 = ~w27362;// level 8
assign po04636 = ~w27365;// level 8
assign po04637 = ~w27368;// level 8
assign po04638 = ~w27371;// level 8
assign po04639 = ~w27374;// level 8
assign po04640 = ~w27377;// level 8
assign po04641 = ~w27380;// level 8
assign po04642 = ~w27383;// level 8
assign po04643 = ~w27386;// level 8
assign po04644 = ~w27389;// level 8
assign po04645 = ~w27392;// level 8
assign po04646 = ~w27395;// level 8
assign po04647 = ~w27398;// level 8
assign po04648 = ~w27401;// level 8
assign po04649 = ~w27404;// level 8
assign po04650 = ~w27407;// level 8
assign po04651 = ~w27410;// level 8
assign po04652 = ~w27413;// level 8
assign po04653 = ~w27416;// level 8
assign po04654 = ~w27419;// level 8
assign po04655 = ~w27422;// level 8
assign po04656 = ~w27425;// level 8
assign po04657 = ~w27428;// level 8
assign po04658 = ~w27431;// level 8
assign po04659 = ~w27435;// level 8
assign po04660 = ~w27438;// level 8
assign po04661 = ~w27441;// level 8
assign po04662 = ~w27444;// level 8
assign po04663 = ~w27447;// level 8
assign po04664 = ~w27450;// level 8
assign po04665 = ~w27453;// level 8
assign po04666 = ~w27456;// level 8
assign po04667 = ~w27459;// level 8
assign po04668 = ~w27462;// level 8
assign po04669 = ~w27465;// level 8
assign po04670 = ~w27468;// level 8
assign po04671 = ~w27471;// level 8
assign po04672 = ~w27474;// level 8
assign po04673 = ~w27477;// level 8
assign po04674 = ~w27480;// level 8
assign po04675 = ~w27483;// level 8
assign po04676 = ~w27486;// level 8
assign po04677 = ~w27489;// level 8
assign po04678 = ~w27492;// level 8
assign po04679 = ~w27495;// level 8
assign po04680 = ~w27498;// level 8
assign po04681 = ~w27501;// level 8
assign po04682 = ~w27504;// level 8
assign po04683 = ~w27507;// level 8
assign po04684 = ~w27510;// level 8
assign po04685 = ~w27513;// level 8
assign po04686 = ~w27516;// level 8
assign po04687 = ~w27519;// level 8
assign po04688 = ~w27522;// level 8
assign po04689 = ~w27525;// level 8
assign po04690 = ~w27528;// level 8
assign po04691 = ~w27531;// level 8
assign po04692 = ~w27534;// level 8
assign po04693 = ~w27537;// level 8
assign po04694 = ~w27540;// level 8
assign po04695 = ~w27543;// level 8
assign po04696 = ~w27546;// level 8
assign po04697 = ~w27549;// level 8
assign po04698 = ~w27552;// level 8
assign po04699 = ~w27555;// level 8
assign po04700 = ~w27558;// level 8
assign po04701 = ~w27561;// level 8
assign po04702 = ~w27564;// level 8
assign po04703 = ~w27567;// level 8
assign po04704 = ~w27570;// level 8
assign po04705 = ~w27573;// level 8
assign po04706 = ~w27576;// level 8
assign po04707 = ~w27579;// level 8
assign po04708 = ~w27582;// level 8
assign po04709 = ~w27585;// level 8
assign po04710 = ~w27588;// level 8
assign po04711 = ~w27591;// level 8
assign po04712 = ~w27594;// level 8
assign po04713 = ~w27598;// level 8
assign po04714 = ~w27601;// level 8
assign po04715 = ~w27604;// level 8
assign po04716 = ~w27607;// level 8
assign po04717 = ~w27610;// level 8
assign po04718 = ~w27613;// level 8
assign po04719 = ~w27616;// level 8
assign po04720 = ~w27619;// level 8
assign po04721 = ~w27622;// level 8
assign po04722 = ~w27625;// level 8
assign po04723 = ~w27628;// level 8
assign po04724 = ~w27631;// level 8
assign po04725 = ~w27634;// level 8
assign po04726 = ~w27637;// level 8
assign po04727 = ~w27640;// level 8
assign po04728 = ~w27643;// level 8
assign po04729 = ~w27646;// level 8
assign po04730 = ~w27649;// level 8
assign po04731 = ~w27652;// level 8
assign po04732 = ~w27655;// level 8
assign po04733 = ~w27658;// level 8
assign po04734 = ~w27661;// level 8
assign po04735 = ~w27664;// level 8
assign po04736 = ~w27667;// level 8
assign po04737 = ~w27670;// level 8
assign po04738 = ~w27673;// level 8
assign po04739 = ~w27676;// level 8
assign po04740 = ~w27679;// level 8
assign po04741 = ~w27682;// level 8
assign po04742 = ~w27685;// level 8
assign po04743 = ~w27688;// level 8
assign po04744 = ~w27691;// level 8
assign po04745 = ~w27694;// level 8
assign po04746 = ~w27697;// level 8
assign po04747 = ~w27700;// level 8
assign po04748 = ~w27703;// level 8
assign po04749 = ~w27706;// level 8
assign po04750 = ~w27709;// level 8
assign po04751 = ~w27712;// level 8
assign po04752 = ~w27715;// level 8
assign po04753 = ~w27718;// level 8
assign po04754 = ~w27721;// level 8
assign po04755 = ~w27724;// level 8
assign po04756 = ~w27727;// level 8
assign po04757 = ~w27730;// level 8
assign po04758 = ~w27733;// level 8
assign po04759 = ~w27736;// level 8
assign po04760 = ~w27739;// level 8
assign po04761 = ~w27742;// level 8
assign po04762 = ~w27745;// level 8
assign po04763 = ~w27748;// level 8
assign po04764 = ~w27751;// level 8
assign po04765 = ~w27754;// level 8
assign po04766 = ~w27757;// level 8
assign po04767 = ~w27760;// level 8
assign po04768 = ~w27763;// level 8
assign po04769 = ~w27766;// level 8
assign po04770 = ~w27769;// level 8
assign po04771 = ~w27772;// level 8
assign po04772 = ~w27775;// level 8
assign po04773 = ~w27778;// level 8
assign po04774 = ~w27781;// level 8
assign po04775 = ~w27784;// level 8
assign po04776 = ~w27787;// level 8
assign po04777 = ~w27790;// level 8
assign po04778 = ~w27793;// level 8
assign po04779 = ~w27796;// level 8
assign po04780 = ~w27799;// level 8
assign po04781 = ~w27802;// level 8
assign po04782 = ~w27805;// level 8
assign po04783 = ~w27808;// level 8
assign po04784 = ~w27811;// level 8
assign po04785 = ~w27814;// level 8
assign po04786 = ~w27817;// level 8
assign po04787 = ~w27820;// level 8
assign po04788 = ~w27823;// level 8
assign po04789 = ~w27826;// level 8
assign po04790 = ~w27829;// level 8
assign po04791 = ~w27832;// level 8
assign po04792 = ~w27835;// level 8
assign po04793 = ~w27838;// level 8
assign po04794 = ~w27841;// level 8
assign po04795 = ~w27844;// level 8
assign po04796 = ~w27847;// level 8
assign po04797 = ~w27850;// level 8
assign po04798 = ~w27853;// level 8
assign po04799 = ~w27856;// level 8
assign po04800 = ~w27859;// level 8
assign po04801 = ~w27862;// level 8
assign po04802 = ~w27865;// level 8
assign po04803 = ~w27868;// level 8
assign po04804 = ~w27871;// level 8
assign po04805 = ~w27874;// level 8
assign po04806 = ~w27877;// level 8
assign po04807 = ~w27880;// level 8
assign po04808 = ~w27883;// level 8
assign po04809 = ~w27886;// level 8
assign po04810 = ~w27889;// level 8
assign po04811 = ~w27892;// level 8
assign po04812 = ~w27895;// level 8
assign po04813 = ~w27898;// level 8
assign po04814 = ~w27901;// level 8
assign po04815 = ~w27904;// level 8
assign po04816 = ~w27907;// level 8
assign po04817 = ~w27910;// level 8
assign po04818 = ~w27913;// level 8
assign po04819 = ~w27916;// level 8
assign po04820 = ~w27919;// level 8
assign po04821 = ~w27922;// level 8
assign po04822 = ~w27925;// level 8
assign po04823 = ~w27928;// level 8
assign po04824 = ~w27931;// level 8
assign po04825 = ~w27934;// level 8
assign po04826 = ~w27937;// level 8
assign po04827 = ~w27940;// level 8
assign po04828 = ~w27943;// level 8
assign po04829 = ~w27946;// level 8
assign po04830 = ~w27949;// level 8
assign po04831 = ~w27952;// level 8
assign po04832 = ~w27955;// level 8
assign po04833 = ~w27958;// level 8
assign po04834 = ~w27961;// level 8
assign po04835 = ~w27964;// level 8
assign po04836 = ~w27967;// level 8
assign po04837 = ~w27970;// level 8
assign po04838 = ~w27973;// level 8
assign po04839 = ~w27976;// level 8
assign po04840 = ~w27979;// level 8
assign po04841 = ~w27982;// level 8
assign po04842 = ~w27985;// level 8
assign po04843 = ~w27988;// level 8
assign po04844 = ~w27991;// level 8
assign po04845 = ~w27994;// level 8
assign po04846 = ~w27997;// level 8
assign po04847 = ~w28000;// level 8
assign po04848 = ~w28003;// level 8
assign po04849 = ~w28006;// level 8
assign po04850 = ~w28009;// level 8
assign po04851 = ~w28012;// level 8
assign po04852 = ~w28015;// level 8
assign po04853 = ~w28018;// level 8
assign po04854 = ~w28021;// level 8
assign po04855 = ~w28024;// level 8
assign po04856 = ~w28027;// level 8
assign po04857 = ~w28030;// level 8
assign po04858 = ~w28033;// level 8
assign po04859 = ~w28036;// level 8
assign po04860 = ~w28039;// level 8
assign po04861 = ~w28042;// level 8
assign po04862 = ~w28045;// level 8
assign po04863 = ~w28048;// level 8
assign po04864 = ~w28051;// level 8
assign po04865 = ~w28054;// level 8
assign po04866 = ~w28057;// level 8
assign po04867 = ~w28060;// level 8
assign po04868 = ~w28063;// level 8
assign po04869 = ~w28066;// level 8
assign po04870 = ~w28069;// level 8
assign po04871 = ~w28072;// level 8
assign po04872 = ~w28075;// level 8
assign po04873 = ~w28078;// level 8
assign po04874 = ~w28081;// level 8
assign po04875 = ~w28084;// level 8
assign po04876 = ~w28087;// level 8
assign po04877 = ~w28090;// level 8
assign po04878 = ~w28093;// level 8
assign po04879 = ~w28096;// level 8
assign po04880 = ~w28099;// level 8
assign po04881 = ~w28102;// level 8
assign po04882 = ~w28105;// level 8
assign po04883 = ~w28108;// level 8
assign po04884 = ~w28111;// level 8
assign po04885 = ~w28114;// level 8
assign po04886 = ~w28117;// level 8
assign po04887 = ~w28120;// level 8
assign po04888 = ~w28123;// level 8
assign po04889 = ~w28126;// level 8
assign po04890 = ~w28129;// level 8
assign po04891 = ~w28132;// level 8
assign po04892 = ~w28135;// level 8
assign po04893 = ~w28138;// level 8
assign po04894 = ~w28141;// level 8
assign po04895 = ~w28144;// level 8
assign po04896 = ~w28147;// level 8
assign po04897 = ~w28150;// level 8
assign po04898 = ~w28153;// level 8
assign po04899 = ~w28156;// level 8
assign po04900 = ~w28159;// level 8
assign po04901 = ~w28162;// level 8
assign po04902 = ~w28165;// level 8
assign po04903 = ~w28168;// level 8
assign po04904 = ~w28171;// level 8
assign po04905 = ~w28174;// level 8
assign po04906 = ~w28177;// level 8
assign po04907 = ~w28180;// level 8
assign po04908 = ~w28183;// level 8
assign po04909 = ~w28186;// level 8
assign po04910 = ~w28189;// level 8
assign po04911 = ~w28192;// level 8
assign po04912 = ~w28195;// level 8
assign po04913 = ~w28198;// level 8
assign po04914 = ~w28201;// level 8
assign po04915 = ~w28204;// level 8
assign po04916 = ~w28207;// level 8
assign po04917 = ~w28210;// level 8
assign po04918 = ~w28213;// level 8
assign po04919 = ~w28216;// level 8
assign po04920 = ~w28219;// level 8
assign po04921 = ~w28222;// level 8
assign po04922 = ~w28225;// level 8
assign po04923 = ~w28228;// level 8
assign po04924 = ~w28231;// level 8
assign po04925 = ~w28235;// level 8
assign po04926 = ~w28238;// level 8
assign po04927 = ~w28241;// level 8
assign po04928 = ~w28244;// level 8
assign po04929 = ~w28247;// level 8
assign po04930 = ~w28250;// level 8
assign po04931 = ~w28253;// level 8
assign po04932 = ~w28256;// level 8
assign po04933 = ~w28259;// level 7
assign po04934 = ~w28262;// level 7
assign po04935 = ~w28265;// level 7
assign po04936 = ~w28268;// level 7
assign po04937 = ~w28271;// level 7
assign po04938 = ~w28274;// level 8
assign po04939 = ~w28277;// level 7
assign po04940 = ~w28280;// level 7
assign po04941 = ~w28283;// level 7
assign po04942 = ~w28286;// level 7
assign po04943 = ~w28289;// level 7
assign po04944 = ~w28292;// level 7
assign po04945 = ~w28295;// level 7
assign po04946 = ~w28298;// level 7
assign po04947 = ~w28301;// level 7
assign po04948 = ~w28304;// level 7
assign po04949 = ~w28307;// level 7
assign po04950 = ~w28310;// level 8
assign po04951 = ~w28313;// level 7
assign po04952 = ~w28316;// level 7
assign po04953 = ~w28319;// level 8
assign po04954 = ~w28322;// level 8
assign po04955 = ~w28325;// level 8
assign po04956 = ~w28328;// level 8
assign po04957 = ~w28331;// level 8
assign po04958 = ~w28334;// level 8
assign po04959 = ~w28337;// level 8
assign po04960 = ~w28341;// level 8
assign po04961 = ~w28344;// level 8
assign po04962 = ~w28347;// level 8
assign po04963 = ~w28350;// level 8
assign po04964 = ~w28353;// level 8
assign po04965 = ~w28356;// level 8
assign po04966 = ~w28360;// level 8
assign po04967 = ~w28363;// level 8
assign po04968 = ~w28366;// level 8
assign po04969 = ~w28369;// level 8
assign po04970 = ~w28372;// level 8
assign po04971 = ~w28375;// level 8
assign po04972 = ~w28378;// level 8
assign po04973 = ~w28382;// level 8
assign po04974 = ~w28385;// level 8
assign po04975 = ~w28388;// level 8
assign po04976 = ~w28391;// level 8
assign po04977 = ~w28394;// level 8
assign po04978 = ~w28397;// level 8
assign po04979 = ~w28401;// level 8
assign po04980 = ~w28404;// level 8
assign po04981 = ~w28407;// level 8
assign po04982 = ~w28410;// level 8
assign po04983 = ~w28413;// level 8
assign po04984 = ~w28416;// level 8
assign po04985 = ~w28419;// level 8
assign po04986 = ~w28423;// level 8
assign po04987 = ~w28426;// level 8
assign po04988 = ~w28429;// level 8
assign po04989 = ~w28432;// level 8
assign po04990 = ~w28435;// level 8
assign po04991 = ~w28438;// level 8
assign po04992 = ~w28442;// level 8
assign po04993 = ~w28445;// level 8
assign po04994 = ~w28448;// level 8
assign po04995 = ~w28451;// level 8
assign po04996 = ~w28454;// level 8
assign po04997 = ~w28457;// level 8
assign po04998 = ~w28460;// level 8
assign po04999 = ~w28463;// level 8
assign po05000 = ~w28467;// level 8
assign po05001 = ~w28470;// level 8
assign po05002 = ~w28473;// level 8
assign po05003 = ~w28476;// level 8
assign po05004 = ~w28479;// level 8
assign po05005 = ~w28482;// level 8
assign po05006 = ~w28486;// level 8
assign po05007 = ~w28489;// level 8
assign po05008 = ~w28492;// level 8
assign po05009 = ~w28495;// level 8
assign po05010 = ~w28498;// level 8
assign po05011 = ~w28501;// level 8
assign po05012 = ~w28504;// level 8
assign po05013 = ~w28508;// level 8
assign po05014 = ~w28511;// level 8
assign po05015 = ~w28514;// level 8
assign po05016 = ~w28517;// level 8
assign po05017 = ~w28520;// level 8
assign po05018 = ~w28523;// level 8
assign po05019 = ~w28527;// level 8
assign po05020 = ~w28530;// level 8
assign po05021 = ~w28533;// level 8
assign po05022 = ~w28536;// level 8
assign po05023 = ~w28539;// level 8
assign po05024 = ~w28542;// level 8
assign po05025 = ~w28545;// level 8
assign po05026 = ~w28549;// level 8
assign po05027 = ~w28552;// level 8
assign po05028 = ~w28555;// level 8
assign po05029 = ~w28558;// level 8
assign po05030 = ~w28561;// level 8
assign po05031 = ~w28564;// level 8
assign po05032 = ~w28568;// level 8
assign po05033 = ~w28571;// level 8
assign po05034 = ~w28574;// level 8
assign po05035 = ~w28577;// level 8
assign po05036 = ~w28580;// level 8
assign po05037 = ~w28583;// level 8
assign po05038 = ~w28586;// level 8
assign po05039 = ~w28590;// level 8
assign po05040 = ~w28593;// level 8
assign po05041 = ~w28596;// level 8
assign po05042 = ~w28599;// level 8
assign po05043 = ~w28602;// level 8
assign po05044 = ~w28605;// level 8
assign po05045 = ~w28609;// level 8
assign po05046 = ~w28612;// level 8
assign po05047 = ~w28615;// level 8
assign po05048 = ~w28618;// level 8
assign po05049 = ~w28621;// level 8
assign po05050 = ~w28624;// level 8
assign po05051 = ~w28627;// level 8
assign po05052 = ~w28631;// level 8
assign po05053 = ~w28634;// level 8
assign po05054 = ~w28637;// level 8
assign po05055 = ~w28640;// level 8
assign po05056 = ~w28643;// level 8
assign po05057 = ~w28646;// level 8
assign po05058 = ~w28650;// level 8
assign po05059 = ~w28653;// level 8
assign po05060 = ~w28656;// level 8
assign po05061 = ~w28659;// level 8
assign po05062 = ~w28662;// level 8
assign po05063 = ~w28665;// level 8
assign po05064 = ~w28668;// level 8
assign po05065 = ~w28672;// level 8
assign po05066 = ~w28675;// level 8
assign po05067 = ~w28678;// level 8
assign po05068 = ~w28681;// level 8
assign po05069 = ~w28684;// level 8
assign po05070 = ~w28687;// level 8
assign po05071 = ~w28691;// level 8
assign po05072 = ~w28694;// level 8
assign po05073 = ~w28697;// level 8
assign po05074 = ~w28700;// level 8
assign po05075 = ~w28703;// level 8
assign po05076 = ~w28706;// level 8
assign po05077 = ~w28709;// level 8
assign po05078 = ~w28713;// level 8
assign po05079 = ~w28716;// level 8
assign po05080 = ~w28719;// level 8
assign po05081 = ~w28722;// level 8
assign po05082 = ~w28725;// level 8
assign po05083 = ~w28728;// level 8
assign po05084 = ~w28732;// level 8
assign po05085 = ~w28735;// level 8
assign po05086 = ~w28738;// level 8
assign po05087 = ~w28741;// level 8
assign po05088 = ~w28744;// level 8
assign po05089 = ~w28747;// level 8
assign po05090 = ~w28750;// level 8
assign po05091 = ~w28754;// level 8
assign po05092 = ~w28757;// level 8
assign po05093 = ~w28760;// level 8
assign po05094 = ~w28763;// level 8
assign po05095 = ~w28766;// level 8
assign po05096 = ~w28769;// level 8
assign po05097 = ~w28773;// level 8
assign po05098 = ~w28776;// level 8
assign po05099 = ~w28779;// level 8
assign po05100 = ~w28782;// level 8
assign po05101 = ~w28785;// level 8
assign po05102 = ~w28788;// level 8
assign po05103 = ~w28791;// level 8
assign po05104 = ~w28795;// level 8
assign po05105 = ~w28798;// level 8
assign po05106 = ~w28801;// level 8
assign po05107 = ~w28804;// level 8
assign po05108 = ~w28807;// level 8
assign po05109 = ~w28810;// level 8
assign po05110 = ~w28814;// level 8
assign po05111 = ~w28817;// level 8
assign po05112 = ~w28820;// level 8
assign po05113 = ~w28823;// level 8
assign po05114 = ~w28826;// level 8
assign po05115 = ~w28829;// level 8
assign po05116 = ~w28832;// level 8
assign po05117 = ~w28836;// level 8
assign po05118 = ~w28839;// level 8
assign po05119 = ~w28842;// level 8
assign po05120 = ~w28845;// level 8
assign po05121 = ~w28848;// level 8
assign po05122 = ~w28851;// level 8
assign po05123 = ~w28855;// level 8
assign po05124 = ~w28858;// level 8
assign po05125 = ~w28861;// level 8
assign po05126 = ~w28864;// level 8
assign po05127 = ~w28867;// level 8
assign po05128 = ~w28870;// level 8
assign po05129 = ~w28873;// level 8
assign po05130 = ~w28877;// level 8
assign po05131 = ~w28880;// level 8
assign po05132 = ~w28883;// level 8
assign po05133 = ~w28886;// level 8
assign po05134 = ~w28889;// level 8
assign po05135 = ~w28892;// level 8
assign po05136 = ~w28896;// level 8
assign po05137 = ~w28899;// level 8
assign po05138 = ~w28902;// level 8
assign po05139 = ~w28905;// level 8
assign po05140 = ~w28908;// level 8
assign po05141 = ~w28911;// level 8
assign po05142 = ~w28914;// level 8
assign po05143 = ~w28917;// level 8
assign po05144 = ~w28921;// level 8
assign po05145 = ~w28924;// level 8
assign po05146 = ~w28927;// level 8
assign po05147 = ~w28930;// level 8
assign po05148 = ~w28933;// level 8
assign po05149 = ~w28936;// level 8
assign po05150 = ~w28940;// level 8
assign po05151 = ~w28943;// level 8
assign po05152 = ~w28946;// level 8
assign po05153 = ~w28949;// level 8
assign po05154 = ~w28952;// level 8
assign po05155 = ~w28955;// level 8
assign po05156 = ~w28958;// level 8
assign po05157 = ~w28962;// level 8
assign po05158 = ~w28965;// level 8
assign po05159 = ~w28968;// level 8
assign po05160 = ~w28971;// level 8
assign po05161 = ~w28974;// level 8
assign po05162 = ~w28977;// level 8
assign po05163 = ~w28980;// level 8
assign po05164 = ~w28983;// level 8
assign po05165 = ~w28986;// level 8
assign po05166 = ~w28989;// level 8
assign po05167 = ~w28992;// level 8
assign po05168 = ~w28995;// level 8
assign po05169 = ~w28998;// level 8
assign po05170 = ~w29001;// level 8
assign po05171 = ~w29004;// level 8
assign po05172 = ~w29007;// level 8
assign po05173 = ~w29010;// level 8
assign po05174 = ~w29013;// level 8
assign po05175 = ~w29016;// level 8
assign po05176 = ~w29019;// level 8
assign po05177 = ~w29022;// level 8
assign po05178 = ~w29025;// level 8
assign po05179 = ~w29028;// level 8
assign po05180 = ~w29031;// level 8
assign po05181 = ~w29034;// level 8
assign po05182 = ~w29037;// level 8
assign po05183 = ~w29040;// level 8
assign po05184 = ~w29043;// level 8
assign po05185 = ~w29046;// level 8
assign po05186 = ~w29049;// level 8
assign po05187 = ~w29052;// level 8
assign po05188 = ~w29055;// level 8
assign po05189 = ~w29058;// level 8
assign po05190 = ~w29061;// level 8
assign po05191 = ~w29064;// level 8
assign po05192 = ~w29067;// level 8
assign po05193 = ~w29070;// level 8
assign po05194 = ~w29073;// level 8
assign po05195 = ~w29076;// level 8
assign po05196 = ~w29079;// level 8
assign po05197 = ~w29082;// level 8
assign po05198 = ~w29085;// level 8
assign po05199 = ~w29088;// level 8
assign po05200 = ~w29091;// level 8
assign po05201 = ~w29094;// level 8
assign po05202 = ~w29097;// level 8
assign po05203 = ~w29100;// level 8
assign po05204 = ~w29103;// level 8
assign po05205 = ~w29106;// level 8
assign po05206 = ~w29109;// level 8
assign po05207 = ~w29112;// level 8
assign po05208 = ~w29115;// level 8
assign po05209 = ~w29118;// level 8
assign po05210 = ~w29121;// level 8
assign po05211 = ~w29124;// level 8
assign po05212 = ~w29127;// level 8
assign po05213 = ~w29130;// level 8
assign po05214 = ~w29133;// level 8
assign po05215 = ~w29136;// level 8
assign po05216 = ~w29139;// level 8
assign po05217 = ~w29142;// level 8
assign po05218 = ~w29145;// level 8
assign po05219 = ~w29148;// level 8
assign po05220 = ~w29151;// level 8
assign po05221 = ~w29154;// level 8
assign po05222 = ~w29157;// level 8
assign po05223 = ~w29160;// level 8
assign po05224 = ~w29163;// level 8
assign po05225 = ~w29166;// level 8
assign po05226 = ~w29169;// level 8
assign po05227 = ~w29172;// level 8
assign po05228 = ~w29175;// level 8
assign po05229 = ~w29178;// level 8
assign po05230 = ~w29181;// level 8
assign po05231 = ~w29184;// level 8
assign po05232 = ~w29187;// level 8
assign po05233 = ~w29190;// level 8
assign po05234 = ~w29193;// level 8
assign po05235 = ~w29196;// level 8
assign po05236 = ~w29199;// level 8
assign po05237 = ~w29202;// level 8
assign po05238 = ~w29206;// level 8
assign po05239 = ~w29209;// level 8
assign po05240 = ~w29212;// level 8
assign po05241 = ~w29215;// level 8
assign po05242 = ~w29218;// level 8
assign po05243 = ~w29221;// level 8
assign po05244 = ~w29224;// level 8
assign po05245 = ~w29227;// level 8
assign po05246 = ~w29230;// level 8
assign po05247 = ~w29233;// level 8
assign po05248 = ~w29236;// level 8
assign po05249 = ~w29239;// level 8
assign po05250 = ~w29242;// level 8
assign po05251 = ~w29245;// level 8
assign po05252 = ~w29248;// level 8
assign po05253 = ~w29251;// level 8
assign po05254 = ~w29254;// level 8
assign po05255 = ~w29257;// level 8
assign po05256 = ~w29260;// level 8
assign po05257 = ~w29263;// level 8
assign po05258 = ~w29266;// level 8
assign po05259 = ~w29269;// level 8
assign po05260 = ~w29272;// level 8
assign po05261 = ~w29275;// level 8
assign po05262 = ~w29278;// level 8
assign po05263 = ~w29281;// level 8
assign po05264 = ~w29284;// level 8
assign po05265 = ~w29287;// level 8
assign po05266 = ~w29290;// level 8
assign po05267 = ~w29293;// level 8
assign po05268 = ~w29296;// level 8
assign po05269 = ~w29299;// level 8
assign po05270 = ~w29302;// level 8
assign po05271 = ~w29305;// level 8
assign po05272 = ~w29308;// level 8
assign po05273 = ~w29311;// level 8
assign po05274 = ~w29314;// level 8
assign po05275 = ~w29317;// level 8
assign po05276 = ~w29320;// level 8
assign po05277 = ~w29323;// level 8
assign po05278 = ~w29326;// level 8
assign po05279 = ~w29329;// level 8
assign po05280 = ~w29332;// level 8
assign po05281 = ~w29335;// level 8
assign po05282 = ~w29338;// level 8
assign po05283 = ~w29341;// level 8
assign po05284 = ~w29344;// level 8
assign po05285 = ~w29347;// level 8
assign po05286 = ~w29350;// level 8
assign po05287 = ~w29353;// level 8
assign po05288 = ~w29356;// level 8
assign po05289 = ~w29359;// level 8
assign po05290 = ~w29362;// level 8
assign po05291 = ~w29365;// level 8
assign po05292 = ~w29368;// level 8
assign po05293 = ~w29371;// level 8
assign po05294 = ~w29374;// level 8
assign po05295 = ~w29377;// level 8
assign po05296 = ~w29380;// level 8
assign po05297 = ~w29383;// level 8
assign po05298 = ~w29386;// level 8
assign po05299 = ~w29389;// level 8
assign po05300 = ~w29392;// level 8
assign po05301 = ~w29395;// level 8
assign po05302 = ~w29398;// level 8
assign po05303 = ~w29401;// level 8
assign po05304 = ~w29404;// level 8
assign po05305 = ~w29407;// level 8
assign po05306 = ~w29410;// level 8
assign po05307 = ~w29413;// level 8
assign po05308 = ~w29416;// level 8
assign po05309 = ~w29419;// level 8
assign po05310 = ~w29422;// level 8
assign po05311 = ~w29425;// level 8
assign po05312 = ~w29428;// level 8
assign po05313 = ~w29431;// level 8
assign po05314 = ~w29434;// level 8
assign po05315 = ~w29437;// level 8
assign po05316 = ~w29440;// level 8
assign po05317 = ~w29443;// level 8
assign po05318 = ~w29446;// level 8
assign po05319 = ~w29449;// level 8
assign po05320 = ~w29452;// level 8
assign po05321 = ~w29455;// level 8
assign po05322 = ~w29458;// level 8
assign po05323 = ~w29461;// level 8
assign po05324 = ~w29464;// level 8
assign po05325 = ~w29467;// level 8
assign po05326 = ~w29470;// level 8
assign po05327 = ~w29473;// level 8
assign po05328 = ~w29476;// level 8
assign po05329 = ~w29479;// level 8
assign po05330 = ~w29482;// level 8
assign po05331 = ~w29485;// level 8
assign po05332 = ~w29488;// level 8
assign po05333 = ~w29491;// level 8
assign po05334 = ~w29494;// level 8
assign po05335 = ~w29497;// level 8
assign po05336 = ~w29500;// level 8
assign po05337 = ~w29503;// level 8
assign po05338 = ~w29506;// level 8
assign po05339 = ~w29509;// level 8
assign po05340 = ~w29512;// level 8
assign po05341 = ~w29515;// level 8
assign po05342 = ~w29518;// level 8
assign po05343 = ~w29521;// level 8
assign po05344 = ~w29524;// level 8
assign po05345 = ~w29527;// level 8
assign po05346 = ~w29530;// level 8
assign po05347 = ~w29533;// level 8
assign po05348 = ~w29536;// level 8
assign po05349 = ~w29539;// level 8
assign po05350 = ~w29542;// level 8
assign po05351 = ~w29545;// level 8
assign po05352 = ~w29548;// level 8
assign po05353 = ~w29551;// level 8
assign po05354 = ~w29554;// level 8
assign po05355 = ~w29557;// level 8
assign po05356 = ~w29560;// level 8
assign po05357 = ~w29563;// level 8
assign po05358 = ~w29566;// level 8
assign po05359 = ~w29569;// level 8
assign po05360 = ~w29572;// level 8
assign po05361 = ~w29575;// level 8
assign po05362 = ~w29578;// level 8
assign po05363 = ~w29581;// level 8
assign po05364 = ~w29584;// level 8
assign po05365 = ~w29587;// level 8
assign po05366 = ~w29590;// level 8
assign po05367 = ~w29593;// level 8
assign po05368 = ~w29596;// level 8
assign po05369 = ~w29599;// level 8
assign po05370 = ~w29602;// level 8
assign po05371 = ~w29605;// level 8
assign po05372 = ~w29608;// level 8
assign po05373 = ~w29611;// level 8
assign po05374 = ~w29614;// level 8
assign po05375 = ~w29617;// level 8
assign po05376 = ~w29620;// level 8
assign po05377 = ~w29623;// level 8
assign po05378 = ~w29626;// level 8
assign po05379 = ~w29629;// level 8
assign po05380 = ~w29632;// level 8
assign po05381 = ~w29635;// level 8
assign po05382 = ~w29638;// level 8
assign po05383 = ~w29641;// level 8
assign po05384 = ~w29644;// level 8
assign po05385 = ~w29647;// level 8
assign po05386 = ~w29650;// level 8
assign po05387 = ~w29653;// level 8
assign po05388 = ~w29656;// level 8
assign po05389 = ~w29659;// level 8
assign po05390 = ~w29662;// level 8
assign po05391 = ~w29665;// level 8
assign po05392 = ~w29668;// level 8
assign po05393 = ~w29671;// level 8
assign po05394 = ~w29674;// level 8
assign po05395 = ~w29677;// level 8
assign po05396 = ~w29680;// level 8
assign po05397 = ~w29683;// level 8
assign po05398 = ~w29686;// level 8
assign po05399 = ~w29689;// level 8
assign po05400 = ~w29692;// level 8
assign po05401 = ~w29695;// level 8
assign po05402 = ~w29698;// level 8
assign po05403 = ~w29701;// level 8
assign po05404 = ~w29704;// level 8
assign po05405 = ~w29707;// level 8
assign po05406 = ~w29710;// level 8
assign po05407 = ~w29713;// level 8
assign po05408 = ~w29716;// level 8
assign po05409 = ~w29719;// level 8
assign po05410 = ~w29722;// level 8
assign po05411 = ~w29725;// level 8
assign po05412 = ~w29728;// level 8
assign po05413 = ~w29731;// level 8
assign po05414 = ~w29734;// level 8
assign po05415 = ~w29737;// level 8
assign po05416 = ~w29740;// level 8
assign po05417 = ~w29743;// level 8
assign po05418 = ~w29746;// level 8
assign po05419 = ~w29749;// level 8
assign po05420 = ~w29752;// level 8
assign po05421 = ~w29755;// level 8
assign po05422 = ~w29758;// level 8
assign po05423 = ~w29761;// level 8
assign po05424 = ~w29764;// level 8
assign po05425 = ~w29767;// level 8
assign po05426 = ~w29770;// level 8
assign po05427 = ~w29773;// level 8
assign po05428 = ~w29776;// level 8
assign po05429 = ~w29779;// level 8
assign po05430 = ~w29782;// level 8
assign po05431 = ~w29785;// level 8
assign po05432 = ~w29788;// level 8
assign po05433 = ~w29791;// level 8
assign po05434 = ~w29794;// level 8
assign po05435 = ~w29797;// level 8
assign po05436 = ~w29800;// level 8
assign po05437 = ~w29803;// level 8
assign po05438 = ~w29806;// level 8
assign po05439 = ~w29809;// level 8
assign po05440 = ~w29812;// level 8
assign po05441 = ~w29815;// level 8
assign po05442 = ~w29818;// level 8
assign po05443 = ~w29821;// level 8
assign po05444 = ~w29824;// level 8
assign po05445 = ~w29827;// level 8
assign po05446 = ~w29830;// level 8
assign po05447 = ~w29833;// level 8
assign po05448 = ~w29836;// level 8
assign po05449 = ~w29839;// level 8
assign po05450 = ~w29842;// level 8
assign po05451 = ~w29845;// level 8
assign po05452 = ~w29848;// level 7
assign po05453 = ~w29851;// level 8
assign po05454 = ~w29854;// level 8
assign po05455 = ~w29857;// level 8
assign po05456 = ~w29860;// level 8
assign po05457 = ~w29863;// level 8
assign po05458 = ~w29866;// level 8
assign po05459 = ~w29869;// level 8
assign po05460 = ~w29872;// level 8
assign po05461 = ~w29875;// level 8
assign po05462 = ~w29878;// level 8
assign po05463 = ~w29881;// level 8
assign po05464 = ~w29884;// level 8
assign po05465 = ~w29887;// level 8
assign po05466 = ~w29890;// level 8
assign po05467 = ~w29893;// level 8
assign po05468 = ~w29896;// level 8
assign po05469 = ~w29899;// level 8
assign po05470 = ~w29902;// level 8
assign po05471 = ~w29905;// level 8
assign po05472 = ~w29908;// level 8
assign po05473 = ~w29911;// level 8
assign po05474 = ~w29914;// level 8
assign po05475 = ~w29917;// level 8
assign po05476 = ~w29920;// level 8
assign po05477 = ~w29923;// level 8
assign po05478 = ~w29926;// level 8
assign po05479 = ~w29929;// level 8
assign po05480 = ~w29932;// level 8
assign po05481 = ~w29935;// level 8
assign po05482 = ~w29938;// level 8
assign po05483 = ~w29941;// level 8
assign po05484 = ~w29944;// level 8
assign po05485 = ~w29947;// level 8
assign po05486 = ~w29950;// level 8
assign po05487 = ~w29953;// level 8
assign po05488 = ~w29956;// level 8
assign po05489 = ~w29959;// level 8
assign po05490 = ~w29962;// level 8
assign po05491 = ~w29965;// level 8
assign po05492 = ~w29968;// level 8
assign po05493 = ~w29971;// level 8
assign po05494 = ~w29974;// level 8
assign po05495 = ~w29977;// level 8
assign po05496 = ~w29980;// level 8
assign po05497 = ~w29983;// level 8
assign po05498 = ~w29986;// level 8
assign po05499 = ~w29990;// level 8
assign po05500 = ~w29993;// level 8
assign po05501 = ~w29996;// level 8
assign po05502 = ~w29999;// level 8
assign po05503 = ~w30002;// level 8
assign po05504 = ~w30005;// level 8
assign po05505 = ~w30008;// level 8
assign po05506 = ~w30011;// level 8
assign po05507 = ~w30014;// level 8
assign po05508 = ~w30017;// level 8
assign po05509 = ~w30020;// level 8
assign po05510 = ~w30023;// level 8
assign po05511 = ~w30026;// level 8
assign po05512 = ~w30029;// level 8
assign po05513 = ~w30032;// level 8
assign po05514 = ~w30035;// level 8
assign po05515 = ~w30038;// level 8
assign po05516 = ~w30041;// level 8
assign po05517 = ~w30044;// level 8
assign po05518 = ~w30047;// level 8
assign po05519 = ~w30050;// level 8
assign po05520 = ~w30053;// level 8
assign po05521 = ~w30056;// level 8
assign po05522 = ~w30059;// level 8
assign po05523 = ~w30062;// level 8
assign po05524 = ~w30065;// level 8
assign po05525 = ~w30068;// level 8
assign po05526 = ~w30071;// level 8
assign po05527 = ~w30074;// level 8
assign po05528 = ~w30077;// level 8
assign po05529 = ~w30080;// level 8
assign po05530 = ~w30083;// level 8
assign po05531 = ~w30086;// level 8
assign po05532 = ~w30089;// level 8
assign po05533 = ~w30092;// level 8
assign po05534 = ~w30095;// level 8
assign po05535 = ~w30098;// level 8
assign po05536 = ~w30101;// level 8
assign po05537 = ~w30104;// level 8
assign po05538 = ~w30107;// level 8
assign po05539 = ~w30110;// level 8
assign po05540 = ~w30113;// level 8
assign po05541 = ~w30116;// level 8
assign po05542 = ~w30119;// level 8
assign po05543 = ~w30122;// level 8
assign po05544 = ~w30125;// level 8
assign po05545 = ~w30128;// level 8
assign po05546 = ~w30131;// level 8
assign po05547 = ~w30134;// level 7
assign po05548 = ~w30137;// level 8
assign po05549 = ~w30140;// level 8
assign po05550 = ~w30143;// level 7
assign po05551 = ~w30146;// level 8
assign po05552 = ~w30149;// level 7
assign po05553 = ~w30152;// level 8
assign po05554 = ~w30156;// level 8
assign po05555 = ~w30159;// level 8
assign po05556 = ~w30162;// level 8
assign po05557 = ~w30165;// level 8
assign po05558 = ~w30168;// level 8
assign po05559 = ~w30171;// level 8
assign po05560 = ~w30174;// level 8
assign po05561 = ~w30177;// level 8
assign po05562 = ~w30181;// level 8
assign po05563 = ~w30184;// level 8
assign po05564 = ~w30187;// level 8
assign po05565 = ~w30190;// level 8
assign po05566 = ~w30193;// level 8
assign po05567 = ~w30196;// level 8
assign po05568 = ~w30199;// level 8
assign po05569 = ~w30203;// level 8
assign po05570 = ~w30206;// level 8
assign po05571 = ~w30209;// level 8
assign po05572 = ~w30212;// level 8
assign po05573 = ~w30215;// level 8
assign po05574 = ~w30218;// level 8
assign po05575 = ~w30221;// level 8
assign po05576 = ~w30225;// level 8
assign po05577 = ~w30228;// level 8
assign po05578 = ~w30231;// level 8
assign po05579 = ~w30234;// level 8
assign po05580 = ~w30237;// level 8
assign po05581 = ~w30240;// level 8
assign po05582 = ~w30243;// level 8
assign po05583 = ~w30247;// level 8
assign po05584 = ~w30250;// level 8
assign po05585 = ~w30253;// level 8
assign po05586 = ~w30256;// level 8
assign po05587 = ~w30259;// level 8
assign po05588 = ~w30262;// level 8
assign po05589 = ~w30266;// level 8
assign po05590 = ~w30269;// level 8
assign po05591 = ~w30272;// level 8
assign po05592 = ~w30275;// level 8
assign po05593 = ~w30278;// level 8
assign po05594 = ~w30281;// level 8
assign po05595 = ~w30284;// level 8
assign po05596 = ~w30288;// level 8
assign po05597 = ~w30291;// level 8
assign po05598 = ~w30294;// level 8
assign po05599 = ~w30297;// level 8
assign po05600 = ~w30300;// level 8
assign po05601 = ~w30303;// level 8
assign po05602 = ~w30306;// level 8
assign po05603 = ~w30310;// level 8
assign po05604 = ~w30313;// level 8
assign po05605 = ~w30316;// level 8
assign po05606 = ~w30319;// level 8
assign po05607 = ~w30322;// level 8
assign po05608 = ~w30325;// level 8
assign po05609 = ~w30328;// level 8
assign po05610 = ~w30332;// level 8
assign po05611 = ~w30335;// level 8
assign po05612 = ~w30338;// level 8
assign po05613 = ~w30341;// level 8
assign po05614 = ~w30344;// level 8
assign po05615 = ~w30347;// level 8
assign po05616 = ~w30351;// level 8
assign po05617 = ~w30354;// level 8
assign po05618 = ~w30357;// level 8
assign po05619 = ~w30360;// level 8
assign po05620 = ~w30363;// level 8
assign po05621 = ~w30366;// level 8
assign po05622 = ~w30369;// level 8
assign po05623 = ~w30373;// level 8
assign po05624 = ~w30376;// level 8
assign po05625 = ~w30379;// level 8
assign po05626 = ~w30382;// level 8
assign po05627 = ~w30385;// level 8
assign po05628 = ~w30388;// level 8
assign po05629 = ~w30392;// level 8
assign po05630 = ~w30395;// level 8
assign po05631 = ~w30398;// level 8
assign po05632 = ~w30401;// level 8
assign po05633 = ~w30404;// level 8
assign po05634 = ~w30407;// level 8
assign po05635 = ~w30410;// level 8
assign po05636 = ~w30414;// level 8
assign po05637 = ~w30417;// level 8
assign po05638 = ~w30420;// level 8
assign po05639 = ~w30423;// level 8
assign po05640 = ~w30426;// level 8
assign po05641 = ~w30429;// level 8
assign po05642 = ~w30433;// level 8
assign po05643 = ~w30436;// level 8
assign po05644 = ~w30439;// level 8
assign po05645 = ~w30442;// level 8
assign po05646 = ~w30445;// level 8
assign po05647 = ~w30448;// level 8
assign po05648 = ~w30451;// level 8
assign po05649 = ~w30455;// level 8
assign po05650 = ~w30458;// level 8
assign po05651 = ~w30461;// level 8
assign po05652 = ~w30464;// level 8
assign po05653 = ~w30467;// level 8
assign po05654 = ~w30470;// level 8
assign po05655 = ~w30474;// level 8
assign po05656 = ~w30477;// level 8
assign po05657 = ~w30480;// level 8
assign po05658 = ~w30483;// level 8
assign po05659 = ~w30486;// level 8
assign po05660 = ~w30489;// level 8
assign po05661 = ~w30492;// level 8
assign po05662 = ~w30496;// level 8
assign po05663 = ~w30499;// level 8
assign po05664 = ~w30502;// level 8
assign po05665 = ~w30505;// level 8
assign po05666 = ~w30508;// level 8
assign po05667 = ~w30511;// level 8
assign po05668 = ~w30515;// level 8
assign po05669 = ~w30518;// level 8
assign po05670 = ~w30521;// level 8
assign po05671 = ~w30524;// level 8
assign po05672 = ~w30527;// level 8
assign po05673 = ~w30530;// level 8
assign po05674 = ~w30533;// level 8
assign po05675 = ~w30537;// level 8
assign po05676 = ~w30540;// level 8
assign po05677 = ~w30543;// level 8
assign po05678 = ~w30546;// level 8
assign po05679 = ~w30549;// level 8
assign po05680 = ~w30552;// level 8
assign po05681 = ~w30556;// level 8
assign po05682 = ~w30559;// level 8
assign po05683 = ~w30562;// level 8
assign po05684 = ~w30565;// level 8
assign po05685 = ~w30568;// level 8
assign po05686 = ~w30571;// level 8
assign po05687 = ~w30574;// level 8
assign po05688 = ~w30578;// level 8
assign po05689 = ~w30581;// level 8
assign po05690 = ~w30584;// level 8
assign po05691 = ~w30587;// level 8
assign po05692 = ~w30590;// level 8
assign po05693 = ~w30593;// level 8
assign po05694 = ~w30597;// level 8
assign po05695 = ~w30600;// level 8
assign po05696 = ~w30603;// level 8
assign po05697 = ~w30606;// level 8
assign po05698 = ~w30609;// level 8
assign po05699 = ~w30612;// level 8
assign po05700 = ~w30615;// level 8
assign po05701 = ~w30619;// level 8
assign po05702 = ~w30622;// level 8
assign po05703 = ~w30625;// level 8
assign po05704 = ~w30628;// level 8
assign po05705 = ~w30631;// level 8
assign po05706 = ~w30634;// level 8
assign po05707 = ~w30638;// level 8
assign po05708 = ~w30641;// level 8
assign po05709 = ~w30644;// level 8
assign po05710 = ~w30647;// level 8
assign po05711 = ~w30650;// level 8
assign po05712 = ~w30653;// level 8
assign po05713 = ~w30656;// level 8
assign po05714 = ~w30659;// level 8
assign po05715 = ~w30662;// level 8
assign po05716 = ~w30665;// level 8
assign po05717 = ~w30668;// level 8
assign po05718 = ~w30671;// level 8
assign po05719 = ~w30674;// level 8
assign po05720 = ~w30677;// level 8
assign po05721 = ~w30680;// level 8
assign po05722 = ~w30683;// level 8
assign po05723 = ~w30686;// level 8
assign po05724 = ~w30689;// level 8
assign po05725 = ~w30692;// level 8
assign po05726 = ~w30695;// level 8
assign po05727 = ~w30698;// level 8
assign po05728 = ~w30701;// level 8
assign po05729 = ~w30704;// level 8
assign po05730 = ~w30707;// level 8
assign po05731 = ~w30710;// level 8
assign po05732 = ~w30713;// level 8
assign po05733 = ~w30716;// level 8
assign po05734 = ~w30719;// level 8
assign po05735 = ~w30722;// level 8
assign po05736 = ~w30725;// level 8
assign po05737 = ~w30728;// level 8
assign po05738 = ~w30731;// level 8
assign po05739 = ~w30734;// level 8
assign po05740 = ~w30737;// level 8
assign po05741 = ~w30740;// level 8
assign po05742 = ~w30743;// level 8
assign po05743 = ~w30746;// level 8
assign po05744 = ~w30749;// level 8
assign po05745 = ~w30752;// level 8
assign po05746 = ~w30755;// level 8
assign po05747 = ~w30758;// level 8
assign po05748 = ~w30761;// level 8
assign po05749 = ~w30764;// level 8
assign po05750 = ~w30767;// level 8
assign po05751 = ~w30770;// level 8
assign po05752 = ~w30773;// level 8
assign po05753 = ~w30776;// level 8
assign po05754 = ~w30779;// level 8
assign po05755 = ~w30782;// level 8
assign po05756 = ~w30785;// level 8
assign po05757 = ~w30788;// level 8
assign po05758 = ~w30791;// level 8
assign po05759 = ~w30794;// level 8
assign po05760 = ~w30797;// level 8
assign po05761 = ~w30800;// level 8
assign po05762 = ~w30803;// level 8
assign po05763 = ~w30806;// level 8
assign po05764 = ~w30809;// level 8
assign po05765 = ~w30812;// level 8
assign po05766 = ~w30815;// level 8
assign po05767 = ~w30818;// level 8
assign po05768 = ~w30821;// level 8
assign po05769 = ~w30824;// level 8
assign po05770 = ~w30827;// level 8
assign po05771 = ~w30830;// level 8
assign po05772 = ~w30833;// level 8
assign po05773 = ~w30836;// level 8
assign po05774 = ~w30839;// level 8
assign po05775 = ~w30842;// level 8
assign po05776 = ~w30845;// level 8
assign po05777 = ~w30848;// level 8
assign po05778 = ~w30851;// level 8
assign po05779 = ~w30854;// level 8
assign po05780 = ~w30857;// level 8
assign po05781 = ~w30860;// level 8
assign po05782 = ~w30863;// level 8
assign po05783 = ~w30866;// level 8
assign po05784 = ~w30869;// level 8
assign po05785 = ~w30872;// level 8
assign po05786 = ~w30875;// level 8
assign po05787 = ~w30878;// level 8
assign po05788 = ~w30881;// level 8
assign po05789 = ~w30884;// level 8
assign po05790 = ~w30887;// level 8
assign po05791 = ~w30890;// level 8
assign po05792 = ~w30893;// level 8
assign po05793 = ~w30896;// level 8
assign po05794 = ~w30900;// level 8
assign po05795 = ~w30903;// level 8
assign po05796 = ~w30906;// level 8
assign po05797 = ~w30909;// level 8
assign po05798 = ~w30912;// level 8
assign po05799 = ~w30915;// level 8
assign po05800 = ~w30918;// level 8
assign po05801 = ~w30921;// level 8
assign po05802 = ~w30924;// level 8
assign po05803 = ~w30927;// level 8
assign po05804 = ~w30930;// level 8
assign po05805 = ~w30933;// level 8
assign po05806 = ~w30936;// level 8
assign po05807 = ~w30939;// level 8
assign po05808 = ~w30942;// level 8
assign po05809 = ~w30945;// level 8
assign po05810 = ~w30948;// level 8
assign po05811 = ~w30951;// level 8
assign po05812 = ~w30954;// level 8
assign po05813 = ~w30957;// level 8
assign po05814 = ~w30960;// level 8
assign po05815 = ~w30963;// level 8
assign po05816 = ~w30966;// level 8
assign po05817 = ~w30969;// level 8
assign po05818 = ~w30972;// level 8
assign po05819 = ~w30975;// level 8
assign po05820 = ~w30978;// level 8
assign po05821 = ~w30981;// level 8
assign po05822 = ~w30984;// level 8
assign po05823 = ~w30987;// level 8
assign po05824 = ~w30990;// level 8
assign po05825 = ~w30993;// level 8
assign po05826 = ~w30996;// level 8
assign po05827 = ~w30999;// level 8
assign po05828 = ~w31002;// level 8
assign po05829 = ~w31005;// level 8
assign po05830 = ~w31008;// level 8
assign po05831 = ~w31011;// level 8
assign po05832 = ~w31014;// level 8
assign po05833 = ~w31017;// level 8
assign po05834 = ~w31020;// level 8
assign po05835 = ~w31023;// level 8
assign po05836 = ~w31026;// level 8
assign po05837 = ~w31029;// level 8
assign po05838 = ~w31033;// level 8
assign po05839 = ~w31036;// level 8
assign po05840 = ~w31039;// level 8
assign po05841 = ~w31042;// level 8
assign po05842 = ~w31045;// level 8
assign po05843 = ~w31048;// level 8
assign po05844 = ~w31051;// level 8
assign po05845 = ~w31054;// level 8
assign po05846 = ~w31057;// level 8
assign po05847 = ~w31060;// level 8
assign po05848 = ~w31064;// level 8
assign po05849 = ~w31067;// level 8
assign po05850 = ~w31070;// level 8
assign po05851 = ~w31073;// level 8
assign po05852 = ~w31076;// level 8
assign po05853 = ~w31079;// level 8
assign po05854 = ~w31082;// level 8
assign po05855 = ~w31085;// level 8
assign po05856 = ~w31088;// level 8
assign po05857 = ~w31091;// level 8
assign po05858 = ~w31094;// level 8
assign po05859 = ~w31097;// level 8
assign po05860 = ~w31100;// level 8
assign po05861 = ~w31103;// level 8
assign po05862 = ~w31106;// level 8
assign po05863 = ~w31109;// level 8
assign po05864 = ~w31112;// level 8
assign po05865 = ~w31115;// level 8
assign po05866 = ~w31118;// level 8
assign po05867 = ~w31121;// level 8
assign po05868 = ~w31124;// level 8
assign po05869 = ~w31127;// level 8
assign po05870 = ~w31130;// level 8
assign po05871 = ~w31133;// level 8
assign po05872 = ~w31136;// level 8
assign po05873 = ~w31139;// level 8
assign po05874 = ~w31142;// level 8
assign po05875 = ~w31145;// level 8
assign po05876 = ~w31148;// level 8
assign po05877 = ~w31151;// level 8
assign po05878 = ~w31154;// level 8
assign po05879 = ~w31157;// level 8
assign po05880 = ~w31160;// level 8
assign po05881 = ~w31163;// level 8
assign po05882 = ~w31166;// level 8
assign po05883 = ~w31169;// level 8
assign po05884 = ~w31172;// level 8
assign po05885 = ~w31175;// level 8
assign po05886 = ~w31178;// level 8
assign po05887 = ~w31181;// level 8
assign po05888 = ~w31184;// level 8
assign po05889 = ~w31187;// level 8
assign po05890 = ~w31190;// level 8
assign po05891 = ~w31193;// level 8
assign po05892 = ~w31196;// level 8
assign po05893 = ~w31199;// level 8
assign po05894 = ~w31202;// level 8
assign po05895 = ~w31205;// level 8
assign po05896 = ~w31208;// level 8
assign po05897 = ~w31211;// level 8
assign po05898 = ~w31214;// level 8
assign po05899 = ~w31217;// level 8
assign po05900 = ~w31220;// level 8
assign po05901 = ~w31223;// level 8
assign po05902 = ~w31226;// level 8
assign po05903 = ~w31229;// level 8
assign po05904 = ~w31232;// level 8
assign po05905 = ~w31235;// level 8
assign po05906 = ~w31238;// level 8
assign po05907 = ~w31241;// level 8
assign po05908 = ~w31244;// level 8
assign po05909 = ~w31247;// level 8
assign po05910 = ~w31250;// level 8
assign po05911 = ~w31253;// level 8
assign po05912 = ~w31256;// level 8
assign po05913 = ~w31259;// level 8
assign po05914 = ~w31262;// level 8
assign po05915 = ~w31265;// level 8
assign po05916 = ~w31268;// level 8
assign po05917 = ~w31272;// level 8
assign po05918 = ~w31275;// level 8
assign po05919 = ~w31278;// level 8
assign po05920 = ~w31281;// level 8
assign po05921 = ~w31284;// level 8
assign po05922 = ~w31287;// level 8
assign po05923 = ~w31290;// level 8
assign po05924 = ~w31293;// level 8
assign po05925 = ~w31296;// level 8
assign po05926 = ~w31299;// level 8
assign po05927 = ~w31302;// level 8
assign po05928 = ~w31305;// level 8
assign po05929 = ~w31308;// level 8
assign po05930 = ~w31311;// level 8
assign po05931 = ~w31314;// level 8
assign po05932 = ~w31317;// level 8
assign po05933 = ~w31320;// level 8
assign po05934 = ~w31323;// level 8
assign po05935 = ~w31326;// level 8
assign po05936 = ~w31329;// level 8
assign po05937 = ~w31332;// level 8
assign po05938 = ~w31335;// level 8
assign po05939 = ~w31338;// level 8
assign po05940 = ~w31341;// level 8
assign po05941 = ~w31344;// level 8
assign po05942 = ~w31347;// level 8
assign po05943 = ~w31351;// level 8
assign po05944 = ~w31354;// level 8
assign po05945 = ~w31357;// level 8
assign po05946 = ~w31360;// level 8
assign po05947 = ~w31363;// level 8
assign po05948 = ~w31366;// level 8
assign po05949 = ~w31369;// level 8
assign po05950 = ~w31372;// level 8
assign po05951 = ~w31375;// level 8
assign po05952 = ~w31378;// level 8
assign po05953 = ~w31381;// level 8
assign po05954 = ~w31384;// level 8
assign po05955 = ~w31387;// level 8
assign po05956 = ~w31390;// level 8
assign po05957 = ~w31393;// level 8
assign po05958 = ~w31396;// level 8
assign po05959 = ~w31399;// level 8
assign po05960 = ~w31402;// level 8
assign po05961 = ~w31405;// level 8
assign po05962 = ~w31408;// level 8
assign po05963 = ~w31411;// level 8
assign po05964 = ~w31414;// level 8
assign po05965 = ~w31417;// level 8
assign po05966 = ~w31420;// level 8
assign po05967 = ~w31423;// level 8
assign po05968 = ~w31426;// level 8
assign po05969 = ~w31429;// level 8
assign po05970 = ~w31432;// level 8
assign po05971 = ~w31435;// level 8
assign po05972 = ~w31438;// level 8
assign po05973 = ~w31441;// level 8
assign po05974 = ~w31444;// level 8
assign po05975 = ~w31447;// level 8
assign po05976 = ~w31451;// level 8
assign po05977 = ~w31454;// level 8
assign po05978 = ~w31457;// level 8
assign po05979 = ~w31460;// level 8
assign po05980 = ~w31463;// level 8
assign po05981 = ~w31466;// level 8
assign po05982 = ~w31469;// level 8
assign po05983 = ~w31472;// level 8
assign po05984 = ~w31476;// level 8
assign po05985 = ~w31480;// level 8
assign po05986 = ~w31483;// level 8
assign po05987 = ~w31486;// level 8
assign po05988 = ~w31489;// level 8
assign po05989 = ~w31492;// level 8
assign po05990 = ~w31495;// level 8
assign po05991 = ~w31498;// level 8
assign po05992 = ~w31501;// level 8
assign po05993 = ~w31504;// level 8
assign po05994 = ~w31508;// level 8
assign po05995 = ~w31511;// level 8
assign po05996 = ~w31514;// level 8
assign po05997 = ~w31517;// level 8
assign po05998 = ~w31520;// level 8
assign po05999 = ~w31523;// level 8
assign po06000 = ~w31526;// level 8
assign po06001 = ~w31529;// level 8
assign po06002 = ~w31533;// level 8
assign po06003 = ~w31536;// level 8
assign po06004 = ~w31540;// level 8
assign po06005 = ~w31543;// level 8
assign po06006 = ~w31546;// level 8
assign po06007 = ~w31549;// level 8
assign po06008 = ~w31552;// level 8
assign po06009 = ~w31555;// level 8
assign po06010 = ~w31558;// level 8
assign po06011 = ~w31561;// level 8
assign po06012 = ~w31564;// level 8
assign po06013 = ~w31567;// level 8
assign po06014 = ~w31571;// level 8
assign po06015 = ~w31574;// level 8
assign po06016 = ~w31577;// level 8
assign po06017 = ~w31580;// level 8
assign po06018 = ~w31583;// level 8
assign po06019 = ~w31586;// level 8
assign po06020 = ~w31589;// level 8
assign po06021 = ~w31592;// level 8
assign po06022 = ~w31596;// level 8
assign po06023 = ~w31599;// level 8
assign po06024 = ~w31602;// level 8
assign po06025 = ~w31605;// level 8
assign po06026 = ~w31608;// level 8
assign po06027 = ~w31611;// level 8
assign po06028 = ~w31614;// level 8
assign po06029 = ~w31618;// level 8
assign po06030 = ~w31621;// level 8
assign po06031 = ~w31624;// level 8
assign po06032 = ~w31627;// level 8
assign po06033 = ~w31630;// level 8
assign po06034 = ~w31633;// level 8
assign po06035 = ~w31637;// level 8
assign po06036 = ~w31640;// level 8
assign po06037 = ~w31643;// level 8
assign po06038 = ~w31646;// level 8
assign po06039 = ~w31649;// level 8
assign po06040 = ~w31652;// level 8
assign po06041 = ~w31655;// level 8
assign po06042 = ~w31659;// level 8
assign po06043 = ~w31662;// level 8
assign po06044 = ~w31665;// level 8
assign po06045 = ~w31668;// level 8
assign po06046 = ~w31671;// level 8
assign po06047 = ~w31675;// level 8
assign po06048 = ~w31679;// level 8
assign po06049 = ~w31683;// level 8
assign po06050 = ~w31686;// level 8
assign po06051 = ~w31689;// level 8
assign po06052 = ~w31692;// level 8
assign po06053 = ~w31695;// level 8
assign po06054 = ~w31698;// level 8
assign po06055 = ~w31701;// level 8
assign po06056 = ~w31704;// level 8
assign po06057 = ~w31707;// level 8
assign po06058 = ~w31710;// level 8
assign po06059 = ~w31713;// level 8
assign po06060 = ~w31716;// level 8
assign po06061 = ~w31719;// level 8
assign po06062 = ~w31723;// level 8
assign po06063 = ~w31726;// level 8
assign po06064 = ~w31729;// level 8
assign po06065 = ~w31732;// level 8
assign po06066 = ~w31735;// level 8
assign po06067 = ~w31738;// level 8
assign po06068 = ~w31741;// level 8
assign po06069 = ~w31744;// level 8
assign po06070 = ~w31747;// level 8
assign po06071 = ~w31750;// level 8
assign po06072 = ~w31753;// level 8
assign po06073 = ~w31756;// level 8
assign po06074 = ~w31759;// level 8
assign po06075 = ~w31762;// level 8
assign po06076 = ~w31765;// level 8
assign po06077 = ~w31768;// level 8
assign po06078 = ~w31771;// level 8
assign po06079 = ~w31774;// level 8
assign po06080 = ~w31777;// level 8
assign po06081 = ~w31780;// level 8
assign po06082 = ~w31783;// level 8
assign po06083 = ~w31786;// level 8
assign po06084 = ~w31789;// level 8
assign po06085 = ~w31792;// level 8
assign po06086 = ~w31795;// level 8
assign po06087 = ~w31798;// level 8
assign po06088 = ~w31801;// level 8
assign po06089 = ~w31804;// level 8
assign po06090 = ~w31807;// level 8
assign po06091 = ~w31810;// level 8
assign po06092 = ~w31813;// level 8
assign po06093 = ~w31816;// level 8
assign po06094 = ~w31819;// level 8
assign po06095 = ~w31822;// level 8
assign po06096 = ~w31825;// level 8
assign po06097 = ~w31828;// level 8
assign po06098 = ~w31831;// level 8
assign po06099 = ~w31834;// level 8
assign po06100 = ~w31837;// level 8
assign po06101 = ~w31840;// level 8
assign po06102 = ~w31843;// level 8
assign po06103 = ~w31846;// level 8
assign po06104 = ~w31849;// level 8
assign po06105 = ~w31852;// level 8
assign po06106 = ~w31855;// level 8
assign po06107 = ~w31858;// level 8
assign po06108 = ~w31861;// level 8
assign po06109 = ~w31864;// level 8
assign po06110 = ~w31867;// level 8
assign po06111 = ~w31870;// level 8
assign po06112 = ~w31873;// level 8
assign po06113 = ~w31876;// level 8
assign po06114 = ~w31880;// level 8
assign po06115 = ~w31883;// level 8
assign po06116 = ~w31886;// level 8
assign po06117 = ~w31889;// level 8
assign po06118 = ~w31892;// level 8
assign po06119 = ~w31895;// level 8
assign po06120 = ~w31898;// level 8
assign po06121 = ~w31901;// level 8
assign po06122 = ~w31904;// level 8
assign po06123 = ~w31907;// level 8
assign po06124 = ~w31910;// level 8
assign po06125 = ~w31913;// level 8
assign po06126 = ~w31916;// level 8
assign po06127 = ~w31919;// level 8
assign po06128 = ~w31922;// level 8
assign po06129 = ~w31925;// level 8
assign po06130 = ~w31928;// level 8
assign po06131 = ~w31931;// level 8
assign po06132 = ~w31934;// level 8
assign po06133 = ~w31937;// level 8
assign po06134 = ~w31940;// level 8
assign po06135 = ~w31943;// level 8
assign po06136 = ~w31946;// level 8
assign po06137 = ~w31949;// level 8
assign po06138 = ~w31952;// level 8
assign po06139 = ~w31955;// level 8
assign po06140 = ~w31958;// level 8
assign po06141 = ~w31961;// level 7
assign po06142 = ~w31964;// level 7
assign po06143 = ~w31967;// level 7
assign po06144 = ~w31970;// level 8
assign po06145 = ~w31973;// level 8
assign po06146 = ~w31976;// level 8
assign po06147 = ~w31979;// level 8
assign po06148 = ~w31982;// level 8
assign po06149 = ~w31985;// level 8
assign po06150 = ~w31988;// level 8
assign po06151 = ~w31991;// level 8
assign po06152 = ~w31994;// level 8
assign po06153 = ~w31997;// level 8
assign po06154 = ~w32000;// level 8
assign po06155 = ~w32003;// level 8
assign po06156 = ~w32006;// level 8
assign po06157 = ~w32009;// level 8
assign po06158 = ~w32012;// level 8
assign po06159 = ~w32015;// level 8
assign po06160 = ~w32018;// level 8
assign po06161 = ~w32021;// level 8
assign po06162 = ~w32024;// level 8
assign po06163 = ~w32027;// level 8
assign po06164 = ~w32030;// level 8
assign po06165 = ~w32033;// level 8
assign po06166 = ~w32036;// level 8
assign po06167 = ~w32039;// level 8
assign po06168 = ~w32042;// level 8
assign po06169 = ~w32045;// level 8
assign po06170 = ~w32048;// level 8
assign po06171 = ~w32051;// level 8
assign po06172 = ~w32054;// level 8
assign po06173 = ~w32057;// level 8
assign po06174 = ~w32060;// level 8
assign po06175 = ~w32063;// level 8
assign po06176 = ~w32066;// level 8
assign po06177 = ~w32069;// level 8
assign po06178 = ~w32072;// level 8
assign po06179 = ~w32075;// level 8
assign po06180 = ~w32078;// level 8
assign po06181 = ~w32081;// level 8
assign po06182 = ~w32084;// level 8
assign po06183 = ~w32087;// level 8
assign po06184 = ~w32090;// level 8
assign po06185 = ~w32093;// level 8
assign po06186 = ~w32096;// level 8
assign po06187 = ~w32099;// level 8
assign po06188 = ~w32102;// level 8
assign po06189 = ~w32105;// level 8
assign po06190 = ~w32108;// level 8
assign po06191 = ~w32111;// level 8
assign po06192 = ~w32114;// level 8
assign po06193 = ~w32117;// level 8
assign po06194 = ~w32120;// level 8
assign po06195 = ~w32123;// level 8
assign po06196 = ~w32126;// level 8
assign po06197 = ~w32129;// level 8
assign po06198 = ~w32132;// level 8
assign po06199 = ~w32135;// level 8
assign po06200 = ~w32138;// level 7
assign po06201 = ~w32141;// level 7
assign po06202 = ~w32144;// level 7
assign po06203 = ~w32148;// level 8
assign po06204 = ~w32151;// level 7
assign po06205 = ~w32154;// level 8
assign po06206 = ~w32157;// level 7
assign po06207 = ~w32160;// level 7
assign po06208 = ~w32163;// level 8
assign po06209 = ~w32166;// level 8
assign po06210 = ~w32169;// level 8
assign po06211 = ~w32172;// level 8
assign po06212 = ~w32175;// level 8
assign po06213 = ~w32178;// level 8
assign po06214 = ~w32181;// level 8
assign po06215 = ~w32184;// level 8
assign po06216 = ~w32187;// level 8
assign po06217 = ~w32190;// level 8
assign po06218 = ~w32193;// level 8
assign po06219 = ~w32196;// level 8
assign po06220 = ~w32199;// level 8
assign po06221 = ~w32202;// level 8
assign po06222 = ~w32205;// level 8
assign po06223 = ~w32208;// level 8
assign po06224 = ~w32211;// level 8
assign po06225 = ~w32214;// level 8
assign po06226 = ~w32217;// level 8
assign po06227 = ~w32220;// level 8
assign po06228 = ~w32223;// level 8
assign po06229 = ~w32226;// level 8
assign po06230 = ~w32229;// level 8
assign po06231 = ~w32232;// level 8
assign po06232 = ~w32235;// level 8
assign po06233 = ~w32238;// level 8
assign po06234 = ~w32242;// level 8
assign po06235 = ~w32245;// level 8
assign po06236 = ~w32248;// level 8
assign po06237 = ~w32251;// level 8
assign po06238 = ~w32254;// level 8
assign po06239 = ~w32257;// level 8
assign po06240 = ~w32260;// level 8
assign po06241 = ~w32263;// level 8
assign po06242 = ~w32266;// level 8
assign po06243 = ~w32269;// level 8
assign po06244 = ~w32272;// level 8
assign po06245 = ~w32275;// level 8
assign po06246 = ~w32278;// level 8
assign po06247 = ~w32281;// level 8
assign po06248 = ~w32284;// level 8
assign po06249 = ~w32287;// level 8
assign po06250 = ~w32291;// level 8
assign po06251 = ~w32294;// level 8
assign po06252 = ~w32297;// level 8
assign po06253 = ~w32300;// level 8
assign po06254 = ~w32303;// level 8
assign po06255 = ~w32306;// level 8
assign po06256 = ~w32309;// level 8
assign po06257 = ~w32312;// level 8
assign po06258 = ~w32315;// level 8
assign po06259 = ~w32318;// level 8
assign po06260 = ~w32321;// level 8
assign po06261 = ~w32324;// level 8
assign po06262 = ~w32327;// level 8
assign po06263 = ~w32330;// level 8
assign po06264 = ~w32333;// level 8
assign po06265 = ~w32336;// level 8
assign po06266 = ~w32339;// level 8
assign po06267 = ~w32342;// level 8
assign po06268 = ~w32345;// level 8
assign po06269 = ~w32348;// level 8
assign po06270 = ~w32351;// level 8
assign po06271 = ~w32354;// level 8
assign po06272 = ~w32357;// level 8
assign po06273 = ~w32360;// level 8
assign po06274 = ~w32363;// level 8
assign po06275 = ~w32366;// level 8
assign po06276 = ~w32369;// level 8
assign po06277 = ~w32372;// level 8
assign po06278 = ~w32375;// level 8
assign po06279 = ~w32378;// level 8
assign po06280 = ~w32381;// level 8
assign po06281 = ~w32384;// level 8
assign po06282 = ~w32387;// level 8
assign po06283 = ~w32390;// level 8
assign po06284 = ~w32393;// level 8
assign po06285 = ~w32396;// level 8
assign po06286 = ~w32399;// level 8
assign po06287 = ~w32402;// level 8
assign po06288 = ~w32405;// level 8
assign po06289 = ~w32408;// level 8
assign po06290 = ~w32411;// level 8
assign po06291 = ~w32414;// level 8
assign po06292 = ~w32418;// level 8
assign po06293 = ~w32421;// level 8
assign po06294 = ~w32425;// level 8
assign po06295 = ~w32428;// level 8
assign po06296 = ~w32431;// level 8
assign po06297 = ~w32434;// level 8
assign po06298 = ~w32437;// level 8
assign po06299 = ~w32440;// level 8
assign po06300 = ~w32443;// level 8
assign po06301 = ~w32446;// level 8
assign po06302 = ~w32449;// level 8
assign po06303 = ~w32452;// level 8
assign po06304 = ~w32455;// level 8
assign po06305 = ~w32459;// level 8
assign po06306 = ~w32462;// level 8
assign po06307 = ~w32465;// level 8
assign po06308 = ~w32469;// level 8
assign po06309 = ~w32472;// level 8
assign po06310 = ~w32475;// level 8
assign po06311 = ~w32478;// level 8
assign po06312 = ~w32481;// level 8
assign po06313 = ~w32484;// level 8
assign po06314 = ~w32487;// level 8
assign po06315 = ~w32490;// level 8
assign po06316 = ~w32493;// level 8
assign po06317 = ~w32496;// level 8
assign po06318 = ~w32500;// level 8
assign po06319 = ~w32503;// level 8
assign po06320 = ~w32507;// level 8
assign po06321 = ~w32510;// level 8
assign po06322 = ~w32513;// level 8
assign po06323 = ~w32516;// level 8
assign po06324 = ~w32519;// level 8
assign po06325 = ~w32522;// level 8
assign po06326 = ~w32525;// level 8
assign po06327 = ~w32528;// level 8
assign po06328 = ~w32531;// level 8
assign po06329 = ~w32534;// level 8
assign po06330 = ~w32537;// level 8
assign po06331 = ~w32541;// level 8
assign po06332 = ~w32544;// level 8
assign po06333 = ~w32547;// level 8
assign po06334 = ~w32550;// level 8
assign po06335 = ~w32553;// level 8
assign po06336 = ~w32556;// level 8
assign po06337 = ~w32559;// level 8
assign po06338 = ~w32562;// level 8
assign po06339 = ~w32565;// level 8
assign po06340 = ~w32569;// level 8
assign po06341 = ~w32572;// level 8
assign po06342 = ~w32575;// level 8
assign po06343 = ~w32578;// level 8
assign po06344 = ~w32581;// level 8
assign po06345 = ~w32584;// level 8
assign po06346 = ~w32587;// level 8
assign po06347 = ~w32590;// level 8
assign po06348 = ~w32593;// level 8
assign po06349 = ~w32596;// level 8
assign po06350 = ~w32599;// level 8
assign po06351 = ~w32602;// level 8
assign po06352 = ~w32605;// level 8
assign po06353 = ~w32608;// level 8
assign po06354 = ~w32611;// level 8
assign po06355 = ~w32614;// level 8
assign po06356 = ~w32617;// level 8
assign po06357 = ~w32620;// level 8
assign po06358 = ~w32623;// level 8
assign po06359 = ~w32626;// level 8
assign po06360 = ~w32629;// level 8
assign po06361 = ~w32632;// level 8
assign po06362 = ~w32635;// level 8
assign po06363 = ~w32638;// level 8
assign po06364 = ~w32641;// level 8
assign po06365 = ~w32644;// level 8
assign po06366 = ~w32647;// level 8
assign po06367 = ~w32650;// level 8
assign po06368 = ~w32653;// level 8
assign po06369 = ~w32656;// level 8
assign po06370 = ~w32659;// level 8
assign po06371 = ~w32662;// level 8
assign po06372 = ~w32665;// level 8
assign po06373 = ~w32668;// level 8
assign po06374 = ~w32671;// level 8
assign po06375 = ~w32674;// level 8
assign po06376 = ~w32677;// level 8
assign po06377 = ~w32680;// level 8
assign po06378 = ~w32683;// level 8
assign po06379 = ~w32686;// level 8
assign po06380 = ~w32689;// level 8
assign po06381 = ~w32692;// level 8
assign po06382 = ~w32695;// level 8
assign po06383 = ~w32698;// level 8
assign po06384 = ~w32701;// level 8
assign po06385 = ~w32704;// level 8
assign po06386 = ~w32707;// level 8
assign po06387 = ~w32710;// level 8
assign po06388 = ~w32713;// level 8
assign po06389 = ~w32716;// level 8
assign po06390 = ~w32719;// level 8
assign po06391 = ~w32722;// level 8
assign po06392 = ~w32725;// level 8
assign po06393 = ~w32728;// level 8
assign po06394 = ~w32731;// level 8
assign po06395 = ~w32734;// level 8
assign po06396 = ~w32737;// level 8
assign po06397 = ~w32740;// level 8
assign po06398 = ~w32743;// level 8
assign po06399 = ~w32746;// level 8
assign po06400 = ~w32749;// level 8
assign po06401 = ~w32752;// level 8
assign po06402 = ~w32755;// level 8
assign po06403 = ~w32758;// level 8
assign po06404 = ~w32761;// level 8
assign po06405 = ~w32764;// level 8
assign po06406 = ~w32767;// level 8
assign po06407 = ~w32770;// level 8
assign po06408 = ~w32773;// level 8
assign po06409 = ~w32776;// level 8
assign po06410 = ~w32779;// level 8
assign po06411 = ~w32782;// level 8
assign po06412 = ~w32785;// level 8
assign po06413 = ~w32788;// level 8
assign po06414 = ~w32791;// level 8
assign po06415 = ~w32794;// level 8
assign po06416 = ~w32797;// level 8
assign po06417 = ~w32800;// level 8
assign po06418 = ~w32803;// level 8
assign po06419 = ~w32806;// level 8
assign po06420 = ~w32809;// level 8
assign po06421 = ~w32812;// level 8
assign po06422 = ~w32815;// level 8
assign po06423 = ~w32818;// level 8
assign po06424 = ~w32821;// level 8
assign po06425 = ~w32824;// level 8
assign po06426 = ~w32827;// level 8
assign po06427 = ~w32830;// level 8
assign po06428 = ~w32833;// level 8
assign po06429 = ~w32836;// level 8
assign po06430 = ~w32839;// level 8
assign po06431 = ~w32842;// level 8
assign po06432 = ~w32845;// level 8
assign po06433 = ~w32848;// level 8
assign po06434 = ~w32851;// level 8
assign po06435 = ~w32854;// level 8
assign po06436 = ~w32857;// level 8
assign po06437 = ~w32860;// level 8
assign po06438 = ~w32863;// level 8
assign po06439 = ~w32866;// level 8
assign po06440 = ~w32869;// level 8
assign po06441 = ~w32872;// level 8
assign po06442 = ~w32875;// level 8
assign po06443 = ~w32878;// level 8
assign po06444 = ~w32881;// level 8
assign po06445 = ~w32884;// level 8
assign po06446 = ~w32887;// level 8
assign po06447 = ~w32890;// level 8
assign po06448 = ~w32893;// level 8
assign po06449 = ~w32896;// level 8
assign po06450 = ~w32899;// level 8
assign po06451 = ~w32903;// level 8
assign po06452 = ~w32906;// level 8
assign po06453 = ~w32909;// level 8
assign po06454 = ~w32912;// level 8
assign po06455 = ~w32915;// level 8
assign po06456 = ~w32918;// level 8
assign po06457 = ~w32921;// level 8
assign po06458 = ~w32924;// level 8
assign po06459 = ~w32927;// level 8
assign po06460 = ~w32930;// level 8
assign po06461 = ~w32933;// level 8
assign po06462 = ~w32936;// level 8
assign po06463 = ~w32939;// level 8
assign po06464 = ~w32942;// level 8
assign po06465 = ~w32945;// level 8
assign po06466 = ~w32948;// level 8
assign po06467 = ~w32951;// level 8
assign po06468 = ~w32954;// level 8
assign po06469 = ~w32957;// level 8
assign po06470 = ~w32960;// level 8
assign po06471 = ~w32963;// level 8
assign po06472 = ~w32966;// level 8
assign po06473 = ~w32969;// level 8
assign po06474 = ~w32972;// level 8
assign po06475 = ~w32975;// level 8
assign po06476 = ~w32978;// level 8
assign po06477 = ~w32981;// level 8
assign po06478 = ~w32984;// level 8
assign po06479 = ~w32987;// level 8
assign po06480 = ~w32990;// level 8
assign po06481 = ~w32993;// level 8
assign po06482 = ~w32996;// level 8
assign po06483 = ~w32999;// level 8
assign po06484 = ~w33002;// level 8
assign po06485 = ~w33005;// level 8
assign po06486 = ~w33008;// level 8
assign po06487 = ~w33011;// level 8
assign po06488 = ~w33014;// level 8
assign po06489 = ~w33017;// level 8
assign po06490 = ~w33020;// level 8
assign po06491 = ~w33023;// level 8
assign po06492 = ~w33026;// level 8
assign po06493 = ~w33029;// level 8
assign po06494 = ~w33032;// level 8
assign po06495 = ~w33035;// level 8
assign po06496 = ~w33038;// level 8
assign po06497 = ~w33041;// level 8
assign po06498 = ~w33044;// level 8
assign po06499 = ~w33047;// level 8
assign po06500 = ~w33050;// level 8
assign po06501 = ~w33053;// level 8
assign po06502 = ~w33056;// level 8
assign po06503 = ~w33059;// level 8
assign po06504 = ~w33062;// level 8
assign po06505 = ~w33065;// level 8
assign po06506 = ~w33068;// level 8
assign po06507 = ~w33071;// level 8
assign po06508 = ~w33074;// level 8
assign po06509 = ~w33077;// level 8
assign po06510 = ~w33080;// level 8
assign po06511 = ~w33083;// level 8
assign po06512 = ~w33086;// level 8
assign po06513 = ~w33089;// level 8
assign po06514 = ~w33092;// level 8
assign po06515 = ~w33095;// level 8
assign po06516 = ~w33098;// level 8
assign po06517 = ~w33101;// level 8
assign po06518 = ~w33104;// level 8
assign po06519 = ~w33107;// level 8
assign po06520 = ~w33110;// level 8
assign po06521 = ~w33113;// level 8
assign po06522 = ~w33116;// level 8
assign po06523 = ~w33119;// level 8
assign po06524 = ~w33122;// level 8
assign po06525 = ~w33125;// level 8
assign po06526 = ~w33128;// level 8
assign po06527 = ~w33131;// level 8
assign po06528 = ~w33134;// level 8
assign po06529 = ~w33137;// level 8
assign po06530 = ~w33140;// level 8
assign po06531 = ~w33143;// level 8
assign po06532 = ~w33146;// level 8
assign po06533 = ~w33149;// level 8
assign po06534 = ~w33152;// level 8
assign po06535 = ~w33155;// level 8
assign po06536 = ~w33158;// level 8
assign po06537 = ~w33161;// level 8
assign po06538 = ~w33164;// level 8
assign po06539 = ~w33167;// level 8
assign po06540 = ~w33170;// level 8
assign po06541 = ~w33173;// level 7
assign po06542 = ~w33176;// level 7
assign po06543 = ~w33179;// level 7
assign po06544 = ~w33182;// level 7
assign po06545 = ~w33185;// level 8
assign po06546 = ~w33189;// level 8
assign po06547 = ~w33193;// level 8
assign po06548 = ~w33197;// level 8
assign po06549 = ~w33200;// level 8
assign po06550 = ~w33203;// level 8
assign po06551 = ~w33206;// level 8
assign po06552 = ~w33209;// level 8
assign po06553 = ~w33212;// level 8
assign po06554 = ~w33215;// level 8
assign po06555 = ~w33218;// level 8
assign po06556 = ~w33221;// level 8
assign po06557 = ~w33224;// level 8
assign po06558 = ~w33227;// level 8
assign po06559 = ~w33231;// level 8
assign po06560 = ~w33234;// level 8
assign po06561 = ~w33237;// level 8
assign po06562 = ~w33240;// level 8
assign po06563 = ~w33243;// level 8
assign po06564 = ~w33246;// level 8
assign po06565 = ~w33249;// level 8
assign po06566 = ~w33252;// level 8
assign po06567 = ~w33255;// level 8
assign po06568 = ~w33259;// level 8
assign po06569 = ~w33262;// level 8
assign po06570 = ~w33265;// level 8
assign po06571 = ~w33268;// level 8
assign po06572 = ~w33271;// level 8
assign po06573 = ~w33274;// level 8
assign po06574 = ~w33278;// level 8
assign po06575 = ~w33281;// level 8
assign po06576 = ~w33284;// level 8
assign po06577 = ~w33287;// level 8
assign po06578 = ~w33290;// level 8
assign po06579 = ~w33293;// level 8
assign po06580 = ~w33296;// level 8
assign po06581 = ~w33300;// level 8
assign po06582 = ~w33303;// level 8
assign po06583 = ~w33306;// level 8
assign po06584 = ~w33309;// level 8
assign po06585 = ~w33312;// level 8
assign po06586 = ~w33315;// level 8
assign po06587 = ~w33318;// level 8
assign po06588 = ~w33321;// level 8
assign po06589 = ~w33324;// level 8
assign po06590 = ~w33327;// level 8
assign po06591 = ~w33330;// level 8
assign po06592 = ~w33333;// level 8
assign po06593 = ~w33337;// level 8
assign po06594 = ~w33340;// level 8
assign po06595 = ~w33343;// level 8
assign po06596 = ~w33346;// level 8
assign po06597 = ~w33349;// level 8
assign po06598 = ~w33352;// level 8
assign po06599 = ~w33355;// level 8
assign po06600 = ~w33358;// level 8
assign po06601 = ~w33361;// level 8
assign po06602 = ~w33364;// level 8
assign po06603 = ~w33367;// level 8
assign po06604 = ~w33370;// level 8
assign po06605 = ~w33373;// level 8
assign po06606 = ~w33376;// level 8
assign po06607 = ~w33379;// level 8
assign po06608 = ~w33382;// level 8
assign po06609 = ~w33385;// level 8
assign po06610 = ~w33388;// level 8
assign po06611 = ~w33391;// level 8
assign po06612 = ~w33394;// level 8
assign po06613 = ~w33397;// level 8
assign po06614 = ~w33400;// level 8
assign po06615 = ~w33403;// level 8
assign po06616 = ~w33406;// level 8
assign po06617 = ~w33409;// level 8
assign po06618 = ~w33412;// level 8
assign po06619 = ~w33415;// level 8
assign po06620 = ~w33418;// level 8
assign po06621 = ~w33421;// level 8
assign po06622 = ~w33424;// level 8
assign po06623 = ~w33427;// level 8
assign po06624 = ~w33430;// level 8
assign po06625 = ~w33433;// level 8
assign po06626 = ~w33437;// level 8
assign po06627 = ~w33440;// level 8
assign po06628 = ~w33443;// level 8
assign po06629 = ~w33446;// level 8
assign po06630 = ~w33449;// level 8
assign po06631 = ~w33452;// level 8
assign po06632 = ~w33455;// level 8
assign po06633 = ~w33458;// level 8
assign po06634 = ~w33461;// level 8
assign po06635 = ~w33464;// level 8
assign po06636 = ~w33467;// level 8
assign po06637 = ~w33470;// level 8
assign po06638 = ~w33473;// level 8
assign po06639 = ~w33476;// level 8
assign po06640 = ~w33479;// level 8
assign po06641 = ~w33482;// level 8
assign po06642 = ~w33485;// level 8
assign po06643 = ~w33488;// level 8
assign po06644 = ~w33491;// level 8
assign po06645 = ~w33494;// level 8
assign po06646 = ~w33497;// level 8
assign po06647 = ~w33500;// level 8
assign po06648 = ~w33503;// level 8
assign po06649 = ~w33506;// level 8
assign po06650 = ~w33509;// level 8
assign po06651 = ~w33512;// level 8
assign po06652 = ~w33515;// level 8
assign po06653 = ~w33518;// level 8
assign po06654 = ~w33521;// level 8
assign po06655 = ~w33524;// level 8
assign po06656 = ~w33527;// level 8
assign po06657 = ~w33530;// level 8
assign po06658 = ~w33533;// level 8
assign po06659 = ~w33536;// level 8
assign po06660 = ~w33539;// level 8
assign po06661 = ~w33542;// level 8
assign po06662 = ~w33545;// level 8
assign po06663 = ~w33548;// level 8
assign po06664 = ~w33551;// level 8
assign po06665 = ~w33554;// level 8
assign po06666 = ~w33557;// level 8
assign po06667 = ~w33560;// level 8
assign po06668 = ~w33563;// level 8
assign po06669 = ~w33566;// level 8
assign po06670 = ~w33569;// level 8
assign po06671 = ~w33572;// level 8
assign po06672 = ~w33575;// level 8
assign po06673 = ~w33578;// level 8
assign po06674 = ~w33581;// level 8
assign po06675 = ~w33584;// level 8
assign po06676 = ~w33587;// level 8
assign po06677 = ~w33590;// level 8
assign po06678 = ~w33593;// level 8
assign po06679 = ~w33596;// level 8
assign po06680 = ~w33599;// level 8
assign po06681 = ~w33602;// level 8
assign po06682 = ~w33605;// level 8
assign po06683 = ~w33608;// level 8
assign po06684 = ~w33611;// level 8
assign po06685 = ~w33614;// level 8
assign po06686 = ~w33617;// level 8
assign po06687 = ~w33620;// level 8
assign po06688 = ~w33623;// level 8
assign po06689 = ~w33626;// level 8
assign po06690 = ~w33629;// level 8
assign po06691 = ~w33632;// level 8
assign po06692 = ~w33635;// level 7
assign po06693 = ~w33638;// level 8
assign po06694 = ~w33641;// level 7
assign po06695 = ~w33644;// level 7
assign po06696 = ~w33647;// level 7
assign po06697 = ~w33650;// level 7
assign po06698 = ~w33653;// level 7
assign po06699 = ~w33656;// level 8
assign po06700 = ~w33659;// level 8
assign po06701 = ~w33662;// level 8
assign po06702 = ~w33665;// level 8
assign po06703 = ~w33668;// level 8
assign po06704 = ~w33671;// level 8
assign po06705 = ~w33674;// level 8
assign po06706 = ~w33677;// level 8
assign po06707 = ~w33680;// level 8
assign po06708 = ~w33683;// level 8
assign po06709 = ~w33686;// level 8
assign po06710 = ~w33689;// level 8
assign po06711 = ~w33692;// level 8
assign po06712 = ~w33695;// level 8
assign po06713 = ~w33698;// level 8
assign po06714 = ~w33701;// level 8
assign po06715 = ~w33704;// level 8
assign po06716 = ~w33707;// level 8
assign po06717 = ~w33710;// level 8
assign po06718 = ~w33713;// level 8
assign po06719 = ~w33716;// level 8
assign po06720 = ~w33719;// level 8
assign po06721 = ~w33722;// level 8
assign po06722 = ~w33725;// level 8
assign po06723 = ~w33728;// level 8
assign po06724 = ~w33731;// level 8
assign po06725 = ~w33734;// level 8
assign po06726 = ~w33737;// level 8
assign po06727 = ~w33740;// level 8
assign po06728 = ~w33743;// level 8
assign po06729 = ~w33746;// level 8
assign po06730 = ~w33750;// level 8
assign po06731 = ~w33753;// level 8
assign po06732 = ~w33756;// level 8
assign po06733 = ~w33759;// level 8
assign po06734 = ~w33762;// level 8
assign po06735 = ~w33765;// level 8
assign po06736 = ~w33768;// level 8
assign po06737 = ~w33771;// level 8
assign po06738 = ~w33774;// level 8
assign po06739 = ~w33777;// level 8
assign po06740 = ~w33780;// level 8
assign po06741 = ~w33783;// level 8
assign po06742 = ~w33786;// level 8
assign po06743 = ~w33789;// level 8
assign po06744 = ~w33792;// level 8
assign po06745 = ~w33795;// level 8
assign po06746 = ~w33798;// level 8
assign po06747 = ~w33801;// level 8
assign po06748 = ~w33804;// level 8
assign po06749 = ~w33807;// level 8
assign po06750 = ~w33810;// level 8
assign po06751 = ~w33813;// level 8
assign po06752 = ~w33816;// level 8
assign po06753 = ~w33819;// level 8
assign po06754 = ~w33822;// level 8
assign po06755 = ~w33825;// level 8
assign po06756 = ~w33828;// level 8
assign po06757 = ~w33832;// level 8
assign po06758 = ~w33835;// level 8
assign po06759 = ~w33838;// level 8
assign po06760 = ~w33841;// level 8
assign po06761 = ~w33844;// level 8
assign po06762 = ~w33847;// level 8
assign po06763 = ~w33850;// level 8
assign po06764 = ~w33853;// level 8
assign po06765 = ~w33856;// level 7
assign po06766 = ~w33859;// level 7
assign po06767 = ~w33862;// level 7
assign po06768 = ~w33865;// level 7
assign po06769 = ~w33868;// level 7
assign po06770 = ~w33871;// level 7
assign po06771 = ~w33874;// level 7
assign po06772 = ~w33877;// level 7
assign po06773 = ~w33880;// level 7
assign po06774 = ~w33883;// level 7
assign po06775 = ~w33886;// level 7
assign po06776 = ~w33889;// level 7
assign po06777 = ~w33892;// level 7
assign po06778 = ~w33895;// level 7
assign po06779 = ~w33898;// level 7
assign po06780 = ~w33901;// level 7
assign po06781 = ~w33904;// level 7
assign po06782 = ~w33907;// level 7
assign po06783 = ~w33910;// level 7
assign po06784 = ~w33913;// level 8
assign po06785 = ~w33917;// level 8
assign po06786 = ~w33920;// level 8
assign po06787 = ~w33923;// level 8
assign po06788 = ~w33926;// level 8
assign po06789 = ~w33929;// level 8
assign po06790 = ~w33932;// level 8
assign po06791 = ~w33935;// level 8
assign po06792 = ~w33939;// level 8
assign po06793 = ~w33942;// level 8
assign po06794 = ~w33945;// level 8
assign po06795 = ~w33948;// level 8
assign po06796 = ~w33951;// level 8
assign po06797 = ~w33954;// level 8
assign po06798 = ~w33958;// level 8
assign po06799 = ~w33961;// level 8
assign po06800 = ~w33964;// level 8
assign po06801 = ~w33967;// level 8
assign po06802 = ~w33971;// level 8
assign po06803 = ~w33974;// level 8
assign po06804 = ~w33977;// level 8
assign po06805 = ~w33980;// level 8
assign po06806 = ~w33983;// level 8
assign po06807 = ~w33987;// level 8
assign po06808 = ~w33990;// level 8
assign po06809 = ~w33993;// level 8
assign po06810 = ~w33996;// level 8
assign po06811 = ~w33999;// level 8
assign po06812 = ~w34002;// level 8
assign po06813 = ~w34005;// level 8
assign po06814 = ~w34008;// level 8
assign po06815 = ~w34011;// level 8
assign po06816 = ~w34015;// level 8
assign po06817 = ~w34018;// level 8
assign po06818 = ~w34021;// level 8
assign po06819 = ~w34024;// level 8
assign po06820 = ~w34027;// level 8
assign po06821 = ~w34030;// level 8
assign po06822 = ~w34033;// level 8
assign po06823 = ~w34036;// level 8
assign po06824 = ~w34039;// level 8
assign po06825 = ~w34042;// level 8
assign po06826 = ~w34045;// level 8
assign po06827 = ~w34048;// level 8
assign po06828 = ~w34051;// level 8
assign po06829 = ~w34054;// level 8
assign po06830 = ~w34057;// level 8
assign po06831 = ~w34060;// level 8
assign po06832 = ~w34063;// level 8
assign po06833 = ~w34066;// level 8
assign po06834 = ~w34069;// level 8
assign po06835 = ~w34073;// level 8
assign po06836 = ~w34076;// level 8
assign po06837 = ~w34079;// level 8
assign po06838 = ~w34082;// level 8
assign po06839 = ~w34085;// level 8
assign po06840 = ~w34088;// level 8
assign po06841 = ~w34091;// level 8
assign po06842 = ~w34094;// level 8
assign po06843 = ~w34097;// level 8
assign po06844 = ~w34100;// level 8
assign po06845 = ~w34103;// level 8
assign po06846 = ~w34106;// level 8
assign po06847 = ~w34109;// level 8
assign po06848 = ~w34112;// level 8
assign po06849 = ~w34115;// level 8
assign po06850 = ~w34118;// level 8
assign po06851 = ~w34121;// level 8
assign po06852 = ~w34124;// level 8
assign po06853 = ~w34127;// level 8
assign po06854 = ~w34130;// level 8
assign po06855 = ~w34133;// level 8
assign po06856 = ~w34136;// level 8
assign po06857 = ~w34139;// level 8
assign po06858 = ~w34142;// level 8
assign po06859 = ~w34145;// level 8
assign po06860 = ~w34148;// level 8
assign po06861 = ~w34151;// level 8
assign po06862 = ~w34154;// level 8
assign po06863 = ~w34157;// level 8
assign po06864 = ~w34160;// level 8
assign po06865 = ~w34163;// level 8
assign po06866 = ~w34166;// level 8
assign po06867 = ~w34169;// level 8
assign po06868 = ~w34172;// level 8
assign po06869 = ~w34175;// level 8
assign po06870 = ~w34178;// level 8
assign po06871 = ~w34181;// level 8
assign po06872 = ~w34184;// level 8
assign po06873 = ~w34187;// level 8
assign po06874 = ~w34190;// level 8
assign po06875 = ~w34193;// level 8
assign po06876 = ~w34196;// level 8
assign po06877 = ~w34199;// level 8
assign po06878 = ~w34202;// level 8
assign po06879 = ~w34205;// level 8
assign po06880 = ~w34208;// level 8
assign po06881 = ~w34211;// level 8
assign po06882 = ~w34214;// level 8
assign po06883 = ~w34217;// level 8
assign po06884 = ~w34220;// level 8
assign po06885 = ~w34223;// level 8
assign po06886 = ~w34226;// level 8
assign po06887 = ~w34229;// level 8
assign po06888 = ~w34232;// level 8
assign po06889 = ~w34235;// level 8
assign po06890 = ~w34238;// level 8
assign po06891 = ~w34241;// level 8
assign po06892 = ~w34244;// level 8
assign po06893 = ~w34247;// level 8
assign po06894 = ~w34250;// level 8
assign po06895 = ~w34253;// level 8
assign po06896 = ~w34256;// level 7
assign po06897 = ~w34259;// level 7
assign po06898 = ~w34262;// level 7
assign po06899 = ~w34265;// level 8
assign po06900 = ~w34268;// level 8
assign po06901 = ~w34271;// level 7
assign po06902 = ~w34275;// level 8
assign po06903 = ~w34278;// level 8
assign po06904 = ~w34281;// level 8
assign po06905 = ~w34284;// level 8
assign po06906 = ~w34287;// level 8
assign po06907 = ~w34290;// level 8
assign po06908 = ~w34293;// level 8
assign po06909 = ~w34296;// level 8
assign po06910 = ~w34299;// level 8
assign po06911 = ~w34302;// level 8
assign po06912 = ~w34305;// level 8
assign po06913 = ~w34308;// level 8
assign po06914 = ~w34311;// level 8
assign po06915 = ~w34315;// level 8
assign po06916 = ~w34318;// level 8
assign po06917 = ~w34321;// level 8
assign po06918 = ~w34324;// level 8
assign po06919 = ~w34327;// level 8
assign po06920 = ~w34330;// level 8
assign po06921 = ~w34333;// level 8
assign po06922 = ~w34336;// level 8
assign po06923 = ~w34339;// level 8
assign po06924 = ~w34342;// level 8
assign po06925 = ~w34345;// level 8
assign po06926 = ~w34348;// level 8
assign po06927 = ~w34351;// level 8
assign po06928 = ~w34354;// level 8
assign po06929 = ~w34357;// level 8
assign po06930 = ~w34360;// level 8
assign po06931 = ~w34363;// level 8
assign po06932 = ~w34366;// level 8
assign po06933 = ~w34369;// level 8
assign po06934 = ~w34372;// level 8
assign po06935 = ~w34375;// level 8
assign po06936 = ~w34378;// level 8
assign po06937 = ~w34381;// level 8
assign po06938 = ~w34384;// level 8
assign po06939 = ~w34387;// level 8
assign po06940 = ~w34390;// level 8
assign po06941 = ~w34393;// level 8
assign po06942 = ~w34396;// level 8
assign po06943 = ~w34399;// level 8
assign po06944 = ~w34402;// level 8
assign po06945 = ~w34405;// level 8
assign po06946 = ~w34408;// level 8
assign po06947 = ~w34411;// level 8
assign po06948 = ~w34414;// level 8
assign po06949 = ~w34417;// level 8
assign po06950 = ~w34420;// level 8
assign po06951 = ~w34423;// level 8
assign po06952 = ~w34426;// level 8
assign po06953 = ~w34429;// level 8
assign po06954 = ~w34433;// level 8
assign po06955 = ~w34436;// level 7
assign po06956 = ~w34439;// level 7
assign po06957 = ~w34442;// level 8
assign po06958 = ~w34445;// level 7
assign po06959 = ~w34448;// level 8
assign po06960 = ~w34451;// level 8
assign po06961 = ~w34454;// level 8
assign po06962 = ~w34457;// level 7
assign po06963 = ~w34460;// level 8
assign po06964 = ~w34463;// level 8
assign po06965 = ~w34466;// level 8
assign po06966 = ~w34469;// level 8
assign po06967 = ~w34472;// level 7
assign po06968 = ~w34475;// level 7
assign po06969 = ~w34478;// level 7
assign po06970 = ~w34481;// level 7
assign po06971 = ~w34484;// level 8
assign po06972 = ~w34487;// level 7
assign po06973 = ~w34490;// level 7
assign po06974 = ~w34494;// level 8
assign po06975 = ~w34497;// level 8
assign po06976 = ~w34500;// level 8
assign po06977 = ~w34503;// level 8
assign po06978 = ~w34506;// level 8
assign po06979 = ~w34509;// level 8
assign po06980 = ~w34513;// level 8
assign po06981 = ~w34517;// level 8
assign po06982 = ~w34520;// level 8
assign po06983 = ~w34523;// level 8
assign po06984 = ~w34526;// level 8
assign po06985 = ~w34529;// level 8
assign po06986 = ~w34532;// level 8
assign po06987 = ~w34535;// level 8
assign po06988 = ~w34538;// level 8
assign po06989 = ~w34541;// level 8
assign po06990 = ~w34544;// level 8
assign po06991 = ~w34547;// level 8
assign po06992 = ~w34550;// level 8
assign po06993 = ~w34554;// level 8
assign po06994 = ~w34557;// level 8
assign po06995 = ~w34560;// level 8
assign po06996 = ~w34563;// level 8
assign po06997 = ~w34566;// level 8
assign po06998 = ~w34569;// level 8
assign po06999 = ~w34572;// level 8
assign po07000 = ~w34576;// level 8
assign po07001 = ~w34579;// level 8
assign po07002 = ~w34582;// level 8
assign po07003 = ~w34585;// level 8
assign po07004 = ~w34588;// level 8
assign po07005 = ~w34591;// level 8
assign po07006 = ~w34595;// level 8
assign po07007 = ~w34598;// level 8
assign po07008 = ~w34601;// level 8
assign po07009 = ~w34604;// level 8
assign po07010 = ~w34607;// level 8
assign po07011 = ~w34610;// level 8
assign po07012 = ~w34613;// level 8
assign po07013 = ~w34616;// level 8
assign po07014 = ~w34619;// level 8
assign po07015 = ~w34622;// level 8
assign po07016 = ~w34625;// level 8
assign po07017 = ~w34628;// level 8
assign po07018 = ~w34632;// level 8
assign po07019 = ~w34635;// level 8
assign po07020 = ~w34638;// level 8
assign po07021 = ~w34641;// level 8
assign po07022 = ~w34644;// level 8
assign po07023 = ~w34647;// level 8
assign po07024 = ~w34650;// level 8
assign po07025 = ~w34653;// level 8
assign po07026 = ~w34656;// level 8
assign po07027 = ~w34659;// level 8
assign po07028 = ~w34662;// level 8
assign po07029 = ~w34665;// level 8
assign po07030 = ~w34668;// level 8
assign po07031 = ~w34671;// level 8
assign po07032 = ~w34674;// level 8
assign po07033 = ~w34677;// level 8
assign po07034 = ~w34680;// level 8
assign po07035 = ~w34683;// level 8
assign po07036 = ~w34686;// level 8
assign po07037 = ~w34689;// level 8
assign po07038 = ~w34692;// level 8
assign po07039 = ~w34695;// level 8
assign po07040 = ~w34698;// level 8
assign po07041 = ~w34701;// level 8
assign po07042 = ~w34704;// level 8
assign po07043 = ~w34707;// level 8
assign po07044 = ~w34710;// level 8
assign po07045 = ~w34713;// level 8
assign po07046 = ~w34716;// level 8
assign po07047 = ~w34719;// level 8
assign po07048 = ~w34722;// level 8
assign po07049 = ~w34725;// level 8
assign po07050 = ~w34728;// level 8
assign po07051 = ~w34731;// level 8
assign po07052 = ~w34734;// level 8
assign po07053 = ~w34737;// level 8
assign po07054 = ~w34740;// level 8
assign po07055 = ~w34743;// level 8
assign po07056 = ~w34746;// level 8
assign po07057 = ~w34749;// level 8
assign po07058 = ~w34752;// level 8
assign po07059 = ~w34755;// level 8
assign po07060 = ~w34758;// level 8
assign po07061 = ~w34761;// level 8
assign po07062 = ~w34764;// level 8
assign po07063 = ~w34767;// level 8
assign po07064 = ~w34770;// level 8
assign po07065 = ~w34773;// level 8
assign po07066 = ~w34776;// level 8
assign po07067 = ~w34779;// level 8
assign po07068 = ~w34782;// level 8
assign po07069 = ~w34785;// level 8
assign po07070 = ~w34788;// level 8
assign po07071 = ~w34791;// level 8
assign po07072 = ~w34794;// level 8
assign po07073 = ~w34797;// level 8
assign po07074 = ~w34800;// level 8
assign po07075 = ~w34803;// level 8
assign po07076 = ~w34806;// level 8
assign po07077 = ~w34809;// level 8
assign po07078 = ~w34812;// level 8
assign po07079 = ~w34815;// level 8
assign po07080 = ~w34818;// level 8
assign po07081 = ~w34821;// level 8
assign po07082 = ~w34824;// level 8
assign po07083 = ~w34827;// level 8
assign po07084 = ~w34830;// level 8
assign po07085 = ~w34833;// level 8
assign po07086 = ~w34836;// level 8
assign po07087 = ~w34839;// level 8
assign po07088 = ~w34842;// level 8
assign po07089 = ~w34845;// level 8
assign po07090 = ~w34848;// level 8
assign po07091 = ~w34851;// level 8
assign po07092 = ~w34854;// level 8
assign po07093 = ~w34857;// level 8
assign po07094 = ~w34860;// level 8
assign po07095 = ~w34863;// level 8
assign po07096 = ~w34866;// level 8
assign po07097 = ~w34869;// level 8
assign po07098 = ~w34872;// level 8
assign po07099 = ~w34875;// level 8
assign po07100 = ~w34878;// level 8
assign po07101 = ~w34881;// level 8
assign po07102 = ~w34884;// level 8
assign po07103 = ~w34887;// level 8
assign po07104 = ~w34890;// level 8
assign po07105 = ~w34893;// level 8
assign po07106 = ~w34896;// level 8
assign po07107 = ~w34899;// level 8
assign po07108 = ~w34902;// level 8
assign po07109 = ~w34905;// level 8
assign po07110 = ~w34908;// level 8
assign po07111 = ~w34911;// level 8
assign po07112 = ~w34914;// level 8
assign po07113 = ~w34917;// level 8
assign po07114 = ~w34920;// level 8
assign po07115 = ~w34923;// level 8
assign po07116 = ~w34926;// level 8
assign po07117 = ~w34929;// level 8
assign po07118 = ~w34932;// level 8
assign po07119 = ~w34935;// level 8
assign po07120 = ~w34938;// level 8
assign po07121 = ~w34941;// level 8
assign po07122 = ~w34944;// level 8
assign po07123 = ~w34947;// level 8
assign po07124 = ~w34950;// level 8
assign po07125 = ~w34953;// level 8
assign po07126 = ~w34956;// level 8
assign po07127 = ~w34959;// level 8
assign po07128 = ~w34962;// level 8
assign po07129 = ~w34965;// level 8
assign po07130 = ~w34968;// level 8
assign po07131 = ~w34971;// level 8
assign po07132 = ~w34974;// level 8
assign po07133 = ~w34977;// level 8
assign po07134 = ~w34980;// level 8
assign po07135 = ~w34983;// level 8
assign po07136 = ~w34986;// level 8
assign po07137 = ~w34989;// level 8
assign po07138 = ~w34992;// level 8
assign po07139 = ~w34995;// level 8
assign po07140 = ~w34998;// level 8
assign po07141 = ~w35001;// level 8
assign po07142 = ~w35004;// level 8
assign po07143 = ~w35008;// level 8
assign po07144 = ~w35011;// level 8
assign po07145 = ~w35014;// level 8
assign po07146 = ~w35017;// level 8
assign po07147 = ~w35020;// level 8
assign po07148 = ~w35023;// level 8
assign po07149 = ~w35026;// level 8
assign po07150 = ~w35029;// level 8
assign po07151 = ~w35032;// level 8
assign po07152 = ~w35035;// level 8
assign po07153 = ~w35038;// level 8
assign po07154 = ~w35041;// level 8
assign po07155 = ~w35045;// level 8
assign po07156 = ~w35048;// level 8
assign po07157 = ~w35051;// level 8
assign po07158 = ~w35054;// level 8
assign po07159 = ~w35057;// level 8
assign po07160 = ~w35060;// level 8
assign po07161 = ~w35063;// level 8
assign po07162 = ~w35067;// level 8
assign po07163 = ~w35070;// level 8
assign po07164 = ~w35073;// level 8
assign po07165 = ~w35076;// level 8
assign po07166 = ~w35079;// level 8
assign po07167 = ~w35082;// level 8
assign po07168 = ~w35085;// level 8
assign po07169 = ~w35089;// level 8
assign po07170 = ~w35092;// level 8
assign po07171 = ~w35095;// level 8
assign po07172 = ~w35098;// level 8
assign po07173 = ~w35101;// level 8
assign po07174 = ~w35105;// level 8
assign po07175 = ~w35108;// level 8
assign po07176 = ~w35111;// level 8
assign po07177 = ~w35115;// level 8
assign po07178 = ~w35118;// level 8
assign po07179 = ~w35121;// level 8
assign po07180 = ~w35124;// level 8
assign po07181 = ~w35127;// level 8
assign po07182 = ~w35130;// level 8
assign po07183 = ~w35133;// level 8
assign po07184 = ~w35136;// level 8
assign po07185 = ~w35139;// level 8
assign po07186 = ~w35142;// level 8
assign po07187 = ~w35145;// level 8
assign po07188 = ~w35148;// level 8
assign po07189 = ~w35151;// level 8
assign po07190 = ~w35154;// level 8
assign po07191 = ~w35157;// level 8
assign po07192 = ~w35160;// level 8
assign po07193 = ~w35163;// level 8
assign po07194 = ~w35166;// level 8
assign po07195 = ~w35169;// level 8
assign po07196 = ~w35172;// level 8
assign po07197 = ~w35175;// level 8
assign po07198 = ~w35178;// level 8
assign po07199 = ~w35181;// level 8
assign po07200 = ~w35184;// level 8
assign po07201 = ~w35187;// level 8
assign po07202 = ~w35190;// level 8
assign po07203 = ~w35193;// level 8
assign po07204 = ~w35196;// level 8
assign po07205 = ~w35199;// level 8
assign po07206 = ~w35202;// level 8
assign po07207 = ~w35205;// level 8
assign po07208 = ~w35208;// level 8
assign po07209 = ~w35211;// level 8
assign po07210 = ~w35214;// level 8
assign po07211 = ~w35217;// level 8
assign po07212 = ~w35220;// level 8
assign po07213 = ~w35223;// level 8
assign po07214 = ~w35226;// level 8
assign po07215 = ~w35229;// level 8
assign po07216 = ~w35232;// level 8
assign po07217 = ~w35235;// level 8
assign po07218 = ~w35238;// level 8
assign po07219 = ~w35241;// level 8
assign po07220 = ~w35244;// level 8
assign po07221 = ~w35247;// level 8
assign po07222 = ~w35250;// level 8
assign po07223 = ~w35253;// level 8
assign po07224 = ~w35256;// level 8
assign po07225 = ~w35259;// level 8
assign po07226 = ~w35262;// level 8
assign po07227 = ~w35265;// level 8
assign po07228 = ~w35268;// level 8
assign po07229 = ~w35271;// level 8
assign po07230 = ~w35274;// level 8
assign po07231 = ~w35277;// level 8
assign po07232 = ~w35280;// level 8
assign po07233 = ~w35283;// level 8
assign po07234 = ~w35286;// level 8
assign po07235 = ~w35289;// level 8
assign po07236 = ~w35292;// level 8
assign po07237 = ~w35295;// level 8
assign po07238 = ~w35298;// level 8
assign po07239 = ~w35301;// level 8
assign po07240 = ~w35304;// level 8
assign po07241 = ~w35307;// level 8
assign po07242 = ~w35310;// level 8
assign po07243 = ~w35313;// level 8
assign po07244 = ~w35316;// level 8
assign po07245 = ~w35319;// level 8
assign po07246 = ~w35322;// level 8
assign po07247 = ~w35325;// level 8
assign po07248 = ~w35328;// level 8
assign po07249 = ~w35331;// level 8
assign po07250 = ~w35334;// level 8
assign po07251 = ~w35337;// level 8
assign po07252 = ~w35340;// level 8
assign po07253 = ~w35343;// level 8
assign po07254 = ~w35346;// level 8
assign po07255 = ~w35349;// level 8
assign po07256 = ~w35352;// level 8
assign po07257 = ~w35355;// level 8
assign po07258 = ~w35358;// level 8
assign po07259 = ~w35361;// level 8
assign po07260 = ~w35364;// level 8
assign po07261 = ~w35367;// level 8
assign po07262 = ~w35370;// level 8
assign po07263 = ~w35373;// level 8
assign po07264 = ~w35376;// level 8
assign po07265 = ~w35379;// level 8
assign po07266 = ~w35382;// level 8
assign po07267 = ~w35385;// level 8
assign po07268 = ~w35388;// level 8
assign po07269 = ~w35391;// level 8
assign po07270 = ~w35394;// level 8
assign po07271 = ~w35397;// level 7
assign po07272 = ~w35400;// level 7
assign po07273 = ~w35403;// level 7
assign po07274 = ~w35406;// level 8
assign po07275 = ~w35409;// level 7
assign po07276 = ~w35412;// level 7
assign po07277 = ~w35415;// level 8
assign po07278 = ~w35418;// level 7
assign po07279 = ~w35422;// level 8
assign po07280 = ~w35425;// level 8
assign po07281 = ~w35428;// level 8
assign po07282 = ~w35431;// level 8
assign po07283 = ~w35434;// level 8
assign po07284 = ~w35437;// level 8
assign po07285 = ~w35440;// level 8
assign po07286 = ~w35444;// level 8
assign po07287 = ~w35447;// level 8
assign po07288 = ~w35450;// level 8
assign po07289 = ~w35453;// level 8
assign po07290 = ~w35456;// level 8
assign po07291 = ~w35459;// level 8
assign po07292 = ~w35462;// level 8
assign po07293 = ~w35466;// level 8
assign po07294 = ~w35469;// level 8
assign po07295 = ~w35472;// level 8
assign po07296 = ~w35476;// level 8
assign po07297 = ~w35479;// level 8
assign po07298 = ~w35482;// level 8
assign po07299 = ~w35485;// level 8
assign po07300 = ~w35488;// level 8
assign po07301 = ~w35491;// level 8
assign po07302 = ~w35494;// level 8
assign po07303 = ~w35497;// level 8
assign po07304 = ~w35500;// level 8
assign po07305 = ~w35504;// level 8
assign po07306 = ~w35507;// level 8
assign po07307 = ~w35510;// level 8
assign po07308 = ~w35513;// level 8
assign po07309 = ~w35516;// level 8
assign po07310 = ~w35519;// level 8
assign po07311 = ~w35522;// level 8
assign po07312 = ~w35525;// level 8
assign po07313 = ~w35528;// level 8
assign po07314 = ~w35531;// level 8
assign po07315 = ~w35534;// level 8
assign po07316 = ~w35537;// level 8
assign po07317 = ~w35540;// level 8
assign po07318 = ~w35543;// level 8
assign po07319 = ~w35546;// level 8
assign po07320 = ~w35549;// level 8
assign po07321 = ~w35552;// level 8
assign po07322 = ~w35555;// level 8
assign po07323 = ~w35558;// level 8
assign po07324 = ~w35561;// level 8
assign po07325 = ~w35564;// level 8
assign po07326 = ~w35567;// level 8
assign po07327 = ~w35570;// level 8
assign po07328 = ~w35573;// level 8
assign po07329 = ~w35576;// level 8
assign po07330 = ~w35579;// level 8
assign po07331 = ~w35582;// level 8
assign po07332 = ~w35585;// level 8
assign po07333 = ~w35588;// level 8
assign po07334 = ~w35591;// level 8
assign po07335 = ~w35594;// level 8
assign po07336 = ~w35597;// level 8
assign po07337 = ~w35600;// level 8
assign po07338 = ~w35603;// level 8
assign po07339 = ~w35606;// level 8
assign po07340 = ~w35609;// level 8
assign po07341 = ~w35612;// level 8
assign po07342 = ~w35615;// level 8
assign po07343 = ~w35618;// level 8
assign po07344 = ~w35622;// level 8
assign po07345 = ~w35625;// level 8
assign po07346 = ~w35628;// level 8
assign po07347 = ~w35631;// level 8
assign po07348 = ~w35634;// level 8
assign po07349 = ~w35637;// level 8
assign po07350 = ~w35640;// level 8
assign po07351 = ~w35643;// level 8
assign po07352 = ~w35646;// level 8
assign po07353 = ~w35649;// level 8
assign po07354 = ~w35652;// level 8
assign po07355 = ~w35655;// level 8
assign po07356 = ~w35658;// level 8
assign po07357 = ~w35661;// level 8
assign po07358 = ~w35664;// level 8
assign po07359 = ~w35668;// level 8
assign po07360 = ~w35671;// level 8
assign po07361 = ~w35674;// level 8
assign po07362 = ~w35677;// level 8
assign po07363 = ~w35680;// level 8
assign po07364 = ~w35683;// level 8
assign po07365 = ~w35686;// level 8
assign po07366 = ~w35689;// level 8
assign po07367 = ~w35692;// level 8
assign po07368 = ~w35695;// level 8
assign po07369 = ~w35698;// level 8
assign po07370 = ~w35701;// level 8
assign po07371 = ~w35704;// level 8
assign po07372 = ~w35707;// level 8
assign po07373 = ~w35710;// level 8
assign po07374 = ~w35713;// level 8
assign po07375 = ~w35716;// level 8
assign po07376 = ~w35719;// level 8
assign po07377 = ~w35722;// level 8
assign po07378 = ~w35725;// level 8
assign po07379 = ~w35728;// level 8
assign po07380 = ~w35731;// level 8
assign po07381 = ~w35734;// level 8
assign po07382 = ~w35737;// level 8
assign po07383 = ~w35740;// level 8
assign po07384 = ~w35743;// level 8
assign po07385 = ~w35746;// level 8
assign po07386 = ~w35749;// level 8
assign po07387 = ~w35752;// level 8
assign po07388 = ~w35755;// level 8
assign po07389 = ~w35758;// level 8
assign po07390 = ~w35761;// level 8
assign po07391 = ~w35764;// level 8
assign po07392 = ~w35767;// level 8
assign po07393 = ~w35770;// level 8
assign po07394 = ~w35773;// level 8
assign po07395 = ~w35776;// level 8
assign po07396 = ~w35779;// level 8
assign po07397 = ~w35782;// level 8
assign po07398 = ~w35785;// level 8
assign po07399 = ~w35788;// level 8
assign po07400 = ~w35791;// level 8
assign po07401 = ~w35794;// level 8
assign po07402 = ~w35797;// level 8
assign po07403 = ~w35800;// level 8
assign po07404 = ~w35803;// level 8
assign po07405 = ~w35806;// level 8
assign po07406 = ~w35809;// level 8
assign po07407 = ~w35812;// level 8
assign po07408 = ~w35815;// level 8
assign po07409 = ~w35818;// level 8
assign po07410 = ~w35821;// level 8
assign po07411 = ~w35824;// level 8
assign po07412 = ~w35828;// level 8
assign po07413 = ~w35831;// level 8
assign po07414 = ~w35834;// level 8
assign po07415 = ~w35837;// level 8
assign po07416 = ~w35840;// level 8
assign po07417 = ~w35843;// level 8
assign po07418 = ~w35846;// level 8
assign po07419 = ~w35849;// level 8
assign po07420 = ~w35852;// level 8
assign po07421 = ~w35855;// level 8
assign po07422 = ~w35858;// level 8
assign po07423 = ~w35861;// level 8
assign po07424 = ~w35864;// level 8
assign po07425 = ~w35867;// level 8
assign po07426 = ~w35870;// level 8
assign po07427 = ~w35873;// level 8
assign po07428 = ~w35876;// level 8
assign po07429 = ~w35879;// level 8
assign po07430 = ~w35882;// level 8
assign po07431 = ~w35885;// level 8
assign po07432 = ~w35888;// level 8
assign po07433 = ~w35891;// level 8
assign po07434 = ~w35894;// level 8
assign po07435 = ~w35897;// level 8
assign po07436 = ~w35900;// level 8
assign po07437 = ~w35903;// level 8
assign po07438 = ~w35906;// level 8
assign po07439 = ~w35909;// level 8
assign po07440 = ~w35912;// level 8
assign po07441 = ~w35915;// level 8
assign po07442 = ~w35918;// level 8
assign po07443 = ~w35922;// level 8
assign po07444 = ~w35925;// level 8
assign po07445 = ~w35928;// level 8
assign po07446 = ~w35932;// level 8
assign po07447 = ~w35935;// level 8
assign po07448 = ~w35938;// level 8
assign po07449 = ~w35941;// level 8
assign po07450 = ~w35944;// level 8
assign po07451 = ~w35947;// level 8
assign po07452 = ~w35950;// level 8
assign po07453 = ~w35953;// level 8
assign po07454 = ~w35956;// level 8
assign po07455 = ~w35959;// level 8
assign po07456 = ~w35962;// level 8
assign po07457 = ~w35965;// level 8
assign po07458 = ~w35969;// level 8
assign po07459 = ~w35972;// level 8
assign po07460 = ~w35975;// level 8
assign po07461 = ~w35978;// level 8
assign po07462 = ~w35981;// level 8
assign po07463 = ~w35984;// level 8
assign po07464 = ~w35987;// level 8
assign po07465 = ~w35990;// level 8
assign po07466 = ~w35993;// level 8
assign po07467 = ~w35996;// level 8
assign po07468 = ~w36000;// level 8
assign po07469 = ~w36003;// level 8
assign po07470 = ~w36006;// level 8
assign po07471 = ~w36009;// level 8
assign po07472 = ~w36012;// level 8
assign po07473 = ~w36015;// level 8
assign po07474 = ~w36018;// level 8
assign po07475 = ~w36021;// level 8
assign po07476 = ~w36024;// level 8
assign po07477 = ~w36027;// level 8
assign po07478 = ~w36030;// level 8
assign po07479 = ~w36033;// level 8
assign po07480 = ~w36036;// level 8
assign po07481 = ~w36039;// level 8
assign po07482 = ~w36042;// level 8
assign po07483 = ~w36045;// level 8
assign po07484 = ~w36048;// level 8
assign po07485 = ~w36051;// level 8
assign po07486 = ~w36054;// level 8
assign po07487 = ~w36057;// level 8
assign po07488 = ~w36060;// level 8
assign po07489 = ~w36063;// level 8
assign po07490 = ~w36066;// level 8
assign po07491 = ~w36069;// level 8
assign po07492 = ~w36072;// level 8
assign po07493 = ~w36075;// level 8
assign po07494 = ~w36078;// level 8
assign po07495 = ~w36081;// level 8
assign po07496 = ~w36084;// level 8
assign po07497 = ~w36087;// level 8
assign po07498 = ~w36091;// level 8
assign po07499 = ~w36094;// level 8
assign po07500 = ~w36097;// level 8
assign po07501 = ~w36100;// level 8
assign po07502 = ~w36103;// level 8
assign po07503 = ~w36106;// level 8
assign po07504 = ~w36109;// level 8
assign po07505 = ~w36112;// level 8
assign po07506 = ~w36115;// level 8
assign po07507 = ~w36118;// level 8
assign po07508 = ~w36121;// level 8
assign po07509 = ~w36124;// level 8
assign po07510 = ~w36127;// level 8
assign po07511 = ~w36130;// level 8
assign po07512 = ~w36133;// level 8
assign po07513 = ~w36136;// level 8
assign po07514 = ~w36139;// level 8
assign po07515 = ~w36142;// level 8
assign po07516 = ~w36145;// level 8
assign po07517 = ~w36148;// level 8
assign po07518 = ~w36151;// level 8
assign po07519 = ~w36154;// level 8
assign po07520 = ~w36157;// level 8
assign po07521 = ~w36160;// level 8
assign po07522 = ~w36163;// level 8
assign po07523 = ~w36166;// level 8
assign po07524 = ~w36169;// level 8
assign po07525 = ~w36172;// level 8
assign po07526 = ~w36175;// level 8
assign po07527 = ~w36178;// level 8
assign po07528 = ~w36181;// level 8
assign po07529 = ~w36184;// level 8
assign po07530 = ~w36187;// level 8
assign po07531 = ~w36190;// level 8
assign po07532 = ~w36193;// level 8
assign po07533 = ~w36196;// level 8
assign po07534 = ~w36199;// level 8
assign po07535 = ~w36202;// level 8
assign po07536 = ~w36205;// level 8
assign po07537 = ~w36209;// level 8
assign po07538 = ~w36212;// level 8
assign po07539 = ~w36215;// level 8
assign po07540 = ~w36218;// level 8
assign po07541 = ~w36221;// level 8
assign po07542 = ~w36224;// level 8
assign po07543 = ~w36227;// level 8
assign po07544 = ~w36230;// level 8
assign po07545 = ~w36233;// level 8
assign po07546 = ~w36236;// level 8
assign po07547 = ~w36239;// level 8
assign po07548 = ~w36242;// level 8
assign po07549 = ~w36245;// level 8
assign po07550 = ~w36248;// level 8
assign po07551 = ~w36251;// level 8
assign po07552 = ~w36254;// level 8
assign po07553 = ~w36257;// level 8
assign po07554 = ~w36260;// level 8
assign po07555 = ~w36263;// level 8
assign po07556 = ~w36266;// level 8
assign po07557 = ~w36269;// level 8
assign po07558 = ~w36272;// level 8
assign po07559 = ~w36275;// level 8
assign po07560 = ~w36278;// level 8
assign po07561 = ~w36281;// level 8
assign po07562 = ~w36284;// level 8
assign po07563 = ~w36287;// level 8
assign po07564 = ~w36290;// level 8
assign po07565 = ~w36293;// level 8
assign po07566 = ~w36296;// level 8
assign po07567 = ~w36299;// level 8
assign po07568 = ~w36302;// level 8
assign po07569 = ~w36305;// level 8
assign po07570 = ~w36308;// level 8
assign po07571 = ~w36311;// level 8
assign po07572 = ~w36314;// level 8
assign po07573 = ~w36317;// level 8
assign po07574 = ~w36320;// level 8
assign po07575 = ~w36323;// level 8
assign po07576 = ~w36326;// level 8
assign po07577 = ~w36329;// level 8
assign po07578 = ~w36332;// level 8
assign po07579 = ~w36335;// level 8
assign po07580 = ~w36338;// level 8
assign po07581 = ~w36341;// level 8
assign po07582 = ~w36344;// level 8
assign po07583 = ~w36347;// level 8
assign po07584 = ~w36350;// level 8
assign po07585 = ~w36353;// level 8
assign po07586 = ~w36356;// level 8
assign po07587 = ~w36360;// level 8
assign po07588 = ~w36363;// level 8
assign po07589 = ~w36366;// level 8
assign po07590 = ~w36369;// level 8
assign po07591 = ~w36372;// level 8
assign po07592 = ~w36375;// level 8
assign po07593 = ~w36378;// level 8
assign po07594 = ~w36381;// level 8
assign po07595 = ~w36384;// level 8
assign po07596 = ~w36387;// level 8
assign po07597 = ~w36390;// level 8
assign po07598 = ~w36394;// level 8
assign po07599 = ~w36397;// level 8
assign po07600 = ~w36400;// level 8
assign po07601 = ~w36403;// level 8
assign po07602 = ~w36406;// level 8
assign po07603 = ~w36409;// level 8
assign po07604 = ~w36412;// level 8
assign po07605 = ~w36415;// level 8
assign po07606 = ~w36419;// level 8
assign po07607 = ~w36422;// level 8
assign po07608 = ~w36425;// level 8
assign po07609 = ~w36428;// level 8
assign po07610 = ~w36431;// level 8
assign po07611 = ~w36434;// level 8
assign po07612 = ~w36437;// level 8
assign po07613 = ~w36440;// level 8
assign po07614 = ~w36443;// level 8
assign po07615 = ~w36446;// level 8
assign po07616 = ~w36449;// level 8
assign po07617 = ~w36453;// level 8
assign po07618 = ~w36456;// level 8
assign po07619 = ~w36459;// level 8
assign po07620 = ~w36462;// level 8
assign po07621 = ~w36465;// level 8
assign po07622 = ~w36468;// level 8
assign po07623 = ~w36471;// level 8
assign po07624 = ~w36475;// level 8
assign po07625 = ~w36478;// level 8
assign po07626 = ~w36481;// level 8
assign po07627 = ~w36484;// level 8
assign po07628 = ~w36487;// level 8
assign po07629 = ~w36490;// level 8
assign po07630 = ~w36493;// level 8
assign po07631 = ~w36496;// level 8
assign po07632 = ~w36499;// level 8
assign po07633 = ~w36502;// level 8
assign po07634 = ~w36505;// level 8
assign po07635 = ~w36508;// level 8
assign po07636 = ~w36511;// level 8
assign po07637 = ~w36514;// level 8
assign po07638 = ~w36517;// level 8
assign po07639 = ~w36520;// level 8
assign po07640 = ~w36523;// level 8
assign po07641 = ~w36526;// level 8
assign po07642 = ~w36529;// level 8
assign po07643 = ~w36532;// level 8
assign po07644 = ~w36535;// level 8
assign po07645 = ~w36538;// level 8
assign po07646 = ~w36541;// level 8
assign po07647 = ~w36544;// level 8
assign po07648 = ~w36547;// level 8
assign po07649 = ~w36550;// level 8
assign po07650 = ~w36553;// level 8
assign po07651 = ~w36556;// level 8
assign po07652 = ~w36559;// level 8
assign po07653 = ~w36562;// level 8
assign po07654 = ~w36565;// level 8
assign po07655 = ~w36568;// level 8
assign po07656 = ~w36571;// level 8
assign po07657 = ~w36574;// level 8
assign po07658 = ~w36577;// level 8
assign po07659 = ~w36580;// level 8
assign po07660 = ~w36583;// level 8
assign po07661 = ~w36586;// level 8
assign po07662 = ~w36589;// level 8
assign po07663 = ~w36592;// level 8
assign po07664 = ~w36595;// level 8
assign po07665 = ~w36598;// level 8
assign po07666 = ~w36601;// level 8
assign po07667 = ~w36604;// level 8
assign po07668 = ~w36607;// level 8
assign po07669 = ~w36610;// level 8
assign po07670 = ~w36613;// level 8
assign po07671 = ~w36616;// level 8
assign po07672 = ~w36619;// level 8
assign po07673 = ~w36622;// level 8
assign po07674 = ~w36625;// level 8
assign po07675 = ~w36628;// level 8
assign po07676 = ~w36631;// level 8
assign po07677 = ~w36634;// level 8
assign po07678 = ~w36637;// level 8
assign po07679 = ~w36640;// level 8
assign po07680 = ~w36643;// level 8
assign po07681 = ~w36646;// level 8
assign po07682 = ~w36649;// level 8
assign po07683 = ~w36652;// level 8
assign po07684 = ~w36655;// level 8
assign po07685 = ~w36658;// level 8
assign po07686 = ~w36661;// level 8
assign po07687 = ~w36664;// level 8
assign po07688 = ~w36667;// level 8
assign po07689 = ~w36670;// level 8
assign po07690 = ~w36673;// level 8
assign po07691 = ~w36676;// level 8
assign po07692 = ~w36679;// level 8
assign po07693 = ~w36682;// level 8
assign po07694 = ~w36685;// level 8
assign po07695 = ~w36689;// level 8
assign po07696 = ~w36692;// level 8
assign po07697 = ~w36695;// level 8
assign po07698 = ~w36698;// level 8
assign po07699 = ~w36701;// level 8
assign po07700 = ~w36704;// level 8
assign po07701 = ~w36707;// level 8
assign po07702 = ~w36710;// level 8
assign po07703 = ~w36713;// level 8
assign po07704 = ~w36716;// level 8
assign po07705 = ~w36719;// level 8
assign po07706 = ~w36722;// level 8
assign po07707 = ~w36725;// level 8
assign po07708 = ~w36728;// level 8
assign po07709 = ~w36731;// level 8
assign po07710 = ~w36734;// level 8
assign po07711 = ~w36737;// level 8
assign po07712 = ~w36740;// level 8
assign po07713 = ~w36743;// level 8
assign po07714 = ~w36746;// level 8
assign po07715 = ~w36749;// level 8
assign po07716 = ~w36752;// level 8
assign po07717 = ~w36755;// level 8
assign po07718 = ~w36758;// level 8
assign po07719 = ~w36761;// level 8
assign po07720 = ~w36764;// level 8
assign po07721 = ~w36767;// level 8
assign po07722 = ~w36770;// level 8
assign po07723 = ~w36773;// level 8
assign po07724 = ~w36776;// level 8
assign po07725 = ~w36779;// level 8
assign po07726 = ~w36782;// level 8
assign po07727 = ~w36785;// level 8
assign po07728 = ~w36788;// level 8
assign po07729 = ~w36791;// level 8
assign po07730 = ~w36794;// level 8
assign po07731 = ~w36797;// level 8
assign po07732 = ~w36800;// level 8
assign po07733 = ~w36803;// level 8
assign po07734 = ~w36806;// level 8
assign po07735 = ~w36809;// level 8
assign po07736 = ~w36812;// level 8
assign po07737 = ~w36815;// level 8
assign po07738 = ~w36818;// level 8
assign po07739 = ~w36821;// level 8
assign po07740 = ~w36824;// level 8
assign po07741 = ~w36827;// level 8
assign po07742 = ~w36830;// level 8
assign po07743 = ~w36833;// level 8
assign po07744 = ~w36836;// level 8
assign po07745 = ~w36839;// level 8
assign po07746 = ~w36842;// level 8
assign po07747 = ~w36845;// level 8
assign po07748 = ~w36848;// level 8
assign po07749 = ~w36851;// level 7
assign po07750 = ~w36854;// level 7
assign po07751 = ~w36857;// level 7
assign po07752 = ~w36860;// level 7
assign po07753 = ~w36863;// level 7
assign po07754 = ~w36866;// level 7
assign po07755 = ~w36869;// level 7
assign po07756 = ~w36872;// level 8
assign po07757 = ~w36875;// level 8
assign po07758 = ~w36878;// level 8
assign po07759 = ~w36881;// level 8
assign po07760 = ~w36884;// level 8
assign po07761 = ~w36887;// level 8
assign po07762 = ~w36891;// level 8
assign po07763 = ~w36895;// level 8
assign po07764 = ~w36898;// level 8
assign po07765 = ~w36901;// level 8
assign po07766 = ~w36904;// level 8
assign po07767 = ~w36907;// level 8
assign po07768 = ~w36910;// level 8
assign po07769 = ~w36913;// level 8
assign po07770 = ~w36916;// level 8
assign po07771 = ~w36919;// level 8
assign po07772 = ~w36923;// level 8
assign po07773 = ~w36926;// level 8
assign po07774 = ~w36929;// level 8
assign po07775 = ~w36932;// level 8
assign po07776 = ~w36935;// level 8
assign po07777 = ~w36938;// level 8
assign po07778 = ~w36941;// level 8
assign po07779 = ~w36944;// level 8
assign po07780 = ~w36947;// level 8
assign po07781 = ~w36950;// level 8
assign po07782 = ~w36953;// level 8
assign po07783 = ~w36957;// level 8
assign po07784 = ~w36960;// level 8
assign po07785 = ~w36963;// level 8
assign po07786 = ~w36966;// level 8
assign po07787 = ~w36969;// level 8
assign po07788 = ~w36972;// level 8
assign po07789 = ~w36975;// level 8
assign po07790 = ~w36978;// level 8
assign po07791 = ~w36981;// level 8
assign po07792 = ~w36984;// level 8
assign po07793 = ~w36987;// level 8
assign po07794 = ~w36990;// level 8
assign po07795 = ~w36993;// level 8
assign po07796 = ~w36996;// level 8
assign po07797 = ~w36999;// level 8
assign po07798 = ~w37002;// level 8
assign po07799 = ~w37005;// level 8
assign po07800 = ~w37008;// level 8
assign po07801 = ~w37011;// level 8
assign po07802 = ~w37014;// level 8
assign po07803 = ~w37017;// level 8
assign po07804 = ~w37020;// level 8
assign po07805 = ~w37023;// level 8
assign po07806 = ~w37026;// level 8
assign po07807 = ~w37029;// level 8
assign po07808 = ~w37032;// level 8
assign po07809 = ~w37035;// level 8
assign po07810 = ~w37038;// level 8
assign po07811 = ~w37041;// level 8
assign po07812 = ~w37044;// level 8
assign po07813 = ~w37047;// level 8
assign po07814 = ~w37050;// level 8
assign po07815 = ~w37053;// level 8
assign po07816 = ~w37056;// level 8
assign po07817 = ~w37059;// level 8
assign po07818 = ~w37062;// level 8
assign po07819 = ~w37065;// level 8
assign po07820 = ~w37068;// level 8
assign po07821 = ~w37071;// level 8
assign po07822 = ~w37074;// level 8
assign po07823 = ~w37077;// level 8
assign po07824 = ~w37080;// level 8
assign po07825 = ~w37083;// level 8
assign po07826 = ~w37086;// level 8
assign po07827 = ~w37089;// level 8
assign po07828 = ~w37092;// level 8
assign po07829 = ~w37095;// level 8
assign po07830 = ~w37098;// level 8
assign po07831 = ~w37101;// level 8
assign po07832 = ~w37104;// level 8
assign po07833 = ~w37107;// level 8
assign po07834 = ~w37110;// level 8
assign po07835 = ~w37113;// level 8
assign po07836 = ~w37116;// level 8
assign po07837 = ~w37119;// level 8
assign po07838 = ~w37122;// level 8
assign po07839 = ~w37125;// level 8
assign po07840 = ~w37128;// level 8
assign po07841 = ~w37131;// level 8
assign po07842 = ~w37134;// level 8
assign po07843 = ~w37137;// level 8
assign po07844 = ~w37140;// level 8
assign po07845 = ~w37143;// level 8
assign po07846 = ~w37146;// level 8
assign po07847 = ~w37149;// level 8
assign po07848 = ~w37152;// level 8
assign po07849 = ~w37155;// level 8
assign po07850 = ~w37158;// level 8
assign po07851 = ~w37161;// level 8
assign po07852 = ~w37164;// level 8
assign po07853 = ~w37167;// level 8
assign po07854 = ~w37170;// level 8
assign po07855 = ~w37173;// level 8
assign po07856 = ~w37176;// level 8
assign po07857 = ~w37179;// level 8
assign po07858 = ~w37182;// level 8
assign po07859 = ~w37185;// level 8
assign po07860 = ~w37188;// level 8
assign po07861 = ~w37191;// level 8
assign po07862 = ~w37194;// level 8
assign po07863 = ~w37197;// level 8
assign po07864 = ~w37200;// level 8
assign po07865 = ~w37203;// level 8
assign po07866 = ~w37206;// level 8
assign po07867 = ~w37209;// level 8
assign po07868 = ~w37212;// level 8
assign po07869 = ~w37215;// level 8
assign po07870 = ~w37218;// level 8
assign po07871 = ~w37221;// level 8
assign po07872 = ~w37224;// level 8
assign po07873 = ~w37227;// level 8
assign po07874 = ~w37230;// level 8
assign po07875 = ~w37233;// level 8
assign po07876 = ~w37236;// level 8
assign po07877 = ~w37239;// level 8
assign po07878 = ~w37242;// level 8
assign po07879 = ~w37245;// level 8
assign po07880 = ~w37248;// level 8
assign po07881 = ~w37251;// level 8
assign po07882 = ~w37254;// level 8
assign po07883 = ~w37257;// level 8
assign po07884 = ~w37260;// level 8
assign po07885 = ~w37263;// level 8
assign po07886 = ~w37266;// level 8
assign po07887 = ~w37269;// level 8
assign po07888 = ~w37272;// level 8
assign po07889 = ~w37275;// level 8
assign po07890 = ~w37278;// level 8
assign po07891 = ~w37281;// level 8
assign po07892 = ~w37284;// level 8
assign po07893 = ~w37287;// level 8
assign po07894 = ~w37290;// level 8
assign po07895 = ~w37293;// level 8
assign po07896 = ~w37296;// level 8
assign po07897 = ~w37299;// level 8
assign po07898 = ~w37302;// level 8
assign po07899 = ~w37305;// level 8
assign po07900 = ~w37308;// level 8
assign po07901 = ~w37311;// level 8
assign po07902 = ~w37314;// level 8
assign po07903 = ~w37317;// level 8
assign po07904 = ~w37320;// level 8
assign po07905 = ~w37323;// level 8
assign po07906 = ~w37326;// level 8
assign po07907 = ~w37329;// level 8
assign po07908 = ~w37332;// level 8
assign po07909 = ~w37335;// level 8
assign po07910 = ~w37338;// level 8
assign po07911 = ~w37341;// level 8
assign po07912 = ~w37344;// level 8
assign po07913 = ~w37347;// level 8
assign po07914 = ~w37350;// level 8
assign po07915 = ~w37353;// level 8
assign po07916 = ~w37356;// level 8
assign po07917 = ~w37359;// level 8
assign po07918 = ~w37362;// level 8
assign po07919 = ~w37365;// level 8
assign po07920 = ~w37368;// level 8
assign po07921 = ~w37371;// level 8
assign po07922 = ~w37374;// level 8
assign po07923 = ~w37377;// level 7
assign po07924 = ~w37380;// level 8
assign po07925 = ~w37383;// level 8
assign po07926 = ~w37386;// level 7
assign po07927 = ~w37389;// level 8
assign po07928 = ~w37392;// level 7
assign po07929 = ~w37395;// level 7
assign po07930 = ~w37398;// level 8
assign po07931 = ~w37401;// level 7
assign po07932 = ~w37405;// level 8
assign po07933 = ~w37408;// level 8
assign po07934 = ~w37411;// level 8
assign po07935 = ~w37414;// level 8
assign po07936 = ~w37417;// level 8
assign po07937 = ~w37420;// level 8
assign po07938 = ~w37424;// level 8
assign po07939 = ~w37427;// level 8
assign po07940 = ~w37430;// level 8
assign po07941 = ~w37433;// level 8
assign po07942 = ~w37436;// level 8
assign po07943 = ~w37439;// level 8
assign po07944 = ~w37442;// level 8
assign po07945 = ~w37445;// level 8
assign po07946 = ~w37448;// level 8
assign po07947 = ~w37451;// level 8
assign po07948 = ~w37454;// level 8
assign po07949 = ~w37457;// level 8
assign po07950 = ~w37460;// level 8
assign po07951 = ~w37463;// level 8
assign po07952 = ~w37466;// level 8
assign po07953 = ~w37469;// level 8
assign po07954 = ~w37472;// level 8
assign po07955 = ~w37475;// level 8
assign po07956 = ~w37478;// level 8
assign po07957 = ~w37481;// level 8
assign po07958 = ~w37484;// level 8
assign po07959 = ~w37487;// level 8
assign po07960 = ~w37490;// level 8
assign po07961 = ~w37493;// level 8
assign po07962 = ~w37496;// level 8
assign po07963 = ~w37499;// level 8
assign po07964 = ~w37502;// level 8
assign po07965 = ~w37505;// level 8
assign po07966 = ~w37508;// level 8
assign po07967 = ~w37511;// level 8
assign po07968 = ~w37514;// level 8
assign po07969 = ~w37517;// level 8
assign po07970 = ~w37520;// level 8
assign po07971 = ~w37523;// level 8
assign po07972 = ~w37526;// level 7
assign po07973 = ~w37529;// level 8
assign po07974 = ~w37532;// level 7
assign po07975 = ~w37535;// level 7
assign po07976 = ~w37538;// level 8
assign po07977 = ~w37541;// level 8
assign po07978 = ~w37545;// level 8
assign po07979 = ~w37548;// level 7
assign po07980 = ~w37551;// level 8
assign po07981 = ~w37554;// level 7
assign po07982 = ~w37557;// level 8
assign po07983 = ~w37560;// level 8
assign po07984 = ~w37563;// level 8
assign po07985 = ~w37566;// level 8
assign po07986 = ~w37569;// level 8
assign po07987 = ~w37572;// level 8
assign po07988 = ~w37575;// level 8
assign po07989 = ~w37578;// level 8
assign po07990 = ~w37581;// level 8
assign po07991 = ~w37584;// level 8
assign po07992 = ~w37587;// level 8
assign po07993 = ~w37590;// level 8
assign po07994 = ~w37593;// level 8
assign po07995 = ~w37596;// level 8
assign po07996 = ~w37599;// level 8
assign po07997 = ~w37602;// level 8
assign po07998 = ~w37605;// level 8
assign po07999 = ~w37608;// level 8
assign po08000 = ~w37611;// level 8
assign po08001 = ~w37614;// level 8
assign po08002 = ~w37617;// level 8
assign po08003 = ~w37620;// level 8
assign po08004 = ~w37623;// level 8
assign po08005 = ~w37626;// level 8
assign po08006 = ~w37629;// level 8
assign po08007 = ~w37632;// level 8
assign po08008 = ~w37635;// level 8
assign po08009 = ~w37638;// level 8
assign po08010 = ~w37641;// level 8
assign po08011 = ~w37644;// level 8
assign po08012 = ~w37647;// level 8
assign po08013 = ~w37650;// level 8
assign po08014 = ~w37653;// level 8
assign po08015 = ~w37656;// level 8
assign po08016 = ~w37659;// level 8
assign po08017 = ~w37663;// level 8
assign po08018 = ~w37666;// level 8
assign po08019 = ~w37669;// level 8
assign po08020 = ~w37672;// level 8
assign po08021 = ~w37675;// level 8
assign po08022 = ~w37678;// level 8
assign po08023 = ~w37681;// level 8
assign po08024 = ~w37684;// level 8
assign po08025 = ~w37687;// level 8
assign po08026 = ~w37690;// level 8
assign po08027 = ~w37693;// level 8
assign po08028 = ~w37696;// level 8
assign po08029 = ~w37699;// level 8
assign po08030 = ~w37702;// level 8
assign po08031 = ~w37705;// level 8
assign po08032 = ~w37708;// level 8
assign po08033 = ~w37711;// level 8
assign po08034 = ~w37714;// level 8
assign po08035 = ~w37717;// level 8
assign po08036 = ~w37720;// level 8
assign po08037 = ~w37723;// level 8
assign po08038 = ~w37726;// level 8
assign po08039 = ~w37729;// level 8
assign po08040 = ~w37732;// level 8
assign po08041 = ~w37735;// level 8
assign po08042 = ~w37738;// level 8
assign po08043 = ~w37741;// level 8
assign po08044 = ~w37744;// level 8
assign po08045 = ~w37747;// level 8
assign po08046 = ~w37750;// level 8
assign po08047 = ~w37753;// level 8
assign po08048 = ~w37756;// level 8
assign po08049 = ~w37759;// level 8
assign po08050 = ~w37762;// level 8
assign po08051 = ~w37765;// level 8
assign po08052 = ~w37768;// level 8
assign po08053 = ~w37771;// level 8
assign po08054 = ~w37774;// level 8
assign po08055 = ~w37777;// level 8
assign po08056 = ~w37780;// level 8
assign po08057 = ~w37783;// level 8
assign po08058 = ~w37787;// level 8
assign po08059 = ~w37790;// level 8
assign po08060 = ~w37793;// level 8
assign po08061 = ~w37796;// level 8
assign po08062 = ~w37799;// level 8
assign po08063 = ~w37802;// level 8
assign po08064 = ~w37805;// level 8
assign po08065 = ~w37808;// level 8
assign po08066 = ~w37811;// level 8
assign po08067 = ~w37814;// level 8
assign po08068 = ~w37817;// level 8
assign po08069 = ~w37820;// level 8
assign po08070 = ~w37823;// level 8
assign po08071 = ~w37826;// level 8
assign po08072 = ~w37829;// level 8
assign po08073 = ~w37832;// level 8
assign po08074 = ~w37835;// level 8
assign po08075 = ~w37838;// level 8
assign po08076 = ~w37841;// level 8
assign po08077 = ~w37844;// level 8
assign po08078 = ~w37847;// level 8
assign po08079 = ~w37850;// level 8
assign po08080 = ~w37853;// level 8
assign po08081 = ~w37856;// level 8
assign po08082 = ~w37859;// level 8
assign po08083 = ~w37862;// level 8
assign po08084 = ~w37865;// level 8
assign po08085 = ~w37868;// level 8
assign po08086 = ~w37871;// level 8
assign po08087 = ~w37874;// level 8
assign po08088 = ~w37877;// level 8
assign po08089 = ~w37880;// level 8
assign po08090 = ~w37883;// level 8
assign po08091 = ~w37886;// level 8
assign po08092 = ~w37889;// level 8
assign po08093 = ~w37892;// level 8
assign po08094 = ~w37895;// level 8
assign po08095 = ~w37898;// level 8
assign po08096 = ~w37901;// level 8
assign po08097 = ~w37905;// level 8
assign po08098 = ~w37908;// level 8
assign po08099 = ~w37911;// level 8
assign po08100 = ~w37914;// level 8
assign po08101 = ~w37917;// level 8
assign po08102 = ~w37920;// level 8
assign po08103 = ~w37923;// level 8
assign po08104 = ~w37926;// level 8
assign po08105 = ~w37929;// level 8
assign po08106 = ~w37932;// level 8
assign po08107 = ~w37935;// level 8
assign po08108 = ~w37938;// level 8
assign po08109 = ~w37941;// level 8
assign po08110 = ~w37944;// level 8
assign po08111 = ~w37947;// level 8
assign po08112 = ~w37950;// level 8
assign po08113 = ~w37953;// level 8
assign po08114 = ~w37956;// level 8
assign po08115 = ~w37959;// level 8
assign po08116 = ~w37962;// level 8
assign po08117 = ~w37965;// level 8
assign po08118 = ~w37968;// level 8
assign po08119 = ~w37971;// level 8
assign po08120 = ~w37974;// level 8
assign po08121 = ~w37977;// level 8
assign po08122 = ~w37980;// level 8
assign po08123 = ~w37983;// level 8
assign po08124 = ~w37986;// level 8
assign po08125 = ~w37989;// level 8
assign po08126 = ~w37992;// level 8
assign po08127 = ~w37995;// level 8
assign po08128 = ~w37998;// level 8
assign po08129 = ~w38001;// level 8
assign po08130 = ~w38004;// level 8
assign po08131 = ~w38007;// level 8
assign po08132 = ~w38010;// level 8
assign po08133 = ~w38013;// level 8
assign po08134 = ~w38016;// level 8
assign po08135 = ~w38019;// level 8
assign po08136 = ~w38022;// level 8
assign po08137 = ~w38025;// level 8
assign po08138 = ~w38028;// level 8
assign po08139 = ~w38031;// level 8
assign po08140 = ~w38034;// level 8
assign po08141 = ~w38037;// level 8
assign po08142 = ~w38040;// level 8
assign po08143 = ~w38043;// level 8
assign po08144 = ~w38046;// level 8
assign po08145 = ~w38049;// level 8
assign po08146 = ~w38052;// level 8
assign po08147 = ~w38055;// level 8
assign po08148 = ~w38058;// level 8
assign po08149 = ~w38061;// level 8
assign po08150 = ~w38064;// level 8
assign po08151 = ~w38067;// level 8
assign po08152 = ~w38070;// level 8
assign po08153 = ~w38073;// level 8
assign po08154 = ~w38076;// level 8
assign po08155 = ~w38079;// level 8
assign po08156 = ~w38082;// level 8
assign po08157 = ~w38085;// level 8
assign po08158 = ~w38088;// level 8
assign po08159 = ~w38091;// level 8
assign po08160 = ~w38094;// level 8
assign po08161 = ~w38097;// level 8
assign po08162 = ~w38100;// level 8
assign po08163 = ~w38103;// level 8
assign po08164 = ~w38106;// level 8
assign po08165 = ~w38109;// level 8
assign po08166 = ~w38112;// level 8
assign po08167 = ~w38115;// level 8
assign po08168 = ~w38118;// level 8
assign po08169 = ~w38121;// level 8
assign po08170 = ~w38124;// level 8
assign po08171 = ~w38127;// level 8
assign po08172 = ~w38130;// level 8
assign po08173 = ~w38133;// level 8
assign po08174 = ~w38136;// level 8
assign po08175 = ~w38139;// level 8
assign po08176 = ~w38142;// level 8
assign po08177 = ~w38145;// level 8
assign po08178 = ~w38148;// level 8
assign po08179 = ~w38151;// level 8
assign po08180 = ~w38154;// level 8
assign po08181 = ~w38157;// level 8
assign po08182 = ~w38160;// level 8
assign po08183 = ~w38163;// level 8
assign po08184 = ~w38166;// level 8
assign po08185 = ~w38169;// level 8
assign po08186 = ~w38172;// level 8
assign po08187 = ~w38175;// level 8
assign po08188 = ~w38178;// level 8
assign po08189 = ~w38181;// level 8
assign po08190 = ~w38184;// level 8
assign po08191 = ~w38187;// level 8
assign po08192 = ~w38190;// level 8
assign po08193 = ~w38193;// level 8
assign po08194 = ~w38196;// level 8
assign po08195 = ~w38199;// level 8
assign po08196 = ~w38202;// level 8
assign po08197 = ~w38205;// level 8
assign po08198 = ~w38208;// level 8
assign po08199 = ~w38211;// level 8
assign po08200 = ~w38214;// level 8
assign po08201 = ~w38217;// level 8
assign po08202 = ~w38220;// level 8
assign po08203 = ~w38223;// level 8
assign po08204 = ~w38226;// level 8
assign po08205 = ~w38229;// level 8
assign po08206 = ~w38232;// level 8
assign po08207 = ~w38235;// level 8
assign po08208 = ~w38238;// level 8
assign po08209 = ~w38241;// level 8
assign po08210 = ~w38244;// level 8
assign po08211 = ~w38247;// level 8
assign po08212 = ~w38250;// level 8
assign po08213 = ~w38253;// level 8
assign po08214 = ~w38256;// level 8
assign po08215 = ~w38259;// level 8
assign po08216 = ~w38262;// level 8
assign po08217 = ~w38265;// level 8
assign po08218 = ~w38268;// level 8
assign po08219 = ~w38271;// level 8
assign po08220 = ~w38274;// level 8
assign po08221 = ~w38277;// level 8
assign po08222 = ~w38280;// level 8
assign po08223 = ~w38283;// level 8
assign po08224 = ~w38286;// level 8
assign po08225 = ~w38289;// level 8
assign po08226 = ~w38292;// level 8
assign po08227 = ~w38295;// level 8
assign po08228 = ~w38298;// level 8
assign po08229 = ~w38301;// level 8
assign po08230 = ~w38304;// level 8
assign po08231 = ~w38307;// level 8
assign po08232 = ~w38310;// level 8
assign po08233 = ~w38314;// level 8
assign po08234 = ~w38317;// level 8
assign po08235 = ~w38320;// level 8
assign po08236 = ~w38323;// level 8
assign po08237 = ~w38326;// level 8
assign po08238 = ~w38329;// level 8
assign po08239 = ~w38332;// level 8
assign po08240 = ~w38335;// level 8
assign po08241 = ~w38338;// level 8
assign po08242 = ~w38341;// level 8
assign po08243 = ~w38344;// level 8
assign po08244 = ~w38347;// level 8
assign po08245 = ~w38350;// level 8
assign po08246 = ~w38353;// level 8
assign po08247 = ~w38356;// level 8
assign po08248 = ~w38359;// level 8
assign po08249 = ~w38362;// level 7
assign po08250 = ~w38365;// level 8
assign po08251 = ~w38368;// level 7
assign po08252 = ~w38371;// level 8
assign po08253 = ~w38374;// level 7
assign po08254 = ~w38377;// level 8
assign po08255 = ~w38380;// level 7
assign po08256 = ~w38383;// level 8
assign po08257 = ~w38386;// level 8
assign po08258 = ~w38389;// level 8
assign po08259 = ~w38392;// level 7
assign po08260 = ~w38395;// level 7
assign po08261 = ~w38398;// level 8
assign po08262 = ~w38401;// level 8
assign po08263 = ~w38404;// level 7
assign po08264 = ~w38407;// level 7
assign po08265 = ~w38410;// level 7
assign po08266 = ~w38413;// level 7
assign po08267 = ~w38416;// level 7
assign po08268 = ~w38419;// level 7
assign po08269 = ~w38423;// level 8
assign po08270 = ~w38426;// level 8
assign po08271 = ~w38429;// level 8
assign po08272 = ~w38432;// level 8
assign po08273 = ~w38435;// level 8
assign po08274 = ~w38438;// level 8
assign po08275 = ~w38441;// level 8
assign po08276 = ~w38444;// level 8
assign po08277 = ~w38447;// level 8
assign po08278 = ~w38451;// level 8
assign po08279 = ~w38454;// level 8
assign po08280 = ~w38457;// level 8
assign po08281 = ~w38460;// level 8
assign po08282 = ~w38463;// level 8
assign po08283 = ~w38466;// level 8
assign po08284 = ~w38470;// level 8
assign po08285 = ~w38473;// level 8
assign po08286 = ~w38476;// level 8
assign po08287 = ~w38479;// level 8
assign po08288 = ~w38482;// level 8
assign po08289 = ~w38485;// level 8
assign po08290 = ~w38488;// level 8
assign po08291 = ~w38491;// level 8
assign po08292 = ~w38494;// level 8
assign po08293 = ~w38497;// level 8
assign po08294 = ~w38500;// level 8
assign po08295 = ~w38503;// level 8
assign po08296 = ~w38506;// level 8
assign po08297 = ~w38509;// level 8
assign po08298 = ~w38512;// level 8
assign po08299 = ~w38515;// level 8
assign po08300 = ~w38518;// level 8
assign po08301 = ~w38521;// level 8
assign po08302 = ~w38524;// level 8
assign po08303 = ~w38527;// level 8
assign po08304 = ~w38530;// level 8
assign po08305 = ~w38533;// level 8
assign po08306 = ~w38536;// level 8
assign po08307 = ~w38539;// level 8
assign po08308 = ~w38542;// level 8
assign po08309 = ~w38545;// level 8
assign po08310 = ~w38548;// level 8
assign po08311 = ~w38551;// level 8
assign po08312 = ~w38554;// level 8
assign po08313 = ~w38557;// level 8
assign po08314 = ~w38560;// level 8
assign po08315 = ~w38563;// level 8
assign po08316 = ~w38566;// level 8
assign po08317 = ~w38569;// level 8
assign po08318 = ~w38572;// level 8
assign po08319 = ~w38575;// level 8
assign po08320 = ~w38578;// level 8
assign po08321 = ~w38581;// level 8
assign po08322 = ~w38584;// level 8
assign po08323 = ~w38587;// level 8
assign po08324 = ~w38590;// level 8
assign po08325 = ~w38593;// level 8
assign po08326 = ~w38596;// level 8
assign po08327 = ~w38599;// level 8
assign po08328 = ~w38602;// level 8
assign po08329 = ~w38605;// level 8
assign po08330 = ~w38608;// level 8
assign po08331 = ~w38611;// level 8
assign po08332 = ~w38614;// level 8
assign po08333 = ~w38617;// level 8
assign po08334 = ~w38620;// level 8
assign po08335 = ~w38623;// level 8
assign po08336 = ~w38626;// level 8
assign po08337 = ~w38629;// level 8
assign po08338 = ~w38632;// level 8
assign po08339 = ~w38635;// level 8
assign po08340 = ~w38638;// level 8
assign po08341 = ~w38641;// level 8
assign po08342 = ~w38644;// level 8
assign po08343 = ~w38647;// level 8
assign po08344 = ~w38650;// level 8
assign po08345 = ~w38653;// level 8
assign po08346 = ~w38656;// level 8
assign po08347 = ~w38659;// level 8
assign po08348 = ~w38662;// level 8
assign po08349 = ~w38665;// level 8
assign po08350 = ~w38668;// level 8
assign po08351 = ~w38671;// level 8
assign po08352 = ~w38674;// level 8
assign po08353 = ~w38677;// level 8
assign po08354 = ~w38680;// level 8
assign po08355 = ~w38683;// level 8
assign po08356 = ~w38686;// level 8
assign po08357 = ~w38689;// level 8
assign po08358 = ~w38692;// level 8
assign po08359 = ~w38695;// level 8
assign po08360 = ~w38698;// level 8
assign po08361 = ~w38701;// level 8
assign po08362 = ~w38704;// level 8
assign po08363 = ~w38707;// level 8
assign po08364 = ~w38710;// level 8
assign po08365 = ~w38713;// level 8
assign po08366 = ~w38716;// level 8
assign po08367 = ~w38719;// level 8
assign po08368 = ~w38722;// level 8
assign po08369 = ~w38725;// level 8
assign po08370 = ~w38728;// level 8
assign po08371 = ~w38731;// level 8
assign po08372 = ~w38734;// level 8
assign po08373 = ~w38737;// level 8
assign po08374 = ~w38740;// level 8
assign po08375 = ~w38743;// level 8
assign po08376 = ~w38746;// level 8
assign po08377 = ~w38749;// level 8
assign po08378 = ~w38752;// level 8
assign po08379 = ~w38755;// level 8
assign po08380 = ~w38758;// level 8
assign po08381 = ~w38761;// level 8
assign po08382 = ~w38764;// level 7
assign po08383 = ~w38767;// level 7
assign po08384 = ~w38770;// level 7
assign po08385 = ~w38773;// level 7
assign po08386 = ~w38776;// level 7
assign po08387 = ~w38779;// level 7
assign po08388 = ~w38782;// level 8
assign po08389 = ~w38785;// level 8
assign po08390 = ~w38788;// level 8
assign po08391 = ~w38791;// level 8
assign po08392 = ~w38794;// level 8
assign po08393 = ~w38797;// level 8
assign po08394 = ~w38800;// level 8
assign po08395 = ~w38803;// level 8
assign po08396 = ~w38806;// level 8
assign po08397 = ~w38809;// level 8
assign po08398 = ~w38812;// level 8
assign po08399 = ~w38815;// level 8
assign po08400 = ~w38818;// level 8
assign po08401 = ~w38821;// level 8
assign po08402 = ~w38824;// level 8
assign po08403 = ~w38827;// level 8
assign po08404 = ~w38830;// level 8
assign po08405 = ~w38833;// level 8
assign po08406 = ~w38836;// level 8
assign po08407 = ~w38839;// level 8
assign po08408 = ~w38842;// level 8
assign po08409 = ~w38845;// level 8
assign po08410 = ~w38848;// level 8
assign po08411 = ~w38851;// level 8
assign po08412 = ~w38854;// level 8
assign po08413 = ~w38857;// level 8
assign po08414 = ~w38861;// level 8
assign po08415 = ~w38864;// level 8
assign po08416 = ~w38867;// level 8
assign po08417 = ~w38870;// level 8
assign po08418 = ~w38873;// level 8
assign po08419 = ~w38876;// level 8
assign po08420 = ~w38879;// level 8
assign po08421 = ~w38882;// level 8
assign po08422 = ~w38885;// level 8
assign po08423 = ~w38888;// level 8
assign po08424 = ~w38891;// level 8
assign po08425 = ~w38894;// level 8
assign po08426 = ~w38897;// level 8
assign po08427 = ~w38900;// level 8
assign po08428 = ~w38903;// level 8
assign po08429 = ~w38906;// level 8
assign po08430 = ~w38909;// level 8
assign po08431 = ~w38912;// level 8
assign po08432 = ~w38915;// level 8
assign po08433 = ~w38918;// level 8
assign po08434 = ~w38921;// level 7
assign po08435 = ~w38924;// level 8
assign po08436 = ~w38927;// level 7
assign po08437 = ~w38930;// level 7
assign po08438 = ~w38933;// level 7
assign po08439 = ~w38936;// level 7
assign po08440 = ~w38939;// level 8
assign po08441 = ~w38942;// level 7
assign po08442 = ~w38945;// level 8
assign po08443 = ~w38948;// level 7
assign po08444 = ~w38951;// level 7
assign po08445 = ~w38954;// level 7
assign po08446 = ~w38957;// level 7
assign po08447 = ~w38960;// level 7
assign po08448 = ~w38963;// level 7
assign po08449 = ~w38966;// level 7
assign po08450 = ~w38969;// level 7
assign po08451 = ~w38972;// level 8
assign po08452 = ~w38975;// level 7
assign po08453 = ~w38979;// level 8
assign po08454 = ~w38982;// level 8
assign po08455 = ~w38985;// level 8
assign po08456 = ~w38988;// level 8
assign po08457 = ~w38991;// level 8
assign po08458 = ~w38994;// level 8
assign po08459 = ~w38997;// level 8
assign po08460 = ~w39000;// level 8
assign po08461 = ~w39003;// level 8
assign po08462 = ~w39006;// level 8
assign po08463 = ~w39009;// level 8
assign po08464 = ~w39012;// level 8
assign po08465 = ~w39015;// level 8
assign po08466 = ~w39018;// level 8
assign po08467 = ~w39021;// level 8
assign po08468 = ~w39024;// level 8
assign po08469 = ~w39027;// level 8
assign po08470 = ~w39030;// level 8
assign po08471 = ~w39033;// level 8
assign po08472 = ~w39036;// level 8
assign po08473 = ~w39039;// level 8
assign po08474 = ~w39042;// level 8
assign po08475 = ~w39045;// level 8
assign po08476 = ~w39048;// level 8
assign po08477 = ~w39051;// level 8
assign po08478 = ~w39054;// level 8
assign po08479 = ~w39057;// level 8
assign po08480 = ~w39060;// level 8
assign po08481 = ~w39063;// level 8
assign po08482 = ~w39066;// level 8
assign po08483 = ~w39069;// level 8
assign po08484 = ~w39072;// level 8
assign po08485 = ~w39075;// level 8
assign po08486 = ~w39078;// level 8
assign po08487 = ~w39081;// level 8
assign po08488 = ~w39084;// level 8
assign po08489 = ~w39087;// level 8
assign po08490 = ~w39090;// level 8
assign po08491 = ~w39093;// level 8
assign po08492 = ~w39096;// level 8
assign po08493 = ~w39099;// level 8
assign po08494 = ~w39102;// level 8
assign po08495 = ~w39105;// level 8
assign po08496 = ~w39108;// level 8
assign po08497 = ~w39111;// level 8
assign po08498 = ~w39114;// level 8
assign po08499 = ~w39117;// level 8
assign po08500 = ~w39120;// level 8
assign po08501 = ~w39123;// level 8
assign po08502 = ~w39126;// level 8
assign po08503 = ~w39129;// level 8
assign po08504 = ~w39132;// level 8
assign po08505 = ~w39135;// level 8
assign po08506 = ~w39138;// level 8
assign po08507 = ~w39141;// level 8
assign po08508 = ~w39144;// level 8
assign po08509 = ~w39147;// level 8
assign po08510 = ~w39150;// level 8
assign po08511 = ~w39153;// level 8
assign po08512 = ~w39156;// level 8
assign po08513 = ~w39159;// level 8
assign po08514 = ~w39162;// level 8
assign po08515 = ~w39165;// level 8
assign po08516 = ~w39168;// level 8
assign po08517 = ~w39171;// level 8
assign po08518 = ~w39174;// level 8
assign po08519 = ~w39177;// level 8
assign po08520 = ~w39180;// level 8
assign po08521 = ~w39183;// level 8
assign po08522 = ~w39186;// level 8
assign po08523 = ~w39189;// level 8
assign po08524 = ~w39192;// level 8
assign po08525 = ~w39195;// level 8
assign po08526 = ~w39198;// level 8
assign po08527 = ~w39201;// level 8
assign po08528 = ~w39204;// level 8
assign po08529 = ~w39207;// level 8
assign po08530 = ~w39210;// level 8
assign po08531 = ~w39213;// level 8
assign po08532 = ~w39216;// level 8
assign po08533 = ~w39219;// level 8
assign po08534 = ~w39222;// level 8
assign po08535 = ~w39225;// level 8
assign po08536 = ~w39228;// level 8
assign po08537 = ~w39231;// level 8
assign po08538 = ~w39234;// level 8
assign po08539 = ~w39237;// level 8
assign po08540 = ~w39240;// level 8
assign po08541 = ~w39243;// level 8
assign po08542 = ~w39246;// level 8
assign po08543 = ~w39249;// level 8
assign po08544 = ~w39252;// level 8
assign po08545 = ~w39255;// level 8
assign po08546 = ~w39258;// level 8
assign po08547 = ~w39261;// level 8
assign po08548 = ~w39264;// level 8
assign po08549 = ~w39267;// level 8
assign po08550 = ~w39270;// level 8
assign po08551 = ~w39273;// level 8
assign po08552 = ~w39276;// level 8
assign po08553 = ~w39279;// level 8
assign po08554 = ~w39282;// level 8
assign po08555 = ~w39285;// level 8
assign po08556 = ~w39288;// level 8
assign po08557 = ~w39291;// level 8
assign po08558 = ~w39294;// level 8
assign po08559 = ~w39297;// level 8
assign po08560 = ~w39300;// level 8
assign po08561 = ~w39303;// level 8
assign po08562 = ~w39306;// level 8
assign po08563 = ~w39309;// level 8
assign po08564 = ~w39312;// level 8
assign po08565 = ~w39315;// level 8
assign po08566 = ~w39318;// level 8
assign po08567 = ~w39321;// level 8
assign po08568 = ~w39324;// level 8
assign po08569 = ~w39327;// level 8
assign po08570 = ~w39330;// level 8
assign po08571 = ~w39333;// level 8
assign po08572 = ~w39336;// level 8
assign po08573 = ~w39339;// level 8
assign po08574 = ~w39342;// level 8
assign po08575 = ~w39345;// level 8
assign po08576 = ~w39348;// level 8
assign po08577 = ~w39351;// level 8
assign po08578 = ~w39354;// level 8
assign po08579 = ~w39357;// level 8
assign po08580 = ~w39360;// level 8
assign po08581 = ~w39363;// level 8
assign po08582 = ~w39366;// level 8
assign po08583 = ~w39369;// level 8
assign po08584 = ~w39372;// level 8
assign po08585 = ~w39375;// level 8
assign po08586 = ~w39378;// level 8
assign po08587 = ~w39381;// level 8
assign po08588 = ~w39384;// level 8
assign po08589 = ~w39387;// level 8
assign po08590 = ~w39390;// level 8
assign po08591 = ~w39393;// level 7
assign po08592 = ~w39396;// level 7
assign po08593 = ~w39399;// level 7
assign po08594 = ~w39402;// level 7
assign po08595 = ~w39405;// level 7
assign po08596 = ~w39408;// level 8
assign po08597 = ~w39411;// level 7
assign po08598 = ~w39414;// level 7
assign po08599 = ~w39417;// level 7
assign po08600 = ~w39420;// level 7
assign po08601 = ~w39423;// level 7
assign po08602 = ~w39426;// level 8
assign po08603 = ~w39429;// level 8
assign po08604 = ~w39432;// level 8
assign po08605 = ~w39435;// level 8
assign po08606 = ~w39438;// level 8
assign po08607 = ~w39441;// level 8
assign po08608 = ~w39444;// level 8
assign po08609 = ~w39447;// level 8
assign po08610 = ~w39450;// level 8
assign po08611 = ~w39453;// level 8
assign po08612 = ~w39456;// level 8
assign po08613 = ~w39459;// level 8
assign po08614 = ~w39462;// level 8
assign po08615 = ~w39465;// level 8
assign po08616 = ~w39468;// level 7
assign po08617 = ~w39471;// level 8
assign po08618 = ~w39474;// level 7
assign po08619 = ~w39477;// level 7
assign po08620 = ~w39480;// level 7
assign po08621 = ~w39483;// level 7
assign po08622 = ~w39486;// level 7
assign po08623 = ~w39489;// level 8
assign po08624 = ~w39492;// level 8
assign po08625 = ~w39495;// level 8
assign po08626 = ~w39498;// level 8
assign po08627 = ~w39501;// level 8
assign po08628 = ~w39504;// level 8
assign po08629 = ~w39507;// level 8
assign po08630 = ~w39510;// level 8
assign po08631 = ~w39513;// level 8
assign po08632 = ~w39516;// level 8
assign po08633 = ~w39519;// level 8
assign po08634 = ~w39522;// level 8
assign po08635 = ~w39525;// level 8
assign po08636 = ~w39528;// level 8
assign po08637 = ~w39531;// level 8
assign po08638 = ~w39534;// level 8
assign po08639 = ~w39537;// level 8
assign po08640 = ~w39540;// level 8
assign po08641 = ~w39543;// level 8
assign po08642 = ~w39546;// level 8
assign po08643 = ~w39549;// level 8
assign po08644 = ~w39552;// level 8
assign po08645 = ~w39555;// level 8
assign po08646 = ~w39558;// level 8
assign po08647 = ~w39561;// level 8
assign po08648 = ~w39564;// level 8
assign po08649 = ~w39567;// level 8
assign po08650 = ~w39570;// level 8
assign po08651 = ~w39573;// level 8
assign po08652 = ~w39576;// level 8
assign po08653 = ~w39579;// level 8
assign po08654 = ~w39582;// level 8
assign po08655 = ~w39585;// level 8
assign po08656 = ~w39588;// level 8
assign po08657 = ~w39591;// level 8
assign po08658 = ~w39594;// level 8
assign po08659 = ~w39597;// level 8
assign po08660 = ~w39600;// level 8
assign po08661 = ~w39603;// level 8
assign po08662 = ~w39606;// level 8
assign po08663 = ~w39609;// level 8
assign po08664 = ~w39612;// level 8
assign po08665 = ~w39615;// level 8
assign po08666 = ~w39618;// level 8
assign po08667 = ~w39621;// level 8
assign po08668 = ~w39624;// level 8
assign po08669 = ~w39627;// level 8
assign po08670 = ~w39630;// level 8
assign po08671 = ~w39633;// level 8
assign po08672 = ~w39636;// level 8
assign po08673 = ~w39639;// level 8
assign po08674 = ~w39642;// level 8
assign po08675 = ~w39645;// level 8
assign po08676 = ~w39648;// level 8
assign po08677 = ~w39651;// level 8
assign po08678 = ~w39654;// level 8
assign po08679 = ~w39657;// level 8
assign po08680 = ~w39660;// level 8
assign po08681 = ~w39663;// level 8
assign po08682 = ~w39666;// level 8
assign po08683 = ~w39669;// level 8
assign po08684 = ~w39672;// level 8
assign po08685 = ~w39675;// level 8
assign po08686 = ~w39678;// level 8
assign po08687 = ~w39681;// level 8
assign po08688 = ~w39684;// level 8
assign po08689 = ~w39687;// level 8
assign po08690 = ~w39690;// level 8
assign po08691 = ~w39693;// level 8
assign po08692 = ~w39696;// level 8
assign po08693 = ~w39699;// level 8
assign po08694 = ~w39702;// level 8
assign po08695 = ~w39705;// level 8
assign po08696 = ~w39708;// level 8
assign po08697 = ~w39711;// level 8
assign po08698 = ~w39714;// level 8
assign po08699 = ~w39717;// level 8
assign po08700 = ~w39720;// level 8
assign po08701 = ~w39723;// level 8
assign po08702 = ~w39726;// level 8
assign po08703 = ~w39729;// level 8
assign po08704 = ~w39732;// level 8
assign po08705 = ~w39735;// level 8
assign po08706 = ~w39738;// level 8
assign po08707 = ~w39741;// level 8
assign po08708 = ~w39744;// level 8
assign po08709 = ~w39747;// level 8
assign po08710 = ~w39750;// level 8
assign po08711 = ~w39753;// level 8
assign po08712 = ~w39756;// level 8
assign po08713 = ~w39759;// level 8
assign po08714 = ~w39762;// level 8
assign po08715 = ~w39765;// level 8
assign po08716 = ~w39768;// level 8
assign po08717 = ~w39771;// level 8
assign po08718 = ~w39774;// level 8
assign po08719 = ~w39777;// level 8
assign po08720 = ~w39780;// level 7
assign po08721 = ~w39783;// level 7
assign po08722 = ~w39786;// level 7
assign po08723 = ~w39789;// level 8
assign po08724 = ~w39792;// level 7
assign po08725 = ~w39795;// level 8
assign po08726 = ~w39798;// level 8
assign po08727 = ~w39801;// level 8
assign po08728 = ~w39804;// level 8
assign po08729 = ~w39807;// level 8
assign po08730 = ~w39810;// level 8
assign po08731 = ~w39813;// level 8
assign po08732 = ~w39816;// level 8
assign po08733 = ~w39819;// level 8
assign po08734 = ~w39822;// level 8
assign po08735 = ~w39825;// level 8
assign po08736 = ~w39828;// level 8
assign po08737 = ~w39831;// level 8
assign po08738 = ~w39834;// level 8
assign po08739 = ~w39837;// level 8
assign po08740 = ~w39840;// level 8
assign po08741 = ~w39843;// level 8
assign po08742 = ~w39846;// level 8
assign po08743 = ~w39849;// level 8
assign po08744 = ~w39852;// level 8
assign po08745 = ~w39855;// level 8
assign po08746 = ~w39858;// level 8
assign po08747 = ~w39861;// level 8
assign po08748 = ~w39864;// level 8
assign po08749 = ~w39867;// level 8
assign po08750 = ~w39870;// level 8
assign po08751 = ~w39873;// level 8
assign po08752 = ~w39876;// level 8
assign po08753 = ~w39879;// level 8
assign po08754 = ~w39882;// level 8
assign po08755 = ~w39885;// level 8
assign po08756 = ~w39888;// level 8
assign po08757 = ~w39891;// level 8
assign po08758 = ~w39894;// level 8
assign po08759 = ~w39897;// level 8
assign po08760 = ~w39900;// level 7
assign po08761 = ~w39903;// level 7
assign po08762 = ~w39906;// level 8
assign po08763 = ~w39909;// level 7
assign po08764 = ~w39912;// level 7
assign po08765 = ~w39915;// level 8
assign po08766 = ~w39918;// level 8
assign po08767 = ~w39921;// level 8
assign po08768 = ~w39924;// level 8
assign po08769 = ~w39927;// level 8
assign po08770 = ~w39930;// level 8
assign po08771 = ~w39933;// level 8
assign po08772 = ~w39936;// level 8
assign po08773 = ~w39939;// level 8
assign po08774 = ~w39942;// level 8
assign po08775 = ~w39945;// level 8
assign po08776 = ~w39948;// level 8
assign po08777 = ~w39951;// level 8
assign po08778 = ~w39954;// level 8
assign po08779 = ~w39957;// level 8
assign po08780 = ~w39960;// level 8
assign po08781 = ~w39963;// level 8
assign po08782 = ~w39966;// level 8
assign po08783 = ~w39969;// level 8
assign po08784 = ~w39972;// level 8
assign po08785 = ~w39975;// level 8
assign po08786 = ~w39978;// level 8
assign po08787 = ~w39981;// level 8
assign po08788 = ~w39984;// level 8
assign po08789 = ~w39987;// level 8
assign po08790 = ~w39990;// level 8
assign po08791 = ~w39993;// level 8
assign po08792 = ~w39996;// level 8
assign po08793 = ~w39999;// level 8
assign po08794 = ~w40002;// level 8
assign po08795 = ~w40005;// level 8
assign po08796 = ~w40008;// level 8
assign po08797 = ~w40011;// level 8
assign po08798 = ~w40014;// level 8
assign po08799 = ~w40017;// level 8
assign po08800 = ~w40020;// level 8
assign po08801 = ~w40023;// level 8
assign po08802 = ~w40026;// level 8
assign po08803 = ~w40029;// level 8
assign po08804 = ~w40032;// level 8
assign po08805 = ~w40035;// level 8
assign po08806 = ~w40038;// level 8
assign po08807 = ~w40041;// level 8
assign po08808 = ~w40044;// level 8
assign po08809 = ~w40047;// level 8
assign po08810 = ~w40050;// level 8
assign po08811 = ~w40053;// level 8
assign po08812 = ~w40056;// level 7
assign po08813 = ~w40059;// level 7
assign po08814 = ~w40062;// level 7
assign po08815 = ~w40065;// level 7
assign po08816 = ~w40068;// level 7
assign po08817 = ~w40071;// level 7
assign po08818 = ~w40074;// level 7
assign po08819 = ~w40077;// level 7
assign po08820 = ~w40080;// level 7
assign po08821 = ~w40083;// level 7
assign po08822 = ~w40086;// level 7
assign po08823 = ~w40089;// level 7
assign po08824 = ~w40092;// level 7
assign po08825 = ~w40095;// level 7
assign po08826 = ~w40098;// level 7
assign po08827 = ~w40101;// level 7
assign po08828 = ~w40104;// level 7
assign po08829 = ~w40107;// level 7
assign po08830 = ~w40111;// level 8
assign po08831 = ~w40114;// level 8
assign po08832 = ~w40117;// level 8
assign po08833 = ~w40120;// level 8
assign po08834 = ~w40123;// level 8
assign po08835 = ~w40126;// level 8
assign po08836 = ~w40129;// level 8
assign po08837 = ~w40132;// level 8
assign po08838 = ~w40135;// level 8
assign po08839 = ~w40138;// level 8
assign po08840 = ~w40141;// level 8
assign po08841 = ~w40144;// level 8
assign po08842 = ~w40147;// level 8
assign po08843 = ~w40150;// level 8
assign po08844 = ~w40153;// level 8
assign po08845 = ~w40156;// level 8
assign po08846 = ~w40159;// level 8
assign po08847 = ~w40162;// level 8
assign po08848 = ~w40165;// level 8
assign po08849 = ~w40168;// level 8
assign po08850 = ~w40171;// level 8
assign po08851 = ~w40174;// level 8
assign po08852 = ~w40177;// level 8
assign po08853 = ~w40180;// level 8
assign po08854 = ~w40183;// level 8
assign po08855 = ~w40186;// level 8
assign po08856 = ~w40189;// level 8
assign po08857 = ~w40192;// level 8
assign po08858 = ~w40195;// level 8
assign po08859 = ~w40198;// level 8
assign po08860 = ~w40201;// level 8
assign po08861 = ~w40204;// level 8
assign po08862 = ~w40207;// level 8
assign po08863 = ~w40210;// level 8
assign po08864 = ~w40213;// level 8
assign po08865 = ~w40216;// level 8
assign po08866 = ~w40219;// level 8
assign po08867 = ~w40222;// level 8
assign po08868 = ~w40225;// level 8
assign po08869 = ~w40228;// level 8
assign po08870 = ~w40231;// level 8
assign po08871 = ~w40234;// level 8
assign po08872 = ~w40237;// level 8
assign po08873 = ~w40240;// level 8
assign po08874 = ~w40243;// level 8
assign po08875 = ~w40246;// level 8
assign po08876 = ~w40249;// level 8
assign po08877 = ~w40252;// level 8
assign po08878 = ~w40255;// level 8
assign po08879 = ~w40258;// level 8
assign po08880 = ~w40261;// level 8
assign po08881 = ~w40264;// level 8
assign po08882 = ~w40267;// level 8
assign po08883 = ~w40270;// level 8
assign po08884 = ~w40273;// level 8
assign po08885 = ~w40276;// level 8
assign po08886 = ~w40279;// level 8
assign po08887 = ~w40282;// level 8
assign po08888 = ~w40285;// level 8
assign po08889 = ~w40288;// level 8
assign po08890 = ~w40291;// level 8
assign po08891 = ~w40294;// level 8
assign po08892 = ~w40297;// level 8
assign po08893 = ~w40300;// level 8
assign po08894 = ~w40303;// level 8
assign po08895 = ~w40306;// level 8
assign po08896 = ~w40309;// level 8
assign po08897 = ~w40312;// level 7
assign po08898 = ~w40315;// level 8
assign po08899 = ~w40318;// level 7
assign po08900 = ~w40321;// level 8
assign po08901 = ~w40324;// level 7
assign po08902 = ~w40327;// level 7
assign po08903 = ~w40330;// level 7
assign po08904 = ~w40333;// level 8
assign po08905 = ~w40336;// level 8
assign po08906 = ~w40339;// level 8
assign po08907 = ~w40342;// level 8
assign po08908 = ~w40345;// level 8
assign po08909 = ~w40348;// level 8
assign po08910 = ~w40351;// level 8
assign po08911 = ~w40354;// level 8
assign po08912 = ~w40357;// level 8
assign po08913 = ~w40360;// level 8
assign po08914 = ~w40363;// level 8
assign po08915 = ~w40366;// level 8
assign po08916 = ~w40369;// level 8
assign po08917 = ~w40372;// level 8
assign po08918 = ~w40375;// level 8
assign po08919 = ~w40378;// level 8
assign po08920 = ~w40381;// level 8
assign po08921 = ~w40384;// level 8
assign po08922 = ~w40387;// level 8
assign po08923 = ~w40390;// level 8
assign po08924 = ~w40393;// level 8
assign po08925 = ~w40396;// level 8
assign po08926 = ~w40399;// level 8
assign po08927 = ~w40402;// level 8
assign po08928 = ~w40405;// level 8
assign po08929 = ~w40408;// level 8
assign po08930 = ~w40411;// level 8
assign po08931 = ~w40414;// level 8
assign po08932 = ~w40417;// level 8
assign po08933 = ~w40420;// level 8
assign po08934 = ~w40423;// level 8
assign po08935 = ~w40426;// level 8
assign po08936 = ~w40429;// level 8
assign po08937 = ~w40432;// level 8
assign po08938 = ~w40435;// level 8
assign po08939 = ~w40438;// level 8
assign po08940 = ~w40441;// level 8
assign po08941 = ~w40444;// level 8
assign po08942 = ~w40447;// level 8
assign po08943 = ~w40450;// level 8
assign po08944 = ~w40453;// level 8
assign po08945 = ~w40456;// level 8
assign po08946 = ~w40459;// level 8
assign po08947 = ~w40462;// level 8
assign po08948 = ~w40465;// level 8
assign po08949 = ~w40468;// level 8
assign po08950 = ~w40471;// level 8
assign po08951 = ~w40474;// level 8
assign po08952 = ~w40477;// level 8
assign po08953 = ~w40480;// level 8
assign po08954 = ~w40483;// level 8
assign po08955 = ~w40486;// level 8
assign po08956 = ~w40489;// level 7
assign po08957 = ~w40492;// level 7
assign po08958 = ~w40495;// level 7
assign po08959 = ~w40498;// level 7
assign po08960 = ~w40501;// level 8
assign po08961 = ~w40504;// level 8
assign po08962 = ~w40507;// level 8
assign po08963 = ~w40510;// level 8
assign po08964 = ~w40513;// level 8
assign po08965 = ~w40516;// level 8
assign po08966 = ~w40519;// level 8
assign po08967 = ~w40522;// level 8
assign po08968 = ~w40525;// level 8
assign po08969 = ~w40528;// level 7
assign po08970 = ~w40531;// level 7
assign po08971 = ~w40534;// level 7
assign po08972 = ~w40537;// level 7
assign po08973 = ~w40540;// level 7
assign po08974 = ~w40543;// level 7
assign po08975 = ~w40546;// level 7
assign po08976 = ~w40549;// level 7
assign po08977 = ~w40552;// level 7
assign po08978 = ~w40555;// level 7
assign po08979 = ~w40558;// level 7
assign po08980 = ~w40561;// level 7
assign po08981 = ~w40564;// level 7
assign po08982 = ~w40567;// level 8
assign po08983 = ~w40570;// level 8
assign po08984 = ~w40573;// level 8
assign po08985 = ~w40576;// level 8
assign po08986 = ~w40579;// level 8
assign po08987 = ~w40582;// level 8
assign po08988 = ~w40585;// level 8
assign po08989 = ~w40588;// level 8
assign po08990 = ~w40591;// level 8
assign po08991 = ~w40594;// level 8
assign po08992 = ~w40597;// level 8
assign po08993 = ~w40600;// level 8
assign po08994 = ~w40603;// level 8
assign po08995 = ~w40606;// level 8
assign po08996 = ~w40609;// level 8
assign po08997 = ~w40612;// level 8
assign po08998 = ~w40615;// level 8
assign po08999 = ~w40618;// level 8
assign po09000 = ~w40621;// level 8
assign po09001 = ~w40624;// level 8
assign po09002 = ~w40627;// level 8
assign po09003 = ~w40630;// level 8
assign po09004 = ~w40633;// level 8
assign po09005 = ~w40636;// level 8
assign po09006 = ~w40639;// level 8
assign po09007 = ~w40642;// level 8
assign po09008 = ~w40645;// level 8
assign po09009 = ~w40648;// level 8
assign po09010 = ~w40651;// level 8
assign po09011 = ~w40654;// level 8
assign po09012 = ~w40657;// level 8
assign po09013 = ~w40660;// level 8
assign po09014 = ~w40663;// level 8
assign po09015 = ~w40666;// level 8
assign po09016 = ~w40669;// level 8
assign po09017 = ~w40672;// level 8
assign po09018 = ~w40675;// level 8
assign po09019 = ~w40678;// level 8
assign po09020 = ~w40681;// level 8
assign po09021 = ~w40684;// level 7
assign po09022 = ~w40687;// level 7
assign po09023 = ~w40690;// level 7
assign po09024 = ~w40693;// level 7
assign po09025 = ~w40696;// level 7
assign po09026 = ~w40699;// level 7
assign po09027 = ~w40702;// level 8
assign po09028 = ~w40705;// level 8
assign po09029 = ~w40708;// level 8
assign po09030 = ~w40711;// level 8
assign po09031 = ~w40714;// level 8
assign po09032 = ~w40717;// level 8
assign po09033 = ~w40720;// level 8
assign po09034 = ~w40723;// level 8
assign po09035 = ~w40726;// level 8
assign po09036 = ~w40729;// level 8
assign po09037 = ~w40732;// level 8
assign po09038 = ~w40735;// level 8
assign po09039 = ~w40738;// level 8
assign po09040 = ~w40741;// level 8
assign po09041 = ~w40744;// level 8
assign po09042 = ~w40747;// level 8
assign po09043 = ~w40750;// level 8
assign po09044 = ~w40753;// level 8
assign po09045 = ~w40756;// level 8
assign po09046 = ~w40759;// level 8
assign po09047 = ~w40762;// level 8
assign po09048 = ~w40765;// level 8
assign po09049 = ~w40768;// level 8
assign po09050 = ~w40771;// level 8
assign po09051 = ~w40774;// level 8
assign po09052 = ~w40777;// level 8
assign po09053 = ~w40780;// level 8
assign po09054 = ~w40783;// level 8
assign po09055 = ~w40786;// level 8
assign po09056 = ~w40789;// level 8
assign po09057 = ~w40792;// level 8
assign po09058 = ~w40795;// level 8
assign po09059 = ~w40798;// level 8
assign po09060 = ~w40801;// level 7
assign po09061 = ~w40804;// level 7
assign po09062 = ~w40807;// level 7
assign po09063 = ~w40810;// level 7
assign po09064 = ~w40813;// level 8
assign po09065 = ~w40816;// level 7
assign po09066 = ~w40819;// level 8
assign po09067 = ~w40822;// level 8
assign po09068 = ~w40825;// level 8
assign po09069 = ~w40828;// level 8
assign po09070 = ~w40831;// level 8
assign po09071 = ~w40834;// level 8
assign po09072 = ~w40837;// level 8
assign po09073 = ~w40840;// level 8
assign po09074 = ~w40843;// level 8
assign po09075 = ~w40846;// level 8
assign po09076 = ~w40849;// level 8
assign po09077 = ~w40852;// level 8
assign po09078 = ~w40855;// level 8
assign po09079 = ~w40858;// level 7
assign po09080 = ~w40861;// level 7
assign po09081 = ~w40864;// level 7
assign po09082 = ~w40867;// level 7
assign po09083 = ~w40870;// level 7
assign po09084 = ~w40873;// level 7
assign po09085 = ~w40876;// level 7
assign po09086 = ~w40879;// level 7
assign po09087 = ~w40882;// level 7
assign po09088 = ~w40885;// level 7
assign po09089 = ~w40888;// level 7
assign po09090 = ~w40891;// level 7
assign po09091 = ~w40894;// level 7
assign po09092 = ~w40897;// level 8
assign po09093 = ~w40900;// level 7
assign po09094 = ~w40903;// level 7
assign po09095 = ~w40906;// level 8
assign po09096 = ~w40909;// level 8
assign po09097 = ~w40912;// level 7
assign po09098 = ~w40915;// level 8
assign po09099 = ~w40918;// level 8
assign po09100 = ~w40921;// level 8
assign po09101 = ~w40924;// level 8
assign po09102 = ~w40927;// level 8
assign po09103 = ~w40930;// level 8
assign po09104 = ~w40933;// level 8
assign po09105 = ~w40936;// level 8
assign po09106 = ~w40939;// level 8
assign po09107 = ~w40942;// level 8
assign po09108 = ~w40945;// level 8
assign po09109 = ~w40948;// level 8
assign po09110 = ~w40951;// level 8
assign po09111 = ~w40954;// level 8
assign po09112 = ~w40957;// level 8
assign po09113 = ~w40960;// level 8
assign po09114 = ~w40963;// level 8
assign po09115 = ~w40966;// level 8
assign po09116 = ~w40969;// level 8
assign po09117 = ~w40972;// level 8
assign po09118 = ~w40975;// level 8
assign po09119 = ~w40978;// level 8
assign po09120 = ~w40981;// level 8
assign po09121 = ~w40984;// level 8
assign po09122 = ~w40987;// level 8
assign po09123 = ~w40990;// level 8
assign po09124 = ~w40993;// level 8
assign po09125 = ~w40996;// level 8
assign po09126 = ~w40999;// level 8
assign po09127 = ~w41002;// level 8
assign po09128 = ~w41005;// level 8
assign po09129 = ~w41008;// level 8
assign po09130 = ~w41011;// level 8
assign po09131 = ~w41014;// level 8
assign po09132 = ~w41017;// level 8
assign po09133 = ~w41020;// level 8
assign po09134 = ~w41023;// level 8
assign po09135 = ~w41026;// level 8
assign po09136 = ~w41029;// level 8
assign po09137 = ~w41032;// level 8
assign po09138 = ~w41035;// level 8
assign po09139 = ~w41038;// level 8
assign po09140 = ~w41041;// level 8
assign po09141 = ~w41044;// level 8
assign po09142 = ~w41047;// level 8
assign po09143 = ~w41050;// level 8
assign po09144 = ~w41053;// level 8
assign po09145 = ~w41056;// level 8
assign po09146 = ~w41059;// level 8
assign po09147 = ~w41062;// level 8
assign po09148 = ~w41065;// level 8
assign po09149 = ~w41068;// level 8
assign po09150 = ~w41071;// level 8
assign po09151 = ~w41074;// level 8
assign po09152 = ~w41077;// level 8
assign po09153 = ~w41080;// level 8
assign po09154 = ~w41083;// level 8
assign po09155 = ~w41086;// level 8
assign po09156 = ~w41089;// level 8
assign po09157 = ~w41092;// level 8
assign po09158 = ~w41095;// level 8
assign po09159 = ~w41098;// level 8
assign po09160 = ~w41101;// level 8
assign po09161 = ~w41104;// level 8
assign po09162 = ~w41107;// level 8
assign po09163 = ~w41110;// level 8
assign po09164 = ~w41113;// level 8
assign po09165 = ~w41116;// level 8
assign po09166 = ~w41119;// level 8
assign po09167 = ~w41122;// level 8
assign po09168 = ~w41125;// level 8
assign po09169 = ~w41128;// level 8
assign po09170 = ~w41131;// level 8
assign po09171 = ~w41134;// level 8
assign po09172 = ~w41137;// level 8
assign po09173 = ~w41140;// level 8
assign po09174 = ~w41143;// level 8
assign po09175 = ~w41146;// level 8
assign po09176 = ~w41149;// level 8
assign po09177 = ~w41152;// level 8
assign po09178 = ~w41155;// level 8
assign po09179 = ~w41158;// level 8
assign po09180 = ~w41161;// level 8
assign po09181 = ~w41164;// level 8
assign po09182 = ~w41167;// level 8
assign po09183 = ~w41170;// level 8
assign po09184 = ~w41173;// level 8
assign po09185 = ~w41176;// level 8
assign po09186 = ~w41179;// level 8
assign po09187 = ~w41182;// level 8
assign po09188 = ~w41185;// level 8
assign po09189 = ~w41188;// level 8
assign po09190 = ~w41191;// level 8
assign po09191 = ~w41194;// level 7
assign po09192 = ~w41197;// level 7
assign po09193 = ~w41200;// level 7
assign po09194 = ~w41203;// level 7
assign po09195 = ~w41206;// level 8
assign po09196 = ~w41209;// level 8
assign po09197 = ~w41212;// level 8
assign po09198 = ~w41215;// level 8
assign po09199 = ~w41218;// level 8
assign po09200 = ~w41221;// level 8
assign po09201 = ~w41224;// level 8
assign po09202 = ~w41227;// level 8
assign po09203 = ~w41230;// level 8
assign po09204 = ~w41233;// level 8
assign po09205 = ~w41236;// level 8
assign po09206 = ~w41239;// level 8
assign po09207 = ~w41242;// level 8
assign po09208 = ~w41245;// level 8
assign po09209 = ~w41248;// level 8
assign po09210 = ~w41251;// level 8
assign po09211 = ~w41254;// level 8
assign po09212 = ~w41257;// level 8
assign po09213 = ~w41260;// level 8
assign po09214 = ~w41263;// level 8
assign po09215 = ~w41266;// level 8
assign po09216 = ~w41269;// level 8
assign po09217 = ~w41272;// level 8
assign po09218 = ~w41275;// level 8
assign po09219 = ~w41278;// level 8
assign po09220 = ~w41281;// level 8
assign po09221 = ~w41284;// level 8
assign po09222 = ~w41287;// level 8
assign po09223 = ~w41290;// level 8
assign po09224 = ~w41293;// level 8
assign po09225 = ~w41296;// level 8
assign po09226 = ~w41299;// level 8
assign po09227 = ~w41302;// level 8
assign po09228 = ~w41305;// level 8
assign po09229 = ~w41308;// level 8
assign po09230 = ~w41311;// level 8
assign po09231 = ~w41314;// level 8
assign po09232 = ~w41317;// level 8
assign po09233 = ~w41320;// level 8
assign po09234 = ~w41323;// level 8
assign po09235 = ~w41326;// level 8
assign po09236 = ~w41329;// level 8
assign po09237 = ~w41332;// level 8
assign po09238 = ~w41335;// level 8
assign po09239 = ~w41338;// level 8
assign po09240 = ~w41341;// level 8
assign po09241 = ~w41344;// level 8
assign po09242 = ~w41347;// level 8
assign po09243 = ~w41350;// level 8
assign po09244 = ~w41353;// level 8
assign po09245 = ~w41356;// level 8
assign po09246 = ~w41359;// level 8
assign po09247 = ~w41362;// level 8
assign po09248 = ~w41365;// level 8
assign po09249 = ~w41368;// level 8
assign po09250 = ~w41371;// level 8
assign po09251 = ~w41374;// level 8
assign po09252 = ~w41377;// level 8
assign po09253 = ~w41380;// level 8
assign po09254 = ~w41383;// level 8
assign po09255 = ~w41386;// level 8
assign po09256 = ~w41389;// level 8
assign po09257 = ~w41392;// level 8
assign po09258 = ~w41395;// level 8
assign po09259 = ~w41398;// level 8
assign po09260 = ~w41401;// level 8
assign po09261 = ~w41404;// level 8
assign po09262 = ~w41407;// level 8
assign po09263 = ~w41410;// level 8
assign po09264 = ~w41413;// level 8
assign po09265 = ~w41416;// level 8
assign po09266 = ~w41419;// level 8
assign po09267 = ~w41422;// level 8
assign po09268 = ~w41425;// level 8
assign po09269 = ~w41429;// level 8
assign po09270 = ~w41432;// level 8
assign po09271 = ~w41435;// level 8
assign po09272 = ~w41438;// level 8
assign po09273 = ~w41441;// level 8
assign po09274 = ~w41444;// level 8
assign po09275 = ~w41447;// level 8
assign po09276 = ~w41450;// level 8
assign po09277 = ~w41453;// level 8
assign po09278 = ~w41456;// level 8
assign po09279 = ~w41459;// level 8
assign po09280 = ~w41462;// level 8
assign po09281 = ~w41465;// level 8
assign po09282 = ~w41468;// level 8
assign po09283 = ~w41471;// level 8
assign po09284 = ~w41474;// level 8
assign po09285 = ~w41477;// level 8
assign po09286 = ~w41480;// level 8
assign po09287 = ~w41483;// level 8
assign po09288 = ~w41486;// level 8
assign po09289 = ~w41489;// level 8
assign po09290 = ~w41492;// level 8
assign po09291 = ~w41495;// level 8
assign po09292 = ~w41498;// level 8
assign po09293 = ~w41501;// level 8
assign po09294 = ~w41504;// level 8
assign po09295 = ~w41507;// level 7
assign po09296 = ~w41510;// level 7
assign po09297 = ~w41513;// level 7
assign po09298 = ~w41516;// level 7
assign po09299 = ~w41519;// level 7
assign po09300 = ~w41522;// level 7
assign po09301 = ~w41526;// level 8
assign po09302 = ~w41529;// level 8
assign po09303 = ~w41532;// level 8
assign po09304 = ~w41535;// level 8
assign po09305 = ~w41538;// level 8
assign po09306 = ~w41541;// level 8
assign po09307 = ~w41544;// level 8
assign po09308 = ~w41547;// level 8
assign po09309 = ~w41550;// level 8
assign po09310 = ~w41553;// level 8
assign po09311 = ~w41556;// level 8
assign po09312 = ~w41559;// level 8
assign po09313 = ~w41562;// level 8
assign po09314 = ~w41565;// level 8
assign po09315 = ~w41568;// level 8
assign po09316 = ~w41571;// level 8
assign po09317 = ~w41574;// level 8
assign po09318 = ~w41577;// level 8
assign po09319 = ~w41580;// level 8
assign po09320 = ~w41583;// level 8
assign po09321 = ~w41586;// level 8
assign po09322 = ~w41589;// level 8
assign po09323 = ~w41592;// level 8
assign po09324 = ~w41595;// level 8
assign po09325 = ~w41598;// level 8
assign po09326 = ~w41601;// level 8
assign po09327 = ~w41604;// level 8
assign po09328 = ~w41607;// level 8
assign po09329 = ~w41610;// level 8
assign po09330 = ~w41613;// level 8
assign po09331 = ~w41616;// level 8
assign po09332 = ~w41619;// level 8
assign po09333 = ~w41622;// level 8
assign po09334 = ~w41625;// level 8
assign po09335 = ~w41628;// level 8
assign po09336 = ~w41631;// level 8
assign po09337 = ~w41634;// level 8
assign po09338 = ~w41637;// level 8
assign po09339 = ~w41640;// level 8
assign po09340 = ~w41643;// level 8
assign po09341 = ~w41646;// level 8
assign po09342 = ~w41649;// level 8
assign po09343 = ~w41652;// level 8
assign po09344 = ~w41655;// level 8
assign po09345 = ~w41658;// level 8
assign po09346 = ~w41661;// level 8
assign po09347 = ~w41664;// level 8
assign po09348 = ~w41667;// level 8
assign po09349 = ~w41670;// level 8
assign po09350 = ~w41673;// level 8
assign po09351 = ~w41676;// level 8
assign po09352 = ~w41679;// level 8
assign po09353 = ~w41682;// level 8
assign po09354 = ~w41685;// level 8
assign po09355 = ~w41688;// level 8
assign po09356 = ~w41691;// level 8
assign po09357 = ~w41694;// level 8
assign po09358 = ~w41697;// level 8
assign po09359 = ~w41700;// level 8
assign po09360 = ~w41703;// level 8
assign po09361 = ~w41706;// level 8
assign po09362 = ~w41709;// level 8
assign po09363 = ~w41712;// level 8
assign po09364 = ~w41715;// level 8
assign po09365 = ~w41718;// level 8
assign po09366 = ~w41721;// level 8
assign po09367 = ~w41724;// level 8
assign po09368 = ~w41727;// level 7
assign po09369 = ~w41730;// level 8
assign po09370 = ~w41733;// level 8
assign po09371 = ~w41736;// level 8
assign po09372 = ~w41739;// level 8
assign po09373 = ~w41742;// level 8
assign po09374 = ~w41745;// level 8
assign po09375 = ~w41748;// level 8
assign po09376 = ~w41751;// level 8
assign po09377 = ~w41754;// level 8
assign po09378 = ~w41757;// level 8
assign po09379 = ~w41760;// level 8
assign po09380 = ~w41763;// level 8
assign po09381 = ~w41766;// level 8
assign po09382 = ~w41769;// level 8
assign po09383 = ~w41772;// level 8
assign po09384 = ~w41775;// level 8
assign po09385 = ~w41778;// level 8
assign po09386 = ~w41781;// level 8
assign po09387 = ~w41784;// level 8
assign po09388 = ~w41787;// level 8
assign po09389 = ~w41790;// level 8
assign po09390 = ~w41793;// level 8
assign po09391 = ~w41796;// level 8
assign po09392 = ~w41799;// level 8
assign po09393 = ~w41802;// level 8
assign po09394 = ~w41805;// level 8
assign po09395 = ~w41808;// level 8
assign po09396 = ~w41811;// level 8
assign po09397 = ~w41814;// level 8
assign po09398 = ~w41817;// level 8
assign po09399 = ~w41820;// level 8
assign po09400 = ~w41823;// level 8
assign po09401 = ~w41826;// level 8
assign po09402 = ~w41829;// level 8
assign po09403 = ~w41832;// level 8
assign po09404 = ~w41835;// level 8
assign po09405 = ~w41838;// level 8
assign po09406 = ~w41841;// level 8
assign po09407 = ~w41844;// level 8
assign po09408 = ~w41847;// level 8
assign po09409 = ~w41850;// level 8
assign po09410 = ~w41853;// level 8
assign po09411 = ~w41856;// level 8
assign po09412 = ~w41859;// level 8
assign po09413 = ~w41862;// level 8
assign po09414 = ~w41865;// level 8
assign po09415 = ~w41868;// level 8
assign po09416 = ~w41871;// level 8
assign po09417 = ~w41874;// level 8
assign po09418 = ~w41877;// level 8
assign po09419 = ~w41880;// level 8
assign po09420 = ~w41883;// level 8
assign po09421 = ~w41886;// level 8
assign po09422 = ~w41889;// level 8
assign po09423 = ~w41892;// level 8
assign po09424 = ~w41895;// level 8
assign po09425 = ~w41898;// level 8
assign po09426 = ~w41901;// level 8
assign po09427 = ~w41904;// level 8
assign po09428 = ~w41907;// level 8
assign po09429 = ~w41910;// level 8
assign po09430 = ~w41913;// level 8
assign po09431 = ~w41916;// level 8
assign po09432 = ~w41919;// level 8
assign po09433 = ~w41922;// level 8
assign po09434 = ~w41925;// level 8
assign po09435 = ~w41928;// level 8
assign po09436 = ~w41931;// level 8
assign po09437 = ~w41934;// level 8
assign po09438 = ~w41937;// level 8
assign po09439 = ~w41940;// level 8
assign po09440 = ~w41943;// level 8
assign po09441 = ~w41946;// level 8
assign po09442 = ~w41949;// level 8
assign po09443 = ~w41952;// level 8
assign po09444 = ~w41955;// level 8
assign po09445 = ~w41958;// level 8
assign po09446 = ~w41961;// level 8
assign po09447 = ~w41964;// level 8
assign po09448 = ~w41967;// level 8
assign po09449 = ~w41970;// level 8
assign po09450 = ~w41973;// level 8
assign po09451 = ~w41976;// level 8
assign po09452 = ~w41979;// level 7
assign po09453 = ~w41982;// level 7
assign po09454 = ~w41985;// level 7
assign po09455 = ~w41988;// level 7
assign po09456 = ~w41991;// level 7
assign po09457 = ~w41994;// level 7
assign po09458 = ~w41997;// level 7
assign po09459 = ~w42000;// level 7
assign po09460 = ~w42003;// level 7
assign po09461 = ~w42006;// level 7
assign po09462 = ~w42009;// level 7
assign po09463 = ~w42012;// level 7
assign po09464 = ~w42015;// level 7
assign po09465 = ~w42018;// level 7
assign po09466 = ~w42021;// level 7
assign po09467 = ~w42024;// level 7
assign po09468 = ~w42027;// level 8
assign po09469 = ~w42030;// level 7
assign po09470 = ~w42033;// level 7
assign po09471 = ~w42037;// level 8
assign po09472 = ~w42040;// level 8
assign po09473 = ~w42043;// level 8
assign po09474 = ~w42046;// level 8
assign po09475 = ~w42049;// level 8
assign po09476 = ~w42052;// level 8
assign po09477 = ~w42055;// level 8
assign po09478 = ~w42058;// level 8
assign po09479 = ~w42061;// level 8
assign po09480 = ~w42064;// level 8
assign po09481 = ~w42067;// level 8
assign po09482 = ~w42070;// level 8
assign po09483 = ~w42073;// level 8
assign po09484 = ~w42076;// level 8
assign po09485 = ~w42079;// level 7
assign po09486 = ~w42082;// level 7
assign po09487 = ~w42085;// level 7
assign po09488 = ~w42088;// level 7
assign po09489 = ~w42091;// level 7
assign po09490 = ~w42094;// level 7
assign po09491 = ~w42097;// level 7
assign po09492 = ~w42100;// level 7
assign po09493 = ~w42103;// level 7
assign po09494 = ~w42106;// level 7
assign po09495 = ~w42109;// level 7
assign po09496 = ~w42112;// level 8
assign po09497 = ~w42115;// level 7
assign po09498 = ~w42118;// level 7
assign po09499 = ~w42121;// level 7
assign po09500 = ~w42124;// level 7
assign po09501 = ~w42127;// level 7
assign po09502 = ~w42130;// level 7
assign po09503 = ~w42133;// level 7
assign po09504 = ~w42136;// level 7
assign po09505 = ~w42139;// level 8
assign po09506 = ~w42142;// level 8
assign po09507 = ~w42145;// level 8
assign po09508 = ~w42148;// level 8
assign po09509 = ~w42151;// level 8
assign po09510 = ~w42154;// level 8
assign po09511 = ~w42157;// level 8
assign po09512 = ~w42160;// level 8
assign po09513 = ~w42163;// level 8
assign po09514 = ~w42166;// level 8
assign po09515 = ~w42169;// level 8
assign po09516 = ~w42172;// level 8
assign po09517 = ~w42175;// level 8
assign po09518 = ~w42178;// level 8
assign po09519 = ~w42181;// level 8
assign po09520 = ~w42184;// level 8
assign po09521 = ~w42187;// level 8
assign po09522 = ~w42190;// level 8
assign po09523 = ~w42193;// level 8
assign po09524 = ~w42196;// level 8
assign po09525 = ~w42199;// level 8
assign po09526 = ~w42202;// level 8
assign po09527 = ~w42205;// level 8
assign po09528 = ~w42208;// level 8
assign po09529 = ~w42211;// level 8
assign po09530 = ~w42214;// level 8
assign po09531 = ~w42217;// level 8
assign po09532 = ~w42220;// level 8
assign po09533 = ~w42223;// level 8
assign po09534 = ~w42226;// level 8
assign po09535 = ~w42229;// level 8
assign po09536 = ~w42232;// level 8
assign po09537 = ~w42235;// level 8
assign po09538 = ~w42238;// level 7
assign po09539 = ~w42241;// level 7
assign po09540 = ~w42244;// level 7
assign po09541 = ~w42247;// level 7
assign po09542 = ~w42250;// level 7
assign po09543 = ~w42253;// level 7
assign po09544 = ~w42256;// level 7
assign po09545 = ~w42259;// level 8
assign po09546 = ~w42262;// level 8
assign po09547 = ~w42265;// level 8
assign po09548 = ~w42268;// level 8
assign po09549 = ~w42271;// level 8
assign po09550 = ~w42274;// level 8
assign po09551 = ~w42277;// level 8
assign po09552 = ~w42280;// level 8
assign po09553 = ~w42283;// level 8
assign po09554 = ~w42286;// level 8
assign po09555 = ~w42289;// level 8
assign po09556 = ~w42292;// level 8
assign po09557 = ~w42295;// level 8
assign po09558 = ~w42298;// level 8
assign po09559 = ~w42301;// level 8
assign po09560 = ~w42304;// level 8
assign po09561 = ~w42307;// level 8
assign po09562 = ~w42310;// level 8
assign po09563 = ~w42313;// level 8
assign po09564 = ~w42316;// level 8
assign po09565 = ~w42319;// level 8
assign po09566 = ~w42322;// level 8
assign po09567 = ~w42325;// level 8
assign po09568 = ~w42328;// level 8
assign po09569 = ~w42331;// level 8
assign po09570 = ~w42334;// level 8
assign po09571 = ~w42337;// level 8
assign po09572 = ~w42340;// level 8
assign po09573 = ~w42343;// level 8
assign po09574 = ~w42346;// level 8
assign po09575 = ~w42349;// level 8
assign po09576 = ~w42352;// level 8
assign po09577 = ~w42355;// level 8
assign po09578 = ~w42358;// level 7
assign po09579 = ~w42361;// level 7
assign po09580 = ~w42364;// level 7
assign po09581 = ~w42367;// level 7
assign po09582 = ~w42370;// level 7
assign po09583 = ~w42373;// level 7
assign po09584 = ~w42376;// level 7
assign po09585 = ~w42379;// level 8
assign po09586 = ~w42382;// level 8
assign po09587 = ~w42385;// level 8
assign po09588 = ~w42388;// level 8
assign po09589 = ~w42391;// level 8
assign po09590 = ~w42394;// level 8
assign po09591 = ~w42397;// level 8
assign po09592 = ~w42400;// level 8
assign po09593 = ~w42403;// level 8
assign po09594 = ~w42406;// level 8
assign po09595 = ~w42409;// level 8
assign po09596 = ~w42412;// level 8
assign po09597 = ~w42415;// level 8
assign po09598 = ~w42418;// level 8
assign po09599 = ~w42421;// level 8
assign po09600 = ~w42424;// level 8
assign po09601 = ~w42427;// level 8
assign po09602 = ~w42430;// level 8
assign po09603 = ~w42433;// level 8
assign po09604 = ~w42436;// level 8
assign po09605 = ~w42439;// level 7
assign po09606 = ~w42442;// level 7
assign po09607 = ~w42445;// level 7
assign po09608 = ~w42448;// level 7
assign po09609 = ~w42451;// level 8
assign po09610 = ~w42454;// level 7
assign po09611 = ~w42457;// level 7
assign po09612 = ~w42460;// level 8
assign po09613 = ~w42463;// level 8
assign po09614 = ~w42466;// level 8
assign po09615 = ~w42469;// level 8
assign po09616 = ~w42472;// level 8
assign po09617 = ~w42475;// level 8
assign po09618 = ~w42478;// level 7
assign po09619 = ~w42481;// level 7
assign po09620 = ~w42484;// level 7
assign po09621 = ~w42487;// level 8
assign po09622 = ~w42490;// level 7
assign po09623 = ~w42493;// level 8
assign po09624 = ~w42496;// level 7
assign po09625 = ~w42499;// level 7
assign po09626 = ~w42502;// level 7
assign po09627 = ~w42505;// level 7
assign po09628 = ~w42508;// level 7
assign po09629 = ~w42511;// level 7
assign po09630 = ~w42514;// level 7
assign po09631 = ~w42517;// level 8
assign po09632 = ~w42521;// level 8
assign po09633 = ~w42524;// level 8
assign po09634 = ~w42527;// level 8
assign po09635 = ~w42530;// level 8
assign po09636 = ~w42533;// level 8
assign po09637 = ~w42536;// level 8
assign po09638 = ~w42539;// level 8
assign po09639 = ~w42542;// level 8
assign po09640 = ~w42545;// level 8
assign po09641 = ~w42548;// level 8
assign po09642 = ~w42551;// level 8
assign po09643 = ~w42554;// level 8
assign po09644 = ~w42557;// level 8
assign po09645 = ~w42565;// level 5
assign po09646 = ~w42568;// level 8
assign po09647 = ~w42571;// level 8
assign po09648 = ~w42574;// level 8
assign po09649 = ~w42577;// level 8
assign po09650 = ~w42580;// level 8
assign po09651 = ~w42583;// level 8
assign po09652 = ~w42586;// level 8
assign po09653 = ~w42589;// level 8
assign po09654 = ~w42592;// level 8
assign po09655 = ~w42595;// level 8
assign po09656 = ~w42598;// level 8
assign po09657 = ~w42601;// level 8
assign po09658 = ~w42604;// level 8
assign po09659 = ~w42607;// level 8
assign po09660 = ~w42610;// level 8
assign po09661 = ~w42613;// level 8
assign po09662 = ~w42616;// level 8
assign po09663 = ~w42619;// level 8
assign po09664 = ~w42622;// level 8
assign po09665 = ~w42625;// level 8
assign po09666 = ~w42628;// level 8
assign po09667 = ~w42631;// level 8
assign po09668 = ~w42634;// level 8
assign po09669 = ~w42637;// level 8
assign po09670 = ~w42640;// level 8
assign po09671 = ~w42643;// level 8
assign po09672 = ~w42646;// level 8
assign po09673 = ~w42649;// level 8
assign po09674 = ~w42652;// level 8
assign po09675 = ~w42655;// level 8
assign po09676 = ~w42658;// level 8
assign po09677 = ~w42661;// level 8
assign po09678 = ~w42664;// level 8
assign po09679 = ~w42667;// level 8
assign po09680 = ~w42670;// level 8
assign po09681 = ~w42673;// level 8
assign po09682 = ~w42676;// level 8
assign po09683 = ~w42679;// level 8
assign po09684 = ~w42682;// level 8
assign po09685 = ~w42685;// level 8
assign po09686 = ~w42688;// level 8
assign po09687 = ~w42691;// level 8
assign po09688 = ~w42694;// level 8
assign po09689 = ~w42697;// level 8
assign po09690 = ~w42700;// level 8
assign po09691 = ~w42703;// level 8
assign po09692 = ~w42706;// level 8
assign po09693 = ~w42709;// level 8
assign po09694 = ~w42712;// level 8
assign po09695 = ~w42715;// level 8
assign po09696 = ~w42718;// level 8
assign po09697 = ~w42721;// level 8
assign po09698 = ~w42724;// level 8
assign po09699 = ~w42727;// level 8
assign po09700 = ~w42730;// level 8
assign po09701 = ~w42733;// level 8
assign po09702 = ~w42736;// level 8
assign po09703 = ~w42739;// level 8
assign po09704 = ~w42742;// level 8
assign po09705 = ~w42745;// level 8
assign po09706 = ~w42748;// level 8
assign po09707 = ~w42751;// level 8
assign po09708 = ~w42754;// level 8
assign po09709 = ~w42757;// level 8
assign po09710 = ~w42760;// level 8
assign po09711 = ~w42763;// level 8
assign po09712 = ~w42766;// level 8
assign po09713 = ~w42769;// level 8
assign po09714 = ~w42772;// level 8
assign po09715 = ~w42775;// level 8
assign po09716 = ~w42778;// level 8
assign po09717 = ~w42781;// level 8
assign po09718 = ~w42784;// level 8
assign po09719 = ~w42787;// level 8
assign po09720 = ~w42790;// level 8
assign po09721 = ~w42793;// level 8
assign po09722 = ~w42796;// level 8
assign po09723 = ~w42799;// level 8
assign po09724 = ~w42802;// level 8
assign po09725 = ~w42805;// level 8
assign po09726 = ~w42808;// level 8
assign po09727 = ~w42811;// level 8
assign po09728 = ~w42814;// level 8
assign po09729 = ~w42817;// level 8
assign po09730 = ~w42820;// level 8
assign po09731 = ~w42823;// level 8
assign po09732 = ~w42826;// level 8
assign po09733 = ~w42829;// level 8
assign po09734 = ~w42832;// level 8
assign po09735 = ~w42835;// level 8
assign po09736 = ~w42838;// level 8
assign po09737 = ~w42841;// level 8
assign po09738 = ~w42844;// level 8
assign po09739 = ~w42847;// level 8
assign po09740 = ~w42850;// level 8
assign po09741 = ~w42853;// level 8
assign po09742 = ~w42856;// level 8
assign po09743 = ~w42859;// level 8
assign po09744 = ~w42862;// level 8
assign po09745 = ~w42865;// level 8
assign po09746 = ~w42868;// level 8
assign po09747 = ~w42871;// level 8
assign po09748 = ~w42874;// level 8
assign po09749 = ~w42877;// level 8
assign po09750 = ~w42880;// level 8
assign po09751 = ~w42883;// level 8
assign po09752 = ~w42886;// level 8
assign po09753 = ~w42889;// level 8
assign po09754 = ~w42892;// level 8
assign po09755 = ~w42895;// level 8
assign po09756 = ~w42898;// level 8
assign po09757 = ~w42901;// level 8
assign po09758 = ~w42904;// level 8
assign po09759 = ~w42907;// level 8
assign po09760 = ~w42910;// level 8
assign po09761 = ~w42913;// level 8
assign po09762 = ~w42916;// level 8
assign po09763 = ~w42919;// level 8
assign po09764 = ~w42922;// level 8
assign po09765 = ~w42925;// level 8
assign po09766 = ~w42928;// level 8
assign po09767 = ~w42931;// level 8
assign po09768 = ~w42934;// level 8
assign po09769 = ~w42937;// level 8
assign po09770 = ~w42940;// level 8
assign po09771 = ~w42943;// level 8
assign po09772 = ~w42946;// level 8
assign po09773 = ~w42949;// level 8
assign po09774 = ~w42952;// level 8
assign po09775 = ~w42955;// level 8
assign po09776 = ~w42958;// level 8
assign po09777 = ~w42961;// level 8
assign po09778 = ~w42964;// level 8
assign po09779 = ~w42967;// level 8
assign po09780 = ~w42970;// level 8
assign po09781 = ~w42973;// level 8
assign po09782 = ~w42976;// level 8
assign po09783 = ~w42979;// level 8
assign po09784 = ~w42982;// level 8
assign po09785 = ~w42985;// level 8
assign po09786 = ~w42988;// level 8
assign po09787 = ~w42991;// level 8
assign po09788 = ~w42994;// level 8
assign po09789 = ~w42997;// level 8
assign po09790 = ~w43000;// level 8
assign po09791 = ~w43003;// level 8
assign po09792 = ~w43006;// level 8
assign po09793 = ~w43009;// level 8
assign po09794 = ~w43012;// level 8
assign po09795 = ~w43015;// level 8
assign po09796 = ~w43018;// level 8
assign po09797 = ~w43021;// level 8
assign po09798 = ~w43024;// level 8
assign po09799 = ~w43027;// level 8
assign po09800 = ~w43030;// level 8
assign po09801 = ~w43033;// level 8
assign po09802 = ~w43036;// level 8
assign po09803 = ~w43039;// level 8
assign po09804 = ~w43042;// level 8
assign po09805 = ~w43045;// level 8
assign po09806 = ~w43048;// level 8
assign po09807 = ~w43051;// level 8
assign po09808 = ~w43054;// level 8
assign po09809 = ~w43057;// level 8
assign po09810 = ~w43060;// level 8
assign po09811 = ~w43063;// level 8
assign po09812 = ~w43066;// level 8
assign po09813 = ~w43069;// level 8
assign po09814 = ~w43072;// level 8
assign po09815 = ~w43075;// level 8
assign po09816 = ~w43078;// level 8
assign po09817 = ~w43081;// level 8
assign po09818 = ~w43084;// level 8
assign po09819 = ~w43087;// level 8
assign po09820 = ~w43090;// level 8
assign po09821 = ~w43093;// level 8
assign po09822 = ~w43096;// level 8
assign po09823 = ~w43099;// level 8
assign po09824 = ~w43102;// level 8
assign po09825 = ~w43105;// level 8
assign po09826 = ~w43108;// level 8
assign po09827 = ~w43111;// level 8
assign po09828 = ~w43114;// level 8
assign po09829 = ~w43117;// level 8
assign po09830 = ~w43120;// level 8
assign po09831 = ~w43123;// level 8
assign po09832 = ~w43126;// level 8
assign po09833 = ~w43129;// level 8
assign po09834 = ~w43132;// level 8
assign po09835 = ~w43135;// level 8
assign po09836 = ~w43138;// level 8
assign po09837 = ~w43141;// level 8
assign po09838 = ~w43144;// level 8
assign po09839 = ~w43147;// level 8
assign po09840 = ~w43150;// level 8
assign po09841 = ~w43153;// level 8
assign po09842 = ~w43156;// level 8
assign po09843 = ~w43159;// level 8
assign po09844 = ~w43162;// level 8
assign po09845 = ~w43165;// level 8
assign po09846 = ~w43168;// level 8
assign po09847 = ~w43171;// level 8
assign po09848 = ~w43174;// level 8
assign po09849 = ~w43177;// level 8
assign po09850 = ~w43180;// level 8
assign po09851 = ~w43183;// level 8
assign po09852 = ~w43186;// level 8
assign po09853 = ~w43189;// level 8
assign po09854 = ~w43192;// level 8
assign po09855 = ~w43195;// level 8
assign po09856 = ~w43198;// level 8
assign po09857 = ~w43201;// level 8
assign po09858 = ~w43204;// level 8
assign po09859 = ~w43207;// level 8
assign po09860 = ~w43210;// level 8
assign po09861 = ~w43213;// level 8
assign po09862 = ~w43216;// level 8
assign po09863 = ~w43219;// level 8
assign po09864 = ~w43222;// level 8
assign po09865 = ~w43225;// level 8
assign po09866 = ~w43228;// level 8
assign po09867 = ~w43231;// level 8
assign po09868 = ~w43234;// level 8
assign po09869 = ~w43237;// level 8
assign po09870 = ~w43240;// level 8
assign po09871 = ~w43243;// level 8
assign po09872 = ~w43246;// level 8
assign po09873 = ~w43249;// level 8
assign po09874 = ~w43252;// level 8
assign po09875 = ~w43255;// level 8
assign po09876 = ~w43258;// level 8
assign po09877 = ~w43261;// level 8
assign po09878 = ~w43264;// level 8
assign po09879 = ~w43267;// level 8
assign po09880 = ~w43270;// level 8
assign po09881 = ~w43273;// level 8
assign po09882 = ~w43276;// level 8
assign po09883 = ~w43279;// level 8
assign po09884 = ~w43282;// level 8
assign po09885 = ~w43285;// level 8
assign po09886 = ~w43288;// level 8
assign po09887 = ~w43291;// level 8
assign po09888 = ~w43294;// level 8
assign po09889 = ~w43297;// level 8
assign po09890 = ~w43300;// level 8
assign po09891 = ~w43303;// level 8
assign po09892 = ~w43306;// level 8
assign po09893 = ~w43309;// level 8
assign po09894 = ~w43312;// level 8
assign po09895 = ~w43315;// level 8
assign po09896 = ~w43318;// level 8
assign po09897 = ~w43321;// level 8
assign po09898 = ~w43324;// level 8
assign po09899 = ~w43327;// level 8
assign po09900 = ~w43330;// level 8
assign po09901 = ~w43333;// level 8
assign po09902 = ~w43336;// level 8
assign po09903 = ~w43339;// level 8
assign po09904 = ~w43342;// level 8
assign po09905 = ~w43345;// level 8
assign po09906 = ~w43348;// level 8
assign po09907 = ~w43351;// level 7
assign po09908 = ~w43354;// level 8
assign po09909 = ~w43357;// level 8
assign po09910 = ~w43360;// level 8
assign po09911 = ~w43363;// level 8
assign po09912 = ~w43366;// level 8
assign po09913 = ~w43369;// level 7
assign po09914 = ~w43372;// level 8
assign po09915 = ~w43375;// level 8
assign po09916 = ~w43378;// level 8
assign po09917 = ~w43381;// level 8
assign po09918 = ~w43384;// level 8
assign po09919 = ~w43387;// level 8
assign po09920 = ~w43390;// level 8
assign po09921 = ~w43393;// level 8
assign po09922 = ~w43396;// level 8
assign po09923 = ~w43399;// level 8
assign po09924 = ~w43403;// level 7
assign po09925 = ~w43407;// level 7
assign po09926 = ~w43410;// level 7
assign po09927 = ~w43414;// level 8
assign po09928 = ~w43419;// level 8
assign po09929 = ~w43423;// level 7
assign po09930 = ~w43426;// level 7
assign po09931 = ~w43430;// level 7
assign po09932 = ~w43448;// level 9
assign po09933 = ~w43466;// level 9
assign po09934 = ~w43469;// level 7
assign po09935 = ~w43472;// level 7
assign po09936 = ~w43476;// level 8
assign po09937 = ~w43479;// level 8
assign po09938 = ~w43484;// level 9
assign po09939 = ~w43488;// level 7
assign po09940 = ~w43491;// level 7
assign po09941 = w43495;// level 8
assign po09942 = ~w43499;// level 7
assign po09943 = ~w43502;// level 7
assign po09944 = ~w43506;// level 5
assign po09945 = w43515;// level 6
assign po09946 = w43523;// level 9
assign po09947 = ~w43524;// level 8
assign po09948 = w43527;// level 8
assign po09949 = ~w43532;// level 7
assign po09950 = w43536;// level 6
assign po09951 = w43539;// level 6
assign po09952 = ~w43542;// level 7
assign po09953 = ~w43545;// level 7
assign po09954 = ~w43548;// level 7
assign po09955 = ~w43551;// level 7
assign po09956 = ~w43554;// level 7
assign po09957 = ~w43557;// level 7
assign po09958 = ~w43560;// level 8
assign po09959 = w43563;// level 8
assign po09960 = w43566;// level 8
assign po09961 = w43569;// level 8
assign po09962 = w43572;// level 8
assign po09963 = w43575;// level 8
assign po09964 = w43578;// level 8
assign po09965 = ~w43580;// level 9
assign po09966 = w43584;// level 7
assign po09967 = w43587;// level 7
assign po09968 = ~w43590;// level 7
assign po09969 = w43593;// level 7
assign po09970 = w43596;// level 7
assign po09971 = w43599;// level 7
assign po09972 = ~w43602;// level 7
assign po09973 = ~w43605;// level 7
assign po09974 = ~w43610;// level 9
assign po09975 = ~w43614;// level 7
assign po09976 = ~w43617;// level 7
assign po09977 = ~w43620;// level 7
assign po09978 = w43623;// level 7
assign po09979 = w43626;// level 7
assign po09980 = ~w43629;// level 8
assign po09981 = ~w43631;// level 6
assign po09982 = w43634;// level 6
assign po09983 = ~w43637;// level 8
assign po09984 = ~w43640;// level 8
assign po09985 = w43643;// level 7
assign po09986 = ~w43646;// level 7
assign po09987 = ~w43649;// level 7
assign po09988 = ~w43652;// level 7
assign po09989 = ~w43656;// level 8
assign po09990 = ~w43659;// level 7
assign po09991 = w43671;// level 7
assign po09992 = w43674;// level 9
assign po09993 = w43677;// level 8
assign po09994 = ~w43680;// level 7
assign po09995 = w43683;// level 7
assign po09996 = w43686;// level 7
assign po09997 = ~w43689;// level 7
assign po09998 = ~w43692;// level 7
assign po09999 = ~w43695;// level 7
assign po10000 = ~w43698;// level 8
assign po10001 = ~w43702;// level 7
assign po10002 = ~w43705;// level 8
assign po10003 = ~w43708;// level 7
assign po10004 = ~w43711;// level 8
assign po10005 = ~w43714;// level 7
assign po10006 = ~w43717;// level 8
assign po10007 = ~w43720;// level 7
assign po10008 = ~w43723;// level 7
assign po10009 = ~w43726;// level 7
assign po10010 = ~w43730;// level 7
assign po10011 = ~w43733;// level 7
assign po10012 = ~w43736;// level 7
assign po10013 = ~w43739;// level 7
assign po10014 = ~w43742;// level 7
assign po10015 = ~w43745;// level 7
assign po10016 = ~w43748;// level 7
assign po10017 = ~w43751;// level 8
assign po10018 = ~w43754;// level 7
assign po10019 = ~w43757;// level 7
assign po10020 = ~w43760;// level 8
assign po10021 = ~w43763;// level 8
assign po10022 = ~w43767;// level 7
assign po10023 = ~w43770;// level 7
assign po10024 = ~w43773;// level 7
assign po10025 = ~w43776;// level 7
assign po10026 = ~w43779;// level 7
assign po10027 = ~w43782;// level 7
assign po10028 = ~w43785;// level 7
assign po10029 = ~w43788;// level 7
assign po10030 = ~w43792;// level 7
assign po10031 = ~w43795;// level 7
assign po10032 = ~w43798;// level 7
assign po10033 = ~w43801;// level 7
assign po10034 = ~w43804;// level 7
assign po10035 = ~w43807;// level 7
assign po10036 = ~w43810;// level 7
assign po10037 = ~w43813;// level 7
assign po10038 = w43816;// level 5
assign po10039 = ~w43819;// level 7
assign po10040 = ~w43822;// level 7
assign po10041 = ~w43825;// level 7
assign po10042 = ~w43828;// level 7
assign po10043 = ~w43831;// level 7
assign po10044 = ~w43834;// level 7
assign po10045 = ~w43837;// level 7
assign po10046 = ~w43854;// level 9
assign po10047 = ~w43871;// level 9
assign po10048 = ~w43888;// level 9
assign po10049 = w43890;// level 5
assign po10050 = w43905;// level 7
assign po10051 = w43911;// level 6
assign po10052 = w43914;// level 4
assign po10053 = w43921;// level 8
assign po10054 = ~w43926;// level 6
assign po10055 = ~w43931;// level 5
assign po10056 = w43934;// level 6
assign po10057 = w66;// level 5
assign po10058 = ~pi10350;// level 0
assign po10059 = ~w43939;// level 5
assign po10060 = ~w43943;// level 8
assign po10061 = ~w43946;// level 8
assign po10062 = ~w43949;// level 8
assign po10063 = ~w43953;// level 8
assign po10064 = ~w43956;// level 8
assign po10065 = ~w43961;// level 8
assign po10066 = ~w43964;// level 8
assign po10067 = ~w43967;// level 8
assign po10068 = ~w43970;// level 8
assign po10069 = ~w43974;// level 8
assign po10070 = ~w43978;// level 8
assign po10071 = ~w43981;// level 8
assign po10072 = ~w43984;// level 8
assign po10073 = ~w43987;// level 8
assign po10074 = ~w43990;// level 8
assign po10075 = ~w43994;// level 8
assign po10076 = ~w43997;// level 8
assign po10077 = ~w44000;// level 8
assign po10078 = ~w44003;// level 8
assign po10079 = w44006;// level 7
assign po10080 = ~w44009;// level 9
assign po10081 = w44014;// level 7
assign po10082 = ~w44017;// level 6
assign po10083 = ~w44020;// level 6
assign po10084 = w44024;// level 8
assign po10085 = w44027;// level 6
assign po10086 = ~w44030;// level 9
assign po10087 = ~w44033;// level 9
assign po10088 = ~w44036;// level 9
assign po10089 = w44040;// level 7
assign po10090 = w21604;// level 8
assign po10091 = ~w44045;// level 6
assign po10092 = ~w44047;// level 8
assign po10093 = ~w44050;// level 8
assign po10094 = ~w44053;// level 8
assign po10095 = ~w44056;// level 8
assign po10096 = ~w44059;// level 8
assign po10097 = ~w44062;// level 8
assign po10098 = ~w44065;// level 8
assign po10099 = ~w44068;// level 8
assign po10100 = ~w44071;// level 8
assign po10101 = ~w44074;// level 8
assign po10102 = ~w44077;// level 8
assign po10103 = ~w44080;// level 8
assign po10104 = ~w44083;// level 8
assign po10105 = ~w44086;// level 8
assign po10106 = ~w44089;// level 8
assign po10107 = ~w44092;// level 8
assign po10108 = ~w44095;// level 8
assign po10109 = ~w44098;// level 8
assign po10110 = ~w44101;// level 8
assign po10111 = ~w44104;// level 8
assign po10112 = ~w44107;// level 8
assign po10113 = ~w44110;// level 8
assign po10114 = ~w44113;// level 8
assign po10115 = ~w44116;// level 8
assign po10116 = ~w44119;// level 8
assign po10117 = ~w44122;// level 8
assign po10118 = ~w44125;// level 8
assign po10119 = ~w44128;// level 8
assign po10120 = ~w44131;// level 8
assign po10121 = ~w44134;// level 8
assign po10122 = ~w44136;// level 8
assign po10123 = w44138;// level 8
assign po10124 = ~w44143;// level 8
assign po10125 = w44146;// level 5
assign po10126 = w44154;// level 5
assign po10127 = w44157;// level 3
assign po10128 = w44160;// level 5
assign po10129 = w44163;// level 7
assign po10130 = w44166;// level 6
assign po10131 = w44169;// level 6
assign po10132 = ~w44174;// level 8
assign po10133 = ~w44178;// level 8
assign po10134 = ~w44181;// level 8
assign po10135 = ~w44184;// level 8
assign po10136 = ~w44187;// level 8
assign po10137 = ~w44190;// level 8
assign po10138 = ~w44194;// level 7
assign po10139 = ~w44198;// level 8
assign po10140 = ~w44201;// level 7
assign po10141 = ~w44204;// level 8
assign po10142 = w44206;// level 6
assign po10143 = ~w44209;// level 8
assign po10144 = ~w44213;// level 7
assign po10145 = ~w44216;// level 7
assign po10146 = pi10368;// level 0
assign po10147 = ~w44220;// level 8
assign po10148 = ~w44223;// level 8
assign po10149 = ~w44226;// level 8
assign po10150 = ~w44230;// level 7
assign po10151 = ~w44233;// level 7
assign po10152 = ~w44236;// level 7
assign po10153 = ~w44239;// level 7
assign po10154 = ~w44242;// level 8
assign po10155 = ~w44245;// level 8
assign po10156 = w44249;// level 5
assign po10157 = w44255;// level 7
assign po10158 = w44258;// level 7
assign po10159 = w44261;// level 7
assign po10160 = w44264;// level 7
assign po10161 = w44267;// level 7
assign po10162 = w44270;// level 7
assign po10163 = w44273;// level 7
assign po10164 = w44276;// level 7
assign po10165 = w44279;// level 7
assign po10166 = w44282;// level 7
assign po10167 = w44285;// level 7
assign po10168 = w44288;// level 7
assign po10169 = w44291;// level 7
assign po10170 = w44294;// level 7
assign po10171 = w44297;// level 7
assign po10172 = w44300;// level 7
assign po10173 = pi10360;// level 0
assign po10174 = w44303;// level 7
assign po10175 = w44306;// level 6
assign po10176 = ~w44312;// level 5
assign po10177 = w44315;// level 6
assign po10178 = w44318;// level 6
assign po10179 = w44321;// level 7
assign po10180 = w44324;// level 7
assign po10181 = w44327;// level 7
assign po10182 = w44330;// level 7
assign po10183 = w44333;// level 7
assign po10184 = w44336;// level 7
assign po10185 = w44339;// level 7
assign po10186 = w44342;// level 7
assign po10187 = w44345;// level 7
assign po10188 = w44348;// level 7
assign po10189 = w44351;// level 7
assign po10190 = w44354;// level 7
assign po10191 = w44357;// level 7
assign po10192 = w44360;// level 7
assign po10193 = w44363;// level 7
assign po10194 = w44366;// level 7
assign po10195 = w44369;// level 7
assign po10196 = w44372;// level 7
assign po10197 = w44375;// level 7
assign po10198 = w44378;// level 7
assign po10199 = w44381;// level 7
assign po10200 = w44384;// level 7
assign po10201 = w44387;// level 7
assign po10202 = w44390;// level 7
assign po10203 = w44393;// level 7
assign po10204 = w44396;// level 7
assign po10205 = w44399;// level 7
assign po10206 = w44402;// level 7
assign po10207 = w44405;// level 7
assign po10208 = w44408;// level 7
assign po10209 = w44411;// level 7
assign po10210 = w44414;// level 7
assign po10211 = w44417;// level 7
assign po10212 = w44420;// level 7
assign po10213 = w44423;// level 7
assign po10214 = w44426;// level 7
assign po10215 = w44429;// level 7
assign po10216 = w44432;// level 7
assign po10217 = w44435;// level 7
assign po10218 = w44438;// level 7
assign po10219 = w44441;// level 7
assign po10220 = w44444;// level 7
assign po10221 = w44447;// level 7
assign po10222 = w44450;// level 7
assign po10223 = w44453;// level 7
assign po10224 = w44456;// level 7
assign po10225 = w44459;// level 7
assign po10226 = w44462;// level 7
assign po10227 = w44465;// level 7
assign po10228 = w44468;// level 7
assign po10229 = w44471;// level 7
assign po10230 = w44474;// level 7
assign po10231 = w44477;// level 7
assign po10232 = w44480;// level 7
assign po10233 = w44483;// level 7
assign po10234 = w44486;// level 7
assign po10235 = w44489;// level 7
assign po10236 = w44492;// level 7
assign po10237 = w44495;// level 7
assign po10238 = w44498;// level 7
assign po10239 = w44501;// level 7
assign po10240 = w44504;// level 7
assign po10241 = w44507;// level 7
assign po10242 = w44510;// level 7
assign po10243 = w44513;// level 7
assign po10244 = w44516;// level 7
assign po10245 = w44519;// level 7
assign po10246 = w44522;// level 7
assign po10247 = w44525;// level 7
assign po10248 = w44528;// level 7
assign po10249 = w44531;// level 7
assign po10250 = w44534;// level 7
assign po10251 = w44537;// level 7
assign po10252 = w44540;// level 7
assign po10253 = w44543;// level 7
assign po10254 = w44546;// level 7
assign po10255 = w44549;// level 7
assign po10256 = w44552;// level 7
assign po10257 = w44555;// level 7
assign po10258 = w44558;// level 7
assign po10259 = w44561;// level 7
assign po10260 = w44564;// level 7
assign po10261 = w44567;// level 7
assign po10262 = w44570;// level 7
assign po10263 = w44573;// level 7
assign po10264 = w44576;// level 7
assign po10265 = w44579;// level 7
assign po10266 = w44582;// level 7
assign po10267 = w44585;// level 7
assign po10268 = w44588;// level 7
assign po10269 = w44591;// level 7
assign po10270 = w44594;// level 7
assign po10271 = w44597;// level 7
assign po10272 = w44600;// level 7
assign po10273 = w44603;// level 7
assign po10274 = w44606;// level 7
assign po10275 = w44609;// level 7
assign po10276 = w44612;// level 7
assign po10277 = w44615;// level 7
assign po10278 = w44618;// level 7
assign po10279 = w44621;// level 6
assign po10280 = w44624;// level 7
assign po10281 = w44627;// level 7
assign po10282 = w44630;// level 7
assign po10283 = w44633;// level 7
assign po10284 = w44636;// level 7
assign po10285 = w44639;// level 7
assign po10286 = w44642;// level 7
assign po10287 = w44645;// level 7
assign po10288 = w44648;// level 7
assign po10289 = w44651;// level 7
assign po10290 = w44654;// level 7
assign po10291 = w44657;// level 7
assign po10292 = w44660;// level 7
assign po10293 = w44663;// level 7
assign po10294 = w44666;// level 7
assign po10295 = w44669;// level 7
assign po10296 = w44672;// level 7
assign po10297 = w44675;// level 7
assign po10298 = w44678;// level 7
assign po10299 = w44681;// level 7
assign po10300 = w44684;// level 7
assign po10301 = w44687;// level 7
assign po10302 = w44690;// level 7
assign po10303 = w44693;// level 7
assign po10304 = w44696;// level 7
assign po10305 = w44699;// level 7
assign po10306 = w44702;// level 7
assign po10307 = w44705;// level 7
assign po10308 = w44708;// level 7
assign po10309 = w44711;// level 7
assign po10310 = w44714;// level 7
assign po10311 = w44717;// level 7
assign po10312 = w44720;// level 7
assign po10313 = w44723;// level 7
assign po10314 = w44726;// level 7
assign po10315 = w44729;// level 7
assign po10316 = w44732;// level 7
assign po10317 = w44735;// level 7
assign po10318 = w44738;// level 7
assign po10319 = w44741;// level 7
assign po10320 = w44744;// level 6
assign po10321 = w44747;// level 6
assign po10322 = w44750;// level 6
assign po10323 = w44753;// level 6
assign po10324 = w44756;// level 6
assign po10325 = w44759;// level 6
assign po10326 = w44762;// level 6
assign po10327 = w44765;// level 6
assign po10328 = w44768;// level 6
assign po10329 = w44771;// level 6
assign po10330 = w44774;// level 7
assign po10331 = w44777;// level 7
assign po10332 = w44780;// level 7
assign po10333 = w44783;// level 7
assign po10334 = w44786;// level 7
assign po10335 = w44789;// level 7
assign po10336 = w44792;// level 7
assign po10337 = w44795;// level 7
assign po10338 = w44798;// level 7
assign po10339 = w44801;// level 7
assign po10340 = w44804;// level 7
assign po10341 = w44807;// level 7
assign po10342 = w44810;// level 7
assign po10343 = w44813;// level 7
assign po10344 = w44816;// level 7
assign po10345 = w44819;// level 7
assign po10346 = w44822;// level 7
assign po10347 = w44825;// level 7
assign po10348 = w44828;// level 7
assign po10349 = w44831;// level 7
assign po10350 = w44834;// level 7
assign po10351 = w44837;// level 7
assign po10352 = w44840;// level 7
assign po10353 = w44843;// level 7
assign po10354 = w44846;// level 7
assign po10355 = w44849;// level 7
assign po10356 = w44852;// level 7
assign po10357 = w44854;// level 6
assign po10358 = ~w44857;// level 8
assign po10359 = ~w44860;// level 7
assign po10360 = ~w44863;// level 7
assign po10361 = ~w44866;// level 7
assign po10362 = ~w44869;// level 7
assign po10363 = ~w44872;// level 7
assign po10364 = ~w44875;// level 8
assign po10365 = ~w44878;// level 8
assign po10366 = ~w44881;// level 8
assign po10367 = ~w44884;// level 8
assign po10368 = ~w44887;// level 8
assign po10369 = ~w44890;// level 7
assign po10370 = ~w44893;// level 7
assign po10371 = ~w44896;// level 7
assign po10372 = ~w44899;// level 7
assign po10373 = ~w44902;// level 7
assign po10374 = ~w44905;// level 7
assign po10375 = ~w44908;// level 8
assign po10376 = ~w44911;// level 8
assign po10377 = ~w44914;// level 8
assign po10378 = ~w44917;// level 8
assign po10379 = ~w44920;// level 8
assign po10380 = ~w44923;// level 7
assign po10381 = ~w44926;// level 7
assign po10382 = ~w44929;// level 7
assign po10383 = ~w44932;// level 7
assign po10384 = ~w44935;// level 7
assign po10385 = ~w44938;// level 8
assign po10386 = ~w44941;// level 8
assign po10387 = ~w44944;// level 8
assign po10388 = w44947;// level 7
assign po10389 = w44975;// level 7
assign po10390 = ~w44978;// level 4
assign po10391 = ~w44981;// level 3
assign po10392 = pi10365;// level 0
assign po10393 = w44984;// level 7
assign po10394 = w44987;// level 7
assign po10395 = w44990;// level 7
assign po10396 = w44993;// level 7
assign po10397 = w44996;// level 7
assign po10398 = w44999;// level 7
assign po10399 = w45002;// level 7
assign po10400 = w45005;// level 7
assign po10401 = w45008;// level 7
assign po10402 = w45011;// level 7
assign po10403 = w45014;// level 7
assign po10404 = w45017;// level 7
assign po10405 = w45020;// level 7
assign po10406 = w45023;// level 7
assign po10407 = w45026;// level 7
assign po10408 = w45029;// level 7
assign po10409 = w45032;// level 7
assign po10410 = w45035;// level 7
assign po10411 = w45038;// level 7
assign po10412 = w45041;// level 7
assign po10413 = w45044;// level 7
assign po10414 = w45047;// level 7
assign po10415 = w45050;// level 7
assign po10416 = w45053;// level 7
assign po10417 = w45056;// level 7
assign po10418 = w45059;// level 7
assign po10419 = w45062;// level 7
assign po10420 = w45065;// level 7
assign po10421 = w45068;// level 7
assign po10422 = w45071;// level 7
assign po10423 = w45074;// level 7
assign po10424 = w45077;// level 7
assign po10425 = w45080;// level 7
assign po10426 = w45083;// level 7
assign po10427 = w45086;// level 7
assign po10428 = w45089;// level 7
assign po10429 = w45092;// level 7
assign po10430 = w45095;// level 7
assign po10431 = w45098;// level 7
assign po10432 = w45101;// level 7
assign po10433 = w45104;// level 7
assign po10434 = w45107;// level 7
assign po10435 = w45110;// level 7
assign po10436 = w45113;// level 7
assign po10437 = w45116;// level 7
assign po10438 = w45119;// level 7
assign po10439 = w45122;// level 7
assign po10440 = w45125;// level 7
assign po10441 = w45128;// level 7
assign po10442 = w45131;// level 7
assign po10443 = w45134;// level 7
assign po10444 = w45137;// level 7
assign po10445 = w45140;// level 7
assign po10446 = w45143;// level 7
assign po10447 = w45146;// level 7
assign po10448 = w45149;// level 7
assign po10449 = w45152;// level 7
assign po10450 = w45155;// level 7
assign po10451 = w45158;// level 7
assign po10452 = w45161;// level 7
assign po10453 = w45164;// level 7
assign po10454 = w45167;// level 7
assign po10455 = w45170;// level 7
assign po10456 = w45173;// level 7
assign po10457 = w45176;// level 7
assign po10458 = w45179;// level 7
assign po10459 = w45182;// level 7
assign po10460 = w45185;// level 7
assign po10461 = w45188;// level 7
assign po10462 = w45191;// level 7
assign po10463 = w45194;// level 7
assign po10464 = w45197;// level 7
assign po10465 = w45200;// level 7
assign po10466 = w45203;// level 7
assign po10467 = w45206;// level 7
assign po10468 = w45209;// level 7
assign po10469 = w45212;// level 7
assign po10470 = w45215;// level 7
assign po10471 = w45221;// level 4
assign po10472 = w45224;// level 7
assign po10473 = w45227;// level 6
assign po10474 = w45228;// level 1
assign po10475 = w45229;// level 1
assign po10476 = pi10375;// level 0
assign po10477 = w45230;// level 1
assign po10478 = w45233;// level 6
assign po10479 = w45236;// level 5
assign po10480 = w14215;// level 5
assign po10481 = w45240;// level 3
assign po10482 = w45242;// level 6
assign po10483 = w45245;// level 3
assign po10484 = w45250;// level 6
assign po10485 = w45251;// level 1
assign po10486 = w45252;// level 5
assign po10487 = w45255;// level 6
assign po10488 = w43916;// level 3
assign po10489 = ~w45260;// level 5
assign po10490 = ~w45265;// level 7
assign po10491 = w43664;// level 3
assign po10492 = pi10429;// level 0
assign po10493 = w44151;// level 3
assign po10494 = w45268;// level 5
assign po10495 = ~w45272;// level 6
assign po10496 = w45273;// level 6
assign po10497 = ~w45275;// level 5
assign po10498 = w44247;// level 3
assign po10499 = ~w45281;// level 7
assign po10500 = pi10399;// level 0
assign po10501 = pi10392;// level 0
assign po10502 = w45283;// level 5
assign po10503 = w45287;// level 4
assign po10504 = w45291;// level 4
assign po10505 = ~w45292;// level 4
assign po10506 = w45298;// level 6
assign po10507 = w45300;// level 4
assign po10508 = pi10464;// level 0
assign po10509 = ~w45305;// level 4
assign po10510 = w45308;// level 5
assign po10511 = w45311;// level 5
assign po10512 = w45313;// level 4
assign po10513 = ~w45315;// level 2
assign po10514 = w45318;// level 2
assign po10515 = w45320;// level 2
assign po10516 = w45323;// level 4
assign po10517 = w1576;// level 4
assign po10518 = ~w45328;// level 4
assign po10519 = w45331;// level 2
assign po10520 = w45334;// level 2
assign po10521 = w45337;// level 2
assign po10522 = ~pi10448;// level 0
assign po10523 = ~pi10461;// level 0
assign po10524 = pi10436;// level 0
assign po10525 = ~pi10455;// level 0
assign po10526 = w45340;// level 2
assign po10527 = w45343;// level 2
assign po10528 = w45346;// level 2
assign po10529 = w45349;// level 2
assign po10530 = w45352;// level 2
assign po10531 = w45355;// level 2
assign po10532 = ~pi10456;// level 0
assign po10533 = ~w45359;// level 6
assign po10534 = w45362;// level 4
assign po10535 = w45365;// level 2
assign po10536 = w45368;// level 2
assign po10537 = w45371;// level 2
assign po10538 = w45374;// level 2
assign po10539 = w45377;// level 2
assign po10540 = w45380;// level 2
assign po10541 = w45383;// level 2
assign po10542 = w45386;// level 2
assign po10543 = ~w45388;// level 3
assign po10544 = w45391;// level 2
assign po10545 = w45401;// level 5
assign po10546 = w45404;// level 2
assign po10547 = w45406;// level 3
assign po10548 = pi10463;// level 0
assign po10549 = pi10460;// level 0
assign po10550 = pi10458;// level 0
assign po10551 = pi10534;// level 0
assign po10552 = pi10459;// level 0
assign po10553 = ~w158;// level 2
assign po10554 = w45408;// level 2
assign po10555 = w45410;// level 5
assign po10556 = ~w45413;// level 2
assign po10557 = w12854;// level 3
assign po10558 = w45417;// level 3
assign po10559 = ~w45420;// level 3
assign po10560 = ~pi10500;// level 0
assign po10561 = w45425;// level 4
assign po10562 = w16783;// level 4
assign po10563 = pi10498;// level 0
assign po10564 = ~w45430;// level 5
assign po10565 = pi10533;// level 0
assign po10566 = pi10485;// level 0
assign po10567 = w45432;// level 2
assign po10568 = ~w45434;// level 3
assign po10569 = pi10502;// level 0
assign po10570 = pi10499;// level 0
assign po10571 = ~w538;// level 3
assign po10572 = pi10529;// level 0
assign po10573 = pi10509;// level 0
assign po10574 = pi10494;// level 0
assign po10575 = pi10512;// level 0
assign po10576 = pi10531;// level 0
assign po10577 = pi10497;// level 0
assign po10578 = pi10530;// level 0
assign po10579 = pi10506;// level 0
assign po10580 = pi10525;// level 0
assign po10581 = pi10508;// level 0
assign po10582 = pi10478;// level 0
assign po10583 = pi10526;// level 0
assign po10584 = pi10487;// level 0
assign po10585 = pi10484;// level 0
assign po10586 = pi10507;// level 0
assign po10587 = pi10491;// level 0
assign po10588 = ~w642;// level 2
assign po10589 = pi10513;// level 0
assign po10590 = pi10501;// level 0
assign po10591 = pi10503;// level 0
assign po10592 = pi10504;// level 0
assign po10593 = pi10532;// level 0
assign po10594 = ~w45437;// level 3
assign po10595 = pi00250;// level 0
assign po10596 = w45439;// level 4
assign po10597 = w11126;// level 1
assign po10598 = w45441;// level 2
assign po10599 = w45443;// level 2
assign po10600 = w45446;// level 2
assign po10601 = pi10479;// level 0
assign po10602 = ~pi00294;// level 0
assign po10603 = pi09966;// level 0
assign po10604 = ~w45448;// level 2
assign po10605 = w45451;// level 2
assign po10606 = ~pi00823;// level 0
assign po10607 = ~pi00052;// level 0
assign po10608 = ~pi09965;// level 0
assign po10609 = ~pi00820;// level 0
assign po10610 = pi00843;// level 0
assign po10611 = pi02665;// level 0
assign po10612 = ~pi00818;// level 0
assign po10613 = ~pi00539;// level 0
assign po10614 = pi10442;// level 0
assign po10615 = ~pi00821;// level 0
assign po10616 = pi10470;// level 0
assign po10617 = pi10441;// level 0
assign po10618 = ~pi00473;// level 0
assign po10619 = pi10468;// level 0
assign po10620 = ~pi00872;// level 0
assign po10621 = w45237;// level 1
assign po10622 = ~pi00207;// level 0
assign po10623 = pi00476;// level 0
assign po10624 = ~pi01170;// level 0
assign po10625 = ~pi10006;// level 0
assign po10626 = ~pi00311;// level 0
assign po10627 = pi10443;// level 0
assign po10628 = ~pi00822;// level 0
assign po10629 = ~pi00102;// level 0
assign po10630 = pi10446;// level 0
assign po10631 = ~pi10420;// level 0
assign po10632 = pi10469;// level 0
assign po10633 = ~pi00436;// level 0
assign po10634 = pi10466;// level 0
assign po10635 = ~pi10382;// level 0
assign po10636 = pi10587;// level 0
assign po10637 = pi10467;// level 0
assign po10638 = pi00869;// level 0
assign po10639 = ~pi00053;// level 0
assign po10640 = ~pi00819;// level 0
assign po10641 = w45454;// level 2
assign po10642 = w45457;// level 2
assign po10643 = ~w45459;// level 2
assign po10644 = w45462;// level 2
assign po10645 = pi01165;// level 0
assign po10646 = pi00842;// level 0
assign po10647 = w12874;// level 1
assign po10648 = w45440;// level 1
assign po10649 = w45463;// level 1
assign po10650 = pi10445;// level 0
assign po10651 = pi10588;// level 0
assign po10652 = pi01168;// level 0
assign po10653 = pi10390;// level 0
assign po10654 = ~w149;// level 2
assign po10655 = ~w45466;// level 2
assign po10656 = w45469;// level 2
assign po10657 = w45472;// level 2
assign po10658 = w45475;// level 2
assign po10659 = pi09839;// level 0
assign po10660 = pi09953;// level 0
assign po10661 = w45478;// level 2
assign po10662 = pi10266;// level 0
assign po10663 = ~pi00025;// level 0
assign po10664 = pi02700;// level 0
assign po10665 = pi02702;// level 0
assign po10666 = pi10553;// level 0
assign po10667 = pi10556;// level 0
assign po10668 = pi02701;// level 0
assign po10669 = pi02696;// level 0
assign po10670 = pi10547;// level 0
assign po10671 = pi02698;// level 0
assign po10672 = pi10381;// level 0
assign po10673 = pi02699;// level 0
assign po10674 = pi02697;// level 0
assign po10675 = pi00437;// level 0
assign po10676 = pi02180;// level 0
assign po10677 = w45990;// level 13
assign po10678 = ~w46502;// level 13
assign po10679 = ~w47014;// level 13
assign po10680 = w47526;// level 13
assign po10681 = ~w3883;// level 5
assign po10682 = ~w48038;// level 13
assign po10683 = w48550;// level 13
assign po10684 = ~w49062;// level 13
assign po10685 = ~w49574;// level 13
assign po10686 = ~w50086;// level 13
assign po10687 = w50598;// level 13
assign po10688 = ~w51110;// level 13
assign po10689 = ~w51622;// level 13
assign po10690 = ~w52134;// level 13
assign po10691 = ~w52646;// level 13
assign po10692 = ~w53158;// level 13
assign po10693 = ~w53670;// level 13
assign po10694 = ~w54182;// level 13
assign po10695 = ~w54694;// level 13
endmodule
