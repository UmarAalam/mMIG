//Written by the Majority Logic Package Thu Apr 30 14:58:08 2015
module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403;
wire one, v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, v16, v17, v18, v19, v20, v21, v22, v23, v24, v25, v26, v27, v28, v29, v30, v31, v32, v33, v34, v35, v36, v37, v38, v39, v40, v41, v42, v43, v44, v45, v46, v47, v48, v49, v50, v51, v52, v53, v54, v55, v56, v57, v58, v59, v60, v61, v62, v63, v64, v65, v66, v67, v68, v69, v70, v71, v72, v73, v74, v75, v76, v77, v78, v79, v80, v81, v82, v83, v84, v85, v86, v87, v88, v89, v90, v91, v92, v93, v94, v95, v96, v97, v98, v99, v100, v101, v102, v103, v104, v105, v106, v107, v108, v109, v110, v111, v112, v113, v114, v115, v116, v117, v118, v119, v120, v121, v122, v123, v124, v125, v126, v127, v128, v129, v130, v131, v132, v133, v134, v135, v136, v137, v138, v139, v140, v141, v142, v143, v144, v145, v146, v147, v148, v149, v150, v151, v152, v153, v154, v155, v156, v157, v158, v159, v160, v161, v162, v163, v164, v165, v166, v167, v168, v169, v170, v171, v172, v173, v174, v175, v176, v177, v178, v179, v180, v181, v182, v183, v184, v185, v186, v187, v188, v189, v190, v191, v192, v193, v194, v195, v196, v197, v198, v199, v200, v201, v202, v203, v204, v205, v206, v207, v208, v209, v210, v211, v212, v213, v214, v215, v216, v217, v218, v219, v220, v221, v222, v223, v224, v225, v226, v227, v228, v229, v230, v231, v232, v233, v234, v235, v236, v237, v238, v239, v240, v241, v242, v243, v244, v245, v246, v247, v248, v249, v250, v251, v252, v253, v254, v255, v256, v257, v258, v259, v260, v261, v262, v263, v264, v265, v266, v267, v268, v269, v270, v271, v272, v273, v274, v275, v276, v277, v278, v279, v280, v281, v282, v283, v284, v285, v286, v287, v288, v289, v290, v291, v292, v293, v294, v295, v296, v297, v298, v299, v300, v301, v302, v303, v304, v305, v306, v307, v308, v309, v310, v311, v312, v313, v314, v315, v316, v317, v318, v319, v320, v321, v322, v323, v324, v325, v326, v327, v328, v329, v330, v331, v332, v333, v334, v335, v336, v337, v338, v339, v340, v341, v342, v343, v344, v345, v346, v347, v348, v349, v350, v351, v352, v353, v354, v355, v356, v357, v358, v359, v360, v361, v362, v363, v364, v365, v366, v367, v368, v369, v370, v371, v372, v373, v374, v375, v376, v377, v378, v379, v380, v381, v382, v383, v384, v385, v386, v387, v388, v389, v390, v391, v392, v393, v394, v395, v396, v397, v398, v399, v400, v401, v402, v403, v404, v405, v406, v407, v408, v409, v410, v411, v412, v413, v414, v415, v416, v417, v418, v419, v420, v421, v422, v423, v424, v425, v426, v427, v428, v429, v430, v431, v432, v433, v434, v435, v436, v437, v438, v439, v440, v441, v442, v443, v444, v445, v446, v447, v448, v449, v450, v451, v452, v453, v454, v455, v456, v457, v458, v459, v460, v461, v462, v463, v464, v465, v466, v467, v468, v469, v470, v471, v472, v473, v474, v475, v476, v477, v478, v479, v480, v481, v482, v483, v484, v485, v486, v487, v488, v489, v490, v491, v492, v493, v494, v495, v496, v497, v498, v499, v500, v501, v502, v503, v504, v505, v506, v507, v508, v509, v510, v511, v512, v513, v514, v515, v516, v517, v518, v519, v520, v521, v522, v523, v524, v525, v526, v527, v528, v529, v530, v531, v532, v533, v534, v535, v536, v537, v538, v539, v540, v541, v542, v543, v544, v545, v546, v547, v548, v549, v550, v551, v552, v553, v554, v555, v556, v557, v558, v559, v560, v561, v562, v563, v564, v565, v566, v567, v568, v569, v570, v571, v572, v573, v574, v575, v576, v577, v578, v579, v580, v581, v582, v583, v584, v585, v586, v587, v588, v589, v590, v591, v592, v593, v594, v595, v596, v597, v598, v599, v600, v601, v602, v603, v604, v605, v606, v607, v608, v609, v610, v611, v612, v613, v614, v615, v616, v617, v618, v619, v620, v621, v622, v623, v624, v625, v626, v627, v628, v629, v630, v631, v632, v633, v634, v635, v636, v637, v638, v639, v640, v641, v642, v643, v644, v645, v646, v647, v648, v649, v650, v651, v652, v653, v654, v655, v656, v657, v658, v659, v660, v661, v662, v663, v664, v665, v666, v667, v668, v669, v670, v671, v672, v673, v674, v675, v676, v677, v678, v679, v680, v681, v682, v683, v684, v685, v686, v687, v688, v689, v690, v691, v692, v693, v694, v695, v696, v697, v698, v699, v700, v701, v702, v703, v704, v705, v706, v707, v708, v709, v710, v711, v712, v713, v714, v715, v716, v717, v718, v719, v720, v721, v722, v723, v724, v725, v726, v727, v728, v729, v730, v731, v732, v733, v734, v735, v736, v737, v738, v739, v740, v741, v742, v743, v744, v745, v746, v747, v748, v749, v750, v751, v752, v753, v754, v755, v756, v757, v758, v759, v760, v761, v762, v763, v764, v765, v766, v767, v768, v769, v770, v771, v772, v773, v774, v775, v776, v777, v778, v779, v780, v781, v782, v783, v784, v785, v786, v787, v788, v789, v790, v791, v792, v793, v794, v795, v796, v797, v798, v799, v800, v801, v802, v803, v804, v805, v806, v807, v808, v809, v810, v811, v812, v813, v814, v815, v816, v817, v818, v819, v820, v821, v822, v823, v824, v825, v826, v827, v828, v829, v830, v831, v832, v833, v834, v835, v836, v837, v838, v839, v840, v841, v842, v843, v844, v845, v846, v847, v848, v849, v850, v851, v852, v853, v854, v855, v856, v857, v858, v859, v860, v861, v862, v863, v864, v865, v866, v867, v868, v869, v870, v871, v872, v873, v874, v875, v876, v877, v878, v879, v880, v881, v882, v883, v884, v885, v886, v887, v888, v889, v890, v891, v892, v893, v894, v895, v896, v897, v898, v899, v900, v901, v902, v903, v904, v905, v906, v907, v908, v909, v910, v911, v912, v913, v914, v915, v916, v917, v918, v919, v920, v921, v922, v923, v924, v925, v926, v927, v928, v929, v930, v931, v932, v933, v934, v935, v936, v937, v938, v939, v940, v941, v942, v943, v944, v945, v946, v947, v948, v949, v950, v951, v952, v953, v954, v955, v956, v957, v958, v959, v960, v961, v962, v963, v964, v965, v966, v967, v968, v969, v970, v971, v972, v973, v974, v975, v976, v977, v978, v979, v980, v981, v982, v983, v984, v985, v986, v987, v988, v989, v990, v991, v992, v993, v994, v995, v996, v997, v998, v999, v1000, v1001, v1002, v1003, v1004, v1005, v1006, v1007, v1008, v1009, v1010, v1011, v1012, v1013, v1014, v1015, v1016, v1017, v1018, v1019, v1020, v1021, v1022, v1023, v1024, v1025, v1026, v1027, v1028, v1029, v1030, v1031, v1032, v1033, v1034, v1035, v1036, v1037, v1038, v1039, v1040, v1041, v1042, v1043, v1044, v1045, v1046, v1047, v1048, v1049, v1050, v1051, v1052, v1053, v1054, v1055, v1056, v1057, v1058, v1059, v1060, v1061, v1062, v1063, v1064, v1065, v1066, v1067, v1068, v1069, v1070, v1071, v1072, v1073, v1074, v1075, v1076, v1077, v1078, v1079, v1080, v1081, v1082, v1083, v1084, v1085, v1086, v1087, v1088, v1089, v1090, v1091, v1092, v1093, v1094, v1095, v1096, v1097, v1098, v1099, v1100, v1101, v1102, v1103, v1104, v1105, v1106, v1107, v1108, v1109, v1110, v1111, v1112, v1113, v1114, v1115, v1116, v1117, v1118, v1119, v1120, v1121, v1122, v1123, v1124, v1125, v1126, v1127, v1128, v1129, v1130, v1131, v1132, v1133, v1134, v1135, v1136, v1137, v1138, v1139, v1140, v1141, v1142, v1143, v1144, v1145, v1146, v1147, v1148, v1149, v1150, v1151, v1152, v1153, v1154, v1155, v1156, v1157, v1158, v1159, v1160, v1161, v1162, v1163, v1164, v1165, v1166, v1167, v1168, v1169, v1170, v1171, v1172, v1173, v1174, v1175, v1176, v1177, v1178, v1179, v1180, v1181, v1182, v1183, v1184, v1185, v1186, v1187, v1188, v1189, v1190, v1191, v1192, v1193, v1194, v1195, v1196, v1197, v1198, v1199, v1200, v1201, v1202, v1203, v1204, v1205, v1206, v1207, v1208, v1209, v1210, v1211, v1212, v1213, v1214, v1215, v1216, v1217, v1218, v1219, v1220, v1221, v1222, v1223, v1224, v1225, v1226, v1227, v1228, v1229, v1230, v1231, v1232, v1233, v1234, v1235, v1236, v1237, v1238, v1239, v1240, v1241, v1242, v1243, v1244, v1245, v1246, v1247, v1248, v1249, v1250, v1251, v1252, v1253, v1254, v1255, v1256, v1257, v1258, v1259, v1260, v1261, v1262, v1263, v1264, v1265, v1266, v1267, v1268, v1269, v1270, v1271, v1272, v1273, v1274, v1275, v1276, v1277, v1278, v1279, v1280, v1281, v1282, v1283, v1284, v1285, v1286, v1287, v1288, v1289, v1290, v1291, v1292, v1293, v1294, v1295, v1296, v1297, v1298, v1299, v1300, v1301, v1302, v1303, v1304, v1305, v1306, v1307, v1308, v1309, v1310, v1311, v1312, v1313, v1314, v1315, v1316, v1317, v1318, v1319, v1320, v1321, v1322, v1323, v1324, v1325, v1326, v1327, v1328, v1329, v1330, v1331, v1332, v1333, v1334, v1335, v1336, v1337, v1338, v1339, v1340, v1341, v1342, v1343, v1344, v1345, v1346, v1347, v1348, v1349, v1350, v1351, v1352, v1353, v1354, v1355, v1356, v1357, v1358, v1359, v1360, v1361, v1362, v1363, v1364, v1365, v1366, v1367, v1368, v1369, v1370, v1371, v1372, v1373, v1374, v1375, v1376, v1377, v1378, v1379, v1380, v1381, v1382, v1383, v1384, v1385, v1386, v1387, v1388, v1389, v1390, v1391, v1392, v1393, v1394, v1395, v1396, v1397, v1398, v1399, v1400, v1401, v1402, v1403, v1404, v1405, v1406, v1407, v1408, v1409, v1410, v1411, v1412, v1413, v1414, v1415, v1416, v1417, v1418, v1419, v1420, v1421, v1422, v1423, v1424, v1425, v1426, v1427, v1428, v1429, v1430, v1431, v1432, v1433, v1434, v1435, v1436, v1437, v1438, v1439, v1440, v1441, v1442, v1443, v1444, v1445, v1446, v1447, v1448, v1449, v1450, v1451, v1452, v1453, v1454, v1455, v1456, v1457, v1458, v1459, v1460, v1461, v1462, v1463, v1464, v1465, v1466, v1467, v1468, v1469, v1470, v1471, v1472, v1473, v1474, v1475, v1476, v1477, v1478, v1479, v1480, v1481, v1482, v1483, v1484, v1485, v1486, v1487, v1488, v1489, v1490, v1491, v1492, v1493, v1494, v1495, v1496, v1497, v1498, v1499, v1500, v1501, v1502, v1503, v1504, v1505, v1506, v1507, v1508, v1509, v1510, v1511, v1512, v1513, v1514, v1515, v1516, v1517, v1518, v1519, v1520, v1521, v1522, v1523, v1524, v1525, v1526, v1527, v1528, v1529, v1530, v1531, v1532, v1533, v1534, v1535, v1536, v1537, v1538, v1539, v1540, v1541, v1542, v1543, v1544, v1545, v1546, v1547, v1548, v1549, v1550, v1551, v1552, v1553, v1554, v1555, v1556, v1557, v1558, v1559, v1560, v1561, v1562, v1563, v1564, v1565, v1566, v1567, v1568, v1569, v1570, v1571, v1572, v1573, v1574, v1575, v1576, v1577, v1578, v1579, v1580, v1581, v1582, v1583, v1584, v1585, v1586, v1587, v1588, v1589, v1590, v1591, v1592, v1593, v1594, v1595, v1596, v1597, v1598, v1599, v1600, v1601, v1602, v1603, v1604, v1605, v1606, v1607, v1608, v1609, v1610, v1611, v1612, v1613, v1614, v1615, v1616, v1617, v1618, v1619, v1620, v1621, v1622, v1623, v1624, v1625, v1626, v1627, v1628, v1629, v1630, v1631, v1632, v1633, v1634, v1635, v1636, v1637, v1638, v1639, v1640, v1641, v1642, v1643, v1644, v1645, v1646, v1647, v1648, v1649, v1650, v1651, v1652, v1653, v1654, v1655, v1656, v1657, v1658, v1659, v1660, v1661, v1662, v1663, v1664, v1665, v1666, v1667, v1668, v1669, v1670, v1671, v1672, v1673, v1674, v1675, v1676, v1677, v1678, v1679, v1680, v1681, v1682, v1683, v1684, v1685, v1686, v1687, v1688, v1689, v1690, v1691, v1692, v1693, v1694, v1695, v1696, v1697, v1698, v1699, v1700, v1701, v1702, v1703, v1704, v1705, v1706, v1707, v1708, v1709, v1710, v1711, v1712, v1713, v1714, v1715, v1716, v1717, v1718, v1719, v1720, v1721, v1722, v1723, v1724, v1725, v1726, v1727, v1728, v1729, v1730, v1731, v1732, v1733, v1734, v1735, v1736, v1737, v1738, v1739, v1740, v1741, v1742, v1743, v1744, v1745, v1746, v1747, v1748, v1749, v1750, v1751, v1752, v1753, v1754, v1755, v1756, v1757, v1758, v1759, v1760, v1761, v1762, v1763, v1764, v1765, v1766, v1767, v1768, v1769, v1770, v1771, v1772, v1773, v1774, v1775, v1776, v1777, v1778, v1779, v1780, v1781, v1782, v1783, v1784, v1785, v1786, v1787, v1788, v1789, v1790, v1791, v1792, v1793, v1794, v1795, v1796, v1797, v1798, v1799, v1800, v1801, v1802, v1803, v1804, v1805, v1806, v1807, v1808, v1809, v1810, v1811, v1812, v1813, v1814, v1815, v1816, v1817, v1818, v1819, v1820, v1821, v1822, v1823, v1824, v1825, v1826, v1827, v1828, v1829, v1830, v1831, v1832, v1833, v1834, v1835, v1836, v1837, v1838, v1839, v1840, v1841, v1842, v1843, v1844, v1845, v1846, v1847, v1848, v1849, v1850, v1851, v1852, v1853, v1854, v1855, v1856, v1857, v1858, v1859, v1860, v1861, v1862, v1863, v1864, v1865, v1866, v1867, v1868, v1869, v1870, v1871, v1872, v1873, v1874, v1875, v1876, v1877, v1878, v1879, v1880, v1881, v1882, v1883, v1884, v1885, v1886, v1887, v1888, v1889, v1890, v1891, v1892, v1893, v1894, v1895, v1896, v1897, v1898, v1899, v1900, v1901, v1902, v1903, v1904, v1905, v1906, v1907, v1908, v1909, v1910, v1911, v1912, v1913, v1914, v1915, v1916, v1917, v1918, v1919, v1920, v1921, v1922, v1923, v1924, v1925, v1926, v1927, v1928, v1929, v1930, v1931, v1932, v1933, v1934, v1935, v1936, v1937, v1938, v1939, v1940, v1941, v1942, v1943, v1944, v1945, v1946, v1947, v1948, v1949, v1950, v1951, v1952, v1953, v1954, v1955, v1956, v1957, v1958, v1959, v1960, v1961, v1962, v1963, v1964, v1965, v1966, v1967, v1968, v1969, v1970, v1971, v1972, v1973, v1974, v1975, v1976, v1977, v1978, v1979, v1980, v1981, v1982, v1983, v1984,
w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396;
assign v0 = ~(pi294 | pi301);
assign w0 = v0;
assign v1 = ~(pi188 | pi190);
assign w1 = v1;
assign w2 = pi189 & w1;
assign w3 = pi291 & ~pi297;
assign w4 = pi299 & w3;
assign w5 = w3 & w47;
assign w6 = ~pi296 & w5;
assign w7 = w2 & w6;
assign w8 = pi188 & ~pi189;
assign w9 = pi190 & w8;
assign w10 = w6 & w9;
assign v2 = ~(pi302 | pi303);
assign w11 = v2;
assign v3 = ~(pi131 | pi298);
assign w12 = v3;
assign w13 = ~pi102 & pi298;
assign v4 = ~(w12 | w13);
assign w14 = v4;
assign w15 = w11 & ~w14;
assign w16 = ~pi298 & pi302;
assign w17 = pi132 & pi303;
assign w18 = w16 & w17;
assign w19 = pi302 & ~pi303;
assign v5 = ~(pi132 | pi298);
assign w20 = v5;
assign w21 = w19 & w20;
assign w22 = ~pi302 & pi303;
assign w23 = w14 & w22;
assign w24 = pi298 & pi302;
assign w25 = pi178 & ~pi303;
assign w26 = ~pi178 & pi303;
assign w27 = w24 & ~w25;
assign w28 = ~w26 & w27;
assign v6 = ~(w18 | w21);
assign w29 = v6;
assign w30 = ~w15 & w29;
assign v7 = ~(w23 | w28);
assign w31 = v7;
assign w32 = w30 & w31;
assign w33 = w10 & ~w32;
assign w34 = (~w7 & w32) | (~w7 & w6125) | (w32 & w6125);
assign w35 = pi188 & pi190;
assign v8 = ~(pi189 | w35);
assign w36 = v8;
assign w37 = ~w1 & w36;
assign v9 = ~(pi195 | pi196);
assign w38 = v9;
assign v10 = ~(pi291 | pi303);
assign w39 = v10;
assign v11 = ~(pi298 | pi299);
assign w40 = v11;
assign w41 = w39 & w40;
assign v12 = ~(pi296 | pi300);
assign w42 = v12;
assign v13 = ~(pi297 | pi302);
assign w43 = v13;
assign w44 = w42 & w43;
assign w45 = w41 & w44;
assign w46 = ~w38 & w45;
assign w47 = pi299 & pi300;
assign w48 = pi291 & pi297;
assign w49 = w47 & w48;
assign w50 = pi296 & w49;
assign v14 = ~(w46 | w50);
assign w51 = v14;
assign w52 = (w37 & w46) | (w37 & w6126) | (w46 & w6126);
assign v15 = ~(w2 | w9);
assign w53 = v15;
assign w54 = pi296 & pi300;
assign w55 = w43 & w54;
assign w56 = ~pi298 & pi299;
assign w57 = pi291 & pi303;
assign w58 = w56 & w57;
assign w59 = w55 & w58;
assign w60 = ~w53 & w59;
assign w61 = ~pi303 & w54;
assign w62 = w4 & w61;
assign w63 = w37 & w62;
assign v16 = ~(w60 | w63);
assign w64 = v16;
assign w65 = pi297 & ~pi302;
assign w66 = w54 & w65;
assign w67 = pi298 & pi299;
assign w68 = w39 & w67;
assign w69 = w66 & w68;
assign w70 = ~pi188 & pi189;
assign w71 = pi190 & w70;
assign w72 = w69 & w71;
assign w73 = ~pi291 & pi297;
assign w74 = pi296 & ~pi300;
assign w75 = ~pi299 & w74;
assign w76 = w73 & w75;
assign w77 = w75 & w6127;
assign v17 = ~(w72 | w77);
assign w78 = v17;
assign w79 = w64 & w78;
assign w80 = ~w52 & w79;
assign w81 = (w0 & ~w80) | (w0 & w6128) | (~w80 & w6128);
assign w82 = w36 & w6239;
assign w83 = ~pi291 & pi298;
assign w84 = ~pi299 & pi300;
assign w85 = w83 & w84;
assign w86 = ~pi297 & w85;
assign w87 = w37 & w86;
assign w88 = pi299 & ~pi300;
assign v18 = ~(w85 | w88);
assign w89 = v18;
assign w90 = w85 & w1185;
assign v19 = ~(w89 | w90);
assign w91 = v19;
assign w92 = w9 & ~w88;
assign w93 = w91 & w92;
assign v20 = ~(w87 | w93);
assign w94 = v20;
assign w95 = (pi301 & w82) | (pi301 & w6240) | (w82 & w6240);
assign w96 = ~w94 & w95;
assign v21 = ~(w81 | w96);
assign w97 = v21;
assign w98 = w4 & w74;
assign w99 = pi301 & w8;
assign w100 = w98 & w99;
assign w101 = ~pi190 & w8;
assign w102 = w86 & w101;
assign w103 = pi297 & w85;
assign w104 = w9 & w103;
assign v22 = ~(w102 | w104);
assign w105 = v22;
assign w106 = (~w100 & w105) | (~w100 & w6129) | (w105 & w6129);
assign w107 = (w105 & w6137) | (w105 & w6138) | (w6137 & w6138);
assign v23 = ~(pi291 | pi297);
assign w108 = v23;
assign w109 = pi299 & w108;
assign w110 = w61 & w109;
assign w111 = w8 & w110;
assign v24 = ~(w9 | w71);
assign w112 = v24;
assign w113 = w69 & ~w112;
assign v25 = ~(w111 | w113);
assign w114 = v25;
assign w115 = ~w52 & w114;
assign w116 = w34 & w115;
assign w117 = ~pi291 & pi303;
assign w118 = w56 & w117;
assign w119 = w55 & w118;
assign v26 = ~(pi296 | pi297);
assign w120 = v26;
assign w121 = w47 & w120;
assign w122 = ~pi291 & w121;
assign v27 = ~(w119 | w122);
assign w123 = v27;
assign w124 = w8 & ~w123;
assign w125 = w64 & ~w124;
assign w126 = w75 & w6241;
assign w127 = w125 & ~w126;
assign w128 = w106 & w127;
assign w129 = (~w107 & ~w128) | (~w107 & w6130) | (~w128 & w6130);
assign w130 = w8 & w6139;
assign w131 = w85 & w130;
assign w132 = w130 & w6131;
assign v28 = ~(w100 | w132);
assign w133 = v28;
assign w134 = ~w0 & w133;
assign w135 = w75 & w6242;
assign w136 = w125 & w6132;
assign w137 = w116 & w136;
assign v29 = ~(w134 | w137);
assign w138 = v29;
assign w139 = w129 & ~w138;
assign w140 = ~pi097 & pi098;
assign w141 = ~pi099 & w140;
assign w142 = pi301 & w87;
assign w143 = w134 & ~w142;
assign w144 = (~w76 & ~w87) | (~w76 & w6243) | (~w87 & w6243);
assign w145 = w125 & w6244;
assign w146 = pi097 & pi098;
assign w147 = ~pi099 & w146;
assign w148 = w82 & w147;
assign w149 = (~w141 & ~w82) | (~w141 & w6245) | (~w82 & w6245);
assign w150 = ~w143 & w7363;
assign w151 = (~w6133 & w6247) | (~w6133 & w6248) | (w6247 & w6248);
assign w152 = w139 & ~w151;
assign v30 = ~(pi313 | pi314);
assign w153 = v30;
assign w154 = w141 & w153;
assign w155 = w82 & w6249;
assign w156 = (~w6133 & w6250) | (~w6133 & w6251) | (w6250 & w6251);
assign w157 = pi298 & ~pi302;
assign w158 = w47 & w157;
assign w159 = pi303 & w0;
assign w160 = w0 & w6252;
assign w161 = w73 & w160;
assign w162 = w161 & w6253;
assign v31 = ~(pi097 | pi098);
assign w163 = v31;
assign w164 = pi099 & w163;
assign w165 = w161 & w6254;
assign v32 = ~(w162 | w165);
assign w166 = v32;
assign w167 = ~pi311 & w166;
assign v33 = ~(pi304 | w166);
assign w168 = v33;
assign v34 = ~(w167 | w168);
assign w169 = v34;
assign w170 = w156 & w169;
assign w171 = ~w152 & w170;
assign w172 = w139 & w6255;
assign w173 = pi304 & ~w156;
assign v35 = ~(w172 | w173);
assign w174 = v35;
assign w175 = ~w171 & w174;
assign v36 = ~(w129 | w156);
assign w176 = v36;
assign w177 = pi309 & ~w165;
assign v37 = ~(w162 | w177);
assign w178 = v37;
assign w179 = (~w6133 & w6256) | (~w6133 & w6257) | (w6256 & w6257);
assign w180 = (w179 & ~w139) | (w179 & w6258) | (~w139 & w6258);
assign v38 = ~(w176 | w180);
assign w181 = v38;
assign v39 = ~(w138 | w156);
assign w182 = v39;
assign v40 = ~(pi312 | w165);
assign w183 = v40;
assign v41 = ~(w162 | w183);
assign w184 = v41;
assign w185 = (~w6133 & w6259) | (~w6133 & w6260) | (w6259 & w6260);
assign w186 = (w185 & ~w139) | (w185 & w6261) | (~w139 & w6261);
assign v42 = ~(w182 | w186);
assign w187 = v42;
assign w188 = ~w181 & w187;
assign w189 = ~w175 & w188;
assign w190 = ~pi010 & w189;
assign v43 = ~(w181 | w187);
assign w191 = v43;
assign w192 = ~w175 & w191;
assign w193 = ~pi009 & w192;
assign w194 = w181 & w187;
assign w195 = w175 & w194;
assign w196 = ~pi008 & w195;
assign w197 = w175 & w188;
assign w198 = ~pi006 & w197;
assign w199 = ~w175 & w194;
assign w200 = ~pi012 & w199;
assign w201 = w181 & ~w187;
assign w202 = ~w175 & w201;
assign w203 = ~pi011 & w202;
assign w204 = w175 & w201;
assign w205 = ~pi007 & w204;
assign w206 = w175 & w191;
assign w207 = ~pi005 & w206;
assign v44 = ~(w190 | w193);
assign w208 = v44;
assign v45 = ~(w196 | w198);
assign w209 = v45;
assign v46 = ~(w200 | w203);
assign w210 = v46;
assign v47 = ~(w205 | w207);
assign w211 = v47;
assign w212 = w210 & w211;
assign w213 = w208 & w209;
assign w214 = w212 & w213;
assign v48 = ~(w97 | w214);
assign w215 = v48;
assign w216 = w97 & w214;
assign v49 = ~(w215 | w216);
assign w217 = v49;
assign w218 = (pi116 & ~w174) | (pi116 & w6142) | (~w174 & w6142);
assign w219 = w188 & w218;
assign w220 = (pi115 & ~w174) | (pi115 & w6143) | (~w174 & w6143);
assign w221 = w194 & w220;
assign w222 = (~pi100 & ~w174) | (~pi100 & w6144) | (~w174 & w6144);
assign w223 = w174 & w6177;
assign w224 = w191 & ~w222;
assign w225 = ~w223 & w224;
assign w226 = w175 & w187;
assign w227 = (~pi111 & w180) | (~pi111 & w6223) | (w180 & w6223);
assign w228 = ~w180 & w6224;
assign w229 = w226 & w6145;
assign w230 = (~pi114 & ~w174) | (~pi114 & w6178) | (~w174 & w6178);
assign w231 = w174 & w6225;
assign w232 = w201 & ~w230;
assign w233 = ~w231 & w232;
assign v50 = ~(w219 | w221);
assign w234 = v50;
assign w235 = ~w225 & w234;
assign v51 = ~(w229 | w233);
assign w236 = v51;
assign w237 = w235 & w236;
assign v52 = ~(w97 | w237);
assign w238 = v52;
assign w239 = (pi109 & ~w174) | (pi109 & w6146) | (~w174 & w6146);
assign w240 = w194 & w239;
assign w241 = (pi107 & ~w174) | (pi107 & w6147) | (~w174 & w6147);
assign w242 = w188 & w241;
assign w243 = (~pi106 & ~w174) | (~pi106 & w6148) | (~w174 & w6148);
assign w244 = w174 & w6179;
assign w245 = w191 & ~w243;
assign w246 = ~w244 & w245;
assign w247 = (~pi108 & ~w174) | (~pi108 & w6149) | (~w174 & w6149);
assign w248 = w174 & w6180;
assign w249 = w201 & ~w247;
assign w250 = ~w248 & w249;
assign w251 = (~pi103 & w180) | (~pi103 & w6181) | (w180 & w6181);
assign w252 = ~w180 & w6182;
assign w253 = w226 & w6150;
assign v53 = ~(w240 | w242);
assign w254 = v53;
assign w255 = ~w246 & w254;
assign v54 = ~(w250 | w253);
assign w256 = v54;
assign w257 = w255 & w256;
assign v55 = ~(w97 | w257);
assign w258 = v55;
assign v56 = ~(w238 | w258);
assign w259 = v56;
assign w260 = (pi151 & ~w174) | (pi151 & w6151) | (~w174 & w6151);
assign w261 = w188 & w260;
assign w262 = (pi153 & ~w174) | (pi153 & w6152) | (~w174 & w6152);
assign w263 = w194 & w262;
assign w264 = (~pi148 & w180) | (~pi148 & w6183) | (w180 & w6183);
assign w265 = ~w180 & w6184;
assign w266 = w226 & w6153;
assign w267 = (~pi175 & ~w174) | (~pi175 & w6185) | (~w174 & w6185);
assign w268 = ~pi147 & w175;
assign w269 = w191 & ~w267;
assign w270 = ~w268 & w269;
assign w271 = (~pi152 & ~w174) | (~pi152 & w6154) | (~w174 & w6154);
assign w272 = ~pi149 & w175;
assign w273 = w201 & ~w271;
assign w274 = ~w272 & w273;
assign v57 = ~(w261 | w263);
assign w275 = v57;
assign w276 = ~w266 & w275;
assign v58 = ~(w270 | w274);
assign w277 = v58;
assign w278 = w276 & w277;
assign v59 = ~(w97 | w278);
assign w279 = v59;
assign w280 = (pi124 & ~w174) | (pi124 & w6155) | (~w174 & w6155);
assign w281 = w194 & w280;
assign w282 = (pi118 & ~w174) | (pi118 & w6156) | (~w174 & w6156);
assign w283 = w188 & w282;
assign w284 = (~pi123 & ~w174) | (~pi123 & w6157) | (~w174 & w6157);
assign w285 = w174 & w6186;
assign w286 = w191 & ~w284;
assign w287 = ~w285 & w286;
assign w288 = (~pi119 & ~w174) | (~pi119 & w6158) | (~w174 & w6158);
assign w289 = w174 & w6187;
assign w290 = w201 & ~w288;
assign w291 = ~w289 & w290;
assign w292 = (~pi121 & w180) | (~pi121 & w6188) | (w180 & w6188);
assign w293 = ~w180 & w6189;
assign w294 = w226 & w6159;
assign v60 = ~(w281 | w283);
assign w295 = v60;
assign w296 = ~w287 & w295;
assign v61 = ~(w291 | w294);
assign w297 = v61;
assign w298 = w296 & w297;
assign v62 = ~(w97 | w298);
assign w299 = v62;
assign v63 = ~(w279 | w299);
assign w300 = v63;
assign w301 = (pi158 & ~w174) | (pi158 & w6160) | (~w174 & w6160);
assign w302 = w188 & w301;
assign w303 = (pi160 & ~w174) | (pi160 & w6161) | (~w174 & w6161);
assign w304 = w194 & w303;
assign w305 = (~pi159 & ~w174) | (~pi159 & w6162) | (~w174 & w6162);
assign w306 = w174 & w6190;
assign w307 = w201 & ~w305;
assign w308 = ~w306 & w307;
assign w309 = (~pi155 & w180) | (~pi155 & w6262) | (w180 & w6262);
assign w310 = ~w180 & w6263;
assign w311 = w226 & w6163;
assign w312 = (~pi127 & ~w174) | (~pi127 & w6191) | (~w174 & w6191);
assign w313 = ~pi154 & w175;
assign w314 = w191 & ~w312;
assign w315 = ~w313 & w314;
assign v64 = ~(w302 | w304);
assign w316 = v64;
assign w317 = ~w308 & w316;
assign v65 = ~(w311 | w315);
assign w318 = v65;
assign w319 = w317 & w318;
assign v66 = ~(w97 | w319);
assign w320 = v66;
assign w321 = w318 & w6164;
assign w322 = pi171 & w199;
assign w323 = pi166 & w197;
assign w324 = pi165 & w206;
assign w325 = pi167 & w204;
assign w326 = pi170 & w189;
assign w327 = pi169 & w192;
assign w328 = pi168 & w195;
assign w329 = pi176 & w202;
assign v67 = ~(w322 | w323);
assign w330 = v67;
assign v68 = ~(w324 | w325);
assign w331 = v68;
assign v69 = ~(w326 | w327);
assign w332 = v69;
assign v70 = ~(w328 | w329);
assign w333 = v70;
assign w334 = w332 & w333;
assign w335 = w330 & w331;
assign w336 = w334 & w335;
assign v71 = ~(w321 | w336);
assign w337 = v71;
assign v72 = ~(w320 | w337);
assign w338 = v72;
assign w339 = w236 & w6165;
assign w340 = w97 & w298;
assign v73 = ~(w339 | w340);
assign w341 = v73;
assign w342 = w277 & w6166;
assign w343 = w97 & w257;
assign v74 = ~(w342 | w343);
assign w344 = v74;
assign w345 = w341 & w344;
assign w346 = ~w338 & w345;
assign w347 = w300 & ~w346;
assign w348 = pi068 & w204;
assign w349 = pi069 & w189;
assign w350 = pi066 & w206;
assign w351 = (~pi067 & w180) | (~pi067 & w6193) | (w180 & w6193);
assign w352 = ~w180 & w6194;
assign w353 = w226 & w6167;
assign w354 = pi073 & w192;
assign w355 = pi070 & w202;
assign w356 = pi071 & w199;
assign v75 = ~(w348 | w349);
assign w357 = v75;
assign v76 = ~(w350 | w353);
assign w358 = v76;
assign v77 = ~(w354 | w355);
assign w359 = v77;
assign w360 = ~w356 & w359;
assign w361 = w357 & w358;
assign w362 = w360 & w361;
assign w363 = w97 & w362;
assign w364 = pi089 & w202;
assign w365 = pi082 & w199;
assign w366 = pi085 & w204;
assign w367 = (~pi084 & w180) | (~pi084 & w6195) | (w180 & w6195);
assign w368 = ~w180 & w6196;
assign w369 = w226 & w6168;
assign w370 = pi088 & w189;
assign w371 = pi083 & w206;
assign w372 = pi087 & w192;
assign v78 = ~(w364 | w365);
assign w373 = v78;
assign v79 = ~(w366 | w369);
assign w374 = v79;
assign v80 = ~(w370 | w371);
assign w375 = v80;
assign w376 = ~w372 & w375;
assign w377 = w373 & w374;
assign w378 = w376 & w377;
assign w379 = w97 & w378;
assign v81 = ~(w363 | w379);
assign w380 = v81;
assign w381 = pi077 & w195;
assign w382 = pi074 & w206;
assign w383 = pi080 & w199;
assign w384 = pi079 & w202;
assign w385 = pi075 & w197;
assign w386 = pi078 & w192;
assign w387 = pi076 & w204;
assign w388 = pi065 & w189;
assign v82 = ~(w381 | w382);
assign w389 = v82;
assign v83 = ~(w383 | w384);
assign w390 = v83;
assign v84 = ~(w385 | w386);
assign w391 = v84;
assign v85 = ~(w387 | w388);
assign w392 = v85;
assign w393 = w391 & w392;
assign w394 = w389 & w390;
assign w395 = w393 & w394;
assign w396 = w97 & w395;
assign w397 = pi096 & w199;
assign w398 = pi090 & w206;
assign w399 = pi081 & w192;
assign w400 = pi094 & w189;
assign w401 = pi092 & w204;
assign w402 = pi091 & w197;
assign w403 = pi095 & w202;
assign w404 = pi093 & w195;
assign v86 = ~(w397 | w398);
assign w405 = v86;
assign v87 = ~(w399 | w400);
assign w406 = v87;
assign v88 = ~(w401 | w402);
assign w407 = v88;
assign v89 = ~(w403 | w404);
assign w408 = v89;
assign w409 = w407 & w408;
assign w410 = w405 & w406;
assign w411 = w409 & w410;
assign w412 = w97 & w411;
assign v90 = ~(w396 | w412);
assign w413 = v90;
assign w414 = w380 & w413;
assign w415 = (w414 & w346) | (w414 & w6264) | (w346 & w6264);
assign w416 = ~pi056 & w202;
assign w417 = ~pi049 & w206;
assign w418 = ~pi050 & w197;
assign w419 = ~pi055 & w189;
assign w420 = ~pi054 & w199;
assign w421 = ~pi051 & w204;
assign w422 = ~pi052 & w195;
assign w423 = ~pi053 & w192;
assign v91 = ~(w416 | w417);
assign w424 = v91;
assign v92 = ~(w418 | w419);
assign w425 = v92;
assign v93 = ~(w420 | w421);
assign w426 = v93;
assign v94 = ~(w422 | w423);
assign w427 = v94;
assign w428 = w426 & w427;
assign w429 = w424 & w425;
assign w430 = w428 & w429;
assign w431 = w97 & w430;
assign w432 = pi026 & w189;
assign w433 = pi023 & w204;
assign w434 = pi021 & w206;
assign w435 = pi022 & w197;
assign w436 = pi024 & w195;
assign w437 = pi025 & w192;
assign w438 = pi028 & w199;
assign w439 = pi027 & w202;
assign v95 = ~(w432 | w433);
assign w440 = v95;
assign v96 = ~(w434 | w435);
assign w441 = v96;
assign v97 = ~(w436 | w437);
assign w442 = v97;
assign v98 = ~(w438 | w439);
assign w443 = v98;
assign w444 = w442 & w443;
assign w445 = w440 & w441;
assign w446 = w444 & w445;
assign w447 = w97 & w446;
assign v99 = ~(w396 | w447);
assign w448 = v99;
assign w449 = ~pi058 & w197;
assign w450 = ~pi060 & w195;
assign w451 = ~pi057 & w206;
assign w452 = ~pi061 & w192;
assign w453 = ~pi063 & w202;
assign w454 = ~pi064 & w199;
assign w455 = ~pi062 & w189;
assign w456 = ~pi059 & w204;
assign v100 = ~(w449 | w450);
assign w457 = v100;
assign v101 = ~(w451 | w452);
assign w458 = v101;
assign v102 = ~(w453 | w454);
assign w459 = v102;
assign v103 = ~(w455 | w456);
assign w460 = v103;
assign w461 = w459 & w460;
assign w462 = w457 & w458;
assign w463 = w461 & w462;
assign w464 = w97 & w463;
assign w465 = ~pi014 & w197;
assign w466 = ~pi019 & w202;
assign w467 = ~pi018 & w189;
assign w468 = ~pi016 & w195;
assign w469 = ~pi017 & w192;
assign w470 = ~pi015 & w204;
assign w471 = ~pi013 & w206;
assign w472 = ~pi020 & w199;
assign v104 = ~(w465 | w466);
assign w473 = v104;
assign v105 = ~(w467 | w468);
assign w474 = v105;
assign v106 = ~(w469 | w470);
assign w475 = v106;
assign v107 = ~(w471 | w472);
assign w476 = v107;
assign w477 = w475 & w476;
assign w478 = w473 & w474;
assign w479 = w477 & w478;
assign w480 = w97 & w479;
assign v108 = ~(w464 | w480);
assign w481 = v108;
assign w482 = w448 & w481;
assign w483 = ~w431 & w482;
assign w484 = w415 & w483;
assign v109 = ~(w97 | w479);
assign w485 = v109;
assign v110 = ~(w97 | w463);
assign w486 = v110;
assign v111 = ~(w97 | w446);
assign w487 = v111;
assign v112 = ~(w97 | w395);
assign w488 = v112;
assign v113 = ~(w487 | w488);
assign w489 = v113;
assign w490 = ~w486 & w489;
assign w491 = w489 & w6226;
assign v114 = ~(w97 | w362);
assign w492 = v114;
assign v115 = ~(w97 | w378);
assign w493 = v115;
assign v116 = ~(w97 | w411);
assign w494 = v116;
assign v117 = ~(w493 | w494);
assign w495 = v117;
assign w496 = ~w492 & w495;
assign v118 = ~(w97 | w430);
assign w497 = v118;
assign w498 = w495 & w6265;
assign w499 = w491 & w498;
assign w500 = ~w484 & w6227;
assign w501 = (w217 & w484) | (w217 & w6228) | (w484 & w6228);
assign v119 = ~(w500 | w501);
assign w502 = v119;
assign v120 = ~(w480 | w485);
assign w503 = v120;
assign v121 = ~(w447 | w464);
assign w504 = v121;
assign w505 = w414 & w504;
assign w506 = ~w347 & w505;
assign w507 = w259 & ~w492;
assign w508 = w495 & w507;
assign w509 = w490 & w508;
assign w510 = ~w506 & w6197;
assign w511 = (w503 & w506) | (w503 & w6198) | (w506 & w6198);
assign v122 = ~(w510 | w511);
assign w512 = v122;
assign v123 = ~(w363 | w492);
assign w513 = v123;
assign w514 = ~w346 & w6229;
assign w515 = (w513 & w346) | (w513 & w6230) | (w346 & w6230);
assign v124 = ~(w514 | w515);
assign w516 = v124;
assign v125 = ~(w279 | w320);
assign w517 = v125;
assign w518 = w337 & ~w342;
assign w519 = w517 & ~w518;
assign v126 = ~(w299 | w340);
assign w520 = v126;
assign w521 = (w520 & w518) | (w520 & w6266) | (w518 & w6266);
assign v127 = ~(w129 | w138);
assign w522 = v127;
assign w523 = w150 & w522;
assign v128 = ~(w412 | w494);
assign w524 = v128;
assign w525 = (w380 & w346) | (w380 & w6199) | (w346 & w6199);
assign w526 = w259 & w6267;
assign w527 = (w524 & w525) | (w524 & w6231) | (w525 & w6231);
assign w528 = ~w525 & w6232;
assign v129 = ~(w527 | w528);
assign w529 = v129;
assign v130 = ~(w238 | w299);
assign w530 = v130;
assign w531 = ~w518 & w6200;
assign v131 = ~(w379 | w412);
assign w532 = v131;
assign w533 = w341 & w6268;
assign w534 = w532 & w533;
assign w535 = ~w531 & w534;
assign w536 = w495 & w6233;
assign v132 = ~(w396 | w488);
assign w537 = v132;
assign w538 = ~w535 & w6201;
assign w539 = (w537 & w535) | (w537 & w6202) | (w535 & w6202);
assign v133 = ~(w538 | w539);
assign w540 = v133;
assign v134 = ~(w431 | w497);
assign w541 = v134;
assign w542 = (~w535 & w6234) | (~w535 & w6235) | (w6234 & w6235);
assign w543 = ~w541 & w542;
assign w544 = w541 & ~w542;
assign v135 = ~(w543 | w544);
assign w545 = v135;
assign w546 = ~w519 & w533;
assign w547 = w259 & w6269;
assign w548 = w448 & w532;
assign w549 = (w548 & w546) | (w548 & w6204) | (w546 & w6204);
assign v136 = ~(w215 | w497);
assign w550 = v136;
assign w551 = w495 & w550;
assign w552 = w491 & w551;
assign v137 = ~(w216 | w431);
assign w553 = v137;
assign w554 = w481 & w553;
assign w555 = pi041 & w206;
assign w556 = pi042 & w197;
assign w557 = pi048 & w199;
assign w558 = pi044 & w195;
assign w559 = pi043 & w204;
assign w560 = pi045 & w192;
assign w561 = pi046 & w189;
assign w562 = pi047 & w202;
assign v138 = ~(w555 | w556);
assign w563 = v138;
assign v139 = ~(w557 | w558);
assign w564 = v139;
assign v140 = ~(w559 | w560);
assign w565 = v140;
assign v141 = ~(w561 | w562);
assign w566 = v141;
assign w567 = w565 & w566;
assign w568 = w563 & w564;
assign w569 = w567 & w568;
assign w570 = w97 & ~w569;
assign w571 = ~w97 & w569;
assign v142 = ~(w570 | w571);
assign w572 = v142;
assign w573 = (w549 & w6270) | (w549 & w6271) | (w6270 & w6271);
assign w574 = (~w549 & w6272) | (~w549 & w6273) | (w6272 & w6273);
assign v143 = ~(w573 | w574);
assign w575 = v143;
assign v144 = ~(w447 | w487);
assign w576 = v144;
assign w577 = w495 & w6274;
assign w578 = (w576 & w415) | (w576 & w6275) | (w415 & w6275);
assign w579 = ~w415 & w6276;
assign v145 = ~(w578 | w579);
assign w580 = v145;
assign v146 = ~(w464 | w486);
assign w581 = v146;
assign w582 = w489 & w495;
assign w583 = (w6278 & w7361) | (w6278 & w7362) | (w7361 & w7362);
assign w584 = w581 & w7364;
assign v147 = ~(w583 | w584);
assign w585 = v147;
assign v148 = ~(w379 | w493);
assign w586 = v148;
assign w587 = (w586 & w546) | (w586 & w6236) | (w546 & w6236);
assign w588 = ~w546 & w6237;
assign v149 = ~(w587 | w588);
assign w589 = v149;
assign v150 = ~(w238 | w339);
assign w590 = v150;
assign v151 = ~(w279 | w342);
assign w591 = v151;
assign w592 = ~w338 & w591;
assign w593 = ~w338 & w6238;
assign w594 = (w590 & w593) | (w590 & w6279) | (w593 & w6279);
assign w595 = ~w593 & w6280;
assign v152 = ~(w594 | w595);
assign w596 = v152;
assign v153 = ~(w258 | w343);
assign w597 = v153;
assign w598 = ~w531 & w6281;
assign w599 = (w597 & w531) | (w597 & w6282) | (w531 & w6282);
assign v154 = ~(w598 | w599);
assign w600 = v154;
assign w601 = w517 & w523;
assign w602 = w521 & w601;
assign w603 = ~w516 & w602;
assign w604 = ~w589 & w6283;
assign w605 = ~w512 & w603;
assign v155 = ~(w529 | w540);
assign w606 = v155;
assign w607 = ~w580 & w604;
assign w608 = ~w585 & w607;
assign w609 = w605 & w6284;
assign w610 = ~w545 & w575;
assign w611 = w609 & w7334;
assign v156 = ~(pi296 | pi303);
assign w612 = v156;
assign w613 = w108 & w612;
assign v157 = ~(pi299 | pi300);
assign w614 = v157;
assign w615 = pi302 & w614;
assign w616 = w614 & w16;
assign w617 = w613 & w616;
assign w618 = w36 & w6285;
assign w619 = w617 & w618;
assign w620 = pi242 & w619;
assign w621 = (pi000 & ~w619) | (pi000 & w6286) | (~w619 & w6286);
assign w622 = pi215 & pi225;
assign w623 = pi184 & ~pi202;
assign w624 = ~w622 & w623;
assign w625 = w624 & w6287;
assign w626 = w624 & w6288;
assign w627 = (pi198 & ~w624) | (pi198 & w6289) | (~w624 & w6289);
assign v158 = ~(w625 | w627);
assign w628 = v158;
assign w629 = pi198 & pi217;
assign v159 = ~(pi215 | pi225);
assign w630 = v159;
assign w631 = ~w630 & w6290;
assign w632 = w629 & w631;
assign w633 = w631 & w6291;
assign v160 = ~(pi198 | pi217);
assign w634 = v160;
assign v161 = ~(w629 | w634);
assign w635 = v161;
assign w636 = pi198 & w631;
assign v162 = ~(pi198 | w631);
assign w637 = v162;
assign v163 = ~(w636 | w637);
assign w638 = v163;
assign v164 = ~(w635 | w638);
assign w639 = v164;
assign w640 = (~pi223 & ~w631) | (~pi223 & w6292) | (~w631 & w6292);
assign v165 = ~(w633 | w640);
assign w641 = v165;
assign w642 = ~w639 & w641;
assign w643 = (~w633 & w639) | (~w633 & w6293) | (w639 & w6293);
assign w644 = ~pi132 & w643;
assign w645 = (pi217 & ~w624) | (pi217 & w6295) | (~w624 & w6295);
assign v166 = ~(w626 | w645);
assign w646 = v166;
assign w647 = (w643 & w6296) | (w643 & w6297) | (w6296 & w6297);
assign v167 = ~(w628 | w635);
assign w648 = v167;
assign w649 = (w648 & ~w643) | (w648 & w6298) | (~w643 & w6298);
assign v168 = ~(w647 | w649);
assign w650 = v168;
assign w651 = pi129 & ~w650;
assign v169 = ~(pi132 | w633);
assign w652 = v169;
assign w653 = w639 & ~w652;
assign w654 = (~pi217 & ~w631) | (~pi217 & w634) | (~w631 & w634);
assign v170 = ~(w632 | w654);
assign w655 = v170;
assign w656 = (w643 & w6300) | (w643 & w6301) | (w6300 & w6301);
assign v171 = ~(pi129 | w653);
assign w657 = v171;
assign w658 = ~w656 & w657;
assign w659 = (~pi197 & w651) | (~pi197 & w6302) | (w651 & w6302);
assign w660 = (~pi184 & w630) | (~pi184 & w6303) | (w630 & w6303);
assign w661 = pi129 & pi225;
assign v172 = ~(pi129 | pi225);
assign w662 = v172;
assign v173 = ~(w661 | w662);
assign w663 = v173;
assign v174 = ~(w660 | w663);
assign w664 = v174;
assign w665 = pi215 & w664;
assign v175 = ~(pi215 | w664);
assign w666 = v175;
assign v176 = ~(w665 | w666);
assign w667 = v176;
assign w668 = pi129 & ~w624;
assign w669 = (~pi129 & w630) | (~pi129 & w6304) | (w630 & w6304);
assign v177 = ~(w668 | w669);
assign w670 = v177;
assign w671 = (pi216 & w668) | (pi216 & w6305) | (w668 & w6305);
assign w672 = ~w668 & w6306;
assign v178 = ~(w671 | w672);
assign w673 = v178;
assign w674 = ~w667 & w673;
assign w675 = pi129 & ~w628;
assign w676 = ~pi129 & w638;
assign v179 = ~(w675 | w676);
assign w677 = v179;
assign w678 = w644 & ~w677;
assign w679 = ~w644 & w677;
assign v180 = ~(w678 | w679);
assign w680 = v180;
assign w681 = (~w648 & ~w643) | (~w648 & w6307) | (~w643 & w6307);
assign w682 = pi223 & ~w626;
assign w683 = ~pi223 & w626;
assign v181 = ~(w682 | w683);
assign w684 = v181;
assign v182 = ~(w681 | w684);
assign w685 = v182;
assign w686 = (pi129 & ~w681) | (pi129 & w6308) | (~w681 & w6308);
assign w687 = ~w685 & w686;
assign w688 = (~w641 & w639) | (~w641 & w6309) | (w639 & w6309);
assign v183 = ~(w642 | w688);
assign w689 = v183;
assign v184 = ~(pi129 | w689);
assign w690 = v184;
assign w691 = (pi202 & w660) | (pi202 & w6310) | (w660 & w6310);
assign w692 = w668 & ~w691;
assign w693 = w623 & ~w630;
assign w694 = pi202 & w630;
assign v185 = ~(pi129 | w693);
assign w695 = v185;
assign w696 = ~w694 & w695;
assign v186 = ~(w692 | w696);
assign w697 = v186;
assign w698 = (~w697 & w687) | (~w697 & w6311) | (w687 & w6311);
assign w699 = pi256 & ~pi257;
assign w700 = ~pi241 & w699;
assign w701 = w699 & w6312;
assign v187 = ~(pi225 | w660);
assign w702 = v187;
assign w703 = pi225 & w660;
assign v188 = ~(w702 | w703);
assign w704 = v188;
assign w705 = w701 & w704;
assign w706 = w674 & w705;
assign w707 = w680 & w706;
assign w708 = w659 & w707;
assign v189 = ~(pi241 | pi257);
assign w709 = v189;
assign w710 = pi241 & pi257;
assign v190 = ~(w709 | w710);
assign w711 = v190;
assign w712 = pi256 & w711;
assign w713 = w711 & w6313;
assign v191 = ~(pi257 | pi271);
assign w714 = v191;
assign w715 = pi257 & ~pi273;
assign v192 = ~(w714 | w715);
assign w716 = v192;
assign v193 = ~(pi257 | pi272);
assign w717 = v193;
assign w718 = pi257 & ~pi275;
assign v194 = ~(w717 | w718);
assign w719 = v194;
assign v195 = ~(w716 | w719);
assign w720 = v195;
assign v196 = ~(pi257 | pi264);
assign w721 = v196;
assign w722 = pi257 & ~pi270;
assign v197 = ~(w721 | w722);
assign w723 = v197;
assign v198 = ~(pi223 | w723);
assign w724 = v198;
assign v199 = ~(pi257 | pi274);
assign w725 = v199;
assign w726 = pi257 & ~pi269;
assign v200 = ~(w725 | w726);
assign w727 = v200;
assign v201 = ~(pi216 | w727);
assign w728 = v201;
assign w729 = w634 & w720;
assign w730 = w724 & w728;
assign w731 = w729 & w730;
assign w732 = w713 & w731;
assign w733 = pi241 & ~w699;
assign w734 = ~w699 & w6314;
assign w735 = pi243 & ~pi256;
assign w736 = w709 & w735;
assign w737 = w0 & w736;
assign v202 = ~(w734 | w737);
assign w738 = v202;
assign w739 = (pi131 & w737) | (pi131 & w6315) | (w737 & w6315);
assign w740 = ~pi298 & w19;
assign w741 = w19 & w6316;
assign w742 = pi272 & pi303;
assign w743 = w16 & w742;
assign w744 = ~pi241 & pi257;
assign w745 = w735 & w744;
assign w746 = pi303 & w157;
assign w747 = w157 & w6317;
assign w748 = w24 & w6318;
assign w749 = ~pi298 & w22;
assign w750 = w22 & w6319;
assign v203 = ~(pi298 | pi302);
assign w751 = v203;
assign w752 = ~pi303 & w751;
assign w753 = w751 & w6320;
assign w754 = w11 & w6321;
assign w755 = pi269 & ~pi303;
assign w756 = w24 & w755;
assign w757 = ~w743 & w745;
assign w758 = ~w756 & w757;
assign v204 = ~(w741 | w747);
assign w759 = v204;
assign v205 = ~(w748 | w750);
assign w760 = v205;
assign v206 = ~(w753 | w754);
assign w761 = v206;
assign w762 = w760 & w761;
assign w763 = w758 & w759;
assign w764 = w762 & w763;
assign v207 = ~(pi225 | pi303);
assign w765 = v207;
assign w766 = ~pi202 & pi303;
assign v208 = ~(w765 | w766);
assign w767 = v208;
assign w768 = pi198 & pi303;
assign w769 = pi202 & ~pi303;
assign v209 = ~(w768 | w769);
assign w770 = v209;
assign w771 = ~w767 & w770;
assign w772 = pi223 & pi303;
assign w773 = w157 & w772;
assign w774 = w22 & w6322;
assign w775 = pi217 & ~pi303;
assign v210 = ~(w18 | w775);
assign w776 = v210;
assign w777 = w776 & w6323;
assign w778 = pi225 & pi303;
assign w779 = w751 & w6324;
assign w780 = w19 & ~w20;
assign v211 = ~(w778 | w780);
assign w781 = v211;
assign w782 = ~w779 & w781;
assign w783 = w777 & w782;
assign w784 = pi215 & pi303;
assign w785 = pi197 & ~pi303;
assign v212 = ~(w784 | w785);
assign w786 = v212;
assign w787 = pi198 & ~pi303;
assign v213 = ~(w772 | w787);
assign w788 = v213;
assign v214 = ~(pi216 | pi303);
assign w789 = v214;
assign w790 = ~pi217 & pi303;
assign v215 = ~(w789 | w790);
assign w791 = v215;
assign w792 = w788 & ~w791;
assign w793 = ~w788 & w791;
assign v216 = ~(w792 | w793);
assign w794 = v216;
assign w795 = pi216 & pi303;
assign w796 = pi215 & ~pi303;
assign v217 = ~(w795 | w796);
assign w797 = v217;
assign w798 = w794 & w797;
assign v218 = ~(w794 | w797);
assign w799 = v218;
assign v219 = ~(w798 | w799);
assign w800 = v219;
assign w801 = w786 & w800;
assign w802 = ~w0 & w736;
assign w803 = w771 & w792;
assign w804 = w802 & w803;
assign w805 = w783 & w804;
assign w806 = w801 & w805;
assign v220 = ~(pi278 | pi344);
assign w807 = v220;
assign v221 = ~(pi131 | w807);
assign w808 = v221;
assign w809 = ~pi241 & pi264;
assign w810 = (~w809 & ~w711) | (~w809 & w6325) | (~w711 & w6325);
assign w811 = (~pi197 & ~w711) | (~pi197 & w6327) | (~w711 & w6327);
assign w812 = pi197 & pi264;
assign w813 = ~w699 & w812;
assign v222 = ~(w810 | w813);
assign w814 = v222;
assign w815 = ~w811 & w814;
assign w816 = pi241 & ~pi264;
assign v223 = ~(w809 | w816);
assign w817 = v223;
assign w818 = pi197 & ~w817;
assign w819 = ~pi197 & w817;
assign v224 = ~(w818 | w819);
assign w820 = v224;
assign w821 = pi132 & ~pi256;
assign w822 = ~w711 & w821;
assign v225 = ~(pi241 | w821);
assign w823 = v225;
assign v226 = ~(w822 | w823);
assign w824 = v226;
assign v227 = ~(w820 | w824);
assign w825 = v227;
assign w826 = w820 & w824;
assign w827 = pi256 & ~w710;
assign v228 = ~(w825 | w827);
assign w828 = v228;
assign w829 = (~w815 & ~w828) | (~w815 & w6328) | (~w828 & w6328);
assign w830 = ~pi241 & pi275;
assign w831 = pi223 & w830;
assign v229 = ~(w712 | w831);
assign w832 = v229;
assign v230 = ~(pi223 | pi275);
assign w833 = v230;
assign w834 = pi223 & pi275;
assign w835 = ~w699 & w834;
assign v231 = ~(w833 | w835);
assign w836 = v231;
assign w837 = ~w832 & w836;
assign w838 = pi241 & ~pi275;
assign v232 = ~(w830 | w838);
assign w839 = v232;
assign w840 = pi223 & ~w839;
assign w841 = ~pi223 & w839;
assign v233 = ~(w840 | w841);
assign w842 = v233;
assign v234 = ~(pi241 | pi273);
assign w843 = v234;
assign w844 = pi241 & pi273;
assign v235 = ~(w843 | w844);
assign w845 = v235;
assign v236 = ~(pi198 | w845);
assign w846 = v236;
assign w847 = pi198 & w845;
assign v237 = ~(w846 | w847);
assign w848 = v237;
assign w849 = ~pi241 & pi270;
assign w850 = pi241 & ~pi270;
assign v238 = ~(w849 | w850);
assign w851 = v238;
assign w852 = pi216 & ~w851;
assign w853 = ~pi216 & w851;
assign v239 = ~(w852 | w853);
assign w854 = v239;
assign w855 = pi241 & ~pi272;
assign w856 = ~pi241 & pi272;
assign v240 = ~(w855 | w856);
assign w857 = v240;
assign w858 = pi202 & ~w857;
assign w859 = ~pi202 & w857;
assign v241 = ~(w858 | w859);
assign w860 = v241;
assign v242 = ~(pi241 | pi274);
assign w861 = v242;
assign w862 = pi241 & pi274;
assign v243 = ~(w861 | w862);
assign w863 = v243;
assign w864 = pi215 & w863;
assign v244 = ~(pi215 | w863);
assign w865 = v244;
assign v245 = ~(w864 | w865);
assign w866 = v245;
assign w867 = ~pi241 & pi271;
assign w868 = pi241 & ~pi271;
assign v246 = ~(w867 | w868);
assign w869 = v246;
assign w870 = pi225 & ~w869;
assign w871 = ~pi225 & w869;
assign w872 = w818 & ~w871;
assign v247 = ~(w870 | w872);
assign w873 = v247;
assign w874 = w866 & ~w873;
assign w875 = (~w864 & w873) | (~w864 & w6205) | (w873 & w6205);
assign w876 = w860 & ~w875;
assign v248 = ~(w870 | w871);
assign w877 = v248;
assign w878 = w826 & w877;
assign w879 = ~w866 & w873;
assign v249 = ~(w874 | w879);
assign w880 = v249;
assign w881 = w878 & w880;
assign w882 = ~w860 & w875;
assign v250 = ~(w876 | w882);
assign w883 = v250;
assign w884 = w881 & w883;
assign w885 = (~w858 & w875) | (~w858 & w6329) | (w875 & w6329);
assign w886 = ~w884 & w885;
assign w887 = (w884 & w6330) | (w884 & w6331) | (w6330 & w6331);
assign w888 = pi241 & ~pi269;
assign w889 = ~pi241 & pi269;
assign v251 = ~(w888 | w889);
assign w890 = v251;
assign w891 = pi217 & ~w890;
assign w892 = ~pi217 & w890;
assign v252 = ~(w891 | w892);
assign w893 = v252;
assign v253 = ~(w847 | w852);
assign w894 = v253;
assign v254 = ~(w846 | w894);
assign w895 = v254;
assign w896 = w893 & w895;
assign v255 = ~(w893 | w895);
assign w897 = v255;
assign v256 = ~(w896 | w897);
assign w898 = v256;
assign w899 = (~w891 & ~w895) | (~w891 & w6332) | (~w895 & w6332);
assign w900 = (w887 & w6336) | (w887 & w6337) | (w6336 & w6337);
assign w901 = (w887 & w6338) | (w887 & w6339) | (w6338 & w6339);
assign w902 = ~w900 & w901;
assign v257 = ~(w837 | w902);
assign w903 = v257;
assign v258 = ~(pi198 | pi273);
assign w904 = v258;
assign w905 = pi198 & pi273;
assign v259 = ~(pi241 | w905);
assign w906 = v259;
assign w907 = w699 & ~w906;
assign w908 = pi256 & w744;
assign w909 = ~w905 & w908;
assign v260 = ~(w907 | w909);
assign w910 = v260;
assign v261 = ~(w904 | w910);
assign w911 = v261;
assign w912 = ~w852 & w7365;
assign w913 = w848 & ~w912;
assign w914 = (~w827 & ~w912) | (~w827 & w6340) | (~w912 & w6340);
assign w915 = ~w913 & w914;
assign v262 = ~(w911 | w915);
assign w916 = v262;
assign w917 = pi202 & w856;
assign v263 = ~(w712 | w917);
assign w918 = v263;
assign v264 = ~(pi202 | pi272);
assign w919 = v264;
assign w920 = pi202 & pi272;
assign w921 = ~w699 & w920;
assign v265 = ~(w919 | w921);
assign w922 = v265;
assign w923 = ~w918 & w922;
assign v266 = ~(w881 | w883);
assign w924 = v266;
assign v267 = ~(w827 | w884);
assign w925 = v267;
assign w926 = (~w923 & ~w925) | (~w923 & w6341) | (~w925 & w6341);
assign w927 = w916 & w926;
assign w928 = (~w867 & ~w711) | (~w867 & w6342) | (~w711 & w6342);
assign w929 = (~pi225 & ~w711) | (~pi225 & w6344) | (~w711 & w6344);
assign w930 = pi225 & pi271;
assign w931 = ~w699 & w930;
assign v268 = ~(w928 | w931);
assign w932 = v268;
assign w933 = ~w929 & w932;
assign w934 = ~w826 & w6345;
assign w935 = (w877 & w826) | (w877 & w6346) | (w826 & w6346);
assign v269 = ~(w827 | w934);
assign w936 = v269;
assign w937 = (~w933 & ~w936) | (~w933 & w6347) | (~w936 & w6347);
assign w938 = pi217 & w889;
assign v270 = ~(w712 | w938);
assign w939 = v270;
assign v271 = ~(pi217 | pi269);
assign w940 = v271;
assign w941 = pi217 & pi269;
assign w942 = ~w699 & w941;
assign v272 = ~(w940 | w942);
assign w943 = v272;
assign w944 = ~w939 & w943;
assign v273 = ~(w887 | w898);
assign w945 = v273;
assign w946 = (~w827 & ~w887) | (~w827 & w6348) | (~w887 & w6348);
assign w947 = ~w945 & w946;
assign w948 = ~w947 & w6349;
assign v274 = ~(pi215 | pi274);
assign w949 = v274;
assign w950 = pi215 & pi274;
assign v275 = ~(pi241 | w950);
assign w951 = v275;
assign w952 = w699 & ~w951;
assign w953 = w908 & ~w950;
assign v276 = ~(w952 | w953);
assign w954 = v276;
assign v277 = ~(w949 | w954);
assign w955 = v277;
assign v278 = ~(w878 | w880);
assign w956 = v278;
assign w957 = (~w827 & ~w880) | (~w827 & w6350) | (~w880 & w6350);
assign w958 = ~w956 & w957;
assign v279 = ~(w955 | w958);
assign w959 = v279;
assign w960 = (~w849 & ~w711) | (~w849 & w6351) | (~w711 & w6351);
assign w961 = (~pi216 & ~w711) | (~pi216 & w6353) | (~w711 & w6353);
assign w962 = pi216 & pi270;
assign w963 = ~w699 & w962;
assign v280 = ~(w960 | w963);
assign w964 = v280;
assign w965 = ~w961 & w964;
assign w966 = ~w884 & w6354;
assign w967 = ~w827 & w7365;
assign w968 = ~w966 & w967;
assign w969 = ~w968 & w6355;
assign w970 = w829 & w969;
assign w971 = w927 & w6356;
assign v281 = ~(pi243 | w808);
assign w972 = v281;
assign w973 = (w971 & w6358) | (w971 & w6359) | (w6358 & w6359);
assign v282 = ~(w732 | w739);
assign w974 = v282;
assign w975 = ~w764 & w974;
assign w976 = ~w806 & w975;
assign w977 = (w976 & ~w708) | (w976 & w6360) | (~w708 & w6360);
assign w978 = (~w621 & ~w522) | (~w621 & w6362) | (~w522 & w6362);
assign w979 = w978 & w7366;
assign v283 = ~(w611 | w979);
assign w980 = v283;
assign w981 = ~pi001 & pi247;
assign w982 = w140 & w6363;
assign w983 = w82 & w982;
assign w984 = (~pi001 & ~w82) | (~pi001 & w6364) | (~w82 & w6364);
assign w985 = pi188 & pi189;
assign w986 = ~pi190 & w985;
assign v284 = ~(w82 | w986);
assign w987 = v284;
assign w988 = (pi099 & w82) | (pi099 & w6365) | (w82 & w6365);
assign w989 = ~w82 & w6366;
assign v285 = ~(w988 | w989);
assign w990 = v285;
assign w991 = w0 & ~w986;
assign w992 = w67 & w117;
assign w993 = w54 & w6367;
assign w994 = w992 & w993;
assign v286 = ~(w76 | w994);
assign w995 = v286;
assign w996 = ~pi296 & w48;
assign w997 = w84 & w996;
assign w998 = pi298 & w19;
assign w999 = w19 & w6368;
assign w1000 = pi299 & w999;
assign w1001 = ~w996 & w1000;
assign w1002 = (~w82 & w1001) | (~w82 & w6369) | (w1001 & w6369);
assign w1003 = w40 & w117;
assign w1004 = w42 & w65;
assign w1005 = w1003 & w1004;
assign w1006 = ~w82 & w1005;
assign v287 = ~(w1002 | w1006);
assign w1007 = v287;
assign w1008 = w69 & w985;
assign w1009 = w995 & ~w1008;
assign w1010 = (w991 & ~w1007) | (w991 & w6370) | (~w1007 & w6370);
assign w1011 = ~w1010 & w6371;
assign w1012 = (pi098 & w1010) | (pi098 & w6372) | (w1010 & w6372);
assign v288 = ~(w1011 | w1012);
assign w1013 = v288;
assign w1014 = pi296 & ~pi298;
assign w1015 = w48 & w88;
assign w1016 = w1014 & w1015;
assign w1017 = pi296 & pi297;
assign w1018 = w85 & w1017;
assign v289 = ~(w1016 | w1018);
assign w1019 = v289;
assign w1020 = (pi301 & ~w985) | (pi301 & w6139) | (~w985 & w6139);
assign w1021 = ~w1019 & w1020;
assign v290 = ~(w50 | w617);
assign w1022 = v290;
assign w1023 = w45 & w6373;
assign w1024 = ~w62 & w123;
assign w1025 = w1022 & ~w1023;
assign w1026 = w1024 & w1025;
assign w1027 = w991 & ~w1026;
assign v291 = ~(w987 | w1021);
assign w1028 = v291;
assign w1029 = ~w1027 & w6374;
assign w1030 = (~pi097 & w1027) | (~pi097 & w6375) | (w1027 & w6375);
assign v292 = ~(w990 | w1029);
assign w1031 = v292;
assign w1032 = ~w1030 & w1031;
assign w1033 = ~w1013 & w1032;
assign w1034 = w82 & w6376;
assign v293 = ~(w984 | w1034);
assign w1035 = v293;
assign w1036 = (w1035 & ~w1032) | (w1035 & w6377) | (~w1032 & w6377);
assign w1037 = pi195 & ~pi196;
assign w1038 = w45 & w1037;
assign w1039 = w45 & w6378;
assign w1040 = ~pi296 & pi297;
assign w1041 = w47 & w1040;
assign w1042 = ~pi291 & w1041;
assign w1043 = ~w32 & w1042;
assign w1044 = w39 & w56;
assign w1045 = w66 & w1044;
assign w1046 = w123 & ~w1045;
assign w1047 = (w9 & w1043) | (w9 & w6379) | (w1043 & w6379);
assign w1048 = pi190 & w100;
assign v294 = ~(pi276 | w7368);
assign w1049 = v294;
assign w1050 = w1032 & w6383;
assign w1051 = w108 & w160;
assign w1052 = w158 & w1051;
assign w1053 = pi277 & pi346;
assign w1054 = w1053 & w6207;
assign w1055 = w1053 & w6208;
assign v295 = ~(pi277 | pi346);
assign w1056 = v295;
assign w1057 = w1056 & w6209;
assign w1058 = ~pi277 & pi346;
assign w1059 = ~pi285 & w1058;
assign w1060 = w1058 & w6210;
assign w1061 = pi277 & ~pi346;
assign w1062 = pi285 & w1061;
assign w1063 = w1061 & w6211;
assign w1064 = ~pi285 & w1056;
assign w1065 = w1056 & w6212;
assign w1066 = pi285 & w1058;
assign w1067 = w1058 & w6213;
assign w1068 = w1061 & w6214;
assign v296 = ~(w1054 | w1055);
assign w1069 = v296;
assign v297 = ~(w1057 | w1060);
assign w1070 = v297;
assign v298 = ~(w1063 | w1065);
assign w1071 = v298;
assign v299 = ~(w1067 | w1068);
assign w1072 = v299;
assign w1073 = w1071 & w1072;
assign w1074 = w1069 & w1070;
assign w1075 = w1073 & w1074;
assign w1076 = w1052 & ~w1075;
assign w1077 = ~w1076 & w7368;
assign w1078 = pi195 & pi331;
assign w1079 = ~pi333 & w1078;
assign w1080 = w9 & w1079;
assign w1081 = w0 & w8;
assign w1082 = pi190 & w1081;
assign w1083 = w50 & w1082;
assign v300 = ~(w6 | w59);
assign w1084 = v300;
assign w1085 = w0 & ~w1084;
assign w1086 = ~w1084 & w6384;
assign v301 = ~(w1083 | w1086);
assign w1087 = v301;
assign w1088 = ~w1086 & w6385;
assign w1089 = pi276 & ~w1088;
assign w1090 = pi188 & ~pi310;
assign w1091 = pi190 & ~pi307;
assign w1092 = pi189 & ~pi308;
assign w1093 = ~pi189 & pi308;
assign w1094 = ~pi190 & pi307;
assign w1095 = ~pi188 & pi310;
assign v302 = ~(w1090 | w1091);
assign w1096 = v302;
assign v303 = ~(w1092 | w1093);
assign w1097 = v303;
assign v304 = ~(w1094 | w1095);
assign w1098 = v304;
assign w1099 = w1097 & w1098;
assign w1100 = w1096 & w1099;
assign w1101 = w1099 & w6386;
assign w1102 = ~w1086 & w6387;
assign v305 = ~(w1089 | w1102);
assign w1103 = v305;
assign w1104 = w996 & w999;
assign w1105 = ~pi299 & w1104;
assign w1106 = w66 & w118;
assign v306 = ~(w1105 | w1106);
assign w1107 = v306;
assign w1108 = (w986 & w1105) | (w986 & w6388) | (w1105 & w6388);
assign w1109 = pi294 & ~pi301;
assign w1110 = w8 & ~w88;
assign v307 = ~(pi190 | w1110);
assign w1111 = v307;
assign w1112 = w112 & w996;
assign w1113 = (w1109 & ~w1112) | (w1109 & w6389) | (~w1112 & w6389);
assign w1114 = pi299 & w57;
assign w1115 = pi298 & w55;
assign w1116 = w1114 & w1115;
assign v308 = ~(w77 | w1116);
assign w1117 = v308;
assign w1118 = w118 & w993;
assign w1119 = w57 & w1017;
assign w1120 = w157 & w1119;
assign w1121 = w75 & w1120;
assign v309 = ~(w1118 | w1121);
assign w1122 = v309;
assign w1123 = w54 & w6390;
assign w1124 = w992 & w1123;
assign w1125 = w993 & w1114;
assign v310 = ~(w1124 | w1125);
assign w1126 = v310;
assign w1127 = pi298 & ~pi299;
assign w1128 = pi291 & ~pi303;
assign w1129 = w65 & w74;
assign w1130 = w1127 & w1128;
assign w1131 = w1129 & w1130;
assign w1132 = w108 & w614;
assign w1133 = ~pi296 & w24;
assign w1134 = w1132 & w1133;
assign w1135 = ~pi303 & w1134;
assign w1136 = w88 & ~w996;
assign w1137 = ~w998 & w1136;
assign w1138 = w614 & w24;
assign w1139 = w1128 & w1138;
assign w1140 = w1138 & w6391;
assign v311 = ~(w1137 | w1140);
assign w1141 = v311;
assign w1142 = w55 & w992;
assign v312 = ~(w1135 | w1142);
assign w1143 = v312;
assign w1144 = w1141 & w1143;
assign w1145 = w44 & w1003;
assign w1146 = w1119 & w1138;
assign v313 = ~(w1131 | w1145);
assign w1147 = v313;
assign w1148 = ~w1146 & w1147;
assign w1149 = w1122 & w1148;
assign w1150 = w1126 & w1149;
assign w1151 = w1144 & w1150;
assign w1152 = pi299 & w82;
assign w1153 = w1138 & w6392;
assign w1154 = ~w37 & w1153;
assign w1155 = (~pi300 & ~w19) | (~pi300 & w6393) | (~w19 & w6393);
assign w1156 = w996 & w1155;
assign w1157 = w1104 & w6394;
assign v314 = ~(w1154 | w1156);
assign w1158 = v314;
assign w1159 = (~w1152 & ~w1158) | (~w1152 & w6395) | (~w1158 & w6395);
assign w1160 = w123 & w1084;
assign w1161 = w3 & w614;
assign w1162 = ~w998 & w1161;
assign w1163 = ~w1116 & w6396;
assign w1164 = w1160 & w1163;
assign w1165 = w1150 & w6397;
assign w1166 = ~w1159 & w1165;
assign w1167 = w996 & w1000;
assign w1168 = w68 & w1123;
assign v315 = ~(w62 | w69);
assign w1169 = v315;
assign v316 = ~(w45 | w110);
assign w1170 = v316;
assign v317 = ~(w994 | w1168);
assign w1171 = v317;
assign w1172 = w1169 & w1170;
assign w1173 = w1172 & w6398;
assign w1174 = w84 & ~w996;
assign w1175 = ~pi291 & w1127;
assign w1176 = w44 & w1175;
assign w1177 = w117 & w120;
assign w1178 = w615 & w1177;
assign v318 = ~(w1176 | w1178);
assign w1179 = v318;
assign v319 = ~(w1106 | w1174);
assign w1180 = v319;
assign w1181 = w1179 & w1180;
assign w1182 = ~w1045 & w1181;
assign w1183 = w1173 & w1182;
assign w1184 = w66 & w992;
assign w1185 = pi296 & ~pi297;
assign w1186 = w614 & w1185;
assign w1187 = w39 & w1186;
assign w1188 = w118 & w1123;
assign w1189 = w1044 & w1123;
assign v320 = ~(w1188 | w1189);
assign w1190 = v320;
assign v321 = ~(w101 | w1190);
assign w1191 = v321;
assign v322 = ~(w1041 | w1184);
assign w1192 = v322;
assign w1193 = ~w1187 & w1192;
assign w1194 = ~w1006 & w1193;
assign w1195 = ~w1191 & w1194;
assign w1196 = w117 & w1040;
assign w1197 = w616 & w1196;
assign w1198 = w73 & w612;
assign w1199 = w616 & w1198;
assign v323 = ~(w1197 | w1199);
assign w1200 = v323;
assign w1201 = w75 & w6399;
assign w1202 = w48 & w614;
assign w1203 = w1014 & w1202;
assign w1204 = w41 & w1004;
assign w1205 = ~w82 & w1204;
assign w1206 = w117 & w1186;
assign v324 = ~(w1203 | w1206);
assign w1207 = v324;
assign w1208 = ~w1205 & w1207;
assign w1209 = w42 & w1175;
assign w1210 = w1175 & w1004;
assign w1211 = w53 & w1210;
assign w1212 = w1138 & w1198;
assign w1213 = w1138 & w1196;
assign v325 = ~(w1212 | w1213);
assign w1214 = v325;
assign v326 = ~(w9 | w1214);
assign w1215 = v326;
assign w1216 = w1022 & ~w1201;
assign w1217 = w1200 & ~w1211;
assign w1218 = w1216 & w1217;
assign w1219 = w1208 & ~w1215;
assign w1220 = w1218 & w1219;
assign w1221 = w1194 & w6400;
assign w1222 = w1220 & w1221;
assign w1223 = w1183 & w1222;
assign w1224 = w1166 & w1223;
assign w1225 = w0 & ~w1224;
assign w1226 = ~w82 & w85;
assign w1227 = w36 & w6401;
assign w1228 = w1226 & ~w1227;
assign w1229 = w88 & w1017;
assign w1230 = w157 & w1229;
assign w1231 = w1229 & w6402;
assign w1232 = ~w8 & w1231;
assign w1233 = w108 & w88;
assign w1234 = ~pi296 & w1233;
assign w1235 = ~w82 & w1234;
assign w1236 = w88 & w1198;
assign v327 = ~(w1235 | w1236);
assign w1237 = v327;
assign v328 = ~(w89 | w98);
assign w1238 = v328;
assign w1239 = ~w1232 & w1238;
assign w1240 = ~w1228 & w1239;
assign w1241 = w1237 & w1240;
assign w1242 = ~w82 & w6131;
assign w1243 = ~pi291 & w1229;
assign w1244 = w53 & w1243;
assign w1245 = pi296 & w1233;
assign w1246 = ~w82 & w1245;
assign w1247 = (w48 & ~w1229) | (w48 & w6403) | (~w1229 & w6403);
assign w1248 = (w88 & w1247) | (w88 & w6404) | (w1247 & w6404);
assign w1249 = w4 & w42;
assign v329 = ~(w1246 | w1249);
assign w1250 = v329;
assign w1251 = ~w1248 & w1250;
assign v330 = ~(w1242 | w1244);
assign w1252 = v330;
assign w1253 = w1251 & w1252;
assign w1254 = w1241 & w1253;
assign w1255 = (~w1113 & w1254) | (~w1113 & w6405) | (w1254 & w6405);
assign w1256 = (~w986 & w1225) | (~w986 & w6406) | (w1225 & w6406);
assign v331 = ~(w1108 | w1256);
assign w1257 = v331;
assign w1258 = pi190 & w985;
assign w1259 = ~w1109 & w1258;
assign w1260 = (~w1259 & w1256) | (~w1259 & w6407) | (w1256 & w6407);
assign w1261 = w1250 & w6408;
assign w1262 = (pi301 & ~w1241) | (pi301 & w6409) | (~w1241 & w6409);
assign v332 = ~(w82 | w1200);
assign w1263 = v332;
assign w1264 = ~w617 & w1181;
assign w1265 = w1264 & w6410;
assign v333 = ~(w1184 | w1188);
assign w1266 = v333;
assign v334 = ~(w1045 | w1210);
assign w1267 = v334;
assign v335 = ~(w1042 | w1213);
assign w1268 = v335;
assign w1269 = w1267 & w1268;
assign v336 = ~(w1187 | w1212);
assign w1270 = v336;
assign v337 = ~(w49 | w1189);
assign w1271 = v337;
assign w1272 = ~w1201 & w1271;
assign w1273 = w1270 & w1272;
assign w1274 = w1266 & w1269;
assign w1275 = w1173 & w1274;
assign w1276 = w1273 & w1275;
assign w1277 = w1007 & w1265;
assign w1278 = w1276 & w1277;
assign w1279 = w1166 & w1278;
assign v338 = ~(w1113 | w1262);
assign w1280 = v338;
assign w1281 = (w1280 & w1279) | (w1280 & w6411) | (w1279 & w6411);
assign w1282 = (~w1108 & w1281) | (~w1108 & w6412) | (w1281 & w6412);
assign v339 = ~(w1259 | w1282);
assign w1283 = v339;
assign v340 = ~(pi305 | w153);
assign w1284 = v340;
assign w1285 = (w1284 & w1282) | (w1284 & w6413) | (w1282 & w6413);
assign v341 = ~(w1260 | w1285);
assign w1286 = v341;
assign w1287 = ~w37 & w98;
assign w1288 = (~pi296 & ~w8) | (~pi296 & w6414) | (~w8 & w6414);
assign w1289 = w86 & w1288;
assign w1290 = w91 & ~w1289;
assign w1291 = ~w101 & w1018;
assign w1292 = ~w82 & w2725;
assign v342 = ~(w1231 | w1287);
assign w1293 = v342;
assign w1294 = ~w1291 & w1293;
assign w1295 = w1237 & w1294;
assign w1296 = w1290 & ~w1292;
assign w1297 = w1295 & w6415;
assign w1298 = w53 & w59;
assign w1299 = w32 & w82;
assign w1300 = w32 & w6416;
assign w1301 = w1214 & w1267;
assign w1302 = ~w50 & w1170;
assign w1303 = w1024 & w1302;
assign v343 = ~(w37 | w1303);
assign w1304 = v343;
assign w1305 = w6 & w34;
assign v344 = ~(w2 | w82);
assign w1306 = v344;
assign w1307 = ~w8 & w69;
assign w1308 = w1306 & w1307;
assign v345 = ~(w997 | w1105);
assign w1309 = v345;
assign w1310 = w38 & w45;
assign v346 = ~(w1000 | w1161);
assign w1311 = v346;
assign v347 = ~(w1116 | w1156);
assign w1312 = v347;
assign v348 = ~(w1168 | w1298);
assign w1313 = v348;
assign w1314 = ~w1310 & w1313;
assign w1315 = w1312 & w6417;
assign w1316 = w1301 & w1314;
assign w1317 = ~w1308 & w1309;
assign w1318 = w1316 & w1317;
assign w1319 = w1195 & w1315;
assign v349 = ~(w1300 | w1304);
assign w1320 = v349;
assign w1321 = w1319 & w1320;
assign w1322 = w1151 & w1318;
assign w1323 = w1265 & ~w1305;
assign w1324 = w1322 & w1323;
assign w1325 = (w0 & ~w1324) | (w0 & w6418) | (~w1324 & w6418);
assign v350 = ~(w985 | w1109);
assign w1326 = v350;
assign w1327 = (w1326 & w1297) | (w1326 & w6419) | (w1297 & w6419);
assign w1328 = ~w1325 & w1327;
assign w1329 = ~w1286 & w6420;
assign w1330 = w1283 & w1328;
assign w1331 = ~w1257 & w1330;
assign w1332 = w1330 & w6421;
assign v351 = ~(w1260 | w1328);
assign w1333 = v351;
assign w1334 = ~w1283 & w1333;
assign w1335 = pi305 & ~w153;
assign w1336 = w1333 & w6422;
assign w1337 = pi276 & w1336;
assign w1338 = w1257 & w1330;
assign w1339 = w1330 & w6423;
assign w1340 = (~w153 & w1325) | (~w153 & w6424) | (w1325 & w6424);
assign w1341 = ~w1283 & w6425;
assign w1342 = w1283 & w1333;
assign w1343 = w1229 & w6426;
assign w1344 = w0 & w1210;
assign v352 = ~(w1343 | w1344);
assign w1345 = v352;
assign w1346 = (w2 & w1344) | (w2 & w6427) | (w1344 & w6427);
assign w1347 = pi282 & w1346;
assign w1348 = (~pi276 & ~w1346) | (~pi276 & w6428) | (~w1346 & w6428);
assign w1349 = w1346 & w1764;
assign v353 = ~(w1348 | w1349);
assign w1350 = v353;
assign w1351 = w1333 & w6429;
assign v354 = ~(w1332 | w1341);
assign w1352 = v354;
assign v355 = ~(w1339 | w1351);
assign w1353 = v355;
assign w1354 = w1352 & w1353;
assign v356 = ~(w1329 | w1337);
assign w1355 = v356;
assign w1356 = w1354 & w1355;
assign w1357 = (w1103 & w1356) | (w1103 & w6430) | (w1356 & w6430);
assign w1358 = (w1077 & w1357) | (w1077 & w6431) | (w1357 & w6431);
assign v357 = ~(pi247 | w1036);
assign w1359 = v357;
assign w1360 = (w1359 & w1358) | (w1359 & w6432) | (w1358 & w6432);
assign w1361 = pi359 & ~w981;
assign w1362 = ~w1360 & w1361;
assign w1363 = ~pi002 & pi247;
assign w1364 = (w1047 & w6433) | (w1047 & w6434) | (w6433 & w6434);
assign w1365 = w1032 & w6435;
assign w1366 = w1056 & w6436;
assign w1367 = w1061 & w6437;
assign w1368 = w1058 & w6438;
assign w1369 = w1056 & w6439;
assign w1370 = w1053 & w6440;
assign w1371 = w1061 & w6441;
assign w1372 = w1053 & w6442;
assign w1373 = w1058 & w6443;
assign v358 = ~(w1366 | w1367);
assign w1374 = v358;
assign v359 = ~(w1368 | w1369);
assign w1375 = v359;
assign v360 = ~(w1370 | w1371);
assign w1376 = v360;
assign v361 = ~(w1372 | w1373);
assign w1377 = v361;
assign w1378 = w1376 & w1377;
assign w1379 = w1374 & w1375;
assign w1380 = w1378 & w1379;
assign w1381 = w1052 & ~w1380;
assign w1382 = ~w1381 & w7368;
assign w1383 = pi268 & ~w1088;
assign v362 = ~(w1102 | w1383);
assign w1384 = v362;
assign w1385 = w1330 & w6444;
assign w1386 = (~pi268 & ~w1346) | (~pi268 & w6445) | (~w1346 & w6445);
assign w1387 = w1346 & w6446;
assign w1388 = w1333 & w6447;
assign v363 = ~(w1336 | w1388);
assign w1389 = v363;
assign v364 = ~(w1386 | w1389);
assign w1390 = v364;
assign w1391 = ~w1283 & w6448;
assign w1392 = w1330 & w6449;
assign w1393 = ~w1286 & w6450;
assign v365 = ~(w1385 | w1391);
assign w1394 = v365;
assign w1395 = w1394 & w6451;
assign w1396 = ~w1390 & w1395;
assign w1397 = (w1384 & w1396) | (w1384 & w6452) | (w1396 & w6452);
assign w1398 = (w1382 & w1397) | (w1382 & w6453) | (w1397 & w6453);
assign w1399 = (~pi002 & ~w82) | (~pi002 & w6454) | (~w82 & w6454);
assign w1400 = w82 & w6455;
assign v366 = ~(w1399 | w1400);
assign w1401 = v366;
assign w1402 = (w1401 & ~w1032) | (w1401 & w6456) | (~w1032 & w6456);
assign v367 = ~(pi247 | w1402);
assign w1403 = v367;
assign w1404 = (w1403 & w1398) | (w1403 & w6457) | (w1398 & w6457);
assign w1405 = pi359 & ~w1363;
assign w1406 = ~w1404 & w1405;
assign w1407 = ~pi003 & pi247;
assign w1408 = (w1047 & w6458) | (w1047 & w6459) | (w6458 & w6459);
assign w1409 = w1032 & w6460;
assign w1410 = w1061 & w6461;
assign w1411 = w1053 & w6462;
assign w1412 = w1056 & w6463;
assign w1413 = w1058 & w6464;
assign w1414 = w1058 & w6465;
assign w1415 = w1053 & w6466;
assign w1416 = w1056 & w6467;
assign w1417 = w1061 & w6468;
assign v368 = ~(w1410 | w1411);
assign w1418 = v368;
assign v369 = ~(w1412 | w1413);
assign w1419 = v369;
assign v370 = ~(w1414 | w1415);
assign w1420 = v370;
assign v371 = ~(w1416 | w1417);
assign w1421 = v371;
assign w1422 = w1420 & w1421;
assign w1423 = w1418 & w1419;
assign w1424 = w1422 & w1423;
assign w1425 = w1052 & ~w1424;
assign w1426 = ~w1425 & w7368;
assign w1427 = pi246 & ~w1088;
assign v372 = ~(w1102 | w1427);
assign w1428 = v372;
assign w1429 = ~w1283 & w6469;
assign w1430 = pi265 & pi268;
assign w1431 = w1346 & w6470;
assign w1432 = w1346 & w6471;
assign w1433 = w1333 & w6472;
assign v373 = ~(w1336 | w1433);
assign w1434 = v373;
assign w1435 = pi246 & ~w1434;
assign w1436 = w1330 & w6473;
assign w1437 = w1346 & w6474;
assign w1438 = ~w1286 & w6475;
assign w1439 = w1330 & w6476;
assign v374 = ~(w1429 | w1437);
assign w1440 = v374;
assign w1441 = ~w1436 & w1440;
assign w1442 = w1441 & w6477;
assign w1443 = ~w1435 & w1442;
assign w1444 = (w1428 & w1443) | (w1428 & w6478) | (w1443 & w6478);
assign w1445 = (w1426 & w1444) | (w1426 & w6479) | (w1444 & w6479);
assign w1446 = (~pi003 & ~w82) | (~pi003 & w6480) | (~w82 & w6480);
assign w1447 = w82 & w6481;
assign v375 = ~(w1446 | w1447);
assign w1448 = v375;
assign w1449 = (w1448 & ~w1032) | (w1448 & w6482) | (~w1032 & w6482);
assign v376 = ~(pi247 | w1449);
assign w1450 = v376;
assign w1451 = (w1450 & w1445) | (w1450 & w6483) | (w1445 & w6483);
assign w1452 = pi359 & ~w1407;
assign w1453 = ~w1451 & w1452;
assign w1454 = ~pi004 & pi247;
assign w1455 = (w1047 & w6484) | (w1047 & w6485) | (w6484 & w6485);
assign w1456 = w1032 & w6486;
assign w1457 = w1061 & w6487;
assign w1458 = w1053 & w6488;
assign w1459 = w1058 & w6489;
assign w1460 = w1058 & w6490;
assign w1461 = w1053 & w6491;
assign w1462 = w1061 & w6492;
assign w1463 = w1056 & w6493;
assign w1464 = w1056 & w6494;
assign v377 = ~(w1457 | w1458);
assign w1465 = v377;
assign v378 = ~(w1459 | w1460);
assign w1466 = v378;
assign v379 = ~(w1461 | w1462);
assign w1467 = v379;
assign v380 = ~(w1463 | w1464);
assign w1468 = v380;
assign w1469 = w1467 & w1468;
assign w1470 = w1465 & w1466;
assign w1471 = w1469 & w1470;
assign w1472 = w1052 & ~w1471;
assign w1473 = ~w1472 & w7368;
assign w1474 = pi233 & ~w1088;
assign v381 = ~(w1102 | w1474);
assign w1475 = v381;
assign w1476 = w1330 & w6495;
assign w1477 = (~pi233 & ~w1346) | (~pi233 & w6497) | (~w1346 & w6497);
assign w1478 = w1346 & w6498;
assign w1479 = w1342 & ~w1478;
assign w1480 = (~w1477 & w1479) | (~w1477 & w6499) | (w1479 & w6499);
assign w1481 = ~w1283 & w6500;
assign w1482 = w1330 & w6501;
assign w1483 = ~w1286 & w6502;
assign v382 = ~(w1476 | w1481);
assign w1484 = v382;
assign w1485 = w1484 & w6503;
assign w1486 = ~w1480 & w1485;
assign w1487 = (w1475 & w1486) | (w1475 & w6504) | (w1486 & w6504);
assign w1488 = (w1473 & w1487) | (w1473 & w6505) | (w1487 & w6505);
assign w1489 = (~pi004 & ~w82) | (~pi004 & w6506) | (~w82 & w6506);
assign w1490 = w82 & w6507;
assign v383 = ~(w1489 | w1490);
assign w1491 = v383;
assign w1492 = (w1491 & ~w1032) | (w1491 & w6508) | (~w1032 & w6508);
assign v384 = ~(pi247 | w1492);
assign w1493 = v384;
assign w1494 = (w1493 & w1488) | (w1493 & w6509) | (w1488 & w6509);
assign w1495 = pi359 & ~w1454;
assign w1496 = ~w1494 & w1495;
assign v385 = ~(pi234 | pi240);
assign w1497 = v385;
assign w1498 = ~pi231 & pi251;
assign w1499 = ~w1497 & w1498;
assign w1500 = pi097 & ~pi098;
assign w1501 = ~pi099 & w1500;
assign w1502 = w1500 & w6510;
assign v386 = ~(pi242 | w1502);
assign w1503 = v386;
assign w1504 = pi256 & w710;
assign w1505 = w710 & w6511;
assign w1506 = pi242 & w1505;
assign v387 = ~(w1503 | w1506);
assign w1507 = v387;
assign w1508 = w1507 & w6512;
assign w1509 = ~w82 & w141;
assign v388 = ~(w148 | w1509);
assign w1510 = v388;
assign w1511 = ~w143 & w7369;
assign w1512 = w129 & w138;
assign w1513 = (~pi361 & ~w82) | (~pi361 & w6514) | (~w82 & w6514);
assign w1514 = w1511 & ~w1513;
assign w1515 = ~w1512 & w1514;
assign w1516 = (~pi247 & w1515) | (~pi247 & w6516) | (w1515 & w6516);
assign w1517 = w206 & w1516;
assign w1518 = pi284 & ~w162;
assign v389 = ~(pi283 | w162);
assign w1519 = v389;
assign v390 = ~(w1518 | w1519);
assign w1520 = v390;
assign w1521 = pi280 & ~w162;
assign w1522 = pi304 & w162;
assign v391 = ~(w1521 | w1522);
assign w1523 = v391;
assign w1524 = w1520 & w1523;
assign w1525 = ~pi006 & w1524;
assign w1526 = ~w162 & w6517;
assign w1527 = w1523 & w1526;
assign w1528 = w1523 & w6518;
assign w1529 = ~w162 & w6519;
assign w1530 = ~w1523 & w1529;
assign w1531 = ~w1523 & w6520;
assign w1532 = ~w162 & w6521;
assign w1533 = w1523 & w1532;
assign w1534 = w1523 & w6522;
assign w1535 = ~w1523 & w1532;
assign w1536 = ~w1523 & w6523;
assign w1537 = w1523 & w1529;
assign w1538 = w1523 & w6524;
assign w1539 = w1520 & ~w1523;
assign w1540 = ~pi010 & w1539;
assign w1541 = ~w1523 & w1526;
assign w1542 = ~w1523 & w6525;
assign v392 = ~(w1525 | w1528);
assign w1543 = v392;
assign v393 = ~(w1531 | w1534);
assign w1544 = v393;
assign v394 = ~(w1536 | w1538);
assign w1545 = v394;
assign v395 = ~(w1540 | w1542);
assign w1546 = v395;
assign w1547 = w1545 & w1546;
assign w1548 = w1543 & w1544;
assign w1549 = w1547 & w1548;
assign w1550 = w162 & ~w1549;
assign v396 = ~(w165 | w1511);
assign w1551 = v396;
assign w1552 = w1136 & w6526;
assign v397 = ~(pi242 | pi347);
assign w1553 = v397;
assign w1554 = w736 & ~w788;
assign w1555 = pi241 & w735;
assign w1556 = (~pi269 & ~w19) | (~pi269 & w6528) | (~w19 & w6528);
assign w1557 = w19 & w6529;
assign w1558 = w1555 & ~w1556;
assign w1559 = ~w1557 & w1558;
assign w1560 = ~w651 & w6530;
assign w1561 = w745 & w756;
assign w1562 = w711 & w6531;
assign w1563 = pi242 & ~w1554;
assign w1564 = ~w1561 & w1563;
assign w1565 = w1564 & w6532;
assign w1566 = ~w1560 & w1565;
assign w1567 = w1566 & w7370;
assign v398 = ~(w1552 | w1553);
assign w1568 = v398;
assign w1569 = pi269 & w1552;
assign w1570 = (~w1569 & w1567) | (~w1569 & w6533) | (w1567 & w6533);
assign w1571 = ~pi250 & w165;
assign w1572 = ~w162 & w7371;
assign v399 = ~(w1550 | w1572);
assign w1573 = v399;
assign w1574 = (w502 & w6535) | (w502 & w6536) | (w6535 & w6536);
assign w1575 = (~pi005 & ~w206) | (~pi005 & w6537) | (~w206 & w6537);
assign v400 = ~(w1574 | w1575);
assign w1576 = v400;
assign w1577 = w197 & w1516;
assign w1578 = (w502 & w6538) | (w502 & w6539) | (w6538 & w6539);
assign w1579 = (~pi006 & ~w197) | (~pi006 & w6540) | (~w197 & w6540);
assign v401 = ~(w1578 | w1579);
assign w1580 = v401;
assign w1581 = w204 & w1516;
assign w1582 = (w502 & w6541) | (w502 & w6542) | (w6541 & w6542);
assign w1583 = (~pi007 & ~w204) | (~pi007 & w6543) | (~w204 & w6543);
assign v402 = ~(w1582 | w1583);
assign w1584 = v402;
assign w1585 = w195 & w1516;
assign w1586 = (w502 & w6544) | (w502 & w6545) | (w6544 & w6545);
assign w1587 = (~pi008 & ~w195) | (~pi008 & w6546) | (~w195 & w6546);
assign v403 = ~(w1586 | w1587);
assign w1588 = v403;
assign w1589 = w192 & w1516;
assign w1590 = (w502 & w6547) | (w502 & w6548) | (w6547 & w6548);
assign w1591 = (~pi009 & ~w192) | (~pi009 & w6549) | (~w192 & w6549);
assign v404 = ~(w1590 | w1591);
assign w1592 = v404;
assign w1593 = w189 & w1516;
assign w1594 = (w502 & w6550) | (w502 & w6551) | (w6550 & w6551);
assign w1595 = (~pi010 & ~w189) | (~pi010 & w6552) | (~w189 & w6552);
assign v405 = ~(w1594 | w1595);
assign w1596 = v405;
assign w1597 = w202 & w1516;
assign w1598 = (w502 & w6553) | (w502 & w6554) | (w6553 & w6554);
assign w1599 = (~pi011 & ~w202) | (~pi011 & w6555) | (~w202 & w6555);
assign v406 = ~(w1598 | w1599);
assign w1600 = v406;
assign w1601 = w199 & w1516;
assign w1602 = (w502 & w6556) | (w502 & w6557) | (w6556 & w6557);
assign v407 = ~(pi012 | w1601);
assign w1603 = v407;
assign v408 = ~(w1602 | w1603);
assign w1604 = v408;
assign v409 = ~(pi242 | pi352);
assign w1605 = v409;
assign w1606 = w736 & ~w770;
assign w1607 = (~pi270 & ~w11) | (~pi270 & w6559) | (~w11 & w6559);
assign w1608 = w11 & w6529;
assign w1609 = w1555 & ~w1607;
assign w1610 = ~w1608 & w1609;
assign w1611 = ~w673 & w701;
assign w1612 = w745 & w754;
assign w1613 = w711 & w6560;
assign w1614 = pi242 & ~w1606;
assign w1615 = ~w1612 & w1614;
assign w1616 = w1615 & w6561;
assign w1617 = ~w1611 & w1616;
assign v410 = ~(w1552 | w1605);
assign w1618 = v410;
assign w1619 = pi270 & w1552;
assign w1620 = ~w1619 & w7372;
assign w1621 = ~pi249 & w165;
assign w1622 = ~w162 & w7373;
assign w1623 = ~pi015 & w1537;
assign w1624 = ~w1523 & w6567;
assign w1625 = ~w1523 & w6568;
assign w1626 = ~pi014 & w1524;
assign w1627 = w1523 & w6569;
assign w1628 = ~pi018 & w1539;
assign w1629 = w1523 & w6570;
assign w1630 = ~w1523 & w6571;
assign v411 = ~(w1623 | w1624);
assign w1631 = v411;
assign v412 = ~(w1625 | w1626);
assign w1632 = v412;
assign v413 = ~(w1627 | w1628);
assign w1633 = v413;
assign v414 = ~(w1629 | w1630);
assign w1634 = v414;
assign w1635 = w1633 & w1634;
assign w1636 = w1631 & w1632;
assign w1637 = w1635 & w1636;
assign w1638 = w162 & ~w1637;
assign v415 = ~(w1622 | w1638);
assign w1639 = v415;
assign w1640 = (w1639 & ~w512) | (w1639 & w6572) | (~w512 & w6572);
assign w1641 = w1517 & ~w1640;
assign w1642 = (~pi013 & ~w206) | (~pi013 & w6573) | (~w206 & w6573);
assign v416 = ~(w1641 | w1642);
assign w1643 = v416;
assign w1644 = (w512 & w6574) | (w512 & w6575) | (w6574 & w6575);
assign w1645 = (~pi014 & ~w197) | (~pi014 & w6576) | (~w197 & w6576);
assign v417 = ~(w1644 | w1645);
assign w1646 = v417;
assign w1647 = (w512 & w6577) | (w512 & w6578) | (w6577 & w6578);
assign w1648 = (~pi015 & ~w204) | (~pi015 & w6579) | (~w204 & w6579);
assign v418 = ~(w1647 | w1648);
assign w1649 = v418;
assign w1650 = (w512 & w6580) | (w512 & w6581) | (w6580 & w6581);
assign w1651 = (~pi016 & ~w195) | (~pi016 & w6582) | (~w195 & w6582);
assign v419 = ~(w1650 | w1651);
assign w1652 = v419;
assign w1653 = (w512 & w6583) | (w512 & w6584) | (w6583 & w6584);
assign w1654 = (~pi017 & ~w192) | (~pi017 & w6585) | (~w192 & w6585);
assign v420 = ~(w1653 | w1654);
assign w1655 = v420;
assign w1656 = (w512 & w6586) | (w512 & w6587) | (w6586 & w6587);
assign w1657 = (~pi018 & ~w189) | (~pi018 & w6588) | (~w189 & w6588);
assign v421 = ~(w1656 | w1657);
assign w1658 = v421;
assign w1659 = (w512 & w6589) | (w512 & w6590) | (w6589 & w6590);
assign w1660 = (~pi019 & ~w202) | (~pi019 & w6591) | (~w202 & w6591);
assign v422 = ~(w1659 | w1660);
assign w1661 = v422;
assign w1662 = (w512 & w6592) | (w512 & w6593) | (w6592 & w6593);
assign w1663 = (~pi020 & ~w199) | (~pi020 & w6594) | (~w199 & w6594);
assign v423 = ~(w1662 | w1663);
assign w1664 = v423;
assign w1665 = pi026 & w1539;
assign w1666 = w1523 & w6595;
assign w1667 = ~w1523 & w6596;
assign w1668 = ~w1523 & w6597;
assign w1669 = w1523 & w6598;
assign w1670 = pi022 & w1524;
assign w1671 = w1523 & w6599;
assign w1672 = ~w1523 & w6600;
assign v424 = ~(w1665 | w1666);
assign w1673 = v424;
assign v425 = ~(w1667 | w1668);
assign w1674 = v425;
assign v426 = ~(w1669 | w1670);
assign w1675 = v426;
assign v427 = ~(w1671 | w1672);
assign w1676 = v427;
assign w1677 = w1675 & w1676;
assign w1678 = w1673 & w1674;
assign w1679 = w1677 & w1678;
assign w1680 = w162 & w1679;
assign v428 = ~(pi242 | pi351);
assign w1681 = v428;
assign w1682 = w736 & w767;
assign w1683 = (~pi274 & ~w19) | (~pi274 & w6601) | (~w19 & w6601);
assign w1684 = w19 & w6602;
assign w1685 = w1555 & ~w1683;
assign w1686 = ~w1684 & w1685;
assign w1687 = w667 & w701;
assign w1688 = w741 & w745;
assign w1689 = w713 & w727;
assign w1690 = pi242 & ~w1682;
assign w1691 = ~w1688 & w1690;
assign w1692 = w1691 & w6604;
assign w1693 = ~w1687 & w1692;
assign v429 = ~(w1552 | w1681);
assign w1694 = v429;
assign w1695 = (w958 & w6607) | (w958 & w6608) | (w6607 & w6608);
assign w1696 = pi274 & w1552;
assign v430 = ~(w1695 | w1696);
assign w1697 = v430;
assign w1698 = w1551 & ~w1697;
assign w1699 = ~pi248 & w165;
assign v431 = ~(w162 | w1699);
assign w1700 = v431;
assign w1701 = (w1700 & w1697) | (w1700 & w6609) | (w1697 & w6609);
assign v432 = ~(w1680 | w1701);
assign w1702 = v432;
assign w1703 = (~w1702 & ~w580) | (~w1702 & w6610) | (~w580 & w6610);
assign w1704 = w1517 & ~w1703;
assign w1705 = (pi021 & ~w206) | (pi021 & w6611) | (~w206 & w6611);
assign v433 = ~(w1704 | w1705);
assign w1706 = v433;
assign w1707 = (w580 & w6612) | (w580 & w6613) | (w6612 & w6613);
assign w1708 = (pi022 & ~w197) | (pi022 & w6614) | (~w197 & w6614);
assign v434 = ~(w1707 | w1708);
assign w1709 = v434;
assign w1710 = (w580 & w6615) | (w580 & w6616) | (w6615 & w6616);
assign w1711 = (pi023 & ~w204) | (pi023 & w6617) | (~w204 & w6617);
assign v435 = ~(w1710 | w1711);
assign w1712 = v435;
assign w1713 = (w580 & w6618) | (w580 & w6619) | (w6618 & w6619);
assign w1714 = (pi024 & ~w195) | (pi024 & w6620) | (~w195 & w6620);
assign v436 = ~(w1713 | w1714);
assign w1715 = v436;
assign w1716 = (w580 & w6621) | (w580 & w6622) | (w6621 & w6622);
assign w1717 = (pi025 & ~w192) | (pi025 & w6623) | (~w192 & w6623);
assign v437 = ~(w1716 | w1717);
assign w1718 = v437;
assign w1719 = (w580 & w6624) | (w580 & w6625) | (w6624 & w6625);
assign w1720 = (pi026 & ~w189) | (pi026 & w6626) | (~w189 & w6626);
assign v438 = ~(w1719 | w1720);
assign w1721 = v438;
assign w1722 = (w580 & w6627) | (w580 & w6628) | (w6627 & w6628);
assign w1723 = (pi027 & ~w202) | (pi027 & w6629) | (~w202 & w6629);
assign v439 = ~(w1722 | w1723);
assign w1724 = v439;
assign w1725 = (w580 & w6630) | (w580 & w6631) | (w6630 & w6631);
assign w1726 = (pi028 & ~w199) | (pi028 & w6632) | (~w199 & w6632);
assign v440 = ~(w1725 | w1726);
assign w1727 = v440;
assign w1728 = pi247 & pi359;
assign w1729 = pi029 & w1728;
assign w1730 = w82 & w6633;
assign w1731 = ~pi247 & pi359;
assign w1732 = ~pi099 & w82;
assign w1733 = w82 & w6634;
assign w1734 = ~pi029 & w1733;
assign w1735 = (w1047 & w6635) | (w1047 & w6636) | (w6635 & w6636);
assign w1736 = w1032 & w6637;
assign w1737 = (pi029 & ~w1032) | (pi029 & w6638) | (~w1032 & w6638);
assign w1738 = w1032 & w6639;
assign w1739 = w1058 & w6640;
assign w1740 = w1061 & w6641;
assign w1741 = w1058 & w6642;
assign w1742 = w1056 & w6643;
assign w1743 = w1056 & w6644;
assign w1744 = w1061 & w6645;
assign w1745 = w1053 & w6646;
assign w1746 = w1053 & w6647;
assign v441 = ~(w1739 | w1740);
assign w1747 = v441;
assign v442 = ~(w1741 | w1742);
assign w1748 = v442;
assign v443 = ~(w1743 | w1744);
assign w1749 = v443;
assign v444 = ~(w1745 | w1746);
assign w1750 = v444;
assign w1751 = w1749 & w1750;
assign w1752 = w1747 & w1748;
assign w1753 = w1751 & w1752;
assign w1754 = w1052 & w1753;
assign w1755 = w1738 & ~w1754;
assign w1756 = w1088 & ~w1101;
assign w1757 = ~w1283 & w6648;
assign w1758 = w1330 & w6649;
assign w1759 = pi229 & w1336;
assign w1760 = ~w1286 & w6650;
assign v445 = ~(pi348 | w1346);
assign w1761 = v445;
assign w1762 = pi233 & pi244;
assign w1763 = pi246 & pi259;
assign w1764 = pi276 & pi282;
assign w1765 = w1763 & w1764;
assign w1766 = w1430 & w1762;
assign w1767 = w1765 & w1766;
assign w1768 = pi238 & w1767;
assign w1769 = w1767 & w6651;
assign w1770 = w1767 & w6652;
assign w1771 = w1767 & w6653;
assign w1772 = (~pi229 & ~w1767) | (~pi229 & w6654) | (~w1767 & w6654);
assign v446 = ~(w1771 | w1772);
assign w1773 = v446;
assign w1774 = w1346 & ~w1773;
assign v447 = ~(w1761 | w1774);
assign w1775 = v447;
assign w1776 = w1333 & w6655;
assign w1777 = w1330 & w6656;
assign v448 = ~(w1757 | w1758);
assign w1778 = v448;
assign v449 = ~(w1776 | w1777);
assign w1779 = v449;
assign w1780 = w1778 & w1779;
assign v450 = ~(w1759 | w1760);
assign w1781 = v450;
assign w1782 = w1780 & w1781;
assign w1783 = (pi229 & w1086) | (pi229 & w6657) | (w1086 & w6657);
assign w1784 = w1080 & ~w1101;
assign w1785 = w1087 & w6658;
assign v451 = ~(w1052 | w1783);
assign w1786 = v451;
assign w1787 = ~w1785 & w1786;
assign w1788 = (w1787 & w1782) | (w1787 & w6659) | (w1782 & w6659);
assign v452 = ~(w1732 | w1736);
assign w1789 = v452;
assign w1790 = ~w1737 & w1789;
assign w1791 = ~w1730 & w1731;
assign w1792 = ~w1734 & w1791;
assign w1793 = w1792 & w7374;
assign v453 = ~(w1729 | w1793);
assign w1794 = v453;
assign w1795 = pi030 & w1728;
assign w1796 = w82 & w6661;
assign w1797 = ~pi030 & w1733;
assign w1798 = (w1047 & w6662) | (w1047 & w6663) | (w6662 & w6663);
assign w1799 = w1032 & w6664;
assign w1800 = (pi030 & ~w1032) | (pi030 & w6665) | (~w1032 & w6665);
assign w1801 = w1061 & w6666;
assign w1802 = w1058 & w6667;
assign w1803 = w1058 & w6668;
assign w1804 = w1053 & w6669;
assign w1805 = w1056 & w6670;
assign w1806 = w1053 & w6671;
assign w1807 = w1056 & w6672;
assign w1808 = w1061 & w6673;
assign v454 = ~(w1801 | w1802);
assign w1809 = v454;
assign v455 = ~(w1803 | w1804);
assign w1810 = v455;
assign v456 = ~(w1805 | w1806);
assign w1811 = v456;
assign v457 = ~(w1807 | w1808);
assign w1812 = v457;
assign w1813 = w1811 & w1812;
assign w1814 = w1809 & w1810;
assign w1815 = w1813 & w1814;
assign w1816 = w1052 & w1815;
assign w1817 = w1738 & ~w1816;
assign w1818 = ~w1283 & w6674;
assign w1819 = w1330 & w6675;
assign w1820 = pi226 & w1336;
assign w1821 = ~w1286 & w6676;
assign v458 = ~(pi352 | w1346);
assign w1822 = v458;
assign w1823 = pi226 & w1771;
assign v459 = ~(pi226 | w1771);
assign w1824 = v459;
assign v460 = ~(w1823 | w1824);
assign w1825 = v460;
assign w1826 = w1346 & ~w1825;
assign v461 = ~(w1822 | w1826);
assign w1827 = v461;
assign w1828 = w1333 & w6677;
assign w1829 = w1330 & w6678;
assign v462 = ~(w1818 | w1819);
assign w1830 = v462;
assign v463 = ~(w1828 | w1829);
assign w1831 = v463;
assign w1832 = w1830 & w1831;
assign v464 = ~(w1820 | w1821);
assign w1833 = v464;
assign w1834 = w1832 & w1833;
assign w1835 = (pi226 & w1086) | (pi226 & w6679) | (w1086 & w6679);
assign w1836 = w1087 & w6680;
assign v465 = ~(w1052 | w1835);
assign w1837 = v465;
assign w1838 = ~w1836 & w1837;
assign w1839 = (w1838 & w1834) | (w1838 & w6681) | (w1834 & w6681);
assign v466 = ~(w1732 | w1799);
assign w1840 = v466;
assign w1841 = ~w1800 & w1840;
assign w1842 = w1731 & ~w1796;
assign w1843 = ~w1797 & w1842;
assign w1844 = w1843 & w7375;
assign v467 = ~(w1795 | w1844);
assign w1845 = v467;
assign w1846 = pi031 & w1728;
assign w1847 = w82 & w6683;
assign w1848 = ~pi031 & w1733;
assign w1849 = (w1047 & w6684) | (w1047 & w6685) | (w6684 & w6685);
assign w1850 = w1032 & w6686;
assign w1851 = (pi031 & ~w1032) | (pi031 & w6687) | (~w1032 & w6687);
assign w1852 = w1053 & w6688;
assign w1853 = w1053 & w6689;
assign w1854 = w1061 & w6690;
assign w1855 = w1058 & w6691;
assign w1856 = w1058 & w6692;
assign w1857 = w1056 & w6693;
assign w1858 = w1056 & w6694;
assign w1859 = w1061 & w6695;
assign v468 = ~(w1852 | w1853);
assign w1860 = v468;
assign v469 = ~(w1854 | w1855);
assign w1861 = v469;
assign v470 = ~(w1856 | w1857);
assign w1862 = v470;
assign v471 = ~(w1858 | w1859);
assign w1863 = v471;
assign w1864 = w1862 & w1863;
assign w1865 = w1860 & w1861;
assign w1866 = w1864 & w1865;
assign w1867 = w1052 & w1866;
assign w1868 = w1738 & ~w1867;
assign w1869 = ~w1283 & w6696;
assign w1870 = w1330 & w6697;
assign w1871 = pi227 & w1336;
assign w1872 = ~w1286 & w6698;
assign v472 = ~(pi353 | w1346);
assign w1873 = v472;
assign w1874 = w1771 & w6699;
assign w1875 = (~pi227 & ~w1771) | (~pi227 & w6700) | (~w1771 & w6700);
assign v473 = ~(w1874 | w1875);
assign w1876 = v473;
assign w1877 = w1346 & ~w1876;
assign v474 = ~(w1873 | w1877);
assign w1878 = v474;
assign w1879 = w1333 & w6701;
assign w1880 = w1330 & w6702;
assign v475 = ~(w1869 | w1870);
assign w1881 = v475;
assign v476 = ~(w1879 | w1880);
assign w1882 = v476;
assign w1883 = w1881 & w1882;
assign v477 = ~(w1871 | w1872);
assign w1884 = v477;
assign w1885 = w1883 & w1884;
assign w1886 = (pi227 & w1086) | (pi227 & w6703) | (w1086 & w6703);
assign w1887 = w1087 & w6704;
assign v478 = ~(w1052 | w1886);
assign w1888 = v478;
assign w1889 = ~w1887 & w1888;
assign w1890 = (w1889 & w1885) | (w1889 & w6705) | (w1885 & w6705);
assign v479 = ~(w1732 | w1850);
assign w1891 = v479;
assign w1892 = ~w1851 & w1891;
assign w1893 = w1731 & ~w1847;
assign w1894 = ~w1848 & w1893;
assign w1895 = w1894 & w7376;
assign v480 = ~(w1846 | w1895);
assign w1896 = v480;
assign w1897 = pi032 & w1728;
assign w1898 = w82 & w6707;
assign w1899 = ~pi032 & w1733;
assign w1900 = (w1047 & w6708) | (w1047 & w6709) | (w6708 & w6709);
assign w1901 = w1032 & w6710;
assign w1902 = (pi032 & ~w1032) | (pi032 & w6711) | (~w1032 & w6711);
assign w1903 = w1056 & w6712;
assign w1904 = w1053 & w6713;
assign w1905 = w1058 & w6714;
assign w1906 = w1061 & w6715;
assign w1907 = w1056 & w6716;
assign w1908 = w1058 & w6717;
assign w1909 = w1053 & w6718;
assign w1910 = w1061 & w6719;
assign v481 = ~(w1903 | w1904);
assign w1911 = v481;
assign v482 = ~(w1905 | w1906);
assign w1912 = v482;
assign v483 = ~(w1907 | w1908);
assign w1913 = v483;
assign v484 = ~(w1909 | w1910);
assign w1914 = v484;
assign w1915 = w1913 & w1914;
assign w1916 = w1911 & w1912;
assign w1917 = w1915 & w1916;
assign w1918 = w1052 & w1917;
assign w1919 = w1738 & ~w1918;
assign w1920 = ~w1283 & w6720;
assign w1921 = w1330 & w6721;
assign w1922 = pi191 & w1336;
assign w1923 = ~w1286 & w6722;
assign v485 = ~(pi347 | w1346);
assign w1924 = v485;
assign w1925 = (~pi191 & ~w1771) | (~pi191 & w6723) | (~w1771 & w6723);
assign w1926 = w1771 & w6724;
assign v486 = ~(w1925 | w1926);
assign w1927 = v486;
assign w1928 = w1346 & ~w1927;
assign v487 = ~(w1924 | w1928);
assign w1929 = v487;
assign w1930 = w1333 & w6725;
assign w1931 = w1330 & w6726;
assign v488 = ~(w1920 | w1921);
assign w1932 = v488;
assign v489 = ~(w1930 | w1931);
assign w1933 = v489;
assign w1934 = w1932 & w1933;
assign v490 = ~(w1922 | w1923);
assign w1935 = v490;
assign w1936 = w1934 & w1935;
assign w1937 = (pi191 & w1086) | (pi191 & w6727) | (w1086 & w6727);
assign w1938 = w1087 & w6728;
assign v491 = ~(w1052 | w1937);
assign w1939 = v491;
assign w1940 = ~w1938 & w1939;
assign w1941 = (w1940 & w1936) | (w1940 & w6729) | (w1936 & w6729);
assign v492 = ~(w1732 | w1901);
assign w1942 = v492;
assign w1943 = ~w1902 & w1942;
assign w1944 = w1731 & ~w1898;
assign w1945 = ~w1899 & w1944;
assign w1946 = w1945 & w7377;
assign v493 = ~(w1897 | w1946);
assign w1947 = v493;
assign w1948 = pi033 & w1728;
assign w1949 = w82 & w6731;
assign w1950 = ~pi033 & w1733;
assign w1951 = (~pi033 & ~w1032) | (~pi033 & w6732) | (~w1032 & w6732);
assign w1952 = (w1047 & w6733) | (w1047 & w6734) | (w6733 & w6734);
assign w1953 = w1032 & w6735;
assign v494 = ~(w1951 | w1953);
assign w1954 = v494;
assign w1955 = w1056 & w6736;
assign w1956 = w1053 & w6737;
assign w1957 = w1053 & w6738;
assign w1958 = w1058 & w6739;
assign w1959 = w1058 & w6740;
assign w1960 = w1056 & w6741;
assign w1961 = w1061 & w6742;
assign w1962 = w1061 & w6743;
assign v495 = ~(w1955 | w1956);
assign w1963 = v495;
assign v496 = ~(w1957 | w1958);
assign w1964 = v496;
assign v497 = ~(w1959 | w1960);
assign w1965 = v497;
assign v498 = ~(w1961 | w1962);
assign w1966 = v498;
assign w1967 = w1965 & w1966;
assign w1968 = w1963 & w1964;
assign w1969 = w1967 & w1968;
assign w1970 = w1052 & w1969;
assign w1971 = w1738 & ~w1970;
assign w1972 = ~w1283 & w6744;
assign w1973 = w1330 & w6745;
assign w1974 = pi222 & w1336;
assign w1975 = ~w1286 & w6746;
assign v499 = ~(pi351 | w1346);
assign w1976 = v499;
assign w1977 = (~pi222 & ~w1767) | (~pi222 & w6747) | (~w1767 & w6747);
assign v500 = ~(w1770 | w1977);
assign w1978 = v500;
assign w1979 = w1346 & ~w1978;
assign v501 = ~(w1976 | w1979);
assign w1980 = v501;
assign w1981 = w1333 & w6748;
assign w1982 = w1330 & w6749;
assign v502 = ~(w1972 | w1973);
assign w1983 = v502;
assign v503 = ~(w1981 | w1982);
assign w1984 = v503;
assign w1985 = w1983 & w1984;
assign v504 = ~(w1974 | w1975);
assign w1986 = v504;
assign w1987 = w1985 & w1986;
assign w1988 = (pi222 & w1086) | (pi222 & w6750) | (w1086 & w6750);
assign w1989 = w1087 & w6751;
assign v505 = ~(w1052 | w1988);
assign w1990 = v505;
assign w1991 = ~w1989 & w1990;
assign w1992 = (w1991 & w1987) | (w1991 & w6752) | (w1987 & w6752);
assign v506 = ~(w1732 | w1954);
assign w1993 = v506;
assign w1994 = w1731 & ~w1949;
assign w1995 = ~w1950 & w1994;
assign w1996 = w1995 & w7378;
assign v507 = ~(w1948 | w1996);
assign w1997 = v507;
assign w1998 = pi034 & w1728;
assign w1999 = w82 & w6754;
assign w2000 = ~pi034 & w1733;
assign w2001 = (w1047 & w6755) | (w1047 & w6756) | (w6755 & w6756);
assign w2002 = w1032 & w6757;
assign w2003 = (pi034 & ~w1032) | (pi034 & w6758) | (~w1032 & w6758);
assign w2004 = w1056 & w6759;
assign w2005 = w1053 & w6760;
assign w2006 = w1058 & w6761;
assign w2007 = w1061 & w6762;
assign w2008 = w1058 & w6763;
assign w2009 = w1053 & w6764;
assign w2010 = w1061 & w6765;
assign w2011 = w1056 & w6766;
assign v508 = ~(w2004 | w2005);
assign w2012 = v508;
assign v509 = ~(w2006 | w2007);
assign w2013 = v509;
assign v510 = ~(w2008 | w2009);
assign w2014 = v510;
assign v511 = ~(w2010 | w2011);
assign w2015 = v511;
assign w2016 = w2014 & w2015;
assign w2017 = w2012 & w2013;
assign w2018 = w2016 & w2017;
assign w2019 = w1052 & w2018;
assign w2020 = w1738 & ~w2019;
assign v512 = ~(w1088 | w1102);
assign w2021 = v512;
assign w2022 = (~w1052 & ~w2021) | (~w1052 & w6767) | (~w2021 & w6767);
assign w2023 = (~pi259 & ~w1346) | (~pi259 & w6768) | (~w1346 & w6768);
assign v513 = ~(w1434 | w2023);
assign w2024 = v513;
assign w2025 = ~w1283 & w6769;
assign w2026 = w1330 & w6770;
assign w2027 = ~w1286 & w6771;
assign w2028 = (~w2025 & ~w1331) | (~w2025 & w6772) | (~w1331 & w6772);
assign w2029 = w2028 & w6773;
assign w2030 = ~w2024 & w2029;
assign w2031 = (w2022 & w2030) | (w2022 & w6774) | (w2030 & w6774);
assign v514 = ~(w1732 | w2002);
assign w2032 = v514;
assign w2033 = ~w2003 & w2032;
assign w2034 = w1731 & ~w1999;
assign w2035 = ~w2000 & w2034;
assign w2036 = w2035 & w7379;
assign v515 = ~(w1998 | w2036);
assign w2037 = v515;
assign w2038 = w82 & w6776;
assign w2039 = (pi035 & ~w82) | (pi035 & w6777) | (~w82 & w6777);
assign v516 = ~(w2038 | w2039);
assign w2040 = v516;
assign w2041 = (~w2040 & ~w1032) | (~w2040 & w6778) | (~w1032 & w6778);
assign w2042 = (w1047 & w6779) | (w1047 & w6780) | (w6779 & w6780);
assign w2043 = w1032 & w6781;
assign w2044 = w1058 & w6782;
assign w2045 = w1053 & w6783;
assign w2046 = w1058 & w6784;
assign w2047 = w1061 & w6785;
assign w2048 = w1053 & w6786;
assign w2049 = w1061 & w6787;
assign w2050 = w1056 & w6788;
assign w2051 = w1056 & w6789;
assign v517 = ~(w2044 | w2045);
assign w2052 = v517;
assign v518 = ~(w2046 | w2047);
assign w2053 = v518;
assign v519 = ~(w2048 | w2049);
assign w2054 = v519;
assign v520 = ~(w2050 | w2051);
assign w2055 = v520;
assign w2056 = w2054 & w2055;
assign w2057 = w2052 & w2053;
assign w2058 = w2056 & w2057;
assign w2059 = w1052 & ~w2058;
assign w2060 = ~w2059 & w7368;
assign w2061 = pi282 & w2021;
assign w2062 = w1330 & w6790;
assign w2063 = ~w1283 & w6791;
assign v521 = ~(pi282 | w1346);
assign w2064 = v521;
assign v522 = ~(w1347 | w2064);
assign w2065 = v522;
assign w2066 = w1333 & w6792;
assign w2067 = pi282 & w1336;
assign w2068 = ~w1286 & w6793;
assign w2069 = w1330 & w6794;
assign v523 = ~(w2062 | w2063);
assign w2070 = v523;
assign v524 = ~(w2066 | w2069);
assign w2071 = v524;
assign w2072 = w2070 & w2071;
assign v525 = ~(w2067 | w2068);
assign w2073 = v525;
assign w2074 = w2072 & w2073;
assign w2075 = (~w2061 & w2074) | (~w2061 & w6795) | (w2074 & w6795);
assign w2076 = (w2060 & w2075) | (w2060 & w6796) | (w2075 & w6796);
assign v526 = ~(pi247 | w2041);
assign w2077 = v526;
assign w2078 = (w2077 & w2076) | (w2077 & w6797) | (w2076 & w6797);
assign w2079 = ~pi035 & pi247;
assign w2080 = pi359 & ~w2079;
assign w2081 = ~w2078 & w2080;
assign w2082 = pi036 & w1728;
assign w2083 = w82 & w6798;
assign w2084 = ~pi036 & w1733;
assign w2085 = (w1047 & w6799) | (w1047 & w6800) | (w6799 & w6800);
assign w2086 = w1032 & w6801;
assign w2087 = (pi036 & ~w1032) | (pi036 & w6802) | (~w1032 & w6802);
assign w2088 = w1061 & w6803;
assign w2089 = w1058 & w6804;
assign w2090 = w1053 & w6805;
assign w2091 = w1056 & w6806;
assign w2092 = w1061 & w6807;
assign w2093 = w1058 & w6808;
assign w2094 = w1056 & w6809;
assign w2095 = w1053 & w6810;
assign v527 = ~(w2088 | w2089);
assign w2096 = v527;
assign v528 = ~(w2090 | w2091);
assign w2097 = v528;
assign v529 = ~(w2092 | w2093);
assign w2098 = v529;
assign v530 = ~(w2094 | w2095);
assign w2099 = v530;
assign w2100 = w2098 & w2099;
assign w2101 = w2096 & w2097;
assign w2102 = w2100 & w2101;
assign w2103 = w1052 & w2102;
assign w2104 = w1738 & ~w2103;
assign w2105 = (~w1052 & ~w2021) | (~w1052 & w6811) | (~w2021 & w6811);
assign w2106 = (~pi265 & ~w1346) | (~pi265 & w6812) | (~w1346 & w6812);
assign w2107 = w1333 & w6813;
assign v531 = ~(w1336 | w2107);
assign w2108 = v531;
assign v532 = ~(w2106 | w2108);
assign w2109 = v532;
assign w2110 = ~w1283 & w6814;
assign w2111 = w1330 & w6815;
assign w2112 = ~w1286 & w6816;
assign w2113 = (~w2110 & ~w1338) | (~w2110 & w6817) | (~w1338 & w6817);
assign w2114 = w2113 & w6818;
assign w2115 = ~w2109 & w2114;
assign w2116 = (w2105 & w2115) | (w2105 & w6819) | (w2115 & w6819);
assign v533 = ~(w1732 | w2086);
assign w2117 = v533;
assign w2118 = ~w2087 & w2117;
assign w2119 = w1731 & ~w2083;
assign w2120 = ~w2084 & w2119;
assign w2121 = w2120 & w7380;
assign v534 = ~(w2082 | w2121);
assign w2122 = v534;
assign w2123 = pi037 & w1728;
assign w2124 = w82 & w6821;
assign w2125 = ~pi037 & w1733;
assign w2126 = (~pi037 & ~w1032) | (~pi037 & w6822) | (~w1032 & w6822);
assign w2127 = (w1047 & w6823) | (w1047 & w6824) | (w6823 & w6824);
assign w2128 = w1032 & w6825;
assign v535 = ~(w2126 | w2128);
assign w2129 = v535;
assign w2130 = w1061 & w6826;
assign w2131 = w1058 & w6827;
assign w2132 = w1056 & w6828;
assign w2133 = w1061 & w6829;
assign w2134 = w1058 & w6830;
assign w2135 = w1053 & w6831;
assign w2136 = w1056 & w6832;
assign w2137 = w1053 & w6833;
assign v536 = ~(w2130 | w2131);
assign w2138 = v536;
assign v537 = ~(w2132 | w2133);
assign w2139 = v537;
assign v538 = ~(w2134 | w2135);
assign w2140 = v538;
assign v539 = ~(w2136 | w2137);
assign w2141 = v539;
assign w2142 = w2140 & w2141;
assign w2143 = w2138 & w2139;
assign w2144 = w2142 & w2143;
assign w2145 = w1052 & w2144;
assign w2146 = ~w1283 & w6834;
assign w2147 = w1330 & w6835;
assign w2148 = ~pi224 & w1336;
assign w2149 = ~w1286 & w6836;
assign v540 = ~(pi350 | w1346);
assign w2150 = v540;
assign w2151 = (pi224 & ~w1771) | (pi224 & w6837) | (~w1771 & w6837);
assign w2152 = w1771 & w6838;
assign v541 = ~(w2151 | w2152);
assign w2153 = v541;
assign w2154 = w1346 & ~w2153;
assign v542 = ~(w2150 | w2154);
assign w2155 = v542;
assign w2156 = w1333 & w6839;
assign w2157 = w1330 & w6840;
assign v543 = ~(w2146 | w2147);
assign w2158 = v543;
assign v544 = ~(w2156 | w2157);
assign w2159 = v544;
assign w2160 = w2158 & w2159;
assign v545 = ~(w2148 | w2149);
assign w2161 = v545;
assign w2162 = w2160 & w2161;
assign w2163 = (~pi224 & w1086) | (~pi224 & w6841) | (w1086 & w6841);
assign w2164 = w1087 & w6842;
assign v546 = ~(w1052 | w2163);
assign w2165 = v546;
assign w2166 = ~w2164 & w2165;
assign w2167 = w1738 & ~w2145;
assign v547 = ~(w1732 | w2129);
assign w2168 = v547;
assign w2169 = w1731 & ~w2124;
assign w2170 = ~w2125 & w2169;
assign w2171 = w2170 & w7381;
assign v548 = ~(w2123 | w2171);
assign w2172 = v548;
assign w2173 = pi038 & w1728;
assign w2174 = w82 & w6848;
assign w2175 = ~pi038 & w1733;
assign w2176 = (w1047 & w6849) | (w1047 & w6850) | (w6849 & w6850);
assign w2177 = w1032 & w6851;
assign w2178 = (pi038 & ~w1032) | (pi038 & w6852) | (~w1032 & w6852);
assign w2179 = w1056 & w6853;
assign w2180 = w1061 & w6854;
assign w2181 = w1056 & w6855;
assign w2182 = w1053 & w6856;
assign w2183 = w1058 & w6857;
assign w2184 = w1053 & w6858;
assign w2185 = w1058 & w6859;
assign w2186 = w1061 & w6860;
assign v549 = ~(w2179 | w2180);
assign w2187 = v549;
assign v550 = ~(w2181 | w2182);
assign w2188 = v550;
assign v551 = ~(w2183 | w2184);
assign w2189 = v551;
assign v552 = ~(w2185 | w2186);
assign w2190 = v552;
assign w2191 = w2189 & w2190;
assign w2192 = w2187 & w2188;
assign w2193 = w2191 & w2192;
assign w2194 = w1052 & w2193;
assign w2195 = w1738 & ~w2194;
assign w2196 = ~w1283 & w6861;
assign w2197 = w1330 & w6862;
assign w2198 = pi238 & w1336;
assign w2199 = ~w1286 & w6863;
assign v553 = ~(pi354 | w1346);
assign w2200 = v553;
assign v554 = ~(pi238 | w1767);
assign w2201 = v554;
assign v555 = ~(w1768 | w2201);
assign w2202 = v555;
assign w2203 = w1346 & ~w2202;
assign v556 = ~(w2200 | w2203);
assign w2204 = v556;
assign w2205 = w1333 & w6864;
assign w2206 = w1330 & w6865;
assign v557 = ~(w2196 | w2197);
assign w2207 = v557;
assign v558 = ~(w2205 | w2206);
assign w2208 = v558;
assign w2209 = w2207 & w2208;
assign v559 = ~(w2198 | w2199);
assign w2210 = v559;
assign w2211 = w2209 & w2210;
assign w2212 = (pi238 & w1086) | (pi238 & w6866) | (w1086 & w6866);
assign w2213 = w1087 & w6867;
assign v560 = ~(w1052 | w2212);
assign w2214 = v560;
assign w2215 = ~w2213 & w2214;
assign w2216 = (w2215 & w2211) | (w2215 & w6868) | (w2211 & w6868);
assign v561 = ~(w1732 | w2177);
assign w2217 = v561;
assign w2218 = ~w2178 & w2217;
assign w2219 = w1731 & ~w2174;
assign w2220 = ~w2175 & w2219;
assign w2221 = w2220 & w7382;
assign v562 = ~(w2173 | w2221);
assign w2222 = v562;
assign w2223 = pi039 & w1728;
assign w2224 = w82 & w6870;
assign w2225 = ~pi039 & w1733;
assign w2226 = w1056 & w6871;
assign w2227 = w1053 & w6872;
assign w2228 = w1058 & w6873;
assign w2229 = w1058 & w6874;
assign w2230 = w1061 & w6875;
assign w2231 = w1053 & w6876;
assign w2232 = w1061 & w6877;
assign w2233 = w1056 & w6878;
assign v563 = ~(w2226 | w2227);
assign w2234 = v563;
assign v564 = ~(w2228 | w2229);
assign w2235 = v564;
assign v565 = ~(w2230 | w2231);
assign w2236 = v565;
assign v566 = ~(w2232 | w2233);
assign w2237 = v566;
assign w2238 = w2236 & w2237;
assign w2239 = w2234 & w2235;
assign w2240 = w2238 & w2239;
assign w2241 = w1052 & w2240;
assign w2242 = w1738 & ~w2241;
assign w2243 = (~w1052 & ~w2021) | (~w1052 & w6879) | (~w2021 & w6879);
assign w2244 = ~pi244 & w1478;
assign w2245 = ~w1283 & w6880;
assign w2246 = (pi244 & w1479) | (pi244 & w6881) | (w1479 & w6881);
assign w2247 = pi135 & w1331;
assign w2248 = ~w1286 & w6882;
assign w2249 = w1330 & w6883;
assign v567 = ~(w2244 | w2245);
assign w2250 = v567;
assign w2251 = ~w2247 & w6884;
assign w2252 = ~w2248 & w2251;
assign w2253 = (w1756 & ~w2252) | (w1756 & w6885) | (~w2252 & w6885);
assign w2254 = (w1047 & w6887) | (w1047 & w6888) | (w6887 & w6888);
assign w2255 = w1032 & w6889;
assign w2256 = (~w1732 & w1033) | (~w1732 & w6890) | (w1033 & w6890);
assign w2257 = ~w2255 & w2256;
assign w2258 = w1731 & ~w2224;
assign w2259 = ~w2225 & w2258;
assign w2260 = (w2253 & w6893) | (w2253 & w6894) | (w6893 & w6894);
assign v568 = ~(w2223 | w2260);
assign w2261 = v568;
assign w2262 = pi040 & w1728;
assign w2263 = w82 & w6895;
assign w2264 = ~pi040 & w1733;
assign w2265 = (w1047 & w6896) | (w1047 & w6897) | (w6896 & w6897);
assign w2266 = w1032 & w6898;
assign w2267 = (pi040 & ~w1032) | (pi040 & w6899) | (~w1032 & w6899);
assign w2268 = w1061 & w6900;
assign w2269 = pi078 & w1059;
assign w2270 = w1053 & w6901;
assign w2271 = pi065 & w1066;
assign w2272 = w1056 & w6902;
assign w2273 = pi074 & w1064;
assign w2274 = w1053 & w6903;
assign w2275 = pi077 & w1062;
assign v569 = ~(w2268 | w2269);
assign w2276 = v569;
assign v570 = ~(w2270 | w2271);
assign w2277 = v570;
assign v571 = ~(w2272 | w2273);
assign w2278 = v571;
assign v572 = ~(w2274 | w2275);
assign w2279 = v572;
assign w2280 = w2278 & w2279;
assign w2281 = w2276 & w2277;
assign w2282 = w2280 & w2281;
assign w2283 = w1052 & w2282;
assign w2284 = w1738 & ~w2283;
assign w2285 = ~w1283 & w6904;
assign w2286 = pi232 & w1336;
assign w2287 = ~w1286 & w6905;
assign v573 = ~(pi349 | w1346);
assign w2288 = v573;
assign w2289 = (~pi232 & ~w1767) | (~pi232 & w6906) | (~w1767 & w6906);
assign v574 = ~(w1769 | w2289);
assign w2290 = v574;
assign w2291 = w1346 & ~w2290;
assign v575 = ~(w2288 | w2291);
assign w2292 = v575;
assign w2293 = w1333 & w6907;
assign w2294 = w1330 & w6908;
assign w2295 = (~w2285 & ~w1331) | (~w2285 & w6909) | (~w1331 & w6909);
assign v576 = ~(w2293 | w2294);
assign w2296 = v576;
assign w2297 = w2295 & w2296;
assign v577 = ~(w2286 | w2287);
assign w2298 = v577;
assign w2299 = w2297 & w2298;
assign w2300 = (pi232 & w1086) | (pi232 & w6910) | (w1086 & w6910);
assign w2301 = w1087 & w6911;
assign v578 = ~(w1052 | w2300);
assign w2302 = v578;
assign w2303 = ~w2301 & w2302;
assign w2304 = (w2303 & w2299) | (w2303 & w6912) | (w2299 & w6912);
assign v579 = ~(w1732 | w2266);
assign w2305 = v579;
assign w2306 = ~w2267 & w2305;
assign w2307 = w1731 & ~w2263;
assign w2308 = ~w2264 & w2307;
assign w2309 = w2308 & w7383;
assign v580 = ~(w2262 | w2309);
assign w2310 = v580;
assign v581 = ~(pi242 | pi350);
assign w2311 = v581;
assign w2312 = w745 & w748;
assign w2313 = w711 & w6914;
assign v582 = ~(w2312 | w2313);
assign w2314 = v582;
assign w2315 = ~w687 & w6915;
assign w2316 = w736 & ~w777;
assign w2317 = (~pi275 & ~w24) | (~pi275 & w3634) | (~w24 & w3634);
assign w2318 = w24 & w6917;
assign w2319 = w1555 & ~w2317;
assign w2320 = (pi242 & ~w2319) | (pi242 & w6918) | (~w2319 & w6918);
assign w2321 = w2314 & w2320;
assign w2322 = ~w2316 & w2321;
assign w2323 = ~w2315 & w2322;
assign w2324 = w2323 & w7384;
assign v583 = ~(w1552 | w2311);
assign w2325 = v583;
assign w2326 = pi275 & w1552;
assign w2327 = (~w2326 & w2324) | (~w2326 & w6919) | (w2324 & w6919);
assign w2328 = ~pi253 & w165;
assign w2329 = (~w2328 & w2327) | (~w2328 & w6920) | (w2327 & w6920);
assign w2330 = (w2327 & w6921) | (w2327 & w6922) | (w6921 & w6922);
assign w2331 = w206 & w7385;
assign w2332 = pi041 & ~w206;
assign v584 = ~(w2331 | w2332);
assign w2333 = v584;
assign w2334 = w197 & w7385;
assign w2335 = pi042 & ~w197;
assign v585 = ~(w2334 | w2335);
assign w2336 = v585;
assign w2337 = pi043 & ~w204;
assign w2338 = w1523 & w6923;
assign w2339 = ~w1523 & w6924;
assign w2340 = w1523 & w6925;
assign w2341 = pi042 & w1524;
assign w2342 = pi046 & w1539;
assign w2343 = ~w1523 & w6926;
assign w2344 = ~w1523 & w6927;
assign w2345 = w1523 & w6928;
assign v586 = ~(w2338 | w2339);
assign w2346 = v586;
assign v587 = ~(w2340 | w2341);
assign w2347 = v587;
assign v588 = ~(w2342 | w2343);
assign w2348 = v588;
assign v589 = ~(w2344 | w2345);
assign w2349 = v589;
assign w2350 = w2348 & w2349;
assign w2351 = w2346 & w2347;
assign w2352 = w2350 & w2351;
assign w2353 = w162 & w2352;
assign w2354 = w204 & ~w2353;
assign w2355 = w2354 & w7385;
assign v590 = ~(w2337 | w2355);
assign w2356 = v590;
assign w2357 = w195 & w7385;
assign w2358 = pi044 & ~w195;
assign v591 = ~(w2357 | w2358);
assign w2359 = v591;
assign w2360 = w192 & w7385;
assign w2361 = pi045 & ~w192;
assign v592 = ~(w2360 | w2361);
assign w2362 = v592;
assign w2363 = w189 & w7385;
assign w2364 = pi046 & ~w189;
assign v593 = ~(w2363 | w2364);
assign w2365 = v593;
assign w2366 = pi047 & ~w202;
assign w2367 = w202 & ~w2353;
assign w2368 = w2367 & w7385;
assign v594 = ~(w2366 | w2368);
assign w2369 = v594;
assign v595 = ~(pi048 | w199);
assign w2370 = v595;
assign w2371 = w199 & w2329;
assign w2372 = (w2371 & w575) | (w2371 & w6929) | (w575 & w6929);
assign v596 = ~(w2370 | w2372);
assign w2373 = v596;
assign w2374 = ~w1523 & w6930;
assign w2375 = w1523 & w6931;
assign w2376 = ~pi055 & w1539;
assign w2377 = ~w1523 & w6932;
assign w2378 = w1523 & w6933;
assign w2379 = w1523 & w6934;
assign w2380 = ~pi050 & w1524;
assign w2381 = ~w1523 & w6935;
assign v597 = ~(w2374 | w2375);
assign w2382 = v597;
assign v598 = ~(w2376 | w2377);
assign w2383 = v598;
assign v599 = ~(w2378 | w2379);
assign w2384 = v599;
assign v600 = ~(w2380 | w2381);
assign w2385 = v600;
assign w2386 = w2384 & w2385;
assign w2387 = w2382 & w2383;
assign w2388 = w2386 & w2387;
assign w2389 = w162 & ~w2388;
assign v601 = ~(pi242 | pi353);
assign w2390 = v601;
assign w2391 = w711 & w6936;
assign w2392 = w736 & w791;
assign v602 = ~(w2391 | w2392);
assign w2393 = v602;
assign w2394 = (w2393 & w680) | (w2393 & w6937) | (w680 & w6937);
assign v603 = ~(pi243 | w916);
assign w2395 = v603;
assign w2396 = w711 & ~w715;
assign w2397 = w746 & ~w2396;
assign w2398 = (w735 & w746) | (w735 & w6938) | (w746 & w6938);
assign w2399 = (pi242 & w2397) | (pi242 & w6939) | (w2397 & w6939);
assign w2400 = w2394 & w2399;
assign v604 = ~(w1552 | w2390);
assign w2401 = v604;
assign w2402 = w2401 & w7386;
assign w2403 = pi273 & w1552;
assign v605 = ~(w2402 | w2403);
assign w2404 = v605;
assign w2405 = ~pi236 & w165;
assign w2406 = (w2402 & w6944) | (w2402 & w6945) | (w6944 & w6945);
assign v606 = ~(w2389 | w2406);
assign w2407 = v606;
assign w2408 = (w545 & w6946) | (w545 & w6947) | (w6946 & w6947);
assign w2409 = (~pi049 & ~w206) | (~pi049 & w6948) | (~w206 & w6948);
assign v607 = ~(w2408 | w2409);
assign w2410 = v607;
assign w2411 = (w545 & w6949) | (w545 & w6950) | (w6949 & w6950);
assign w2412 = (~pi050 & ~w197) | (~pi050 & w6951) | (~w197 & w6951);
assign v608 = ~(w2411 | w2412);
assign w2413 = v608;
assign w2414 = (w545 & w6952) | (w545 & w6953) | (w6952 & w6953);
assign w2415 = (~pi051 & ~w204) | (~pi051 & w6954) | (~w204 & w6954);
assign v609 = ~(w2414 | w2415);
assign w2416 = v609;
assign w2417 = (w545 & w6955) | (w545 & w6956) | (w6955 & w6956);
assign w2418 = (~pi052 & ~w195) | (~pi052 & w6957) | (~w195 & w6957);
assign v610 = ~(w2417 | w2418);
assign w2419 = v610;
assign w2420 = (w545 & w6958) | (w545 & w6959) | (w6958 & w6959);
assign w2421 = (~pi053 & ~w192) | (~pi053 & w6960) | (~w192 & w6960);
assign v611 = ~(w2420 | w2421);
assign w2422 = v611;
assign w2423 = (w545 & w6961) | (w545 & w6962) | (w6961 & w6962);
assign w2424 = (~pi054 & ~w199) | (~pi054 & w6963) | (~w199 & w6963);
assign v612 = ~(w2423 | w2424);
assign w2425 = v612;
assign w2426 = (w545 & w6964) | (w545 & w6965) | (w6964 & w6965);
assign w2427 = (~pi055 & ~w189) | (~pi055 & w6966) | (~w189 & w6966);
assign v613 = ~(w2426 | w2427);
assign w2428 = v613;
assign w2429 = (w545 & w6967) | (w545 & w6968) | (w6967 & w6968);
assign v614 = ~(pi056 | w1597);
assign w2430 = v614;
assign v615 = ~(w2429 | w2430);
assign w2431 = v615;
assign w2432 = w1523 & w6969;
assign w2433 = ~w1523 & w6970;
assign w2434 = ~w1523 & w6971;
assign w2435 = w1523 & w6972;
assign w2436 = ~pi062 & w1539;
assign w2437 = w1523 & w6973;
assign w2438 = ~pi058 & w1524;
assign w2439 = ~w1523 & w6974;
assign v616 = ~(w2432 | w2433);
assign w2440 = v616;
assign v617 = ~(w2434 | w2435);
assign w2441 = v617;
assign v618 = ~(w2436 | w2437);
assign w2442 = v618;
assign v619 = ~(w2438 | w2439);
assign w2443 = v619;
assign w2444 = w2442 & w2443;
assign w2445 = w2440 & w2441;
assign w2446 = w2444 & w2445;
assign w2447 = w2444 & w6975;
assign w2448 = ~pi245 & w165;
assign v620 = ~(pi242 | pi348);
assign w2449 = v620;
assign w2450 = pi303 & w16;
assign w2451 = (~pi272 & ~w16) | (~pi272 & w6976) | (~w16 & w6976);
assign w2452 = w16 & w6917;
assign w2453 = w1555 & ~w2451;
assign w2454 = ~w2452 & w2453;
assign w2455 = w713 & w719;
assign w2456 = w736 & ~w797;
assign w2457 = w697 & w701;
assign v621 = ~(w2455 | w2456);
assign w2458 = v621;
assign w2459 = ~w2457 & w2458;
assign v622 = ~(pi243 | w926);
assign w2460 = v622;
assign w2461 = w743 & w745;
assign v623 = ~(w2454 | w2461);
assign w2462 = v623;
assign w2463 = ~w2457 & w6977;
assign w2464 = (w2463 & w926) | (w2463 & w6978) | (w926 & w6978);
assign w2465 = ~w2449 & w7387;
assign w2466 = ~pi272 & w1552;
assign w2467 = (~w2466 & w2465) | (~w2466 & w6981) | (w2465 & w6981);
assign w2468 = (~w162 & ~w2467) | (~w162 & w6982) | (~w2467 & w6982);
assign w2469 = ~w2448 & w2468;
assign w2470 = (w585 & w6983) | (w585 & w6984) | (w6983 & w6984);
assign w2471 = w1517 & ~w2470;
assign w2472 = (pi057 & ~w206) | (pi057 & w6985) | (~w206 & w6985);
assign v624 = ~(w2471 | w2472);
assign w2473 = v624;
assign w2474 = w1577 & ~w2470;
assign w2475 = (pi058 & ~w197) | (pi058 & w6986) | (~w197 & w6986);
assign v625 = ~(w2474 | w2475);
assign w2476 = v625;
assign w2477 = w1581 & ~w2470;
assign w2478 = (pi059 & ~w204) | (pi059 & w6987) | (~w204 & w6987);
assign v626 = ~(w2477 | w2478);
assign w2479 = v626;
assign w2480 = w1585 & ~w2470;
assign w2481 = (pi060 & ~w195) | (pi060 & w6988) | (~w195 & w6988);
assign v627 = ~(w2480 | w2481);
assign w2482 = v627;
assign w2483 = w1589 & ~w2470;
assign w2484 = (pi061 & ~w192) | (pi061 & w6989) | (~w192 & w6989);
assign v628 = ~(w2483 | w2484);
assign w2485 = v628;
assign w2486 = w1593 & ~w2470;
assign w2487 = (pi062 & ~w189) | (pi062 & w6990) | (~w189 & w6990);
assign v629 = ~(w2486 | w2487);
assign w2488 = v629;
assign w2489 = w1597 & ~w2470;
assign w2490 = (pi063 & ~w202) | (pi063 & w6991) | (~w202 & w6991);
assign v630 = ~(w2489 | w2490);
assign w2491 = v630;
assign w2492 = w1601 & ~w2470;
assign w2493 = (pi064 & ~w199) | (pi064 & w6992) | (~w199 & w6992);
assign v631 = ~(w2492 | w2493);
assign w2494 = v631;
assign w2495 = pi065 & w1539;
assign w2496 = w1523 & w6993;
assign w2497 = ~w1523 & w6994;
assign w2498 = ~w1523 & w6995;
assign w2499 = ~w1523 & w6996;
assign w2500 = w1523 & w6997;
assign w2501 = pi075 & w1524;
assign w2502 = w1523 & w6998;
assign v632 = ~(w2495 | w2496);
assign w2503 = v632;
assign v633 = ~(w2497 | w2498);
assign w2504 = v633;
assign v634 = ~(w2499 | w2500);
assign w2505 = v634;
assign v635 = ~(w2501 | w2502);
assign w2506 = v635;
assign w2507 = w2505 & w2506;
assign w2508 = w2503 & w2504;
assign w2509 = w2507 & w2508;
assign w2510 = w162 & w2509;
assign w2511 = w713 & w716;
assign w2512 = (~pi271 & ~w22) | (~pi271 & w6999) | (~w22 & w6999);
assign w2513 = w22 & w6602;
assign w2514 = w1555 & ~w2512;
assign w2515 = ~w2513 & w2514;
assign w2516 = w745 & w750;
assign w2517 = w736 & ~w786;
assign w2518 = w701 & ~w704;
assign v636 = ~(w2516 | w2517);
assign w2519 = v636;
assign w2520 = ~w2511 & w2519;
assign w2521 = ~w2515 & w2520;
assign w2522 = ~w2518 & w2521;
assign w2523 = (w2522 & w937) | (w2522 & w7000) | (w937 & w7000);
assign w2524 = ~pi242 & pi349;
assign w2525 = (~w2524 & w2523) | (~w2524 & w7001) | (w2523 & w7001);
assign w2526 = pi271 & w1552;
assign w2527 = (~w2526 & w2525) | (~w2526 & w7002) | (w2525 & w7002);
assign w2528 = ~pi255 & w165;
assign v637 = ~(w162 | w2528);
assign w2529 = v637;
assign w2530 = (w2529 & w2527) | (w2529 & w7003) | (w2527 & w7003);
assign v638 = ~(w2510 | w2530);
assign w2531 = v638;
assign w2532 = (~w2531 & ~w540) | (~w2531 & w7004) | (~w540 & w7004);
assign w2533 = w1593 & ~w2532;
assign w2534 = (pi065 & ~w189) | (pi065 & w7005) | (~w189 & w7005);
assign v639 = ~(w2533 | w2534);
assign w2535 = v639;
assign w2536 = w1507 & w7006;
assign w2537 = ~w1515 & w7007;
assign v640 = ~(pi247 | w2537);
assign w2538 = v640;
assign w2539 = w206 & w2538;
assign w2540 = w1523 & w7008;
assign w2541 = ~w1523 & w7009;
assign w2542 = pi069 & w1539;
assign w2543 = pi067 & w1524;
assign w2544 = w1523 & w7010;
assign w2545 = ~w1523 & w7011;
assign w2546 = w1523 & w7012;
assign w2547 = ~w1523 & w7013;
assign v641 = ~(w2540 | w2541);
assign w2548 = v641;
assign v642 = ~(w2542 | w2543);
assign w2549 = v642;
assign v643 = ~(w2544 | w2545);
assign w2550 = v643;
assign v644 = ~(w2546 | w2547);
assign w2551 = v644;
assign w2552 = w2550 & w2551;
assign w2553 = w2548 & w2549;
assign w2554 = w2552 & w2553;
assign w2555 = w2553 & w7014;
assign w2556 = ~pi263 & w165;
assign w2557 = w516 & w1511;
assign v645 = ~(w162 | w2556);
assign w2558 = v645;
assign w2559 = (w2558 & w1570) | (w2558 & w7015) | (w1570 & w7015);
assign w2560 = (~w2555 & w2557) | (~w2555 & w7016) | (w2557 & w7016);
assign w2561 = w2539 & ~w2560;
assign w2562 = (~pi066 & ~w206) | (~pi066 & w7017) | (~w206 & w7017);
assign v646 = ~(w2561 | w2562);
assign w2563 = v646;
assign w2564 = w197 & w2538;
assign w2565 = w2564 & ~w2560;
assign w2566 = (~pi067 & ~w197) | (~pi067 & w7018) | (~w197 & w7018);
assign v647 = ~(w2565 | w2566);
assign w2567 = v647;
assign w2568 = w204 & w2538;
assign w2569 = w2568 & ~w2560;
assign w2570 = (~pi068 & ~w204) | (~pi068 & w7019) | (~w204 & w7019);
assign v648 = ~(w2569 | w2570);
assign w2571 = v648;
assign w2572 = w189 & w2538;
assign w2573 = w2572 & ~w2560;
assign w2574 = (~pi069 & ~w189) | (~pi069 & w7020) | (~w189 & w7020);
assign v649 = ~(w2573 | w2574);
assign w2575 = v649;
assign w2576 = w202 & w2538;
assign w2577 = w2576 & ~w2560;
assign w2578 = (~pi070 & ~w202) | (~pi070 & w7021) | (~w202 & w7021);
assign v650 = ~(w2577 | w2578);
assign w2579 = v650;
assign w2580 = w199 & w2538;
assign w2581 = w2580 & ~w2560;
assign w2582 = (~pi071 & ~w199) | (~pi071 & w7022) | (~w199 & w7022);
assign v651 = ~(w2581 | w2582);
assign w2583 = v651;
assign w2584 = w195 & w2538;
assign w2585 = w2584 & ~w2560;
assign w2586 = (~pi072 & ~w195) | (~pi072 & w7023) | (~w195 & w7023);
assign v652 = ~(w2585 | w2586);
assign w2587 = v652;
assign w2588 = w192 & w2538;
assign w2589 = w2588 & ~w2560;
assign w2590 = (~pi073 & ~w192) | (~pi073 & w7024) | (~w192 & w7024);
assign v653 = ~(w2589 | w2590);
assign w2591 = v653;
assign w2592 = (w540 & w7025) | (w540 & w7026) | (w7025 & w7026);
assign w2593 = (pi074 & ~w206) | (pi074 & w7027) | (~w206 & w7027);
assign v654 = ~(w2592 | w2593);
assign w2594 = v654;
assign w2595 = (w540 & w7028) | (w540 & w7029) | (w7028 & w7029);
assign w2596 = (pi075 & ~w197) | (pi075 & w7030) | (~w197 & w7030);
assign v655 = ~(w2595 | w2596);
assign w2597 = v655;
assign w2598 = (w540 & w7031) | (w540 & w7032) | (w7031 & w7032);
assign w2599 = (pi076 & ~w204) | (pi076 & w7033) | (~w204 & w7033);
assign v656 = ~(w2598 | w2599);
assign w2600 = v656;
assign w2601 = (w540 & w7034) | (w540 & w7035) | (w7034 & w7035);
assign w2602 = (pi077 & ~w195) | (pi077 & w7036) | (~w195 & w7036);
assign v657 = ~(w2601 | w2602);
assign w2603 = v657;
assign w2604 = (w540 & w7037) | (w540 & w7038) | (w7037 & w7038);
assign w2605 = (pi078 & ~w192) | (pi078 & w7039) | (~w192 & w7039);
assign v658 = ~(w2604 | w2605);
assign w2606 = v658;
assign w2607 = (w540 & w7040) | (w540 & w7041) | (w7040 & w7041);
assign w2608 = (pi079 & ~w202) | (pi079 & w7042) | (~w202 & w7042);
assign v659 = ~(w2607 | w2608);
assign w2609 = v659;
assign w2610 = (w540 & w7043) | (w540 & w7044) | (w7043 & w7044);
assign w2611 = (pi080 & ~w199) | (pi080 & w7045) | (~w199 & w7045);
assign v660 = ~(w2610 | w2611);
assign w2612 = v660;
assign w2613 = ~w1523 & w7046;
assign w2614 = pi091 & w1524;
assign w2615 = ~w1523 & w7047;
assign w2616 = w1523 & w7048;
assign w2617 = pi094 & w1539;
assign w2618 = ~w1523 & w7049;
assign w2619 = w1523 & w7050;
assign w2620 = w1523 & w7051;
assign v661 = ~(w2613 | w2614);
assign w2621 = v661;
assign v662 = ~(w2615 | w2616);
assign w2622 = v662;
assign v663 = ~(w2617 | w2618);
assign w2623 = v663;
assign v664 = ~(w2619 | w2620);
assign w2624 = v664;
assign w2625 = w2623 & w2624;
assign w2626 = w2621 & w2622;
assign w2627 = w2625 & w2626;
assign w2628 = w162 & w2627;
assign w2629 = ~pi258 & w165;
assign v665 = ~(pi242 | pi354);
assign w2630 = v665;
assign w2631 = w745 & w753;
assign w2632 = (w736 & ~w781) | (w736 & w7052) | (~w781 & w7052);
assign w2633 = pi197 & w701;
assign w2634 = w713 & w723;
assign v666 = ~(pi243 | w829);
assign w2635 = v666;
assign w2636 = (~pi264 & ~w751) | (~pi264 & w7053) | (~w751 & w7053);
assign w2637 = w751 & w7054;
assign w2638 = w1555 & ~w2636;
assign w2639 = ~w2637 & w2638;
assign w2640 = pi242 & ~w2631;
assign w2641 = ~w2633 & w2640;
assign v667 = ~(w2632 | w2634);
assign w2642 = v667;
assign w2643 = ~w2639 & w2642;
assign w2644 = w2641 & w2643;
assign v668 = ~(w1552 | w2630);
assign w2645 = v668;
assign w2646 = (w2645 & w2635) | (w2645 & w7055) | (w2635 & w7055);
assign w2647 = pi264 & w1552;
assign v669 = ~(w2646 | w2647);
assign w2648 = v669;
assign w2649 = w1551 & ~w2648;
assign v670 = ~(w162 | w2649);
assign w2650 = v670;
assign w2651 = ~w2649 & w7056;
assign w2652 = (w2651 & ~w529) | (w2651 & w7057) | (~w529 & w7057);
assign w2653 = (w1589 & w2652) | (w1589 & w7058) | (w2652 & w7058);
assign w2654 = (~pi081 & ~w192) | (~pi081 & w7059) | (~w192 & w7059);
assign v671 = ~(w2653 | w2654);
assign w2655 = v671;
assign w2656 = w589 & w1511;
assign w2657 = ~pi254 & w165;
assign w2658 = (~w2657 & w2327) | (~w2657 & w7060) | (w2327 & w7060);
assign w2659 = w1523 & w7061;
assign w2660 = ~w1523 & w7062;
assign w2661 = pi084 & w1524;
assign w2662 = pi088 & w1539;
assign w2663 = ~w1523 & w7063;
assign w2664 = w1523 & w7064;
assign w2665 = ~w1523 & w7065;
assign w2666 = w1523 & w7066;
assign v672 = ~(w2659 | w2660);
assign w2667 = v672;
assign v673 = ~(w2661 | w2662);
assign w2668 = v673;
assign v674 = ~(w2663 | w2664);
assign w2669 = v674;
assign v675 = ~(w2665 | w2666);
assign w2670 = v675;
assign w2671 = w2669 & w2670;
assign w2672 = w2667 & w2668;
assign w2673 = w2671 & w2672;
assign w2674 = (w162 & ~w2672) | (w162 & w7067) | (~w2672 & w7067);
assign w2675 = (~w2674 & w2658) | (~w2674 & w7068) | (w2658 & w7068);
assign w2676 = (w2580 & w2656) | (w2580 & w7069) | (w2656 & w7069);
assign w2677 = (pi082 & ~w199) | (pi082 & w7070) | (~w199 & w7070);
assign v676 = ~(w2676 | w2677);
assign w2678 = v676;
assign w2679 = (w2539 & w2656) | (w2539 & w7071) | (w2656 & w7071);
assign w2680 = (pi083 & ~w206) | (pi083 & w7072) | (~w206 & w7072);
assign v677 = ~(w2679 | w2680);
assign w2681 = v677;
assign w2682 = (w2564 & w2656) | (w2564 & w7073) | (w2656 & w7073);
assign w2683 = (pi084 & ~w197) | (pi084 & w7074) | (~w197 & w7074);
assign v678 = ~(w2682 | w2683);
assign w2684 = v678;
assign w2685 = (w2568 & w2656) | (w2568 & w7075) | (w2656 & w7075);
assign w2686 = (pi085 & ~w204) | (pi085 & w7076) | (~w204 & w7076);
assign v679 = ~(w2685 | w2686);
assign w2687 = v679;
assign w2688 = (w2584 & w2656) | (w2584 & w7077) | (w2656 & w7077);
assign w2689 = (pi086 & ~w195) | (pi086 & w7078) | (~w195 & w7078);
assign v680 = ~(w2688 | w2689);
assign w2690 = v680;
assign w2691 = (w2588 & w2656) | (w2588 & w7079) | (w2656 & w7079);
assign w2692 = (pi087 & ~w192) | (pi087 & w7080) | (~w192 & w7080);
assign v681 = ~(w2691 | w2692);
assign w2693 = v681;
assign w2694 = (w2572 & w2656) | (w2572 & w7081) | (w2656 & w7081);
assign w2695 = (pi088 & ~w189) | (pi088 & w7082) | (~w189 & w7082);
assign v682 = ~(w2694 | w2695);
assign w2696 = v682;
assign w2697 = (w2576 & w2656) | (w2576 & w7083) | (w2656 & w7083);
assign w2698 = pi089 & ~w2576;
assign v683 = ~(w2697 | w2698);
assign w2699 = v683;
assign w2700 = (pi090 & ~w206) | (pi090 & w7084) | (~w206 & w7084);
assign w2701 = ~w2652 & w7085;
assign v684 = ~(w2700 | w2701);
assign w2702 = v684;
assign w2703 = (w1577 & w2652) | (w1577 & w7086) | (w2652 & w7086);
assign w2704 = (~pi091 & ~w197) | (~pi091 & w7087) | (~w197 & w7087);
assign v685 = ~(w2703 | w2704);
assign w2705 = v685;
assign w2706 = (w1581 & w2652) | (w1581 & w7088) | (w2652 & w7088);
assign w2707 = (~pi092 & ~w204) | (~pi092 & w7089) | (~w204 & w7089);
assign v686 = ~(w2706 | w2707);
assign w2708 = v686;
assign w2709 = (w1585 & w2652) | (w1585 & w7090) | (w2652 & w7090);
assign w2710 = (~pi093 & ~w195) | (~pi093 & w7091) | (~w195 & w7091);
assign v687 = ~(w2709 | w2710);
assign w2711 = v687;
assign w2712 = (w1593 & w2652) | (w1593 & w7092) | (w2652 & w7092);
assign w2713 = (~pi094 & ~w189) | (~pi094 & w7093) | (~w189 & w7093);
assign v688 = ~(w2712 | w2713);
assign w2714 = v688;
assign w2715 = (w1597 & w2652) | (w1597 & w7094) | (w2652 & w7094);
assign w2716 = (~pi095 & ~w202) | (~pi095 & w7095) | (~w202 & w7095);
assign v689 = ~(w2715 | w2716);
assign w2717 = v689;
assign w2718 = (w1601 & w2652) | (w1601 & w7096) | (w2652 & w7096);
assign v690 = ~(pi096 | w1601);
assign w2719 = v690;
assign v691 = ~(w2718 | w2719);
assign w2720 = v691;
assign w2721 = w1032 & w7097;
assign w2722 = ~w38 & w82;
assign w2723 = w82 & w7098;
assign w2724 = w130 & w1018;
assign w2725 = w85 & w1040;
assign w2726 = w8 & w7099;
assign w2727 = (w2726 & w2725) | (w2726 & w7100) | (w2725 & w7100);
assign w2728 = w1082 & ~w1190;
assign v692 = ~(w2724 | w2727);
assign w2729 = v692;
assign w2730 = ~w2728 & w2729;
assign w2731 = (~w2723 & w2730) | (~w2723 & w7101) | (w2730 & w7101);
assign w2732 = ~pi361 & w141;
assign w2733 = pi247 & pi356;
assign w2734 = (~w2733 & ~w141) | (~w2733 & w7102) | (~w141 & w7102);
assign w2735 = (w2734 & ~w1032) | (w2734 & w7103) | (~w1032 & w7103);
assign w2736 = w2735 & w7104;
assign w2737 = (~pi097 & ~w2735) | (~pi097 & w7105) | (~w2735 & w7105);
assign v693 = ~(w2736 | w2737);
assign w2738 = v693;
assign v694 = ~(w2721 | w2738);
assign w2739 = v694;
assign w2740 = pi359 & ~w2739;
assign w2741 = (w2730 & w7106) | (w2730 & w7107) | (w7106 & w7107);
assign w2742 = w2735 & w2741;
assign w2743 = (~pi098 & ~w2735) | (~pi098 & w7108) | (~w2735 & w7108);
assign w2744 = pi359 & ~w2721;
assign w2745 = ~w2742 & w2744;
assign w2746 = ~w2743 & w2745;
assign w2747 = (~w2741 & w2735) | (~w2741 & w7110) | (w2735 & w7110);
assign w2748 = pi356 & w1033;
assign w2749 = (~w2733 & ~w1033) | (~w2733 & w7111) | (~w1033 & w7111);
assign w2750 = pi099 & w2749;
assign w2751 = ~w2747 & w2750;
assign w2752 = (w2735 & w7112) | (w2735 & w7113) | (w7112 & w7113);
assign w2753 = ~w2751 & w2752;
assign w2754 = ~w1523 & w7114;
assign w2755 = ~w1523 & w7115;
assign w2756 = w1523 & w7116;
assign w2757 = ~w1523 & w7117;
assign w2758 = w1523 & w7118;
assign w2759 = w1523 & w7119;
assign w2760 = pi111 & w1524;
assign w2761 = pi116 & w1539;
assign v695 = ~(w2754 | w2755);
assign w2762 = v695;
assign v696 = ~(w2756 | w2757);
assign w2763 = v696;
assign v697 = ~(w2758 | w2759);
assign w2764 = v697;
assign v698 = ~(w2760 | w2761);
assign w2765 = v698;
assign w2766 = w2764 & w2765;
assign w2767 = w2762 & w2763;
assign w2768 = w2766 & w2767;
assign w2769 = w2766 & w7120;
assign w2770 = ~pi266 & w165;
assign w2771 = w596 & w1511;
assign v699 = ~(w162 | w2770);
assign w2772 = v699;
assign w2773 = (w2772 & w1620) | (w2772 & w7121) | (w1620 & w7121);
assign w2774 = (~w2769 & w2771) | (~w2769 & w7122) | (w2771 & w7122);
assign w2775 = w2588 & ~w2774;
assign w2776 = (~pi100 & ~w192) | (~pi100 & w7123) | (~w192 & w7123);
assign v700 = ~(w2775 | w2776);
assign w2777 = v700;
assign w2778 = ~w1523 & w7124;
assign w2779 = w1523 & w7125;
assign w2780 = pi107 & w1539;
assign w2781 = ~w1523 & w7126;
assign w2782 = ~w1523 & w7127;
assign w2783 = w1523 & w7128;
assign w2784 = pi103 & w1524;
assign w2785 = w1523 & w7129;
assign v701 = ~(w2778 | w2779);
assign w2786 = v701;
assign v702 = ~(w2780 | w2781);
assign w2787 = v702;
assign v703 = ~(w2782 | w2783);
assign w2788 = v703;
assign v704 = ~(w2784 | w2785);
assign w2789 = v704;
assign w2790 = w2788 & w2789;
assign w2791 = w2786 & w2787;
assign w2792 = w2790 & w2791;
assign w2793 = w162 & w2792;
assign w2794 = ~pi262 & w165;
assign w2795 = ~w600 & w1511;
assign v705 = ~(w162 | w2794);
assign w2796 = v705;
assign w2797 = w2796 & w7388;
assign w2798 = (~w2793 & w2795) | (~w2793 & w7130) | (w2795 & w7130);
assign w2799 = w2539 & ~w2798;
assign w2800 = (~pi101 & ~w206) | (~pi101 & w7131) | (~w206 & w7131);
assign v706 = ~(w2799 | w2800);
assign w2801 = v706;
assign w2802 = ~pi231 & pi234;
assign w2803 = ~pi251 & w2802;
assign w2804 = w2802 & w7132;
assign w2805 = w1507 & w7133;
assign w2806 = ~w1695 & w7134;
assign w2807 = w86 & w130;
assign w2808 = w86 & w7135;
assign w2809 = pi242 & ~w619;
assign w2810 = (~w745 & w619) | (~w745 & w7136) | (w619 & w7136);
assign w2811 = ~pi102 & pi344;
assign w2812 = (w887 & w7137) | (w887 & w7138) | (w7137 & w7138);
assign w2813 = ~w840 & w7389;
assign v707 = ~(w827 | w2812);
assign w2814 = v707;
assign w2815 = (~w926 & w915) | (~w926 & w7139) | (w915 & w7139);
assign v708 = ~(w927 | w2815);
assign w2816 = v708;
assign w2817 = (~w937 & w947) | (~w937 & w7140) | (w947 & w7140);
assign v709 = ~(w948 | w2817);
assign w2818 = v709;
assign w2819 = w2816 & ~w2818;
assign w2820 = ~w2816 & w2818;
assign v710 = ~(w2819 | w2820);
assign w2821 = v710;
assign w2822 = (~w959 & w968) | (~w959 & w7141) | (w968 & w7141);
assign v711 = ~(w969 | w2822);
assign w2823 = v711;
assign w2824 = ~w829 & w2823;
assign w2825 = w829 & ~w2823;
assign v712 = ~(w2824 | w2825);
assign w2826 = v712;
assign w2827 = ~w903 & w2826;
assign w2828 = w903 & ~w2826;
assign v713 = ~(w2827 | w2828);
assign w2829 = v713;
assign w2830 = w2821 & w2829;
assign v714 = ~(w2821 | w2829);
assign w2831 = v714;
assign w2832 = w827 & ~w2830;
assign w2833 = ~w2831 & w2832;
assign w2834 = (~pi344 & ~w2814) | (~pi344 & w7142) | (~w2814 & w7142);
assign v715 = ~(pi243 | w2811);
assign w2835 = v715;
assign v716 = ~(w786 | w800);
assign w2836 = v716;
assign v717 = ~(w801 | w2836);
assign w2837 = v717;
assign w2838 = w767 & ~w770;
assign v718 = ~(w771 | w2838);
assign w2839 = v718;
assign v719 = ~(w777 | w782);
assign w2840 = v719;
assign v720 = ~(w783 | w2840);
assign w2841 = v720;
assign w2842 = w2839 & ~w2841;
assign w2843 = ~w2839 & w2841;
assign v721 = ~(w2842 | w2843);
assign w2844 = v721;
assign v722 = ~(w2837 | w2844);
assign w2845 = v722;
assign w2846 = w2837 & w2844;
assign w2847 = w802 & ~w2845;
assign w2848 = ~w2846 & w2847;
assign w2849 = (pi102 & w737) | (pi102 & w7144) | (w737 & w7144);
assign w2850 = pi223 & w723;
assign v723 = ~(w724 | w2850);
assign w2851 = v723;
assign w2852 = pi216 & w727;
assign v724 = ~(w728 | w2852);
assign w2853 = v724;
assign w2854 = w2851 & ~w2853;
assign w2855 = ~w2851 & w2853;
assign v725 = ~(w2854 | w2855);
assign w2856 = v725;
assign w2857 = w716 & w719;
assign v726 = ~(w720 | w2857);
assign w2858 = v726;
assign w2859 = w635 & ~w2858;
assign w2860 = ~w635 & w2858;
assign v727 = ~(w2859 | w2860);
assign w2861 = v727;
assign w2862 = w2856 & ~w2861;
assign w2863 = ~w2856 & w2861;
assign w2864 = w713 & ~w2862;
assign w2865 = ~w687 & w7145;
assign v728 = ~(w698 | w2865);
assign w2866 = v728;
assign w2867 = ~w704 & w2866;
assign w2868 = w704 & ~w2866;
assign v729 = ~(w2867 | w2868);
assign w2869 = v729;
assign w2870 = ~w651 & w7146;
assign v730 = ~(w659 | w2870);
assign w2871 = v730;
assign w2872 = w667 & ~w673;
assign v731 = ~(w674 | w2872);
assign w2873 = v731;
assign w2874 = (w681 & w7147) | (w681 & w7148) | (w7147 & w7148);
assign w2875 = w677 & ~w2874;
assign w2876 = w680 & w2874;
assign w2877 = (w2873 & w2876) | (w2873 & w7149) | (w2876 & w7149);
assign w2878 = ~w2876 & w7150;
assign v732 = ~(w2877 | w2878);
assign w2879 = v732;
assign w2880 = w2871 & w2879;
assign v733 = ~(w2871 | w2879);
assign w2881 = v733;
assign v734 = ~(w2880 | w2881);
assign w2882 = v734;
assign w2883 = w2869 & w2882;
assign w2884 = (w701 & w2882) | (w701 & w7151) | (w2882 & w7151);
assign w2885 = ~w2883 & w2884;
assign w2886 = (~w2849 & ~w763) | (~w2849 & w7152) | (~w763 & w7152);
assign w2887 = (w2886 & ~w2864) | (w2886 & w7153) | (~w2864 & w7153);
assign w2888 = ~w2848 & w2887;
assign w2889 = ~w2885 & w2888;
assign w2890 = w2889 & w7390;
assign w2891 = w1234 & w2726;
assign w2892 = w1032 & w7154;
assign w2893 = pi301 & w1015;
assign w2894 = w1015 & w7155;
assign w2895 = w1015 & w7156;
assign w2896 = w147 & w1014;
assign w2897 = w2893 & w2896;
assign w2898 = ~w2895 & w2897;
assign w2899 = w2897 & w7157;
assign w2900 = w159 & w1145;
assign w2901 = ~w1732 & w2900;
assign w2902 = pi323 & w2901;
assign w2903 = pi102 & ~w2901;
assign v735 = ~(w2898 | w2902);
assign w2904 = v735;
assign w2905 = w2810 & ~w2899;
assign w2906 = (w2905 & ~w2904) | (w2905 & w7158) | (~w2904 & w7158);
assign v736 = ~(w2892 | w2906);
assign w2907 = v736;
assign w2908 = (w2907 & w2890) | (w2907 & w7159) | (w2890 & w7159);
assign v737 = ~(pi351 | pi352);
assign w2909 = v737;
assign w2910 = pi351 & pi352;
assign v738 = ~(w2909 | w2910);
assign w2911 = v738;
assign v739 = ~(pi347 | pi349);
assign w2912 = v739;
assign w2913 = pi347 & pi349;
assign v740 = ~(w2912 | w2913);
assign w2914 = v740;
assign w2915 = w2911 & ~w2914;
assign w2916 = ~w2911 & w2914;
assign v741 = ~(w2915 | w2916);
assign w2917 = v741;
assign v742 = ~(pi353 | pi354);
assign w2918 = v742;
assign w2919 = pi353 & pi354;
assign v743 = ~(w2918 | w2919);
assign w2920 = v743;
assign v744 = ~(pi348 | pi350);
assign w2921 = v744;
assign w2922 = pi348 & pi350;
assign v745 = ~(w2921 | w2922);
assign w2923 = v745;
assign w2924 = w2920 & ~w2923;
assign w2925 = ~w2920 & w2923;
assign v746 = ~(w2924 | w2925);
assign w2926 = v746;
assign w2927 = w2917 & w2926;
assign v747 = ~(w2917 | w2926);
assign w2928 = v747;
assign v748 = ~(w2927 | w2928);
assign w2929 = v748;
assign w2930 = (~w2807 & ~w2892) | (~w2807 & w7160) | (~w2892 & w7160);
assign v749 = ~(w2805 | w2808);
assign w2931 = v749;
assign v750 = ~(pi247 | w2806);
assign w2932 = v750;
assign w2933 = w2932 & w7391;
assign w2934 = pi102 & pi247;
assign w2935 = pi359 & ~w2934;
assign w2936 = ~w2933 & w2935;
assign w2937 = w2564 & ~w2798;
assign w2938 = (~pi103 & ~w197) | (~pi103 & w7162) | (~w197 & w7162);
assign v751 = ~(w2937 | w2938);
assign w2939 = v751;
assign w2940 = w2568 & ~w2798;
assign w2941 = (~pi104 & ~w204) | (~pi104 & w7163) | (~w204 & w7163);
assign v752 = ~(w2940 | w2941);
assign w2942 = v752;
assign w2943 = w2584 & ~w2798;
assign w2944 = (~pi105 & ~w195) | (~pi105 & w7164) | (~w195 & w7164);
assign v753 = ~(w2943 | w2944);
assign w2945 = v753;
assign w2946 = w2588 & ~w2798;
assign w2947 = (~pi106 & ~w192) | (~pi106 & w7165) | (~w192 & w7165);
assign v754 = ~(w2946 | w2947);
assign w2948 = v754;
assign w2949 = w2572 & ~w2798;
assign w2950 = (~pi107 & ~w189) | (~pi107 & w7166) | (~w189 & w7166);
assign v755 = ~(w2949 | w2950);
assign w2951 = v755;
assign w2952 = w2576 & ~w2798;
assign w2953 = (~pi108 & ~w202) | (~pi108 & w7167) | (~w202 & w7167);
assign v756 = ~(w2952 | w2953);
assign w2954 = v756;
assign w2955 = w2580 & ~w2798;
assign w2956 = (~pi109 & ~w199) | (~pi109 & w7168) | (~w199 & w7168);
assign v757 = ~(w2955 | w2956);
assign w2957 = v757;
assign w2958 = w2539 & ~w2774;
assign w2959 = (~pi110 & ~w206) | (~pi110 & w7169) | (~w206 & w7169);
assign v758 = ~(w2958 | w2959);
assign w2960 = v758;
assign w2961 = w2564 & ~w2774;
assign w2962 = (~pi111 & ~w197) | (~pi111 & w7170) | (~w197 & w7170);
assign v759 = ~(w2961 | w2962);
assign w2963 = v759;
assign w2964 = w2568 & ~w2774;
assign w2965 = (~pi112 & ~w204) | (~pi112 & w7171) | (~w204 & w7171);
assign v760 = ~(w2964 | w2965);
assign w2966 = v760;
assign w2967 = w2584 & ~w2774;
assign w2968 = (~pi113 & ~w195) | (~pi113 & w7172) | (~w195 & w7172);
assign v761 = ~(w2967 | w2968);
assign w2969 = v761;
assign w2970 = w2576 & ~w2774;
assign w2971 = (~pi114 & ~w202) | (~pi114 & w7173) | (~w202 & w7173);
assign v762 = ~(w2970 | w2971);
assign w2972 = v762;
assign w2973 = w2580 & ~w2774;
assign w2974 = (~pi115 & ~w199) | (~pi115 & w7174) | (~w199 & w7174);
assign v763 = ~(w2973 | w2974);
assign w2975 = v763;
assign w2976 = w2572 & ~w2774;
assign w2977 = (~pi116 & ~w189) | (~pi116 & w7175) | (~w189 & w7175);
assign v764 = ~(w2976 | w2977);
assign w2978 = v764;
assign w2979 = ~pi117 & w1728;
assign w2980 = w146 & w7176;
assign w2981 = ~w81 & w6169;
assign v765 = ~(w2980 | w2981);
assign w2982 = v765;
assign w2983 = (pi117 & ~w146) | (pi117 & w7177) | (~w146 & w7177);
assign w2984 = (~w2983 & w1917) | (~w2983 & w7178) | (w1917 & w7178);
assign w2985 = ~w2982 & w2984;
assign w2986 = ~w2981 & w7179;
assign v766 = ~(w2985 | w2986);
assign w2987 = v766;
assign w2988 = (pi185 & ~w146) | (pi185 & w7180) | (~w146 & w7180);
assign w2989 = (~w2988 & w2282) | (~w2988 & w7181) | (w2282 & w7181);
assign w2990 = ~w2982 & w2989;
assign w2991 = (pi187 & ~w146) | (pi187 & w7182) | (~w146 & w7182);
assign w2992 = (~w2991 & w2193) | (~w2991 & w7183) | (w2193 & w7183);
assign w2993 = ~w2982 & w2992;
assign w2994 = w146 & w7184;
assign v767 = ~(w2981 | w2994);
assign w2995 = v767;
assign w2996 = (pi144 & ~w146) | (pi144 & w7185) | (~w146 & w7185);
assign w2997 = (~w2996 & w1424) | (~w2996 & w7186) | (w1424 & w7186);
assign w2998 = w2995 & ~w2997;
assign w2999 = w146 & w7187;
assign w3000 = (pi130 & ~w146) | (pi130 & w7188) | (~w146 & w7188);
assign w3001 = (~w3000 & w1075) | (~w3000 & w7189) | (w1075 & w7189);
assign w3002 = (w3001 & w2981) | (w3001 & w6170) | (w2981 & w6170);
assign w3003 = ~w2981 & w6171;
assign v768 = ~(w3002 | w3003);
assign w3004 = v768;
assign w3005 = (pi174 & ~w146) | (pi174 & w7190) | (~w146 & w7190);
assign w3006 = w146 & w7191;
assign w3007 = (~w3005 & w2058) | (~w3005 & w7192) | (w2058 & w7192);
assign w3008 = w3004 & w3007;
assign w3009 = (~w3002 & ~w3004) | (~w3002 & w6219) | (~w3004 & w6219);
assign w3010 = w146 & w7193;
assign v769 = ~(w2981 | w3010);
assign w3011 = v769;
assign w3012 = (pi172 & ~w146) | (pi172 & w7194) | (~w146 & w7194);
assign w3013 = (~w3012 & w1380) | (~w3012 & w7195) | (w1380 & w7195);
assign w3014 = ~w3011 & w3013;
assign w3015 = w3009 & ~w3014;
assign w3016 = w146 & w7196;
assign w3017 = (pi173 & ~w146) | (pi173 & w7197) | (~w146 & w7197);
assign w3018 = (~w3017 & w2102) | (~w3017 & w7198) | (w2102 & w7198);
assign w3019 = ~w2981 & w7335;
assign w3020 = ~w2981 & w7199;
assign v770 = ~(w3019 | w3020);
assign w3021 = v770;
assign w3022 = ~w3015 & w3021;
assign w3023 = (w3018 & w2981) | (w3018 & w7200) | (w2981 & w7200);
assign w3024 = w146 & w7201;
assign w3025 = (pi146 & ~w146) | (pi146 & w7202) | (~w146 & w7202);
assign w3026 = (~w3025 & w2018) | (~w3025 & w7203) | (w2018 & w7203);
assign w3027 = (w3026 & w2981) | (w3026 & w7336) | (w2981 & w7336);
assign v771 = ~(w3023 | w3027);
assign w3028 = v771;
assign w3029 = (w3028 & w3015) | (w3028 & w7204) | (w3015 & w7204);
assign w3030 = ~w2981 & w7205;
assign v772 = ~(w3030 | w3029);
assign w3031 = v772;
assign w3032 = (w2997 & w2981) | (w2997 & w7206) | (w2981 & w7206);
assign v773 = ~(w2998 | w3032);
assign w3033 = v773;
assign w3034 = (w3033 & w3029) | (w3033 & w7207) | (w3029 & w7207);
assign v774 = ~(w2998 | w3034);
assign w3035 = v774;
assign w3036 = (pi135 & ~w146) | (pi135 & w7208) | (~w146 & w7208);
assign w3037 = (~w3036 & w2240) | (~w3036 & w7209) | (w2240 & w7209);
assign w3038 = ~w2982 & w3037;
assign w3039 = w146 & w7210;
assign v775 = ~(w2981 | w3039);
assign w3040 = v775;
assign w3041 = (pi137 & ~w146) | (pi137 & w7211) | (~w146 & w7211);
assign w3042 = (~w3041 & w1471) | (~w3041 & w7212) | (w1471 & w7212);
assign w3043 = ~w3040 & w3042;
assign v776 = ~(w3038 | w3043);
assign w3044 = v776;
assign w3045 = ~w3035 & w3044;
assign w3046 = ~w2981 & w7213;
assign w3047 = ~w2981 & w7214;
assign w3048 = (~w3046 & w3038) | (~w3046 & w7215) | (w3038 & w7215);
assign w3049 = ~w3045 & w3048;
assign v777 = ~(w2990 | w2993);
assign w3050 = v777;
assign w3051 = ~w2981 & w7217;
assign w3052 = ~w2981 & w7218;
assign v778 = ~(w3051 | w3052);
assign w3053 = v778;
assign w3054 = w3053 & w7392;
assign w3055 = (pi183 & ~w146) | (pi183 & w7221) | (~w146 & w7221);
assign w3056 = (~w3055 & w1866) | (~w3055 & w7222) | (w1866 & w7222);
assign w3057 = ~w2982 & w3056;
assign w3058 = (pi186 & ~w146) | (pi186 & w7223) | (~w146 & w7223);
assign w3059 = (~w3058 & w1753) | (~w3058 & w7224) | (w1753 & w7224);
assign w3060 = ~w2982 & w3059;
assign w3061 = (pi177 & ~w146) | (pi177 & w7225) | (~w146 & w7225);
assign w3062 = (~w3061 & w1815) | (~w3061 & w7226) | (w1815 & w7226);
assign w3063 = ~w2982 & w3062;
assign v779 = ~(w3060 | w3063);
assign w3064 = v779;
assign w3065 = ~w3057 & w3064;
assign w3066 = (pi182 & ~w146) | (pi182 & w7227) | (~w146 & w7227);
assign w3067 = (~w3066 & w1969) | (~w3066 & w7228) | (w1969 & w7228);
assign w3068 = ~w2982 & w3067;
assign w3069 = w3064 & w7229;
assign w3070 = ~w2981 & w7232;
assign w3071 = ~w2981 & w7233;
assign w3072 = ~w2981 & w7234;
assign w3073 = ~w2981 & w7235;
assign v780 = ~(w3072 | w3073);
assign w3074 = v780;
assign w3075 = ~w3071 & w3074;
assign w3076 = w3074 & w7236;
assign w3077 = w3076 & w7393;
assign w3078 = w2987 & w3077;
assign v781 = ~(w2987 | w3077);
assign w3079 = v781;
assign v782 = ~(w3078 | w3079);
assign w3080 = v782;
assign w3081 = (~w982 & ~w82) | (~w982 & w7237) | (~w82 & w7237);
assign w3082 = ~pi117 & w3081;
assign w3083 = w24 & w47;
assign w3084 = w1051 & w3083;
assign v783 = ~(w3082 | w3084);
assign w3085 = v783;
assign w3086 = w1512 & w3085;
assign w3087 = w1512 & ~w3081;
assign w3088 = (~w3084 & ~w1512) | (~w3084 & w7238) | (~w1512 & w7238);
assign w3089 = pi117 & w3088;
assign w3090 = (~w1732 & w1917) | (~w1732 & w7239) | (w1917 & w7239);
assign w3091 = ~w3089 & w3090;
assign w3092 = pi240 & w2803;
assign w3093 = w1507 & w7241;
assign w3094 = ~pi117 & w1732;
assign v784 = ~(w3093 | w3094);
assign w3095 = v784;
assign w3096 = w3095 & w7394;
assign w3097 = (w1731 & w1570) | (w1731 & w7242) | (w1570 & w7242);
assign w3098 = ~w3096 & w3097;
assign v785 = ~(w2979 | w3098);
assign w3099 = v785;
assign w3100 = ~w1523 & w7243;
assign w3101 = w1523 & w7244;
assign w3102 = w1523 & w7245;
assign w3103 = pi121 & w1524;
assign w3104 = pi118 & w1539;
assign w3105 = ~w1523 & w7246;
assign w3106 = w1523 & w7247;
assign w3107 = ~w1523 & w7248;
assign v786 = ~(w3100 | w3101);
assign w3108 = v786;
assign v787 = ~(w3102 | w3103);
assign w3109 = v787;
assign v788 = ~(w3104 | w3105);
assign w3110 = v788;
assign v789 = ~(w3106 | w3107);
assign w3111 = v789;
assign w3112 = w3110 & w3111;
assign w3113 = w3108 & w3109;
assign w3114 = w3112 & w3113;
assign w3115 = w162 & w3114;
assign w3116 = ~pi267 & w165;
assign w3117 = ~w518 & w7249;
assign w3118 = ~w521 & w1511;
assign w3119 = ~w3116 & w2468;
assign w3120 = (w3119 & ~w3118) | (w3119 & w7250) | (~w3118 & w7250);
assign w3121 = (w2572 & w3120) | (w2572 & w7251) | (w3120 & w7251);
assign w3122 = (~pi118 & ~w189) | (~pi118 & w7252) | (~w189 & w7252);
assign v790 = ~(w3121 | w3122);
assign w3123 = v790;
assign w3124 = (w2576 & w3120) | (w2576 & w7253) | (w3120 & w7253);
assign w3125 = (~pi119 & ~w202) | (~pi119 & w7254) | (~w202 & w7254);
assign v791 = ~(w3124 | w3125);
assign w3126 = v791;
assign w3127 = (w2539 & w3120) | (w2539 & w7255) | (w3120 & w7255);
assign w3128 = (~pi120 & ~w206) | (~pi120 & w7256) | (~w206 & w7256);
assign v792 = ~(w3127 | w3128);
assign w3129 = v792;
assign w3130 = (w2564 & w3120) | (w2564 & w7257) | (w3120 & w7257);
assign w3131 = (~pi121 & ~w197) | (~pi121 & w7258) | (~w197 & w7258);
assign v793 = ~(w3130 | w3131);
assign w3132 = v793;
assign w3133 = (w2584 & w3120) | (w2584 & w7259) | (w3120 & w7259);
assign w3134 = (~pi122 & ~w195) | (~pi122 & w7260) | (~w195 & w7260);
assign v794 = ~(w3133 | w3134);
assign w3135 = v794;
assign w3136 = (w2588 & w3120) | (w2588 & w7261) | (w3120 & w7261);
assign w3137 = (~pi123 & ~w192) | (~pi123 & w7262) | (~w192 & w7262);
assign v795 = ~(w3136 | w3137);
assign w3138 = v795;
assign w3139 = (w2580 & w3120) | (w2580 & w7263) | (w3120 & w7263);
assign w3140 = (~pi124 & ~w199) | (~pi124 & w7264) | (~w199 & w7264);
assign v796 = ~(w3139 | w3140);
assign w3141 = v796;
assign w3142 = (w2568 & w3120) | (w2568 & w7265) | (w3120 & w7265);
assign v797 = ~(pi125 | w2568);
assign w3143 = v797;
assign v798 = ~(w3142 | w3143);
assign w3144 = v798;
assign w3145 = pi126 & pi247;
assign w3146 = w1497 & w1498;
assign w3147 = w1507 & w7266;
assign w3148 = ~w2646 & w7267;
assign w3149 = w2450 & w2894;
assign v799 = ~(w2895 | w3149);
assign w3150 = v799;
assign w3151 = ~w3149 & w7268;
assign w3152 = w2894 & w7269;
assign w3153 = (w2897 & w3151) | (w2897 & w7270) | (w3151 & w7270);
assign w3154 = pi326 & w2901;
assign w3155 = w0 & w614;
assign w3156 = w1120 & w3155;
assign w3157 = w1032 & w7271;
assign v800 = ~(w2901 | w3157);
assign w3158 = v800;
assign w3159 = ~w3157 & w7272;
assign w3160 = (~w3154 & ~w3157) | (~w3154 & w7273) | (~w3157 & w7273);
assign w3161 = ~w3159 & w3160;
assign v801 = ~(w3147 | w3153);
assign w3162 = v801;
assign v802 = ~(pi247 | w3148);
assign w3163 = v802;
assign w3164 = w3163 & w7395;
assign w3165 = pi359 & ~w3145;
assign w3166 = ~w3164 & w3165;
assign w3167 = pi155 & w1524;
assign w3168 = pi158 & w1539;
assign w3169 = ~w1523 & w7275;
assign w3170 = w1523 & w7276;
assign w3171 = w1523 & w7277;
assign w3172 = ~w1523 & w7278;
assign w3173 = ~w1523 & w7279;
assign w3174 = w1523 & w7280;
assign v803 = ~(w3167 | w3168);
assign w3175 = v803;
assign v804 = ~(w3169 | w3170);
assign w3176 = v804;
assign v805 = ~(w3171 | w3172);
assign w3177 = v805;
assign v806 = ~(w3173 | w3174);
assign w3178 = v806;
assign w3179 = w3177 & w3178;
assign w3180 = w3175 & w3176;
assign w3181 = w3179 & w3180;
assign w3182 = w3180 & w7281;
assign w3183 = ~pi260 & w165;
assign v807 = ~(w320 | w321);
assign w3184 = v807;
assign w3185 = w336 & w1511;
assign w3186 = w3184 & w3185;
assign w3187 = ~w336 & w1511;
assign w3188 = ~w3184 & w3187;
assign v808 = ~(w162 | w3183);
assign w3189 = v808;
assign w3190 = (w3189 & w2527) | (w3189 & w7282) | (w2527 & w7282);
assign w3191 = ~w3186 & w3190;
assign w3192 = (~w3182 & ~w3191) | (~w3182 & w7283) | (~w3191 & w7283);
assign w3193 = w2588 & ~w3192;
assign w3194 = (~pi127 & ~w192) | (~pi127 & w7284) | (~w192 & w7284);
assign v809 = ~(w3193 | w3194);
assign w3195 = v809;
assign w3196 = w1507 & w7285;
assign w3197 = (w1502 & ~w1507) | (w1502 & w7286) | (~w1507 & w7286);
assign w3198 = w1 & w7287;
assign w3199 = w1231 & w3198;
assign w3200 = (~pi273 & ~w1231) | (~pi273 & w7288) | (~w1231 & w7288);
assign w3201 = ~pi271 & pi303;
assign v810 = ~(w765 | w3201);
assign w3202 = v810;
assign w3203 = w1231 & w7289;
assign v811 = ~(w3200 | w3203);
assign w3204 = v811;
assign w3205 = w3197 & w3204;
assign w3206 = (~w3205 & w2404) | (~w3205 & w7290) | (w2404 & w7290);
assign w3207 = w1731 & ~w3206;
assign w3208 = (~w1502 & ~w1507) | (~w1502 & w7291) | (~w1507 & w7291);
assign w3209 = (pi359 & w3208) | (pi359 & w1728) | (w3208 & w1728);
assign w3210 = pi128 & w3209;
assign v812 = ~(w3207 | w3210);
assign w3211 = v812;
assign w3212 = ~pi129 & w1728;
assign w3213 = w2805 & ~w2527;
assign v813 = ~(w701 | w733);
assign w3214 = v813;
assign w3215 = ~pi129 & pi243;
assign v814 = ~(w3214 | w3215);
assign w3216 = v814;
assign w3217 = ~w2810 & w3216;
assign w3218 = ~pi320 & w2901;
assign w3219 = ~w3157 & w7292;
assign w3220 = w0 & w1140;
assign w3221 = w0 & w1146;
assign v815 = ~(w3220 | w3221);
assign w3222 = v815;
assign w3223 = w1032 & w7293;
assign w3224 = w2810 & ~w3218;
assign w3225 = ~w3223 & w3224;
assign w3226 = ~w3219 & w3225;
assign w3227 = w6131 & w7294;
assign v816 = ~(w2805 | w3227);
assign w3228 = v816;
assign w3229 = ~w2892 & w3228;
assign w3230 = (w3229 & w3226) | (w3229 & w7295) | (w3226 & w7295);
assign w3231 = w1731 & ~w3213;
assign w3232 = ~w3230 & w3231;
assign v817 = ~(w3212 | w3232);
assign w3233 = v817;
assign w3234 = pi130 & pi247;
assign w3235 = w1507 & w7296;
assign w3236 = w82 & w7297;
assign v818 = ~(w3004 | w3007);
assign w3237 = v818;
assign v819 = ~(w3008 | w3237);
assign w3238 = v819;
assign w3239 = ~pi130 & w3088;
assign w3240 = (~w1732 & ~w1075) | (~w1732 & w7239) | (~w1075 & w7239);
assign w3241 = ~w3239 & w3240;
assign w3242 = (w3241 & ~w3238) | (w3241 & w7298) | (~w3238 & w7298);
assign v820 = ~(w3235 | w3236);
assign w3243 = v820;
assign w3244 = ~w3242 & w3243;
assign w3245 = (~pi247 & ~w2527) | (~pi247 & w7299) | (~w2527 & w7299);
assign w3246 = ~w3244 & w3245;
assign w3247 = pi359 & ~w3234;
assign w3248 = ~w3246 & w3247;
assign w3249 = pi131 & pi247;
assign v821 = ~(pi131 | w2901);
assign w3250 = v821;
assign w3251 = ~pi325 & w2901;
assign w3252 = w2810 & ~w3250;
assign w3253 = ~w3251 & w3252;
assign v822 = ~(w2892 | w3253);
assign w3254 = v822;
assign w3255 = w2909 & w2912;
assign w3256 = w2918 & w2921;
assign w3257 = w3255 & w3256;
assign w3258 = w2892 & ~w3257;
assign w3259 = (w973 & w7305) | (w973 & w7306) | (w7305 & w7306);
assign v823 = ~(w2805 | w3259);
assign w3260 = v823;
assign w3261 = ~pi247 & w7396;
assign w3262 = ~w3260 & w3261;
assign w3263 = pi359 & ~w3249;
assign w3264 = ~w3262 & w3263;
assign w3265 = pi132 & pi247;
assign w3266 = ~w2646 & w7307;
assign w3267 = pi132 & pi243;
assign w3268 = ~w709 & w3267;
assign w3269 = (w701 & ~w643) | (w701 & w7308) | (~w643 & w7308);
assign v824 = ~(pi335 | w2810);
assign w3270 = v824;
assign v825 = ~(pi223 | pi303);
assign w3271 = v825;
assign w3272 = ~pi197 & pi303;
assign v826 = ~(w3271 | w3272);
assign w3273 = v826;
assign w3274 = w736 & w3273;
assign v827 = ~(w840 | w2812);
assign w3275 = v827;
assign v828 = ~(pi241 | pi256);
assign w3276 = v828;
assign v829 = ~(w3275 | w3276);
assign w3277 = v829;
assign w3278 = ~w733 & w3275;
assign v830 = ~(pi243 | w3277);
assign w3279 = v830;
assign w3280 = ~w3278 & w3279;
assign v831 = ~(w3268 | w3274);
assign w3281 = v831;
assign w3282 = w3270 & w3281;
assign w3283 = ~w3269 & w3282;
assign w3284 = ~w3280 & w3283;
assign w3285 = pi322 & w2901;
assign v832 = ~(w1732 | w2900);
assign w3286 = v832;
assign w3287 = w1033 & w3221;
assign w3288 = pi132 & ~w3287;
assign w3289 = pi132 & ~w3220;
assign w3290 = w3223 & ~w3289;
assign v833 = ~(w3288 | w3290);
assign w3291 = v833;
assign w3292 = w3286 & ~w3291;
assign w3293 = pi132 & w1732;
assign v834 = ~(w3285 | w3293);
assign w3294 = v834;
assign w3295 = ~w3270 & w3294;
assign w3296 = ~w3292 & w3295;
assign v835 = ~(w3284 | w3296);
assign w3297 = v835;
assign v836 = ~(w2805 | w3297);
assign w3298 = v836;
assign v837 = ~(pi247 | w3266);
assign w3299 = v837;
assign w3300 = ~w3298 & w3299;
assign w3301 = pi359 & ~w3265;
assign w3302 = ~w3300 & w3301;
assign w3303 = pi133 & pi247;
assign w3304 = w2327 & w3147;
assign w3305 = pi339 & w3150;
assign w3306 = pi332 & w3149;
assign v838 = ~(w3305 | w3306);
assign w3307 = v838;
assign w3308 = w2897 & ~w3307;
assign w3309 = pi330 & w2901;
assign w3310 = ~pi133 & w3157;
assign w3311 = pi133 & w3158;
assign v839 = ~(w3309 | w3310);
assign w3312 = v839;
assign w3313 = ~w3311 & w3312;
assign v840 = ~(w2898 | w3313);
assign w3314 = v840;
assign v841 = ~(w3147 | w3308);
assign w3315 = v841;
assign w3316 = ~w3314 & w3315;
assign v842 = ~(pi247 | w3316);
assign w3317 = v842;
assign w3318 = ~w3304 & w3317;
assign w3319 = pi359 & ~w3303;
assign w3320 = ~w3318 & w3319;
assign w3321 = ~w2327 & w3196;
assign v843 = ~(pi275 | w3199);
assign w3322 = v843;
assign v844 = ~(w742 | w769);
assign w3323 = v844;
assign w3324 = w3199 & w3323;
assign v845 = ~(w3322 | w3324);
assign w3325 = v845;
assign w3326 = w3197 & w3325;
assign v846 = ~(w3321 | w3326);
assign w3327 = v846;
assign w3328 = w1731 & ~w3327;
assign w3329 = pi134 & w3209;
assign v847 = ~(w3328 | w3329);
assign w3330 = v847;
assign w3331 = pi135 & pi247;
assign w3332 = w2327 & w3235;
assign v848 = ~(w1732 | w3088);
assign w3333 = v848;
assign w3334 = pi135 & ~w3333;
assign w3335 = ~w2240 & w3084;
assign v849 = ~(w3038 | w3046);
assign w3336 = v849;
assign v850 = ~(w3032 | w3043);
assign w3337 = v850;
assign w3338 = ~w3031 & w3337;
assign w3339 = w2998 & ~w3043;
assign v851 = ~(w3047 | w3339);
assign w3340 = v851;
assign w3341 = ~w3338 & w3340;
assign w3342 = w3336 & ~w3341;
assign w3343 = ~w3336 & w3341;
assign v852 = ~(w3342 | w3343);
assign w3344 = v852;
assign w3345 = w3087 & w3344;
assign v853 = ~(w3335 | w3345);
assign w3346 = v853;
assign v854 = ~(w1732 | w3346);
assign w3347 = v854;
assign v855 = ~(w3235 | w3334);
assign w3348 = v855;
assign w3349 = ~w3347 & w3348;
assign v856 = ~(pi247 | w3332);
assign w3350 = v856;
assign w3351 = ~w3349 & w3350;
assign w3352 = pi359 & ~w3331;
assign w3353 = ~w3351 & w3352;
assign w3354 = ~w1570 & w3196;
assign v857 = ~(pi269 | w3199);
assign w3355 = v857;
assign w3356 = pi274 & pi303;
assign v858 = ~(w796 | w3356);
assign w3357 = v858;
assign w3358 = w3199 & w3357;
assign v859 = ~(w3355 | w3358);
assign w3359 = v859;
assign w3360 = w3197 & w3359;
assign v860 = ~(w3354 | w3360);
assign w3361 = v860;
assign w3362 = w1731 & ~w3361;
assign w3363 = pi136 & w3209;
assign v861 = ~(w3362 | w3363);
assign w3364 = v861;
assign w3365 = pi137 & pi247;
assign w3366 = w1570 & w3235;
assign w3367 = ~w1471 & w3084;
assign v862 = ~(w3043 | w3047);
assign w3368 = v862;
assign w3369 = w3035 & w3368;
assign v863 = ~(w3035 | w3368);
assign w3370 = v863;
assign v864 = ~(w3369 | w3370);
assign w3371 = v864;
assign w3372 = w3087 & ~w3371;
assign v865 = ~(w3367 | w3372);
assign w3373 = v865;
assign v866 = ~(w1732 | w3373);
assign w3374 = v866;
assign w3375 = pi137 & ~w3333;
assign v867 = ~(w3235 | w3375);
assign w3376 = v867;
assign w3377 = ~w3374 & w3376;
assign v868 = ~(pi247 | w3366);
assign w3378 = v868;
assign w3379 = ~w3377 & w3378;
assign w3380 = pi359 & ~w3365;
assign w3381 = ~w3379 & w3380;
assign w3382 = pi138 & pi247;
assign w3383 = ~w2467 & w3147;
assign w3384 = pi343 & w3150;
assign w3385 = pi288 & w3149;
assign v869 = ~(w3384 | w3385);
assign w3386 = v869;
assign w3387 = w2897 & ~w3386;
assign w3388 = pi316 & w2901;
assign w3389 = ~pi138 & w3157;
assign w3390 = pi138 & w3158;
assign v870 = ~(w3388 | w3389);
assign w3391 = v870;
assign w3392 = ~w3390 & w3391;
assign v871 = ~(w2898 | w3392);
assign w3393 = v871;
assign v872 = ~(w3147 | w3387);
assign w3394 = v872;
assign w3395 = ~w3393 & w3394;
assign v873 = ~(pi247 | w3383);
assign w3396 = v873;
assign w3397 = ~w3395 & w3396;
assign w3398 = pi359 & ~w3382;
assign w3399 = ~w3397 & w3398;
assign w3400 = pi139 & pi247;
assign w3401 = w2404 & w3147;
assign w3402 = pi336 & w3150;
assign w3403 = pi287 & w3149;
assign v874 = ~(w3402 | w3403);
assign w3404 = v874;
assign w3405 = w2897 & ~w3404;
assign w3406 = pi317 & w2901;
assign w3407 = ~pi139 & w3157;
assign w3408 = pi139 & w3158;
assign v875 = ~(w3406 | w3407);
assign w3409 = v875;
assign w3410 = ~w3408 & w3409;
assign v876 = ~(w2898 | w3410);
assign w3411 = v876;
assign v877 = ~(w3147 | w3405);
assign w3412 = v877;
assign w3413 = ~w3411 & w3412;
assign v878 = ~(pi247 | w3413);
assign w3414 = v878;
assign w3415 = ~w3401 & w3414;
assign w3416 = pi359 & ~w3400;
assign w3417 = ~w3415 & w3416;
assign w3418 = pi140 & pi247;
assign w3419 = w1570 & w3147;
assign w3420 = pi340 & w3150;
assign w3421 = pi286 & w3149;
assign v879 = ~(w3420 | w3421);
assign w3422 = v879;
assign w3423 = w2897 & ~w3422;
assign w3424 = pi329 & w2901;
assign w3425 = ~pi140 & w3157;
assign w3426 = pi140 & w3158;
assign v880 = ~(w3424 | w3425);
assign w3427 = v880;
assign w3428 = ~w3426 & w3427;
assign v881 = ~(w2898 | w3428);
assign w3429 = v881;
assign v882 = ~(w3147 | w3423);
assign w3430 = v882;
assign w3431 = ~w3429 & w3430;
assign v883 = ~(pi247 | w3431);
assign w3432 = v883;
assign w3433 = ~w3419 & w3432;
assign w3434 = pi359 & ~w3418;
assign w3435 = ~w3433 & w3434;
assign w3436 = pi141 & pi247;
assign w3437 = w1697 & w3147;
assign w3438 = pi337 & w3150;
assign w3439 = pi289 & w3149;
assign v884 = ~(w3438 | w3439);
assign w3440 = v884;
assign w3441 = w2897 & ~w3440;
assign w3442 = pi327 & w2901;
assign w3443 = ~pi141 & w3157;
assign w3444 = pi141 & w3158;
assign v885 = ~(w3442 | w3443);
assign w3445 = v885;
assign w3446 = ~w3444 & w3445;
assign v886 = ~(w2898 | w3446);
assign w3447 = v886;
assign v887 = ~(w3147 | w3441);
assign w3448 = v887;
assign w3449 = ~w3447 & w3448;
assign v888 = ~(pi247 | w3437);
assign w3450 = v888;
assign w3451 = ~w3449 & w3450;
assign w3452 = pi359 & ~w3436;
assign w3453 = ~w3451 & w3452;
assign w3454 = pi142 & pi247;
assign w3455 = w2527 & w3147;
assign w3456 = pi342 & w3150;
assign w3457 = pi295 & w3149;
assign v889 = ~(w3456 | w3457);
assign w3458 = v889;
assign w3459 = w2897 & ~w3458;
assign w3460 = pi319 & w2901;
assign w3461 = ~pi142 & w3157;
assign w3462 = pi142 & w3158;
assign v890 = ~(w3460 | w3461);
assign w3463 = v890;
assign w3464 = ~w3462 & w3463;
assign v891 = ~(w2898 | w3464);
assign w3465 = v891;
assign v892 = ~(w3147 | w3459);
assign w3466 = v892;
assign w3467 = ~w3465 & w3466;
assign v893 = ~(pi247 | w3455);
assign w3468 = v893;
assign w3469 = ~w3467 & w3468;
assign w3470 = pi359 & ~w3454;
assign w3471 = ~w3469 & w3470;
assign w3472 = pi143 & pi247;
assign w3473 = w1620 & w3147;
assign w3474 = pi338 & w3150;
assign w3475 = pi290 & w3149;
assign v894 = ~(w3474 | w3475);
assign w3476 = v894;
assign w3477 = w2897 & ~w3476;
assign w3478 = pi328 & w2901;
assign w3479 = ~pi143 & w3157;
assign w3480 = pi143 & w3158;
assign v895 = ~(w3478 | w3479);
assign w3481 = v895;
assign w3482 = ~w3480 & w3481;
assign v896 = ~(w2898 | w3482);
assign w3483 = v896;
assign v897 = ~(w3147 | w3477);
assign w3484 = v897;
assign w3485 = ~w3483 & w3484;
assign v898 = ~(pi247 | w3473);
assign w3486 = v898;
assign w3487 = ~w3485 & w3486;
assign w3488 = pi359 & ~w3472;
assign w3489 = ~w3487 & w3488;
assign w3490 = pi144 & pi247;
assign w3491 = w2404 & w3235;
assign w3492 = ~w1424 & w3084;
assign w3493 = w3031 & ~w3033;
assign v899 = ~(w3034 | w3493);
assign w3494 = v899;
assign w3495 = w3087 & w3494;
assign v900 = ~(w3492 | w3495);
assign w3496 = v900;
assign v901 = ~(w1732 | w3496);
assign w3497 = v901;
assign w3498 = pi144 & ~w3333;
assign v902 = ~(w3235 | w3498);
assign w3499 = v902;
assign w3500 = ~w3497 & w3499;
assign v903 = ~(pi247 | w3491);
assign w3501 = v903;
assign w3502 = ~w3500 & w3501;
assign w3503 = pi359 & ~w3490;
assign w3504 = ~w3502 & w3503;
assign w3505 = ~w1620 & w3196;
assign v904 = ~(pi270 | w3199);
assign w3506 = v904;
assign w3507 = pi264 & pi303;
assign v905 = ~(w785 | w3507);
assign w3508 = v905;
assign w3509 = w3199 & w3508;
assign v906 = ~(w3506 | w3509);
assign w3510 = v906;
assign w3511 = w3197 & w3510;
assign v907 = ~(w3505 | w3511);
assign w3512 = v907;
assign w3513 = w1731 & ~w3512;
assign w3514 = pi145 & w3209;
assign v908 = ~(w3513 | w3514);
assign w3515 = v908;
assign w3516 = pi146 & pi247;
assign w3517 = w1620 & w3235;
assign w3518 = pi146 & ~w3333;
assign w3519 = ~w2018 & w3084;
assign v909 = ~(w3027 | w3030);
assign w3520 = v909;
assign v910 = ~(w3022 | w3023);
assign w3521 = v910;
assign w3522 = w3520 & w3521;
assign v911 = ~(w3520 | w3521);
assign w3523 = v911;
assign v912 = ~(w3522 | w3523);
assign w3524 = v912;
assign w3525 = w3087 & w3524;
assign v913 = ~(w3519 | w3525);
assign w3526 = v913;
assign v914 = ~(w1732 | w3526);
assign w3527 = v914;
assign v915 = ~(w3235 | w3518);
assign w3528 = v915;
assign w3529 = ~w3527 & w3528;
assign v916 = ~(pi247 | w3517);
assign w3530 = v916;
assign w3531 = ~w3529 & w3530;
assign w3532 = pi359 & ~w3516;
assign w3533 = ~w3531 & w3532;
assign w3534 = pi152 & w1530;
assign w3535 = pi150 & w1527;
assign w3536 = pi153 & w1541;
assign w3537 = pi149 & w1537;
assign w3538 = pi148 & w1524;
assign w3539 = pi147 & w1533;
assign w3540 = pi175 & w1535;
assign w3541 = pi151 & w1539;
assign v917 = ~(w3534 | w3535);
assign w3542 = v917;
assign v918 = ~(w3536 | w3537);
assign w3543 = v918;
assign v919 = ~(w3538 | w3539);
assign w3544 = v919;
assign v920 = ~(w3540 | w3541);
assign w3545 = v920;
assign w3546 = w3544 & w3545;
assign w3547 = w3542 & w3543;
assign w3548 = w3546 & w3547;
assign w3549 = w162 & w3548;
assign w3550 = ~pi261 & w165;
assign w3551 = w338 & ~w591;
assign w3552 = ~w592 & w1511;
assign w3553 = ~w3551 & w3552;
assign v921 = ~(w162 | w3550);
assign w3554 = v921;
assign w3555 = ~w1698 & w3554;
assign w3556 = ~w3553 & w3555;
assign v922 = ~(w3549 | w3556);
assign w3557 = v922;
assign w3558 = w2539 & ~w3557;
assign v923 = ~(pi147 | w2539);
assign w3559 = v923;
assign v924 = ~(w3558 | w3559);
assign w3560 = v924;
assign w3561 = w2564 & ~w3557;
assign v925 = ~(pi148 | w2564);
assign w3562 = v925;
assign v926 = ~(w3561 | w3562);
assign w3563 = v926;
assign w3564 = w2568 & ~w3557;
assign v927 = ~(pi149 | w2568);
assign w3565 = v927;
assign v928 = ~(w3564 | w3565);
assign w3566 = v928;
assign w3567 = w2584 & ~w3557;
assign v929 = ~(pi150 | w2584);
assign w3568 = v929;
assign v930 = ~(w3567 | w3568);
assign w3569 = v930;
assign w3570 = w2572 & ~w3557;
assign v931 = ~(pi151 | w2572);
assign w3571 = v931;
assign v932 = ~(w3570 | w3571);
assign w3572 = v932;
assign w3573 = w2576 & ~w3557;
assign v933 = ~(pi152 | w2576);
assign w3574 = v933;
assign v934 = ~(w3573 | w3574);
assign w3575 = v934;
assign w3576 = w2580 & ~w3557;
assign v935 = ~(pi153 | w2580);
assign w3577 = v935;
assign v936 = ~(w3576 | w3577);
assign w3578 = v936;
assign w3579 = w2539 & ~w3192;
assign v937 = ~(pi154 | w2539);
assign w3580 = v937;
assign v938 = ~(w3579 | w3580);
assign w3581 = v938;
assign w3582 = w2564 & ~w3192;
assign v939 = ~(pi155 | w2564);
assign w3583 = v939;
assign v940 = ~(w3582 | w3583);
assign w3584 = v940;
assign w3585 = w2568 & ~w3192;
assign v941 = ~(pi156 | w2568);
assign w3586 = v941;
assign v942 = ~(w3585 | w3586);
assign w3587 = v942;
assign w3588 = w2584 & ~w3192;
assign v943 = ~(pi157 | w2584);
assign w3589 = v943;
assign v944 = ~(w3588 | w3589);
assign w3590 = v944;
assign w3591 = w2572 & ~w3192;
assign v945 = ~(pi158 | w2572);
assign w3592 = v945;
assign v946 = ~(w3591 | w3592);
assign w3593 = v946;
assign w3594 = w2576 & ~w3192;
assign v947 = ~(pi159 | w2576);
assign w3595 = v947;
assign v948 = ~(w3594 | w3595);
assign w3596 = v948;
assign w3597 = w2580 & ~w3192;
assign v949 = ~(pi160 | w2580);
assign w3598 = v949;
assign v950 = ~(w3597 | w3598);
assign w3599 = v950;
assign w3600 = pi161 & w3209;
assign w3601 = ~w2648 & w3196;
assign v951 = ~(pi264 | w3199);
assign w3602 = v951;
assign v952 = ~(pi270 | pi303);
assign w3603 = v952;
assign v953 = ~(w3272 | w3603);
assign w3604 = v953;
assign w3605 = w3199 & ~w3604;
assign v954 = ~(w3602 | w3605);
assign w3606 = v954;
assign w3607 = w3197 & w3606;
assign v955 = ~(w3601 | w3607);
assign w3608 = v955;
assign w3609 = w1731 & ~w3608;
assign v956 = ~(w3600 | w3609);
assign w3610 = v956;
assign w3611 = ~w2527 & w3196;
assign v957 = ~(pi271 | w3199);
assign w3612 = v957;
assign w3613 = pi273 & ~pi303;
assign v958 = ~(w778 | w3613);
assign w3614 = v958;
assign w3615 = w3199 & w3614;
assign v959 = ~(w3612 | w3615);
assign w3616 = v959;
assign w3617 = w3197 & w3616;
assign v960 = ~(w3611 | w3617);
assign w3618 = v960;
assign w3619 = w1731 & ~w3618;
assign w3620 = pi162 & w3209;
assign v961 = ~(w3619 | w3620);
assign w3621 = v961;
assign w3622 = ~w1697 & w3196;
assign v962 = ~(pi274 | w3199);
assign w3623 = v962;
assign v963 = ~(w755 | w784);
assign w3624 = v963;
assign w3625 = w3199 & w3624;
assign v964 = ~(w3623 | w3625);
assign w3626 = v964;
assign w3627 = w3197 & w3626;
assign v965 = ~(w3622 | w3627);
assign w3628 = v965;
assign w3629 = w1731 & ~w3628;
assign w3630 = pi163 & w3209;
assign v966 = ~(w3629 | w3630);
assign w3631 = v966;
assign w3632 = w2467 & w3196;
assign v967 = ~(pi272 | w3199);
assign w3633 = v967;
assign v968 = ~(pi275 | pi303);
assign w3634 = v968;
assign v969 = ~(w766 | w3634);
assign w3635 = v969;
assign w3636 = w3199 & ~w3635;
assign v970 = ~(w3633 | w3636);
assign w3637 = v970;
assign w3638 = w3197 & w3637;
assign v971 = ~(w3632 | w3638);
assign w3639 = v971;
assign w3640 = w1731 & ~w3639;
assign w3641 = pi164 & w3209;
assign v972 = ~(w3640 | w3641);
assign w3642 = v972;
assign w3643 = pi166 & w1524;
assign w3644 = pi170 & w1539;
assign w3645 = pi168 & w1527;
assign w3646 = pi171 & w1541;
assign w3647 = pi165 & w1533;
assign w3648 = pi169 & w1535;
assign w3649 = pi167 & w1537;
assign w3650 = pi176 & w1530;
assign v973 = ~(w3643 | w3644);
assign w3651 = v973;
assign v974 = ~(w3645 | w3646);
assign w3652 = v974;
assign v975 = ~(w3647 | w3648);
assign w3653 = v975;
assign v976 = ~(w3649 | w3650);
assign w3654 = v976;
assign w3655 = w3653 & w3654;
assign w3656 = w3651 & w3652;
assign w3657 = w3655 & w3656;
assign w3658 = w162 & w3657;
assign w3659 = ~pi235 & w165;
assign w3660 = w2650 & ~w3659;
assign w3661 = ~w3185 & w3660;
assign v977 = ~(w3658 | w3661);
assign w3662 = v977;
assign w3663 = w2539 & ~w3662;
assign v978 = ~(pi165 | w2539);
assign w3664 = v978;
assign v979 = ~(w3663 | w3664);
assign w3665 = v979;
assign w3666 = w2564 & ~w3662;
assign v980 = ~(pi166 | w2564);
assign w3667 = v980;
assign v981 = ~(w3666 | w3667);
assign w3668 = v981;
assign w3669 = w2568 & ~w3662;
assign v982 = ~(pi167 | w2568);
assign w3670 = v982;
assign v983 = ~(w3669 | w3670);
assign w3671 = v983;
assign w3672 = w2584 & ~w3662;
assign v984 = ~(pi168 | w2584);
assign w3673 = v984;
assign v985 = ~(w3672 | w3673);
assign w3674 = v985;
assign w3675 = w2588 & ~w3662;
assign v986 = ~(pi169 | w2588);
assign w3676 = v986;
assign v987 = ~(w3675 | w3676);
assign w3677 = v987;
assign w3678 = w2572 & ~w3662;
assign v988 = ~(pi170 | w2572);
assign w3679 = v988;
assign v989 = ~(w3678 | w3679);
assign w3680 = v989;
assign w3681 = w2580 & ~w3662;
assign v990 = ~(pi171 | w2580);
assign w3682 = v990;
assign v991 = ~(w3681 | w3682);
assign w3683 = v991;
assign w3684 = pi172 & pi247;
assign w3685 = w1697 & w3235;
assign w3686 = pi172 & w1732;
assign w3687 = w1380 & w3084;
assign v992 = ~(w3014 | w3020);
assign w3688 = v992;
assign v993 = ~(w3009 | w3688);
assign w3689 = v993;
assign w3690 = w3009 & w3688;
assign v994 = ~(w3689 | w3690);
assign w3691 = v994;
assign w3692 = w3087 & ~w3691;
assign w3693 = ~pi172 & w3088;
assign v995 = ~(w1732 | w3687);
assign w3694 = v995;
assign w3695 = ~w3693 & w3694;
assign w3696 = ~w3692 & w3695;
assign v996 = ~(w3235 | w3686);
assign w3697 = v996;
assign w3698 = ~w3696 & w3697;
assign v997 = ~(pi247 | w3685);
assign w3699 = v997;
assign w3700 = ~w3698 & w3699;
assign w3701 = pi359 & ~w3684;
assign w3702 = ~w3700 & w3701;
assign w3703 = pi173 & pi247;
assign w3704 = ~w2467 & w3235;
assign w3705 = pi173 & w1732;
assign w3706 = w2102 & w3084;
assign v998 = ~(w3015 | w3020);
assign w3707 = v998;
assign v999 = ~(w3019 | w3023);
assign w3708 = v999;
assign w3709 = w3707 & w3708;
assign v1000 = ~(w3707 | w3708);
assign w3710 = v1000;
assign v1001 = ~(w3709 | w3710);
assign w3711 = v1001;
assign w3712 = w3087 & w3711;
assign w3713 = ~pi173 & w3088;
assign v1002 = ~(w1732 | w3706);
assign w3714 = v1002;
assign w3715 = ~w3713 & w3714;
assign w3716 = ~w3712 & w3715;
assign v1003 = ~(w3235 | w3705);
assign w3717 = v1003;
assign w3718 = ~w3716 & w3717;
assign v1004 = ~(pi247 | w3704);
assign w3719 = v1004;
assign w3720 = ~w3718 & w3719;
assign w3721 = pi359 & ~w3703;
assign w3722 = ~w3720 & w3721;
assign w3723 = pi174 & pi247;
assign w3724 = w2648 & w3235;
assign w3725 = w2058 & w3084;
assign w3726 = ~pi354 & w147;
assign w3727 = w2058 & w3726;
assign w3728 = w3007 & ~w3727;
assign w3729 = w3087 & ~w3728;
assign v1005 = ~(w3725 | w3729);
assign w3730 = v1005;
assign v1006 = ~(w1732 | w3730);
assign w3731 = v1006;
assign v1007 = ~(pi174 | w3333);
assign w3732 = v1007;
assign v1008 = ~(w3731 | w3732);
assign w3733 = v1008;
assign v1009 = ~(w3235 | w3733);
assign w3734 = v1009;
assign v1010 = ~(pi247 | w3724);
assign w3735 = v1010;
assign w3736 = ~w3734 & w3735;
assign w3737 = pi359 & ~w3723;
assign w3738 = ~w3736 & w3737;
assign w3739 = w2588 & ~w3557;
assign v1011 = ~(pi175 | w2588);
assign w3740 = v1011;
assign v1012 = ~(w3739 | w3740);
assign w3741 = v1012;
assign w3742 = w2576 & ~w3662;
assign v1013 = ~(pi176 | w2576);
assign w3743 = v1013;
assign v1014 = ~(w3742 | w3743);
assign w3744 = v1014;
assign v1015 = ~(w3063 | w3073);
assign w3745 = v1015;
assign v1016 = ~(w3060 | w3068);
assign w3746 = v1016;
assign w3747 = ~w3054 & w3746;
assign v1017 = ~(w3070 | w3072);
assign w3748 = v1017;
assign w3749 = ~w3747 & w3748;
assign w3750 = w3745 & ~w3749;
assign w3751 = ~w3745 & w3749;
assign v1018 = ~(w3750 | w3751);
assign w3752 = v1018;
assign w3753 = w3087 & w3752;
assign w3754 = ~w1815 & w3084;
assign w3755 = pi177 & w3088;
assign v1019 = ~(w1732 | w3754);
assign w3756 = v1019;
assign w3757 = ~w3755 & w3756;
assign w3758 = ~w3753 & w3757;
assign w3759 = ~pi177 & w1732;
assign v1020 = ~(w3093 | w3759);
assign w3760 = v1020;
assign w3761 = ~w3758 & w3760;
assign w3762 = ~w1620 & w3093;
assign w3763 = w1731 & ~w3762;
assign w3764 = ~w3761 & w3763;
assign w3765 = ~pi177 & w1728;
assign v1021 = ~(w3764 | w3765);
assign w3766 = v1021;
assign w3767 = pi178 & pi247;
assign w3768 = w2327 & w2805;
assign w3769 = pi350 & w2892;
assign w3770 = pi178 & ~w2901;
assign w3771 = pi318 & w2901;
assign w3772 = w2810 & ~w3770;
assign w3773 = ~w3771 & w3772;
assign w3774 = ~pi178 & pi344;
assign w3775 = ~pi344 & w903;
assign v1022 = ~(pi243 | w3774);
assign w3776 = v1022;
assign w3777 = ~w3775 & w3776;
assign w3778 = ~w777 & w802;
assign w3779 = pi178 & ~w738;
assign w3780 = w2314 & ~w3779;
assign w3781 = ~w3778 & w3780;
assign w3782 = ~w2810 & w3781;
assign w3783 = ~w2315 & w3782;
assign w3784 = ~w3777 & w3783;
assign v1023 = ~(w2892 | w3773);
assign w3785 = v1023;
assign w3786 = ~w3784 & w3785;
assign v1024 = ~(w2805 | w3769);
assign w3787 = v1024;
assign w3788 = ~w3786 & w3787;
assign v1025 = ~(pi247 | w3768);
assign w3789 = v1025;
assign w3790 = ~w3788 & w3789;
assign w3791 = pi359 & ~w3767;
assign w3792 = ~w3790 & w3791;
assign w3793 = pi179 & w3081;
assign v1026 = ~(w2993 | w3038);
assign w3794 = v1026;
assign v1027 = ~(w2990 | w3068);
assign w3795 = v1027;
assign w3796 = w3794 & w3795;
assign w3797 = ~w3341 & w3796;
assign v1028 = ~(w3046 | w3052);
assign w3798 = v1028;
assign v1029 = ~(w3051 | w3070);
assign w3799 = v1029;
assign w3800 = w3798 & w3799;
assign w3801 = ~w3797 & w3800;
assign w3802 = ~w2985 & w3065;
assign w3803 = ~w3801 & w3802;
assign w3804 = ~w2986 & w3075;
assign w3805 = ~w3803 & w3804;
assign w3806 = w147 & ~w2144;
assign w3807 = pi179 & ~w147;
assign v1030 = ~(w3806 | w3807);
assign w3808 = v1030;
assign w3809 = w2982 & ~w3808;
assign w3810 = ~w2982 & w3808;
assign v1031 = ~(w3809 | w3810);
assign w3811 = v1031;
assign w3812 = w3805 & w3811;
assign v1032 = ~(w3805 | w3811);
assign w3813 = v1032;
assign v1033 = ~(w3812 | w3813);
assign w3814 = v1033;
assign w3815 = w1512 & w3814;
assign v1034 = ~(pi179 | w1512);
assign w3816 = v1034;
assign v1035 = ~(w3081 | w3816);
assign w3817 = v1035;
assign w3818 = ~w3815 & w3817;
assign v1036 = ~(w3084 | w3793);
assign w3819 = v1036;
assign w3820 = ~w3818 & w3819;
assign w3821 = w2144 & w3084;
assign v1037 = ~(w1732 | w3821);
assign w3822 = v1037;
assign w3823 = ~w3820 & w3822;
assign w3824 = pi179 & w1732;
assign v1038 = ~(w3093 | w3824);
assign w3825 = v1038;
assign w3826 = ~w3823 & w3825;
assign w3827 = w2327 & w3093;
assign v1039 = ~(pi247 | w3827);
assign w3828 = v1039;
assign w3829 = ~w3826 & w3828;
assign w3830 = pi179 & pi247;
assign w3831 = pi359 & ~w3830;
assign w3832 = ~w3829 & w3831;
assign w3833 = ~pi180 & pi247;
assign w3834 = ~w2467 & w2805;
assign w3835 = ~pi272 & w1504;
assign v1040 = ~(w1505 | w2460);
assign w3836 = v1040;
assign v1041 = ~(w3835 | w3836);
assign w3837 = v1041;
assign w3838 = w745 & ~w996;
assign w3839 = pi272 & w3838;
assign w3840 = ~pi180 & w734;
assign v1042 = ~(w3839 | w3840);
assign w3841 = v1042;
assign w3842 = ~w2810 & w3841;
assign w3843 = w2459 & w3842;
assign w3844 = ~w3837 & w3843;
assign w3845 = ~pi180 & w1732;
assign w3846 = pi321 & w2901;
assign v1043 = ~(w3157 | w3223);
assign w3847 = v1043;
assign w3848 = pi180 & w3847;
assign w3849 = pi138 & ~w3156;
assign w3850 = ~pi138 & w3222;
assign v1044 = ~(w3849 | w3850);
assign w3851 = v1044;
assign w3852 = w1033 & w3851;
assign w3853 = w3286 & ~w3852;
assign w3854 = ~w3848 & w3853;
assign w3855 = w2810 & ~w3845;
assign w3856 = ~w3846 & w3855;
assign w3857 = ~w3854 & w3856;
assign v1045 = ~(w3844 | w3857);
assign w3858 = v1045;
assign v1046 = ~(w3227 | w3858);
assign w3859 = v1046;
assign w3860 = w2464 & w3227;
assign v1047 = ~(w3859 | w3860);
assign w3861 = v1047;
assign v1048 = ~(w2805 | w3861);
assign w3862 = v1048;
assign v1049 = ~(pi247 | w3834);
assign w3863 = v1049;
assign w3864 = ~w3862 & w3863;
assign w3865 = pi359 & ~w3833;
assign w3866 = ~w3864 & w3865;
assign w3867 = ~pi181 & pi247;
assign w3868 = w2404 & w2805;
assign w3869 = ~pi273 & w1504;
assign v1050 = ~(w1505 | w2395);
assign w3870 = v1050;
assign v1051 = ~(w3869 | w3870);
assign w3871 = v1051;
assign w3872 = ~pi181 & w734;
assign w3873 = pi273 & w3838;
assign v1052 = ~(w3872 | w3873);
assign w3874 = v1052;
assign w3875 = ~w2810 & w3874;
assign w3876 = w2394 & w3875;
assign w3877 = ~w3871 & w3876;
assign w3878 = ~pi181 & w1732;
assign w3879 = ~pi139 & w3222;
assign w3880 = pi139 & ~w3156;
assign v1053 = ~(w3879 | w3880);
assign w3881 = v1053;
assign w3882 = w1033 & w3881;
assign w3883 = pi181 & w3847;
assign w3884 = w3286 & ~w3882;
assign w3885 = ~w3883 & w3884;
assign w3886 = pi315 & w2901;
assign w3887 = w2810 & ~w3878;
assign w3888 = ~w3886 & w3887;
assign w3889 = ~w3885 & w3888;
assign v1054 = ~(w3877 | w3889);
assign w3890 = v1054;
assign v1055 = ~(w3227 | w3890);
assign w3891 = v1055;
assign w3892 = w2523 & w3227;
assign v1056 = ~(w3891 | w3892);
assign w3893 = v1056;
assign v1057 = ~(w2805 | w3893);
assign w3894 = v1057;
assign v1058 = ~(pi247 | w3868);
assign w3895 = v1058;
assign w3896 = ~w3894 & w3895;
assign w3897 = pi359 & ~w3867;
assign w3898 = ~w3896 & w3897;
assign v1059 = ~(w3068 | w3070);
assign w3899 = v1059;
assign w3900 = ~w3054 & w3899;
assign w3901 = w3054 & ~w3899;
assign v1060 = ~(w3900 | w3901);
assign w3902 = v1060;
assign w3903 = w3087 & ~w3902;
assign w3904 = w1969 & w3084;
assign v1061 = ~(w3903 | w3904);
assign w3905 = v1061;
assign v1062 = ~(w1732 | w3905);
assign w3906 = v1062;
assign v1063 = ~(pi182 | w3333);
assign w3907 = v1063;
assign v1064 = ~(w3906 | w3907);
assign w3908 = v1064;
assign v1065 = ~(w3093 | w3908);
assign w3909 = v1065;
assign w3910 = w1697 & w3093;
assign v1066 = ~(pi247 | w3910);
assign w3911 = v1066;
assign w3912 = ~w3909 & w3911;
assign w3913 = pi182 & pi247;
assign w3914 = pi359 & ~w3913;
assign w3915 = ~w3912 & w3914;
assign w3916 = pi183 & w3081;
assign v1067 = ~(w3057 | w3071);
assign w3917 = v1067;
assign w3918 = w3064 & ~w3801;
assign w3919 = w3074 & ~w3918;
assign w3920 = w3917 & ~w3919;
assign w3921 = ~w3917 & w3919;
assign v1068 = ~(w3920 | w3921);
assign w3922 = v1068;
assign w3923 = w1512 & ~w3922;
assign v1069 = ~(pi183 | w1512);
assign w3924 = v1069;
assign v1070 = ~(w3081 | w3924);
assign w3925 = v1070;
assign w3926 = ~w3923 & w3925;
assign v1071 = ~(w3084 | w3916);
assign w3927 = v1071;
assign w3928 = ~w3926 & w3927;
assign w3929 = w1866 & w3084;
assign v1072 = ~(w1732 | w3929);
assign w3930 = v1072;
assign w3931 = ~w3928 & w3930;
assign w3932 = pi183 & w1732;
assign v1073 = ~(w3093 | w3932);
assign w3933 = v1073;
assign w3934 = ~w3931 & w3933;
assign w3935 = w2404 & w3093;
assign v1074 = ~(pi247 | w3935);
assign w3936 = v1074;
assign w3937 = ~w3934 & w3936;
assign w3938 = pi183 & pi247;
assign w3939 = pi359 & ~w3938;
assign w3940 = ~w3937 & w3939;
assign w3941 = ~pi184 & w1728;
assign w3942 = ~w1620 & w2805;
assign w3943 = ~pi184 & w1732;
assign v1075 = ~(pi184 | w3157);
assign w3944 = v1075;
assign w3945 = ~w3287 & w3944;
assign v1076 = ~(w3290 | w3945);
assign w3946 = v1076;
assign v1077 = ~(w2900 | w3946);
assign w3947 = v1077;
assign w3948 = ~pi324 & w2901;
assign v1078 = ~(w3943 | w3948);
assign w3949 = v1078;
assign w3950 = ~w3947 & w3949;
assign w3951 = w2810 & ~w3950;
assign w3952 = pi184 & w734;
assign w3953 = pi243 & ~w670;
assign w3954 = w700 & ~w3953;
assign w3955 = ~w733 & w886;
assign v1079 = ~(w886 | w3276);
assign w3956 = v1079;
assign v1080 = ~(pi243 | w3955);
assign w3957 = v1080;
assign w3958 = ~w3956 & w3957;
assign v1081 = ~(w745 | w3952);
assign w3959 = v1081;
assign w3960 = w2809 & w3959;
assign w3961 = ~w3954 & w3960;
assign w3962 = ~w3958 & w3961;
assign w3963 = w3229 & ~w3962;
assign w3964 = ~w3951 & w3963;
assign w3965 = w1731 & ~w3942;
assign w3966 = ~w3964 & w3965;
assign v1082 = ~(w3941 | w3966);
assign w3967 = v1082;
assign w3968 = pi185 & pi247;
assign w3969 = w2527 & w3093;
assign w3970 = pi185 & ~w3333;
assign w3971 = ~w2282 & w3084;
assign w3972 = ~w3341 & w3794;
assign w3973 = w3798 & ~w3972;
assign v1083 = ~(w2990 | w3051);
assign w3974 = v1083;
assign w3975 = w3973 & w3974;
assign v1084 = ~(w3973 | w3974);
assign w3976 = v1084;
assign v1085 = ~(w3975 | w3976);
assign w3977 = v1085;
assign w3978 = w3087 & ~w3977;
assign v1086 = ~(w3971 | w3978);
assign w3979 = v1086;
assign v1087 = ~(w1732 | w3979);
assign w3980 = v1087;
assign v1088 = ~(w3093 | w3970);
assign w3981 = v1088;
assign w3982 = ~w3980 & w3981;
assign v1089 = ~(pi247 | w3969);
assign w3983 = v1089;
assign w3984 = ~w3982 & w3983;
assign w3985 = pi359 & ~w3968;
assign w3986 = ~w3984 & w3985;
assign w3987 = pi186 & pi247;
assign w3988 = ~w2467 & w3093;
assign v1090 = ~(pi186 | w3333);
assign w3989 = v1090;
assign w3990 = w1753 & w3084;
assign v1091 = ~(w3060 | w3072);
assign w3991 = v1091;
assign w3992 = ~w3801 & w3991;
assign w3993 = w3801 & ~w3991;
assign v1092 = ~(w3992 | w3993);
assign w3994 = v1092;
assign w3995 = w3087 & ~w3994;
assign v1093 = ~(w3990 | w3995);
assign w3996 = v1093;
assign v1094 = ~(w1732 | w3996);
assign w3997 = v1094;
assign v1095 = ~(w3989 | w3997);
assign w3998 = v1095;
assign v1096 = ~(w3093 | w3998);
assign w3999 = v1096;
assign v1097 = ~(pi247 | w3988);
assign w4000 = v1097;
assign w4001 = ~w3999 & w4000;
assign w4002 = pi359 & ~w3987;
assign w4003 = ~w4001 & w4002;
assign w4004 = pi187 & pi247;
assign w4005 = w2648 & w3093;
assign w4006 = pi187 & ~w3333;
assign w4007 = ~w2193 & w3084;
assign v1098 = ~(w2993 | w3052);
assign w4008 = v1098;
assign w4009 = w3049 & w4008;
assign v1099 = ~(w3049 | w4008);
assign w4010 = v1099;
assign v1100 = ~(w4009 | w4010);
assign w4011 = v1100;
assign w4012 = w3087 & ~w4011;
assign v1101 = ~(w4007 | w4012);
assign w4013 = v1101;
assign v1102 = ~(w1732 | w4013);
assign w4014 = v1102;
assign v1103 = ~(w3093 | w4006);
assign w4015 = v1103;
assign w4016 = ~w4014 & w4015;
assign v1104 = ~(pi247 | w4005);
assign w4017 = v1104;
assign w4018 = ~w4016 & w4017;
assign w4019 = pi359 & ~w4004;
assign w4020 = ~w4018 & w4019;
assign w4021 = pi188 & pi356;
assign w4022 = w1728 & w4021;
assign w4023 = pi359 & ~w2733;
assign v1105 = ~(pi188 | w1033);
assign w4024 = v1105;
assign w4025 = ~pi190 & w1109;
assign w4026 = w985 & ~w4025;
assign w4027 = ~pi356 & w4026;
assign w4028 = pi213 & pi214;
assign v1106 = ~(pi213 | pi214);
assign w4029 = v1106;
assign v1107 = ~(w4028 | w4029);
assign w4030 = v1107;
assign w4031 = w4027 & w4030;
assign w4032 = w82 & ~w1107;
assign v1108 = ~(w1334 | w4032);
assign w4033 = v1108;
assign w4034 = w1284 & ~w4033;
assign w4035 = w1033 & ~w4034;
assign v1109 = ~(w2748 | w4035);
assign w4036 = v1109;
assign v1110 = ~(pi356 | w4026);
assign w4037 = v1110;
assign w4038 = pi000 & w101;
assign w4039 = w619 & w4038;
assign w4040 = pi345 & ~w1100;
assign w4041 = ~w4039 & w4040;
assign w4042 = w4037 & w4041;
assign v1111 = ~(w1 | w35);
assign w4043 = v1111;
assign w4044 = w4042 & w4043;
assign v1112 = ~(w4021 | w4031);
assign w4045 = v1112;
assign w4046 = ~w4044 & w4045;
assign w4047 = ~w4036 & w4046;
assign w4048 = w4023 & ~w4024;
assign w4049 = ~w4047 & w4048;
assign v1113 = ~(w4022 | w4049);
assign w4050 = v1113;
assign v1114 = ~(pi189 | w1033);
assign w4051 = v1114;
assign w4052 = pi201 & ~w4029;
assign w4053 = ~pi201 & w4029;
assign v1115 = ~(w4052 | w4053);
assign w4054 = v1115;
assign w4055 = w4027 & w4054;
assign w4056 = ~w36 & w4042;
assign v1116 = ~(w4055 | w4056);
assign w4057 = v1116;
assign w4058 = ~w4036 & w4057;
assign w4059 = w4023 & ~w4051;
assign w4060 = ~w4058 & w4059;
assign w4061 = pi189 & pi356;
assign w4062 = pi359 & w4061;
assign v1117 = ~(w4060 | w4062);
assign w4063 = v1117;
assign w4064 = ~pi190 & w2744;
assign w4065 = pi213 & w985;
assign w4066 = pi190 & w4041;
assign v1118 = ~(w4026 | w4066);
assign w4067 = v1118;
assign v1119 = ~(w4065 | w4067);
assign w4068 = v1119;
assign v1120 = ~(w4034 | w4068);
assign w4069 = v1120;
assign w4070 = pi359 & w2721;
assign w4071 = ~w4069 & w4070;
assign v1121 = ~(w4064 | w4071);
assign w4072 = v1121;
assign w4073 = pi191 & w1728;
assign w4074 = w147 & w986;
assign w4075 = w982 & w1083;
assign v1122 = ~(w4074 | w4075);
assign w4076 = v1122;
assign w4077 = pi191 & w4076;
assign w4078 = ~w3080 & w4074;
assign w4079 = ~w1085 & w1345;
assign w4080 = w9 & w147;
assign w4081 = ~w4079 & w4080;
assign v1123 = ~(w4077 | w4081);
assign w4082 = v1123;
assign w4083 = ~w4078 & w4082;
assign w4084 = ~pi347 & w4081;
assign w4085 = w1731 & ~w4084;
assign w4086 = ~w4083 & w4085;
assign v1124 = ~(w4073 | w4086);
assign w4087 = v1124;
assign w4088 = w47 & w751;
assign w4089 = w161 & w4088;
assign w4090 = w5 & w160;
assign w4091 = ~w751 & w4090;
assign v1125 = ~(w4089 | w4091);
assign w4092 = v1125;
assign w4093 = pi355 & w4092;
assign w4094 = w161 & w3083;
assign w4095 = ~pi192 & pi358;
assign w4096 = ~w4094 & w4095;
assign w4097 = w4092 & w4096;
assign v1126 = ~(w4093 | w4097);
assign w4098 = v1126;
assign w4099 = w4037 & ~w4041;
assign w4100 = w4035 & w4099;
assign w4101 = ~w4098 & w4100;
assign w4102 = w141 & w1048;
assign w4103 = pi193 & w4102;
assign w4104 = w0 & w147;
assign w4105 = w1168 & w4104;
assign w4106 = pi359 & ~w4105;
assign w4107 = w141 & w4094;
assign w4108 = pi192 & ~w4102;
assign w4109 = ~w4107 & w4108;
assign w4110 = ~w4103 & w4106;
assign w4111 = ~w4109 & w4110;
assign w4112 = ~w4101 & w4111;
assign w4113 = pi193 & ~w4107;
assign w4114 = ~pi355 & w4097;
assign w4115 = w4100 & w4114;
assign w4116 = w4106 & ~w4113;
assign w4117 = ~w4115 & w4116;
assign w4118 = ~pi099 & w163;
assign v1127 = ~(pi194 | w983);
assign w4119 = v1127;
assign v1128 = ~(w4118 | w4119);
assign w4120 = v1128;
assign w4121 = ~w4100 & w4120;
assign w4122 = pi359 & ~w4121;
assign w4123 = pi195 & ~w4100;
assign v1129 = ~(w4115 | w4123);
assign w4124 = v1129;
assign w4125 = pi359 & ~w4124;
assign w4126 = ~w4093 & w4100;
assign v1130 = ~(pi196 | w4100);
assign w4127 = v1130;
assign w4128 = pi359 & ~w4126;
assign w4129 = ~w4127 & w4128;
assign w4130 = w70 & w1229;
assign w4131 = w117 & w4130;
assign w4132 = w24 & w4131;
assign v1131 = ~(w1249 | w4132);
assign w4133 = v1131;
assign w4134 = pi301 & ~w4133;
assign w4135 = ~pi190 & w110;
assign v1132 = ~(w1187 | w4135);
assign w4136 = v1132;
assign w4137 = w24 & w1081;
assign w4138 = ~w4136 & w4137;
assign v1133 = ~(w4134 | w4138);
assign w4139 = v1133;
assign w4140 = w9 & w1231;
assign v1134 = ~(w102 | w4140);
assign w4141 = v1134;
assign w4142 = ~w1249 & w4141;
assign w4143 = pi297 & pi298;
assign w4144 = w101 & ~w998;
assign w4145 = w1234 & w4144;
assign v1135 = ~(w4131 | w4145);
assign w4146 = v1135;
assign w4147 = pi302 & ~w4143;
assign w4148 = ~w4146 & w4147;
assign w4149 = w4142 & ~w4148;
assign w4150 = pi301 & ~w4149;
assign v1136 = ~(w1131 | w1203);
assign w4151 = v1136;
assign w4152 = w101 & w996;
assign w4153 = pi300 & w4152;
assign w4154 = ~w1174 & w4151;
assign w4155 = ~w4153 & w4154;
assign w4156 = w101 & w1153;
assign v1137 = ~(w1162 | w4156);
assign w4157 = v1137;
assign w4158 = w101 & w1156;
assign v1138 = ~(w1137 | w4158);
assign w4159 = v1138;
assign w4160 = w4157 & w4159;
assign w4161 = w8 & w1187;
assign w4162 = ~pi298 & w4161;
assign v1139 = ~(w111 | w4162);
assign w4163 = v1139;
assign w4164 = w4160 & w4163;
assign w4165 = pi302 & ~w4164;
assign w4166 = w4155 & ~w4165;
assign w4167 = w0 & ~w4166;
assign w4168 = pi297 & w1109;
assign v1140 = ~(w4150 | w4168);
assign w4169 = v1140;
assign w4170 = ~w4167 & w4169;
assign w4171 = pi296 & w1109;
assign w4172 = pi190 & ~w24;
assign w4173 = ~pi190 & w24;
assign v1141 = ~(w4172 | w4173);
assign w4174 = v1141;
assign w4175 = w4131 & w4174;
assign w4176 = w4141 & ~w4175;
assign w4177 = pi301 & ~w4176;
assign w4178 = w1040 & w1136;
assign w4179 = pi303 & w1234;
assign v1142 = ~(w4178 | w4179);
assign w4180 = v1142;
assign w4181 = w2726 & ~w4180;
assign w4182 = w111 & ~w4172;
assign w4183 = w4161 & w4174;
assign w4184 = w69 & w101;
assign w4185 = ~w1161 & w4159;
assign w4186 = pi303 & ~w4185;
assign w4187 = pi303 & w1210;
assign w4188 = w70 & w4187;
assign w4189 = w8 & w1206;
assign v1143 = ~(w4188 | w4189);
assign w4190 = v1143;
assign v1144 = ~(pi190 | w4190);
assign w4191 = v1144;
assign v1145 = ~(w4182 | w4184);
assign w4192 = v1145;
assign w4193 = ~w4183 & w4192;
assign w4194 = w4155 & w4193;
assign w4195 = ~w4186 & w4194;
assign w4196 = ~w4191 & w4195;
assign w4197 = w0 & ~w4196;
assign v1146 = ~(w4171 | w4181);
assign w4198 = v1146;
assign w4199 = ~w4177 & w4198;
assign w4200 = ~w4197 & w4199;
assign v1147 = ~(w4170 | w4200);
assign w4201 = v1147;
assign w4202 = w8 & w4178;
assign v1148 = ~(w4140 | w4202);
assign w4203 = v1148;
assign w4204 = pi296 & pi302;
assign w4205 = pi298 & ~w4204;
assign w4206 = ~w4146 & w4205;
assign w4207 = ~w102 & w4203;
assign w4208 = ~w4206 & w4207;
assign w4209 = pi301 & ~w4208;
assign w4210 = pi291 & w1109;
assign w4211 = w4155 & ~w4189;
assign w4212 = pi298 & ~w4160;
assign v1149 = ~(w111 | w4161);
assign w4213 = v1149;
assign w4214 = pi190 & pi298;
assign w4215 = w110 & w4214;
assign v1150 = ~(w157 | w4215);
assign w4216 = v1150;
assign v1151 = ~(w4213 | w4216);
assign w4217 = v1151;
assign v1152 = ~(w2 | w101);
assign w4218 = v1152;
assign w4219 = w69 & ~w4218;
assign v1153 = ~(w4188 | w4219);
assign w4220 = v1153;
assign w4221 = w4211 & ~w4217;
assign w4222 = w4220 & w4221;
assign w4223 = ~w4212 & w4222;
assign w4224 = w0 & ~w4223;
assign v1154 = ~(w4209 | w4210);
assign w4225 = v1154;
assign w4226 = ~w4224 & w4225;
assign w4227 = ~w4201 & w4226;
assign v1155 = ~(w4139 | w4227);
assign w4228 = v1155;
assign v1156 = ~(pi247 | w4228);
assign w4229 = v1156;
assign w4230 = pi197 & ~w4229;
assign v1157 = ~(w4170 | w4226);
assign w4231 = v1157;
assign w4232 = ~w4200 & w4231;
assign w4233 = pi126 & w4232;
assign w4234 = w411 & w4200;
assign w4235 = w4139 & ~w4231;
assign w4236 = w336 & ~w4200;
assign w4237 = ~w4234 & w4235;
assign w4238 = ~w4236 & w4237;
assign w4239 = w4200 & w4231;
assign w4240 = pi354 & w4239;
assign w4241 = ~w4139 & w4170;
assign w4242 = ~w4200 & w4241;
assign w4243 = pi187 & w4242;
assign w4244 = w4200 & w4241;
assign w4245 = pi174 & w4244;
assign v1158 = ~(w4233 | w4240);
assign w4246 = v1158;
assign v1159 = ~(w4243 | w4245);
assign w4247 = v1159;
assign w4248 = w4246 & w4247;
assign w4249 = ~w4238 & w4248;
assign v1160 = ~(pi247 | w4249);
assign w4250 = v1160;
assign v1161 = ~(w4230 | w4250);
assign w4251 = v1161;
assign w4252 = pi198 & ~w4229;
assign w4253 = pi139 & w4232;
assign w4254 = w430 & w4200;
assign w4255 = w257 & ~w4200;
assign w4256 = w4235 & ~w4255;
assign w4257 = ~w4254 & w4256;
assign w4258 = pi353 & w4239;
assign w4259 = pi183 & w4242;
assign w4260 = pi144 & w4244;
assign v1162 = ~(w4253 | w4258);
assign w4261 = v1162;
assign v1163 = ~(w4259 | w4260);
assign w4262 = v1163;
assign w4263 = w4261 & w4262;
assign w4264 = ~w4257 & w4263;
assign v1164 = ~(pi247 | w4264);
assign w4265 = v1164;
assign v1165 = ~(w4252 | w4265);
assign w4266 = v1165;
assign w4267 = ~pi199 & pi247;
assign w4268 = w613 & w615;
assign w4269 = w1179 & ~w4268;
assign w4270 = (w1082 & ~w1179) | (w1082 & w6134) | (~w1179 & w6134);
assign v1166 = ~(pi228 | w4270);
assign w4271 = v1166;
assign w4272 = ~pi350 & w4270;
assign v1167 = ~(w4271 | w4272);
assign w4273 = v1167;
assign v1168 = ~(pi199 | w4273);
assign w4274 = v1168;
assign w4275 = pi199 & w4273;
assign v1169 = ~(w4274 | w4275);
assign w4276 = v1169;
assign w4277 = pi200 & w4273;
assign v1170 = ~(pi212 | w4273);
assign w4278 = v1170;
assign v1171 = ~(pi200 | w4273);
assign w4279 = v1171;
assign w4280 = ~pi347 & w4270;
assign v1172 = ~(w4271 | w4280);
assign w4281 = v1172;
assign v1173 = ~(pi211 | w4281);
assign w4282 = v1173;
assign w4283 = ~pi353 & w4270;
assign v1174 = ~(w4271 | w4283);
assign w4284 = v1174;
assign v1175 = ~(pi210 | w4284);
assign w4285 = v1175;
assign w4286 = ~pi348 & w4270;
assign v1176 = ~(w4271 | w4286);
assign w4287 = v1176;
assign w4288 = pi208 & w4287;
assign v1177 = ~(pi208 | w4287);
assign w4289 = v1177;
assign v1178 = ~(w4288 | w4289);
assign w4290 = v1178;
assign w4291 = ~pi351 & w4270;
assign v1179 = ~(w4271 | w4291);
assign w4292 = v1179;
assign w4293 = pi207 & w4292;
assign v1180 = ~(pi207 | w4292);
assign w4294 = v1180;
assign v1181 = ~(w4293 | w4294);
assign w4295 = v1181;
assign w4296 = ~pi349 & w4270;
assign v1182 = ~(w4271 | w4296);
assign w4297 = v1182;
assign w4298 = pi206 & w4297;
assign w4299 = pi354 & w4270;
assign v1183 = ~(w4271 | w4299);
assign w4300 = v1183;
assign w4301 = pi220 & ~w4300;
assign v1184 = ~(pi206 | w4297);
assign w4302 = v1184;
assign v1185 = ~(w4298 | w4302);
assign w4303 = v1185;
assign w4304 = w4301 & w4303;
assign w4305 = (~w4298 & ~w4303) | (~w4298 & w6135) | (~w4303 & w6135);
assign w4306 = w4295 & ~w4305;
assign w4307 = (~w4293 & w4305) | (~w4293 & w6172) | (w4305 & w6172);
assign w4308 = w4290 & ~w4307;
assign w4309 = (~w4288 & w4307) | (~w4288 & w6220) | (w4307 & w6220);
assign w4310 = ~pi352 & w4270;
assign v1186 = ~(w4271 | w4310);
assign w4311 = v1186;
assign v1187 = ~(pi209 | w4311);
assign w4312 = v1187;
assign v1188 = ~(w4312 | w4309);
assign w4313 = v1188;
assign w4314 = pi210 & w4284;
assign w4315 = pi209 & w4311;
assign v1189 = ~(w4314 | w4315);
assign w4316 = v1189;
assign w4317 = (~w4285 & w4313) | (~w4285 & w7337) | (w4313 & w7337);
assign w4318 = pi211 & w4281;
assign v1190 = ~(w4282 | w4318);
assign w4319 = v1190;
assign w4320 = ~w4317 & w4319;
assign v1191 = ~(w4282 | w4320);
assign w4321 = v1191;
assign w4322 = ~w4279 & w4321;
assign w4323 = ~w4278 & w4322;
assign w4324 = pi212 & w4273;
assign v1192 = ~(w4277 | w4324);
assign w4325 = v1192;
assign w4326 = ~w4323 & w4325;
assign w4327 = ~w4276 & w4326;
assign w4328 = w4276 & ~w4326;
assign v1193 = ~(w4327 | w4328);
assign w4329 = v1193;
assign w4330 = w0 & w1167;
assign w4331 = pi230 & w38;
assign w4332 = ~w4330 & w4331;
assign w4333 = ~w1086 & w4332;
assign w4334 = w7368 & w4333;
assign w4335 = w982 & w4334;
assign w4336 = ~w4329 & w4335;
assign v1194 = ~(pi199 | w4335);
assign w4337 = v1194;
assign w4338 = w1732 & ~w4337;
assign w4339 = ~w4336 & w4338;
assign w4340 = w99 & w1243;
assign w4341 = ~w1105 & w1259;
assign w4342 = w985 & ~w4341;
assign w4343 = w2 & w1038;
assign v1195 = ~(w84 | w88);
assign w4344 = v1195;
assign w4345 = w4152 & w4344;
assign v1196 = ~(pi190 | w1190);
assign w4346 = v1196;
assign w4347 = w1084 & w1270;
assign w4348 = w4269 & w4347;
assign w4349 = w1269 & ~w4346;
assign w4350 = w4348 & w4349;
assign w4351 = w8 & ~w4350;
assign v1197 = ~(w4343 | w4345);
assign w4352 = v1197;
assign w4353 = ~w4351 & w4352;
assign w4354 = w0 & ~w4353;
assign v1198 = ~(pi228 | w4340);
assign w4355 = v1198;
assign w4356 = ~w4342 & w4355;
assign w4357 = ~w4354 & w4356;
assign w4358 = w982 & ~w4357;
assign w4359 = ~w4329 & w4358;
assign w4360 = pi199 & w1756;
assign w4361 = w2303 & ~w4360;
assign w4362 = w2284 & ~w4361;
assign w4363 = pi199 & ~w1033;
assign v1199 = ~(w2266 | w4358);
assign w4364 = v1199;
assign w4365 = ~w4363 & w4364;
assign w4366 = ~w4362 & w4365;
assign v1200 = ~(w1732 | w4366);
assign w4367 = v1200;
assign w4368 = ~w4359 & w4367;
assign v1201 = ~(pi247 | w4339);
assign w4369 = v1201;
assign w4370 = ~w4368 & w4369;
assign w4371 = pi359 & ~w4267;
assign w4372 = ~w4370 & w4371;
assign w4373 = ~pi200 & pi247;
assign v1202 = ~(w4277 | w4279);
assign w4374 = v1202;
assign w4375 = ~w4321 & w4374;
assign w4376 = w4321 & ~w4374;
assign v1203 = ~(w4375 | w4376);
assign w4377 = v1203;
assign w4378 = w4335 & w4377;
assign v1204 = ~(pi200 | w4335);
assign w4379 = v1204;
assign w4380 = w1732 & ~w4379;
assign w4381 = ~w4378 & w4380;
assign w4382 = pi200 & ~w1033;
assign w4383 = pi200 & w1756;
assign w4384 = w2243 & ~w4383;
assign w4385 = w2242 & ~w4384;
assign v1205 = ~(w2255 | w4358);
assign w4386 = v1205;
assign w4387 = ~w4382 & w4386;
assign w4388 = ~w4385 & w4387;
assign w4389 = w4358 & w4377;
assign v1206 = ~(w1732 | w4388);
assign w4390 = v1206;
assign w4391 = ~w4389 & w4390;
assign v1207 = ~(pi247 | w4381);
assign w4392 = v1207;
assign w4393 = ~w4391 & w4392;
assign w4394 = pi359 & ~w4373;
assign w4395 = ~w4393 & w4394;
assign w4396 = w2721 & w4034;
assign w4397 = ~pi189 & w4396;
assign w4398 = pi201 & ~w4396;
assign w4399 = pi359 & ~w4397;
assign w4400 = ~w4398 & w4399;
assign w4401 = pi202 & ~w4229;
assign w4402 = pi138 & w4232;
assign w4403 = w463 & w4200;
assign w4404 = w298 & ~w4200;
assign w4405 = w4235 & ~w4404;
assign w4406 = ~w4403 & w4405;
assign w4407 = pi186 & w4242;
assign w4408 = pi173 & w4244;
assign w4409 = pi348 & w4239;
assign v1208 = ~(w4402 | w4407);
assign w4410 = v1208;
assign v1209 = ~(w4408 | w4409);
assign w4411 = v1209;
assign w4412 = w4410 & w4411;
assign w4413 = ~w4406 & w4412;
assign v1210 = ~(pi247 | w4413);
assign w4414 = v1210;
assign v1211 = ~(w4401 | w4414);
assign w4415 = v1211;
assign w4416 = ~pi203 & pi247;
assign v1212 = ~(pi203 | w4273);
assign w4417 = v1212;
assign w4418 = pi203 & w4273;
assign v1213 = ~(w4417 | w4418);
assign w4419 = v1213;
assign v1214 = ~(pi221 | w4273);
assign w4420 = v1214;
assign v1215 = ~(w4274 | w4278);
assign w4421 = v1215;
assign w4422 = ~w4420 & w4421;
assign w4423 = w4322 & w4422;
assign v1216 = ~(w4275 | w4324);
assign w4424 = v1216;
assign w4425 = pi221 & w4273;
assign v1217 = ~(w4277 | w4425);
assign w4426 = v1217;
assign w4427 = w4424 & w4426;
assign w4428 = ~w4423 & w4427;
assign w4429 = ~w4419 & w4428;
assign w4430 = w4419 & ~w4428;
assign v1218 = ~(w4429 | w4430);
assign w4431 = v1218;
assign w4432 = w4335 & ~w4431;
assign v1219 = ~(pi203 | w4335);
assign w4433 = v1219;
assign w4434 = w1732 & ~w4433;
assign w4435 = ~w4432 & w4434;
assign w4436 = pi203 & w1756;
assign w4437 = w1787 & ~w4436;
assign w4438 = w1755 & ~w4437;
assign w4439 = pi203 & ~w1033;
assign v1220 = ~(w1736 | w4358);
assign w4440 = v1220;
assign w4441 = ~w4439 & w4440;
assign w4442 = ~w4438 & w4441;
assign w4443 = w4358 & ~w4431;
assign v1221 = ~(w1732 | w4442);
assign w4444 = v1221;
assign w4445 = ~w4443 & w4444;
assign v1222 = ~(pi247 | w4435);
assign w4446 = v1222;
assign w4447 = ~w4445 & w4446;
assign w4448 = pi359 & ~w4416;
assign w4449 = ~w4447 & w4448;
assign w4450 = ~pi204 & pi247;
assign w4451 = pi204 & w4273;
assign v1223 = ~(pi204 | w4273);
assign w4452 = v1223;
assign v1224 = ~(w4451 | w4452);
assign w4453 = v1224;
assign v1225 = ~(w4279 | w4282);
assign w4454 = v1225;
assign w4455 = w4317 & w4454;
assign w4456 = ~w4279 & w4318;
assign v1226 = ~(w4277 | w4456);
assign w4457 = v1226;
assign w4458 = ~w4455 & w4457;
assign w4459 = w4421 & ~w4458;
assign w4460 = w4424 & ~w4459;
assign v1227 = ~(w4417 | w4420);
assign w4461 = v1227;
assign w4462 = ~w4460 & w4461;
assign v1228 = ~(w4418 | w4425);
assign w4463 = v1228;
assign w4464 = ~w4462 & w4463;
assign w4465 = w4453 & ~w4464;
assign w4466 = ~w4453 & w4464;
assign v1229 = ~(w4465 | w4466);
assign w4467 = v1229;
assign w4468 = w4335 & ~w4467;
assign v1230 = ~(pi204 | w4335);
assign w4469 = v1230;
assign w4470 = w1732 & ~w4469;
assign w4471 = ~w4468 & w4470;
assign w4472 = pi204 & w1756;
assign w4473 = w1838 & ~w4472;
assign w4474 = w1817 & ~w4473;
assign w4475 = pi204 & ~w1033;
assign v1231 = ~(w1799 | w4358);
assign w4476 = v1231;
assign w4477 = ~w4475 & w4476;
assign w4478 = ~w4474 & w4477;
assign w4479 = w4358 & ~w4467;
assign v1232 = ~(w1732 | w4478);
assign w4480 = v1232;
assign w4481 = ~w4479 & w4480;
assign v1233 = ~(pi247 | w4471);
assign w4482 = v1233;
assign w4483 = ~w4481 & w4482;
assign w4484 = pi359 & ~w4450;
assign w4485 = ~w4483 & w4484;
assign w4486 = ~pi205 & pi247;
assign v1234 = ~(pi247 | w1732);
assign w4487 = v1234;
assign w4488 = pi205 & w4273;
assign v1235 = ~(pi205 | w4273);
assign w4489 = v1235;
assign v1236 = ~(w4488 | w4489);
assign w4490 = v1236;
assign v1237 = ~(w4418 | w4451);
assign w4491 = v1237;
assign v1238 = ~(w4417 | w4428);
assign w4492 = v1238;
assign w4493 = ~w4452 & w4492;
assign w4494 = w4491 & ~w4493;
assign w4495 = ~w4490 & w4494;
assign w4496 = w4490 & ~w4494;
assign v1239 = ~(w4495 | w4496);
assign w4497 = v1239;
assign w4498 = w4358 & ~w4497;
assign w4499 = pi205 & ~w1033;
assign w4500 = pi205 & w1756;
assign w4501 = w1889 & ~w4500;
assign w4502 = w1868 & ~w4501;
assign v1240 = ~(w1850 | w4358);
assign w4503 = v1240;
assign w4504 = ~w4499 & w4503;
assign w4505 = ~w4502 & w4504;
assign v1241 = ~(w4498 | w4505);
assign w4506 = v1241;
assign w4507 = w4487 & ~w4506;
assign v1242 = ~(pi205 | w4334);
assign w4508 = v1242;
assign w4509 = w4334 & ~w4497;
assign w4510 = w982 & ~w4508;
assign w4511 = ~w4509 & w4510;
assign w4512 = pi205 & ~w982;
assign v1243 = ~(pi247 | w4512);
assign w4513 = v1243;
assign w4514 = w1732 & w4513;
assign w4515 = ~w4511 & w4514;
assign w4516 = pi359 & ~w4486;
assign w4517 = ~w4507 & w4516;
assign w4518 = ~w4515 & w4517;
assign w4519 = ~pi206 & pi247;
assign v1244 = ~(w4301 | w4303);
assign w4520 = v1244;
assign v1245 = ~(w4304 | w4520);
assign w4521 = v1245;
assign w4522 = w4335 & ~w4521;
assign v1246 = ~(pi206 | w4335);
assign w4523 = v1246;
assign w4524 = w1732 & ~w4522;
assign w4525 = ~w4523 & w4524;
assign w4526 = w4358 & ~w4521;
assign w4527 = pi206 & ~w1033;
assign w4528 = pi206 & w1088;
assign w4529 = w1103 & ~w4528;
assign v1247 = ~(w1052 | w4529);
assign w4530 = v1247;
assign w4531 = w1077 & ~w4530;
assign w4532 = w1050 & ~w4531;
assign v1248 = ~(w4358 | w4527);
assign w4533 = v1248;
assign w4534 = ~w4532 & w4533;
assign v1249 = ~(w1732 | w4526);
assign w4535 = v1249;
assign w4536 = ~w4534 & w4535;
assign v1250 = ~(pi247 | w4525);
assign w4537 = v1250;
assign w4538 = ~w4536 & w4537;
assign w4539 = pi359 & ~w4519;
assign w4540 = ~w4538 & w4539;
assign w4541 = ~pi207 & pi247;
assign w4542 = ~w4295 & w4305;
assign v1251 = ~(w4306 | w4542);
assign w4543 = v1251;
assign w4544 = w4335 & ~w4543;
assign v1252 = ~(pi207 | w4335);
assign w4545 = v1252;
assign w4546 = w1732 & ~w4545;
assign w4547 = ~w4544 & w4546;
assign w4548 = w4358 & ~w4543;
assign w4549 = pi207 & ~w1033;
assign w4550 = pi207 & w1088;
assign w4551 = w1384 & ~w4550;
assign v1253 = ~(w1052 | w4551);
assign w4552 = v1253;
assign w4553 = w1382 & ~w4552;
assign w4554 = w1365 & ~w4553;
assign v1254 = ~(w4358 | w4549);
assign w4555 = v1254;
assign w4556 = ~w4554 & w4555;
assign v1255 = ~(w1732 | w4548);
assign w4557 = v1255;
assign w4558 = ~w4556 & w4557;
assign v1256 = ~(pi247 | w4547);
assign w4559 = v1256;
assign w4560 = ~w4558 & w4559;
assign w4561 = pi359 & ~w4541;
assign w4562 = ~w4560 & w4561;
assign w4563 = pi208 & w1728;
assign v1257 = ~(pi208 | w4335);
assign w4564 = v1257;
assign w4565 = ~w4290 & w4307;
assign v1258 = ~(w4308 | w4565);
assign w4566 = v1258;
assign w4567 = w4335 & ~w4566;
assign w4568 = w1732 & ~w4564;
assign w4569 = ~w4567 & w4568;
assign w4570 = pi208 & ~w1033;
assign w4571 = pi208 & w1756;
assign w4572 = w2105 & ~w4571;
assign w4573 = w2104 & ~w4572;
assign v1259 = ~(w2086 | w4358);
assign w4574 = v1259;
assign w4575 = ~w4570 & w4574;
assign w4576 = ~w4573 & w4575;
assign w4577 = w4358 & ~w4566;
assign v1260 = ~(w1732 | w4577);
assign w4578 = v1260;
assign w4579 = ~w4576 & w4578;
assign v1261 = ~(w4569 | w4579);
assign w4580 = v1261;
assign w4581 = w1731 & ~w4580;
assign v1262 = ~(w4563 | w4581);
assign w4582 = v1262;
assign w4583 = ~pi209 & pi247;
assign v1263 = ~(w4312 | w4315);
assign w4584 = v1263;
assign w4585 = w4309 & ~w4584;
assign w4586 = ~w4309 & w4584;
assign v1264 = ~(w4585 | w4586);
assign w4587 = v1264;
assign w4588 = w4335 & ~w4587;
assign v1265 = ~(pi209 | w4335);
assign w4589 = v1265;
assign w4590 = w1732 & ~w4589;
assign w4591 = ~w4588 & w4590;
assign w4592 = pi209 & w1756;
assign w4593 = w2022 & ~w4592;
assign w4594 = w2020 & ~w4593;
assign w4595 = pi209 & ~w1033;
assign v1266 = ~(w2002 | w4358);
assign w4596 = v1266;
assign w4597 = ~w4595 & w4596;
assign w4598 = ~w4594 & w4597;
assign w4599 = w4358 & ~w4587;
assign v1267 = ~(w1732 | w4598);
assign w4600 = v1267;
assign w4601 = ~w4599 & w4600;
assign v1268 = ~(pi247 | w4591);
assign w4602 = v1268;
assign w4603 = ~w4601 & w4602;
assign w4604 = pi359 & ~w4583;
assign w4605 = ~w4603 & w4604;
assign w4606 = ~pi210 & pi247;
assign v1269 = ~(w4285 | w4314);
assign w4607 = v1269;
assign v1270 = ~(w4313 | w4315);
assign w4608 = v1270;
assign w4609 = ~w4607 & w4608;
assign w4610 = w4607 & ~w4608;
assign v1271 = ~(w4609 | w4610);
assign w4611 = v1271;
assign w4612 = w4358 & ~w4611;
assign w4613 = pi210 & w1088;
assign w4614 = w1428 & ~w4613;
assign v1272 = ~(w1052 | w4614);
assign w4615 = v1272;
assign w4616 = w1426 & ~w4615;
assign w4617 = w1409 & ~w4616;
assign w4618 = pi210 & ~w1033;
assign v1273 = ~(w4358 | w4618);
assign w4619 = v1273;
assign v1274 = ~(w1732 | w4619);
assign w4620 = v1274;
assign v1275 = ~(w4617 | w4620);
assign w4621 = v1275;
assign v1276 = ~(w4612 | w4621);
assign w4622 = v1276;
assign v1277 = ~(pi210 | w4335);
assign w4623 = v1277;
assign w4624 = w4335 & ~w4611;
assign w4625 = w1732 & ~w4623;
assign w4626 = ~w4624 & w4625;
assign v1278 = ~(pi247 | w4622);
assign w4627 = v1278;
assign w4628 = ~w4626 & w4627;
assign w4629 = pi359 & ~w4606;
assign w4630 = ~w4628 & w4629;
assign w4631 = ~pi211 & pi247;
assign w4632 = w4317 & ~w4319;
assign v1279 = ~(w4320 | w4632);
assign w4633 = v1279;
assign w4634 = w4358 & w4633;
assign w4635 = pi211 & w1088;
assign w4636 = w1475 & ~w4635;
assign v1280 = ~(w1052 | w4636);
assign w4637 = v1280;
assign w4638 = w1473 & ~w4637;
assign w4639 = w1456 & ~w4638;
assign w4640 = pi211 & ~w1033;
assign v1281 = ~(w4358 | w4640);
assign w4641 = v1281;
assign v1282 = ~(w1732 | w4641);
assign w4642 = v1282;
assign v1283 = ~(w4639 | w4642);
assign w4643 = v1283;
assign v1284 = ~(w4634 | w4643);
assign w4644 = v1284;
assign v1285 = ~(pi211 | w4335);
assign w4645 = v1285;
assign w4646 = w4335 & w4633;
assign w4647 = w1732 & ~w4645;
assign w4648 = ~w4646 & w4647;
assign v1286 = ~(pi247 | w4644);
assign w4649 = v1286;
assign w4650 = ~w4648 & w4649;
assign w4651 = pi359 & ~w4631;
assign w4652 = ~w4650 & w4651;
assign w4653 = ~pi212 & pi247;
assign v1287 = ~(w4278 | w4324);
assign w4654 = v1287;
assign w4655 = ~w4458 & w4654;
assign w4656 = w4458 & ~w4654;
assign v1288 = ~(w4655 | w4656);
assign w4657 = v1288;
assign w4658 = w4335 & ~w4657;
assign v1289 = ~(pi212 | w4335);
assign w4659 = v1289;
assign w4660 = w1732 & ~w4659;
assign w4661 = ~w4658 & w4660;
assign w4662 = pi212 & w1756;
assign w4663 = w2215 & ~w4662;
assign w4664 = w2195 & ~w4663;
assign w4665 = pi212 & ~w1033;
assign v1290 = ~(w2177 | w4358);
assign w4666 = v1290;
assign w4667 = ~w4665 & w4666;
assign w4668 = ~w4664 & w4667;
assign w4669 = w4358 & ~w4657;
assign v1291 = ~(w1732 | w4668);
assign w4670 = v1291;
assign w4671 = ~w4669 & w4670;
assign v1292 = ~(pi247 | w4661);
assign w4672 = v1292;
assign w4673 = ~w4671 & w4672;
assign w4674 = pi359 & ~w4653;
assign w4675 = ~w4673 & w4674;
assign w4676 = ~pi190 & w4396;
assign w4677 = pi213 & ~w4396;
assign w4678 = pi359 & ~w4676;
assign w4679 = ~w4677 & w4678;
assign w4680 = ~pi188 & w4396;
assign w4681 = pi214 & ~w4396;
assign w4682 = pi359 & ~w4680;
assign w4683 = ~w4681 & w4682;
assign w4684 = pi215 & ~w4229;
assign w4685 = pi141 & w4232;
assign w4686 = w446 & w4200;
assign w4687 = w278 & ~w4200;
assign w4688 = w4235 & ~w4687;
assign w4689 = ~w4686 & w4688;
assign w4690 = pi172 & w4244;
assign w4691 = pi351 & w4239;
assign w4692 = pi182 & w4242;
assign v1293 = ~(w4685 | w4690);
assign w4693 = v1293;
assign v1294 = ~(w4691 | w4692);
assign w4694 = v1294;
assign w4695 = w4693 & w4694;
assign w4696 = ~w4689 & w4695;
assign v1295 = ~(pi247 | w4696);
assign w4697 = v1295;
assign v1296 = ~(w4684 | w4697);
assign w4698 = v1296;
assign w4699 = pi216 & ~w4229;
assign w4700 = pi143 & w4232;
assign w4701 = w479 & w4200;
assign w4702 = w237 & ~w4200;
assign w4703 = w4235 & ~w4702;
assign w4704 = ~w4701 & w4703;
assign w4705 = pi146 & w4244;
assign w4706 = pi352 & w4239;
assign w4707 = pi177 & w4242;
assign v1297 = ~(w4700 | w4705);
assign w4708 = v1297;
assign v1298 = ~(w4706 | w4707);
assign w4709 = v1298;
assign w4710 = w4708 & w4709;
assign w4711 = ~w4704 & w4710;
assign v1299 = ~(pi247 | w4711);
assign w4712 = v1299;
assign v1300 = ~(w4699 | w4712);
assign w4713 = v1300;
assign w4714 = pi217 & ~w4229;
assign w4715 = pi140 & w4232;
assign w4716 = w214 & w4200;
assign w4717 = w362 & ~w4200;
assign w4718 = w4235 & ~w4716;
assign w4719 = ~w4717 & w4718;
assign w4720 = pi347 & w4239;
assign w4721 = pi137 & w4244;
assign w4722 = pi117 & w4242;
assign v1301 = ~(w4715 | w4720);
assign w4723 = v1301;
assign v1302 = ~(w4721 | w4722);
assign w4724 = v1302;
assign w4725 = w4723 & w4724;
assign w4726 = ~w4719 & w4725;
assign v1303 = ~(pi247 | w4726);
assign w4727 = v1303;
assign v1304 = ~(w4714 | w4727);
assign w4728 = v1304;
assign v1305 = ~(pi219 | w4273);
assign w4729 = v1305;
assign v1306 = ~(w4452 | w4489);
assign w4730 = v1306;
assign w4731 = ~w4729 & w4730;
assign w4732 = w4492 & w4731;
assign w4733 = pi219 & w4273;
assign v1307 = ~(w4488 | w4733);
assign w4734 = v1307;
assign w4735 = w4491 & w4734;
assign w4736 = ~w4732 & w4735;
assign w4737 = pi218 & ~w4273;
assign w4738 = ~pi218 & w4273;
assign v1308 = ~(w4737 | w4738);
assign w4739 = v1308;
assign w4740 = w4736 & ~w4739;
assign w4741 = w1732 & ~w4334;
assign w4742 = ~w1732 & w4357;
assign w4743 = w982 & ~w4741;
assign w4744 = ~w4742 & w4743;
assign w4745 = ~w4736 & w4739;
assign w4746 = ~pi247 & w4744;
assign w4747 = ~w4740 & w4746;
assign w4748 = ~w4745 & w4747;
assign w4749 = pi218 & w1756;
assign w4750 = w2166 & ~w4749;
assign w4751 = w7368 & ~w2145;
assign w4752 = ~w4750 & w4751;
assign w4753 = w4487 & ~w4752;
assign w4754 = w2128 & w4753;
assign v1309 = ~(w1033 | w4744);
assign w4755 = v1309;
assign v1310 = ~(pi247 | w4755);
assign w4756 = v1310;
assign v1311 = ~(pi218 | w4756);
assign w4757 = v1311;
assign w4758 = pi359 & ~w4754;
assign w4759 = ~w4757 & w4758;
assign w4760 = ~w4748 & w4759;
assign v1312 = ~(w4729 | w4733);
assign w4761 = v1312;
assign w4762 = ~w4451 & w4464;
assign w4763 = w4730 & ~w4762;
assign v1313 = ~(w4488 | w4763);
assign w4764 = v1313;
assign w4765 = ~w4761 & w4764;
assign w4766 = w4761 & ~w4764;
assign v1314 = ~(w4765 | w4766);
assign w4767 = v1314;
assign w4768 = w4335 & ~w4767;
assign v1315 = ~(pi219 | w4335);
assign w4769 = v1315;
assign w4770 = w1732 & ~w4769;
assign w4771 = ~w4768 & w4770;
assign w4772 = w4358 & ~w4767;
assign w4773 = pi219 & w1756;
assign w4774 = w1940 & ~w4773;
assign w4775 = w1919 & ~w4774;
assign w4776 = pi219 & ~w1033;
assign v1316 = ~(w1901 | w4358);
assign w4777 = v1316;
assign w4778 = ~w4776 & w4777;
assign w4779 = ~w4775 & w4778;
assign v1317 = ~(w1732 | w4779);
assign w4780 = v1317;
assign w4781 = ~w4772 & w4780;
assign v1318 = ~(pi247 | w4771);
assign w4782 = v1318;
assign w4783 = ~w4781 & w4782;
assign w4784 = ~pi219 & pi247;
assign w4785 = pi359 & ~w4784;
assign w4786 = ~w4783 & w4785;
assign w4787 = ~pi220 & pi247;
assign v1319 = ~(pi220 | w4335);
assign w4788 = v1319;
assign w4789 = ~pi220 & w4300;
assign v1320 = ~(w4301 | w4789);
assign w4790 = v1320;
assign w4791 = w4335 & ~w4790;
assign w4792 = w1732 & ~w4788;
assign w4793 = ~w4791 & w4792;
assign w4794 = w4358 & ~w4790;
assign w4795 = pi220 & ~w1033;
assign w4796 = pi220 & w1756;
assign v1321 = ~(w2061 | w4796);
assign w4797 = v1321;
assign v1322 = ~(w1052 | w4797);
assign w4798 = v1322;
assign w4799 = w2060 & ~w4798;
assign w4800 = w2043 & ~w4799;
assign v1323 = ~(w4358 | w4795);
assign w4801 = v1323;
assign w4802 = ~w4800 & w4801;
assign v1324 = ~(w1732 | w4794);
assign w4803 = v1324;
assign w4804 = ~w4802 & w4803;
assign v1325 = ~(pi247 | w4793);
assign w4805 = v1325;
assign w4806 = ~w4804 & w4805;
assign w4807 = pi359 & ~w4787;
assign w4808 = ~w4806 & w4807;
assign w4809 = pi221 & w1756;
assign w4810 = w1991 & ~w4809;
assign w4811 = w1971 & ~w4810;
assign w4812 = w1953 & ~w4811;
assign v1326 = ~(w4420 | w4425);
assign w4813 = v1326;
assign v1327 = ~(w4460 | w4813);
assign w4814 = v1327;
assign w4815 = w4460 & w4813;
assign w4816 = w4744 & ~w4814;
assign w4817 = ~w4815 & w4816;
assign w4818 = ~pi221 & w4755;
assign w4819 = w1731 & ~w4818;
assign w4820 = ~w4812 & w4819;
assign w4821 = ~w4817 & w4820;
assign w4822 = pi221 & w1728;
assign v1328 = ~(w4821 | w4822);
assign w4823 = v1328;
assign w4824 = pi222 & w1728;
assign w4825 = ~pi351 & w4081;
assign w4826 = pi222 & w4076;
assign w4827 = w3902 & w4074;
assign v1329 = ~(w4081 | w4826);
assign w4828 = v1329;
assign w4829 = ~w4827 & w4828;
assign w4830 = w1731 & ~w4825;
assign w4831 = ~w4829 & w4830;
assign v1330 = ~(w4824 | w4831);
assign w4832 = v1330;
assign w4833 = pi223 & ~w4229;
assign w4834 = pi133 & w4232;
assign w4835 = w569 & w4200;
assign w4836 = w378 & ~w4200;
assign w4837 = w4235 & ~w4835;
assign w4838 = ~w4836 & w4837;
assign w4839 = pi135 & w4244;
assign w4840 = pi179 & w4242;
assign w4841 = pi350 & w4239;
assign v1331 = ~(w4834 | w4839);
assign w4842 = v1331;
assign v1332 = ~(w4840 | w4841);
assign w4843 = v1332;
assign w4844 = w4842 & w4843;
assign w4845 = ~w4838 & w4844;
assign v1333 = ~(pi247 | w4845);
assign w4846 = v1333;
assign v1334 = ~(w4833 | w4846);
assign w4847 = v1334;
assign w4848 = ~pi224 & w1728;
assign w4849 = ~pi350 & w4081;
assign w4850 = ~pi224 & w4076;
assign w4851 = ~w3814 & w4074;
assign v1335 = ~(w4081 | w4850);
assign w4852 = v1335;
assign w4853 = ~w4851 & w4852;
assign w4854 = w1731 & ~w4849;
assign w4855 = ~w4853 & w4854;
assign v1336 = ~(w4848 | w4855);
assign w4856 = v1336;
assign w4857 = pi225 & ~w4229;
assign w4858 = pi142 & w4232;
assign w4859 = w395 & w4200;
assign w4860 = w319 & ~w4200;
assign w4861 = w4235 & ~w4860;
assign w4862 = ~w4859 & w4861;
assign w4863 = pi130 & w4244;
assign w4864 = pi185 & w4242;
assign w4865 = pi349 & w4239;
assign v1337 = ~(w4858 | w4863);
assign w4866 = v1337;
assign v1338 = ~(w4864 | w4865);
assign w4867 = v1338;
assign w4868 = w4866 & w4867;
assign w4869 = ~w4862 & w4868;
assign v1339 = ~(pi247 | w4869);
assign w4870 = v1339;
assign v1340 = ~(w4857 | w4870);
assign w4871 = v1340;
assign w4872 = pi226 & w1728;
assign w4873 = pi226 & w4076;
assign w4874 = w3752 & w4074;
assign v1341 = ~(w4081 | w4873);
assign w4875 = v1341;
assign w4876 = ~w4874 & w4875;
assign w4877 = ~pi352 & w4081;
assign w4878 = w1731 & ~w4877;
assign w4879 = ~w4876 & w4878;
assign v1342 = ~(w4872 | w4879);
assign w4880 = v1342;
assign w4881 = pi227 & w1728;
assign w4882 = ~pi353 & w4081;
assign w4883 = pi227 & w4076;
assign w4884 = w3922 & w4074;
assign v1343 = ~(w4081 | w4883);
assign w4885 = v1343;
assign w4886 = ~w4884 & w4885;
assign w4887 = w1731 & ~w4882;
assign w4888 = ~w4886 & w4887;
assign v1344 = ~(w4881 | w4888);
assign w4889 = v1344;
assign w4890 = ~pi247 & w1033;
assign w4891 = pi228 & ~w4890;
assign w4892 = pi345 & w131;
assign w4893 = w4890 & w4892;
assign v1345 = ~(w4891 | w4893);
assign w4894 = v1345;
assign w4895 = pi359 & ~w4894;
assign w4896 = pi229 & w1728;
assign w4897 = ~pi348 & w4081;
assign w4898 = pi229 & w4076;
assign w4899 = w3994 & w4074;
assign v1346 = ~(w4081 | w4898);
assign w4900 = v1346;
assign w4901 = ~w4899 & w4900;
assign w4902 = w1731 & ~w4897;
assign w4903 = ~w4901 & w4902;
assign v1347 = ~(w4896 | w4903);
assign w4904 = v1347;
assign w4905 = ~pi230 & w38;
assign w4906 = w2734 & w4330;
assign w4907 = w1033 & w4906;
assign v1348 = ~(w4905 | w4907);
assign w4908 = v1348;
assign w4909 = pi359 & ~w4908;
assign w4910 = ~pi231 & w1728;
assign w4911 = w1033 & w1731;
assign w4912 = pi301 & ~w1249;
assign w4913 = w2 & w1213;
assign v1349 = ~(w1005 | w1197);
assign w4914 = v1349;
assign w4915 = w101 & ~w4914;
assign w4916 = w9 & w1188;
assign v1350 = ~(pi301 | w4913);
assign w4917 = v1350;
assign w4918 = ~w4916 & w4917;
assign w4919 = ~w4915 & w4918;
assign v1351 = ~(w1109 | w4912);
assign w4920 = v1351;
assign w4921 = ~w4919 & w4920;
assign w4922 = w82 & ~w996;
assign v1352 = ~(w4152 | w4922);
assign w4923 = v1352;
assign w4924 = w1109 & ~w4923;
assign w4925 = ~w88 & w4924;
assign w4926 = w82 & w617;
assign w4927 = w4157 & ~w4926;
assign w4928 = w4211 & w4927;
assign w4929 = w4159 & w4213;
assign w4930 = w4220 & w4929;
assign w4931 = w4928 & w4930;
assign w4932 = w0 & ~w4931;
assign w4933 = w82 & w103;
assign w4934 = w4146 & ~w4933;
assign w4935 = w4203 & w4934;
assign w4936 = pi301 & ~w4935;
assign v1353 = ~(w4921 | w4925);
assign w4937 = v1353;
assign w4938 = ~w4936 & w4937;
assign w4939 = ~w4932 & w4938;
assign w4940 = w4911 & ~w4939;
assign v1354 = ~(w4910 | w4940);
assign w4941 = v1354;
assign w4942 = pi232 & w1728;
assign w4943 = ~pi349 & w4081;
assign w4944 = pi232 & w4076;
assign w4945 = ~w3977 & w4074;
assign v1355 = ~(w4081 | w4944);
assign w4946 = v1355;
assign w4947 = ~w4945 & w4946;
assign w4948 = w1731 & ~w4943;
assign w4949 = ~w4947 & w4948;
assign v1356 = ~(w4942 | w4949);
assign w4950 = v1356;
assign w4951 = pi233 & w1728;
assign v1357 = ~(w98 | w1243);
assign w4952 = v1357;
assign w4953 = w2726 & ~w4952;
assign w4954 = w1038 & ~w1306;
assign w4955 = ~w1042 & w1160;
assign w4956 = w1301 & w4955;
assign w4957 = w101 & ~w4956;
assign v1358 = ~(w4954 | w4957);
assign w4958 = v1358;
assign w4959 = w0 & ~w4958;
assign v1359 = ~(w4953 | w4959);
assign w4960 = v1359;
assign w4961 = w147 & ~w4960;
assign w4962 = ~pi347 & w4961;
assign w4963 = pi233 & w4076;
assign w4964 = ~w3371 & w4074;
assign v1360 = ~(w4961 | w4963);
assign w4965 = v1360;
assign w4966 = ~w4964 & w4965;
assign w4967 = w1731 & ~w4962;
assign w4968 = ~w4966 & w4967;
assign v1361 = ~(w4951 | w4968);
assign w4969 = v1361;
assign w4970 = ~pi234 & w1728;
assign w4971 = w4226 & ~w4921;
assign w4972 = w4911 & ~w4971;
assign v1362 = ~(w4970 | w4972);
assign w4973 = v1362;
assign v1363 = ~(pi247 | w336);
assign w4974 = v1363;
assign w4975 = ~pi235 & pi247;
assign v1364 = ~(w4974 | w4975);
assign w4976 = v1364;
assign v1365 = ~(pi247 | w430);
assign w4977 = v1365;
assign w4978 = ~pi236 & pi247;
assign v1366 = ~(w4977 | w4978);
assign w4979 = v1366;
assign w4980 = pi252 & pi359;
assign w4981 = pi238 & w1728;
assign w4982 = ~pi354 & w4081;
assign w4983 = pi238 & w4076;
assign w4984 = ~w4011 & w4074;
assign v1367 = ~(w4081 | w4983);
assign w4985 = v1367;
assign w4986 = ~w4984 & w4985;
assign w4987 = w1731 & ~w4982;
assign w4988 = ~w4986 & w4987;
assign v1368 = ~(w4981 | w4988);
assign w4989 = v1368;
assign w4990 = ~pi239 & w1728;
assign w4991 = w4200 & ~w4921;
assign w4992 = w4911 & ~w4991;
assign v1369 = ~(w4990 | w4992);
assign w4993 = v1369;
assign w4994 = ~pi240 & w1728;
assign w4995 = w4170 & ~w4921;
assign w4996 = w4911 & ~w4995;
assign v1370 = ~(w4994 | w4996);
assign w4997 = v1370;
assign w4998 = pi241 & w1728;
assign w4999 = w90 & w101;
assign v1371 = ~(w1249 | w4933);
assign w5000 = v1371;
assign w5001 = ~w4999 & w5000;
assign v1372 = ~(pi303 | w4203);
assign w5002 = v1372;
assign w5003 = pi302 & w1016;
assign w5004 = pi302 & ~w612;
assign w5005 = ~w1014 & w5004;
assign w5006 = w1015 & w5005;
assign w5007 = w4952 & ~w5006;
assign w5008 = w1290 & w5007;
assign w5009 = ~w5003 & w5008;
assign w5010 = ~pi296 & w1015;
assign w5011 = w19 & w5010;
assign v1373 = ~(w1233 | w4178);
assign w5012 = v1373;
assign w5013 = w8 & ~w1233;
assign v1374 = ~(w5012 | w5013);
assign w5014 = v1374;
assign v1375 = ~(w103 | w1236);
assign w5015 = v1375;
assign w5016 = ~w5011 & w5015;
assign w5017 = ~w5014 & w5016;
assign w5018 = w5009 & w5017;
assign w5019 = pi302 & ~w5018;
assign w5020 = w5001 & ~w5002;
assign w5021 = ~w5019 & w5020;
assign w5022 = pi301 & ~w5021;
assign v1376 = ~(pi300 | w4923);
assign w5023 = v1376;
assign w5024 = ~pi302 & w4923;
assign w5025 = w1109 & ~w5023;
assign w5026 = ~w5024 & w5025;
assign w5027 = w1153 & w1288;
assign w5028 = ~w8 & w1206;
assign w5029 = ~pi303 & w1210;
assign v1377 = ~(w59 | w5029);
assign w5030 = v1377;
assign v1378 = ~(w1199 | w1204);
assign w5031 = v1378;
assign w5032 = ~w1001 & w5031;
assign w5033 = w123 & ~w1146;
assign w5034 = ~w1156 & w5033;
assign w5035 = w1117 & w1268;
assign w5036 = w4914 & w5035;
assign w5037 = w1309 & w5034;
assign w5038 = w5030 & w5032;
assign w5039 = w5037 & w5038;
assign w5040 = w1273 & w5036;
assign w5041 = w5039 & w5040;
assign w5042 = w1183 & w5041;
assign w5043 = ~w5028 & w5042;
assign w5044 = ~w6 & w1126;
assign w5045 = w1266 & ~w4187;
assign w5046 = w5044 & w5045;
assign v1379 = ~(w1118 | w4268);
assign w5047 = v1379;
assign w5048 = w1141 & w5047;
assign w5049 = ~w5027 & w5048;
assign w5050 = w5046 & w5049;
assign w5051 = w5043 & w5050;
assign w5052 = pi302 & ~w5051;
assign w5053 = pi296 & w1161;
assign v1380 = ~(w4926 | w5053);
assign w5054 = v1380;
assign w5055 = ~w5052 & w5054;
assign w5056 = w0 & ~w5055;
assign v1381 = ~(w5022 | w5026);
assign w5057 = v1381;
assign w5058 = ~w5056 & w5057;
assign w5059 = w4911 & ~w5058;
assign v1382 = ~(w4998 | w5059);
assign w5060 = v1382;
assign w5061 = pi242 & w1728;
assign w5062 = w4203 & w5001;
assign w5063 = pi301 & ~w5062;
assign w5064 = w0 & ~w4928;
assign v1383 = ~(w4925 | w5063);
assign w5065 = v1383;
assign w5066 = ~w5064 & w5065;
assign w5067 = w4911 & ~w5066;
assign v1384 = ~(w5061 | w5067);
assign w5068 = v1384;
assign w5069 = pi243 & w1728;
assign w5070 = w0 & ~w4151;
assign w5071 = w130 & w1231;
assign v1385 = ~(w5070 | w5071);
assign w5072 = v1385;
assign w5073 = ~w4924 & w5072;
assign w5074 = w4911 & ~w5073;
assign v1386 = ~(w5069 | w5074);
assign w5075 = v1386;
assign w5076 = pi244 & w1728;
assign w5077 = ~pi350 & w4961;
assign w5078 = pi244 & w4076;
assign w5079 = w3344 & w4074;
assign v1387 = ~(w4961 | w5078);
assign w5080 = v1387;
assign w5081 = ~w5079 & w5080;
assign w5082 = w1731 & ~w5077;
assign w5083 = ~w5081 & w5082;
assign v1388 = ~(w5076 | w5083);
assign w5084 = v1388;
assign v1389 = ~(pi247 | w463);
assign w5085 = v1389;
assign w5086 = ~pi245 & pi247;
assign v1390 = ~(w5085 | w5086);
assign w5087 = v1390;
assign w5088 = pi246 & w1728;
assign w5089 = ~pi353 & w4961;
assign w5090 = ~w3494 & w4074;
assign w5091 = pi246 & ~w4075;
assign w5092 = pi298 & w4075;
assign v1391 = ~(w4074 | w5091);
assign w5093 = v1391;
assign w5094 = ~w5092 & w5093;
assign v1392 = ~(w1732 | w5094);
assign w5095 = v1392;
assign w5096 = ~w5090 & w5095;
assign w5097 = pi246 & w1732;
assign v1393 = ~(w4961 | w5097);
assign w5098 = v1393;
assign w5099 = ~w5096 & w5098;
assign w5100 = w1731 & ~w5089;
assign w5101 = ~w5099 & w5100;
assign v1394 = ~(w5088 | w5101);
assign w5102 = v1394;
assign w5103 = pi359 & ~w2749;
assign v1395 = ~(pi247 | w446);
assign w5104 = v1395;
assign w5105 = pi247 & ~pi248;
assign v1396 = ~(w5104 | w5105);
assign w5106 = v1396;
assign v1397 = ~(pi247 | w479);
assign w5107 = v1397;
assign w5108 = pi247 & ~pi249;
assign v1398 = ~(w5107 | w5108);
assign w5109 = v1398;
assign v1399 = ~(pi247 | w214);
assign w5110 = v1399;
assign w5111 = pi247 & ~pi250;
assign v1400 = ~(w5110 | w5111);
assign w5112 = v1400;
assign w5113 = ~pi251 & w1728;
assign v1401 = ~(w4139 | w4921);
assign w5114 = v1401;
assign w5115 = w4911 & w5114;
assign v1402 = ~(w5113 | w5115);
assign w5116 = v1402;
assign w5117 = ~w2722 & w2730;
assign w5118 = pi359 & ~w5117;
assign w5119 = ~w1033 & w5118;
assign v1403 = ~(pi247 | w569);
assign w5120 = v1403;
assign w5121 = pi247 & ~pi253;
assign v1404 = ~(w5120 | w5121);
assign w5122 = v1404;
assign v1405 = ~(pi247 | w378);
assign w5123 = v1405;
assign w5124 = pi247 & ~pi254;
assign v1406 = ~(w5123 | w5124);
assign w5125 = v1406;
assign v1407 = ~(pi247 | w395);
assign w5126 = v1407;
assign w5127 = pi247 & ~pi255;
assign v1408 = ~(w5126 | w5127);
assign w5128 = v1408;
assign w5129 = pi256 & w1728;
assign w5130 = pi301 & w4999;
assign w5131 = pi297 & w1226;
assign w5132 = ~pi302 & w5010;
assign v1409 = ~(w5011 | w5132);
assign w5133 = v1409;
assign w5134 = ~w1231 & w5133;
assign w5135 = ~w5014 & w5134;
assign w5136 = w5008 & w5135;
assign w5137 = pi298 & ~w5136;
assign v1410 = ~(w5131 | w5137);
assign w5138 = v1410;
assign w5139 = pi301 & ~w5138;
assign w5140 = pi298 & w1109;
assign w5141 = w4923 & w5140;
assign w5142 = ~w101 & w1153;
assign w5143 = w1122 & ~w5142;
assign w5144 = w5046 & w5143;
assign w5145 = w1144 & w5144;
assign w5146 = w5043 & w5145;
assign w5147 = pi298 & ~w5146;
assign v1411 = ~(w1131 | w5147);
assign w5148 = v1411;
assign w5149 = w0 & ~w5148;
assign v1412 = ~(w5071 | w5130);
assign w5150 = v1412;
assign w5151 = ~w5141 & w5150;
assign w5152 = ~w5139 & w5151;
assign w5153 = ~w5149 & w5152;
assign w5154 = w4911 & ~w5153;
assign v1413 = ~(w5129 | w5154);
assign w5155 = v1413;
assign w5156 = pi257 & w1728;
assign w5157 = w1114 & w1129;
assign v1414 = ~(pi303 | w4202);
assign w5158 = v1414;
assign w5159 = w5012 & ~w5132;
assign w5160 = ~w5131 & w5159;
assign w5161 = w5009 & w5160;
assign v1415 = ~(w5158 | w5161);
assign w5162 = v1415;
assign v1416 = ~(w4999 | w5157);
assign w5163 = v1416;
assign w5164 = ~w5162 & w5163;
assign w5165 = pi301 & ~w5164;
assign w5166 = ~pi303 & w4923;
assign w5167 = w4344 & ~w4923;
assign w5168 = w1109 & ~w5166;
assign w5169 = ~w5167 & w5168;
assign w5170 = ~w101 & w1206;
assign v1417 = ~(w1136 | w1142);
assign w5171 = v1417;
assign w5172 = ~w1145 & w5171;
assign w5173 = ~w5170 & w5172;
assign w5174 = w5144 & w5173;
assign w5175 = w5042 & w5174;
assign w5176 = w159 & ~w5175;
assign v1418 = ~(w5165 | w5169);
assign w5177 = v1418;
assign w5178 = ~w5176 & w5177;
assign w5179 = w4911 & ~w5178;
assign v1419 = ~(w5156 | w5179);
assign w5180 = v1419;
assign v1420 = ~(pi247 | w411);
assign w5181 = v1420;
assign w5182 = pi247 & ~pi258;
assign v1421 = ~(w5181 | w5182);
assign w5183 = v1421;
assign w5184 = pi259 & w1728;
assign w5185 = ~pi352 & w4961;
assign w5186 = pi259 & w1732;
assign w5187 = ~w3524 & w4074;
assign w5188 = pi259 & ~w4075;
assign w5189 = pi302 & w4075;
assign v1422 = ~(w4074 | w5188);
assign w5190 = v1422;
assign w5191 = ~w5189 & w5190;
assign v1423 = ~(w1732 | w5191);
assign w5192 = v1423;
assign w5193 = ~w5187 & w5192;
assign v1424 = ~(w4961 | w5186);
assign w5194 = v1424;
assign w5195 = ~w5193 & w5194;
assign w5196 = w1731 & ~w5185;
assign w5197 = ~w5195 & w5196;
assign v1425 = ~(w5184 | w5197);
assign w5198 = v1425;
assign v1426 = ~(pi247 | w319);
assign w5199 = v1426;
assign w5200 = pi247 & ~pi260;
assign v1427 = ~(w5199 | w5200);
assign w5201 = v1427;
assign v1428 = ~(pi247 | w278);
assign w5202 = v1428;
assign w5203 = pi247 & ~pi261;
assign v1429 = ~(w5202 | w5203);
assign w5204 = v1429;
assign v1430 = ~(pi247 | w257);
assign w5205 = v1430;
assign w5206 = pi247 & ~pi262;
assign v1431 = ~(w5205 | w5206);
assign w5207 = v1431;
assign v1432 = ~(pi247 | w362);
assign w5208 = v1432;
assign w5209 = pi247 & ~pi263;
assign v1433 = ~(w5208 | w5209);
assign w5210 = v1433;
assign v1434 = ~(w63 | w4189);
assign w5211 = v1434;
assign w5212 = w4137 & ~w5211;
assign v1435 = ~(w52 | w60);
assign w5213 = v1435;
assign w5214 = w34 & w5213;
assign w5215 = w4927 & w5214;
assign w5216 = w0 & ~w5215;
assign w5217 = w39 & w1229;
assign w5218 = ~w53 & w5217;
assign v1436 = ~(w4202 | w5218);
assign w5219 = v1436;
assign w5220 = w24 & ~w5219;
assign w5221 = w36 & w4214;
assign w5222 = w1245 & w5221;
assign w5223 = w19 & w5222;
assign v1437 = ~(w4933 | w5223);
assign w5224 = v1437;
assign w5225 = ~w5220 & w5224;
assign w5226 = pi301 & ~w5225;
assign v1438 = ~(w5212 | w5226);
assign w5227 = v1438;
assign w5228 = ~w5216 & w5227;
assign v1439 = ~(w985 | w5228);
assign w5229 = v1439;
assign w5230 = ~pi297 & w985;
assign w5231 = pi190 & w4204;
assign w5232 = w1233 & w5231;
assign v1440 = ~(w103 | w5232);
assign w5233 = v1440;
assign w5234 = w37 & ~w5233;
assign w5235 = w16 & ~w5219;
assign w5236 = w4142 & ~w5234;
assign w5237 = ~w5235 & w5236;
assign w5238 = pi301 & ~w5237;
assign w5239 = w9 & w1212;
assign w5240 = w82 & ~w5031;
assign w5241 = w101 & w1189;
assign v1441 = ~(w5239 | w5241);
assign w5242 = v1441;
assign w5243 = ~w5240 & w5242;
assign w5244 = w101 & w1105;
assign v1442 = ~(w4153 | w5244);
assign w5245 = v1442;
assign w5246 = ~w1002 & w1136;
assign v1443 = ~(w1174 | w5246);
assign w5247 = v1443;
assign w5248 = w5245 & w5247;
assign w5249 = pi297 & ~w5248;
assign v1444 = ~(w16 | w19);
assign w5250 = v1444;
assign v1445 = ~(w5211 | w5250);
assign w5251 = v1445;
assign w5252 = w5243 & ~w5251;
assign w5253 = w4927 & w5252;
assign w5254 = ~w5249 & w5253;
assign w5255 = w0 & ~w5254;
assign v1446 = ~(w985 | w4168);
assign w5256 = v1446;
assign w5257 = ~w5238 & w5256;
assign w5258 = ~w5255 & w5257;
assign v1447 = ~(w5230 | w5258);
assign w5259 = v1447;
assign v1448 = ~(w53 | w5030);
assign w5260 = v1448;
assign v1449 = ~(w52 | w5260);
assign w5261 = v1449;
assign w5262 = pi291 & ~w5247;
assign v1450 = ~(w157 | w5221);
assign w5263 = v1450;
assign v1451 = ~(w5211 | w5263);
assign w5264 = v1451;
assign v1452 = ~(w4219 | w5264);
assign w5265 = v1452;
assign w5266 = w34 & w5265;
assign w5267 = w5243 & w5245;
assign w5268 = w5266 & w5267;
assign w5269 = w5261 & w5268;
assign w5270 = ~w5262 & w5269;
assign w5271 = w0 & ~w5270;
assign w5272 = w157 & ~w5219;
assign w5273 = w4142 & ~w5222;
assign w5274 = ~w5272 & w5273;
assign w5275 = pi301 & ~w5274;
assign w5276 = w103 & w2726;
assign v1453 = ~(w985 | w4210);
assign w5277 = v1453;
assign w5278 = ~w5276 & w5277;
assign w5279 = ~w5275 & w5278;
assign w5280 = ~w5271 & w5279;
assign w5281 = w5229 & w5280;
assign w5282 = w5259 & w5281;
assign w5283 = pi132 & w5282;
assign w5284 = w5229 & w5258;
assign w5285 = ~w5280 & w5284;
assign w5286 = pi220 & w5285;
assign w5287 = w5280 & w5284;
assign w5288 = pi174 & w5287;
assign w5289 = ~pi291 & w985;
assign v1454 = ~(w5280 | w5289);
assign w5290 = v1454;
assign w5291 = w5259 & w5290;
assign w5292 = ~w5229 & w5291;
assign w5293 = pi354 & w5292;
assign v1455 = ~(pi296 | w1326);
assign w5294 = v1455;
assign w5295 = pi303 & w82;
assign w5296 = w1245 & w5295;
assign w5297 = w4174 & w4202;
assign w5298 = ~w4174 & w5218;
assign w5299 = w4912 & ~w5298;
assign w5300 = ~w5296 & w5299;
assign w5301 = ~w5297 & w5300;
assign w5302 = w4174 & ~w5211;
assign w5303 = w101 & ~w1169;
assign w5304 = pi296 & ~w5247;
assign w5305 = pi190 & ~w5261;
assign w5306 = w0 & ~w5303;
assign w5307 = ~w33 & w5306;
assign w5308 = ~w5302 & w5307;
assign w5309 = w5243 & w5308;
assign w5310 = ~w5305 & w5309;
assign w5311 = ~w5304 & w5310;
assign v1456 = ~(w5301 | w5311);
assign w5312 = v1456;
assign v1457 = ~(w985 | w5312);
assign w5313 = v1457;
assign v1458 = ~(w5294 | w5313);
assign w5314 = v1458;
assign v1459 = ~(w5229 | w5291);
assign w5315 = v1459;
assign w5316 = ~w2627 & w5315;
assign v1460 = ~(w5282 | w5314);
assign w5317 = v1460;
assign w5318 = ~w5286 & w5317;
assign w5319 = ~w5288 & w5318;
assign v1461 = ~(w5293 | w5316);
assign w5320 = v1461;
assign w5321 = w5319 & w5320;
assign w5322 = ~w3657 & w5315;
assign w5323 = pi187 & w5287;
assign w5324 = pi212 & w5285;
assign w5325 = pi126 & w5292;
assign w5326 = w5314 & ~w5323;
assign w5327 = ~w5324 & w5326;
assign v1462 = ~(w5322 | w5325);
assign w5328 = v1462;
assign w5329 = w5327 & w5328;
assign v1463 = ~(w5321 | w5329);
assign w5330 = v1463;
assign v1464 = ~(w5283 | w5330);
assign w5331 = v1464;
assign v1465 = ~(pi247 | w5331);
assign w5332 = v1465;
assign w5333 = pi247 & pi264;
assign v1466 = ~(w5332 | w5333);
assign w5334 = v1466;
assign w5335 = pi265 & w1728;
assign w5336 = ~pi348 & w4961;
assign w5337 = pi265 & w1732;
assign w5338 = w3711 & w4074;
assign w5339 = pi265 & ~w4075;
assign w5340 = pi303 & w4075;
assign v1467 = ~(w4074 | w5339);
assign w5341 = v1467;
assign w5342 = ~w5340 & w5341;
assign v1468 = ~(w1732 | w5342);
assign w5343 = v1468;
assign w5344 = ~w5338 & w5343;
assign v1469 = ~(w4961 | w5337);
assign w5345 = v1469;
assign w5346 = ~w5344 & w5345;
assign w5347 = w1731 & ~w5336;
assign w5348 = ~w5346 & w5347;
assign v1470 = ~(w5335 | w5348);
assign w5349 = v1470;
assign v1471 = ~(pi247 | w237);
assign w5350 = v1471;
assign w5351 = pi247 & ~pi266;
assign v1472 = ~(w5350 | w5351);
assign w5352 = v1472;
assign v1473 = ~(pi247 | w298);
assign w5353 = v1473;
assign w5354 = pi247 & ~pi267;
assign v1474 = ~(w5353 | w5354);
assign w5355 = v1474;
assign w5356 = pi268 & w1728;
assign w5357 = ~pi351 & w4961;
assign w5358 = pi268 & w4076;
assign w5359 = w3691 & w4074;
assign v1475 = ~(w4961 | w5358);
assign w5360 = v1475;
assign w5361 = ~w5359 & w5360;
assign w5362 = w1731 & ~w5357;
assign w5363 = ~w5361 & w5362;
assign v1476 = ~(w5356 | w5363);
assign w5364 = v1476;
assign w5365 = pi247 & ~pi269;
assign w5366 = w5292 & ~w5314;
assign w5367 = pi347 & w5366;
assign w5368 = w5287 & ~w5314;
assign w5369 = pi137 & w5368;
assign w5370 = w5285 & ~w5314;
assign w5371 = pi211 & w5370;
assign w5372 = w5285 & w5314;
assign w5373 = pi219 & w5372;
assign w5374 = w5287 & w5314;
assign w5375 = pi117 & w5374;
assign w5376 = w5282 & w5314;
assign w5377 = pi131 & w5376;
assign w5378 = w5292 & w5314;
assign w5379 = pi140 & w5378;
assign w5380 = w1549 & ~w5314;
assign w5381 = w2554 & w5314;
assign v1477 = ~(w5380 | w5381);
assign w5382 = v1477;
assign w5383 = w5315 & w5382;
assign v1478 = ~(pi247 | w5369);
assign w5384 = v1478;
assign v1479 = ~(w5371 | w5373);
assign w5385 = v1479;
assign v1480 = ~(w5375 | w5377);
assign w5386 = v1480;
assign w5387 = ~w5383 & w5386;
assign w5388 = w5384 & w5385;
assign v1481 = ~(w5367 | w5379);
assign w5389 = v1481;
assign w5390 = w5388 & w5389;
assign w5391 = w5387 & w5390;
assign v1482 = ~(w5365 | w5391);
assign w5392 = v1482;
assign w5393 = pi247 & ~pi270;
assign w5394 = pi143 & w5378;
assign w5395 = pi209 & w5370;
assign w5396 = pi146 & w5368;
assign w5397 = pi177 & w5374;
assign w5398 = pi204 & w5372;
assign w5399 = pi184 & w5376;
assign w5400 = pi352 & w5366;
assign w5401 = w1637 & ~w5314;
assign w5402 = w2768 & w5314;
assign v1483 = ~(w5401 | w5402);
assign w5403 = v1483;
assign w5404 = w5315 & w5403;
assign v1484 = ~(pi247 | w5395);
assign w5405 = v1484;
assign v1485 = ~(w5396 | w5397);
assign w5406 = v1485;
assign v1486 = ~(w5398 | w5399);
assign w5407 = v1486;
assign w5408 = ~w5404 & w5407;
assign w5409 = w5405 & w5406;
assign v1487 = ~(w5394 | w5400);
assign w5410 = v1487;
assign w5411 = w5409 & w5410;
assign w5412 = w5408 & w5411;
assign v1488 = ~(w5393 | w5412);
assign w5413 = v1488;
assign w5414 = pi247 & ~pi271;
assign w5415 = pi349 & w5366;
assign w5416 = pi130 & w5368;
assign w5417 = pi199 & w5372;
assign w5418 = pi206 & w5370;
assign w5419 = pi185 & w5374;
assign w5420 = pi129 & w5376;
assign w5421 = pi142 & w5378;
assign w5422 = w2509 & ~w5314;
assign w5423 = w3181 & w5314;
assign v1489 = ~(w5422 | w5423);
assign w5424 = v1489;
assign w5425 = w5315 & w5424;
assign v1490 = ~(pi247 | w5416);
assign w5426 = v1490;
assign v1491 = ~(w5417 | w5418);
assign w5427 = v1491;
assign v1492 = ~(w5419 | w5420);
assign w5428 = v1492;
assign w5429 = ~w5425 & w5428;
assign w5430 = w5426 & w5427;
assign v1493 = ~(w5415 | w5421);
assign w5431 = v1493;
assign w5432 = w5430 & w5431;
assign w5433 = w5429 & w5432;
assign v1494 = ~(w5414 | w5433);
assign w5434 = v1494;
assign w5435 = pi247 & ~pi272;
assign w5436 = pi348 & w5366;
assign w5437 = pi173 & w5368;
assign w5438 = pi186 & w5374;
assign w5439 = pi208 & w5370;
assign w5440 = pi203 & w5372;
assign w5441 = ~pi180 & w5376;
assign w5442 = pi138 & w5378;
assign w5443 = w2446 & ~w5314;
assign w5444 = w3114 & w5314;
assign v1495 = ~(w5443 | w5444);
assign w5445 = v1495;
assign w5446 = w5315 & w5445;
assign v1496 = ~(pi247 | w5437);
assign w5447 = v1496;
assign v1497 = ~(w5438 | w5439);
assign w5448 = v1497;
assign v1498 = ~(w5440 | w5441);
assign w5449 = v1498;
assign w5450 = ~w5446 & w5449;
assign w5451 = w5447 & w5448;
assign v1499 = ~(w5436 | w5442);
assign w5452 = v1499;
assign w5453 = w5451 & w5452;
assign w5454 = w5450 & w5453;
assign v1500 = ~(w5435 | w5454);
assign w5455 = v1500;
assign w5456 = pi247 & ~pi273;
assign w5457 = pi353 & w5366;
assign w5458 = pi210 & w5370;
assign w5459 = pi144 & w5368;
assign w5460 = pi183 & w5374;
assign w5461 = pi205 & w5372;
assign w5462 = ~pi181 & w5376;
assign w5463 = pi139 & w5378;
assign w5464 = w2388 & ~w5314;
assign w5465 = w2792 & w5314;
assign v1501 = ~(w5464 | w5465);
assign w5466 = v1501;
assign w5467 = w5315 & w5466;
assign v1502 = ~(pi247 | w5458);
assign w5468 = v1502;
assign v1503 = ~(w5459 | w5460);
assign w5469 = v1503;
assign v1504 = ~(w5461 | w5462);
assign w5470 = v1504;
assign w5471 = ~w5467 & w5470;
assign w5472 = w5468 & w5469;
assign v1505 = ~(w5457 | w5463);
assign w5473 = v1505;
assign w5474 = w5472 & w5473;
assign w5475 = w5471 & w5474;
assign v1506 = ~(w5456 | w5475);
assign w5476 = v1506;
assign w5477 = pi247 & ~pi274;
assign w5478 = pi141 & w5378;
assign w5479 = pi172 & w5368;
assign w5480 = pi221 & w5372;
assign w5481 = pi207 & w5370;
assign w5482 = pi182 & w5374;
assign w5483 = pi102 & w5376;
assign w5484 = pi351 & w5366;
assign w5485 = w1679 & ~w5314;
assign w5486 = w3548 & w5314;
assign v1507 = ~(w5485 | w5486);
assign w5487 = v1507;
assign w5488 = w5315 & w5487;
assign v1508 = ~(pi247 | w5479);
assign w5489 = v1508;
assign v1509 = ~(w5480 | w5481);
assign w5490 = v1509;
assign v1510 = ~(w5482 | w5483);
assign w5491 = v1510;
assign w5492 = ~w5488 & w5491;
assign w5493 = w5489 & w5490;
assign v1511 = ~(w5478 | w5484);
assign w5494 = v1511;
assign w5495 = w5493 & w5494;
assign w5496 = w5492 & w5495;
assign v1512 = ~(w5477 | w5496);
assign w5497 = v1512;
assign w5498 = pi247 & ~pi275;
assign w5499 = pi350 & w5366;
assign w5500 = pi135 & w5368;
assign w5501 = pi218 & w5372;
assign w5502 = pi179 & w5374;
assign w5503 = pi200 & w5370;
assign w5504 = pi178 & w5376;
assign w5505 = pi133 & w5378;
assign w5506 = w2352 & ~w5314;
assign w5507 = w2673 & w5314;
assign v1513 = ~(w5506 | w5507);
assign w5508 = v1513;
assign w5509 = w5315 & w5508;
assign v1514 = ~(pi247 | w5500);
assign w5510 = v1514;
assign v1515 = ~(w5501 | w5502);
assign w5511 = v1515;
assign v1516 = ~(w5503 | w5504);
assign w5512 = v1516;
assign w5513 = ~w5509 & w5512;
assign w5514 = w5510 & w5511;
assign v1517 = ~(w5499 | w5505);
assign w5515 = v1517;
assign w5516 = w5514 & w5515;
assign w5517 = w5513 & w5516;
assign v1518 = ~(w5498 | w5517);
assign w5518 = v1518;
assign w5519 = pi276 & w1728;
assign w5520 = ~pi349 & w4961;
assign w5521 = pi276 & w4076;
assign w5522 = ~w3238 & w4074;
assign v1519 = ~(w4961 | w5521);
assign w5523 = v1519;
assign w5524 = ~w5522 & w5523;
assign w5525 = w1731 & ~w5520;
assign w5526 = ~w5524 & w5525;
assign v1520 = ~(w5519 | w5526);
assign w5527 = v1520;
assign w5528 = pi247 & ~pi277;
assign v1521 = ~(w1052 | w3084);
assign w5529 = v1521;
assign w5530 = ~w986 & w5529;
assign w5531 = ~pi247 & w5530;
assign w5532 = w1328 & w5531;
assign v1522 = ~(w5528 | w5532);
assign w5533 = v1522;
assign w5534 = pi278 & w1728;
assign w5535 = ~pi294 & w1731;
assign w5536 = w130 & w5535;
assign w5537 = ~w5178 & w5536;
assign w5538 = w5153 & w5537;
assign v1523 = ~(w5534 | w5538);
assign w5539 = v1523;
assign v1524 = ~(w1501 | w2732);
assign w5540 = v1524;
assign v1525 = ~(pi195 | w5540);
assign w5541 = v1525;
assign w5542 = w82 & ~w5541;
assign w5543 = ~w5540 & w5542;
assign w5544 = w2730 & ~w5543;
assign w5545 = w996 & w1109;
assign w5546 = w92 & w5545;
assign w5547 = w2 & w1212;
assign v1526 = ~(pi190 | w5032);
assign w5548 = v1526;
assign v1527 = ~(w1105 | w1189);
assign w5549 = v1527;
assign w5550 = ~w1153 & w5549;
assign w5551 = pi190 & ~w5550;
assign w5552 = w51 & ~w62;
assign w5553 = ~w5548 & w5552;
assign w5554 = ~w5551 & w5553;
assign w5555 = w8 & ~w5554;
assign w5556 = ~w6 & w5030;
assign w5557 = w70 & ~w5556;
assign v1528 = ~(w113 | w5547);
assign w5558 = v1528;
assign w5559 = ~w5557 & w5558;
assign w5560 = ~w5555 & w5559;
assign w5561 = w0 & ~w5560;
assign w5562 = w39 & w4130;
assign v1529 = ~(w93 | w5562);
assign w5563 = v1529;
assign w5564 = pi301 & ~w5563;
assign w5565 = w1245 & w2726;
assign v1530 = ~(w3199 | w5546);
assign w5566 = v1530;
assign w5567 = ~w5565 & w5566;
assign w5568 = ~w5564 & w5567;
assign w5569 = ~w5561 & w5568;
assign v1531 = ~(pi189 | w1185);
assign w5570 = v1531;
assign w5571 = w85 & ~w5570;
assign w5572 = ~w53 & w5571;
assign w5573 = w57 & w101;
assign w5574 = w1230 & w5573;
assign v1532 = ~(w5572 | w5574);
assign w5575 = v1532;
assign w5576 = ~w4202 & w5575;
assign w5577 = pi301 & ~w5576;
assign w5578 = w1081 & w1206;
assign v1533 = ~(w5540 | w5578);
assign w5579 = v1533;
assign w5580 = ~w4270 & w5579;
assign w5581 = ~w4341 & w5580;
assign w5582 = ~w5577 & w5581;
assign w5583 = w5569 & w5582;
assign v1534 = ~(w82 | w5583);
assign w5584 = v1534;
assign w5585 = pi359 & ~w5584;
assign w5586 = pi359 & w1509;
assign w5587 = ~w5569 & w5586;
assign v1535 = ~(w5585 | w5587);
assign w5588 = v1535;
assign v1536 = ~(w5544 | w5588);
assign w5589 = v1536;
assign w5590 = w1284 & w5290;
assign w5591 = ~w5259 & w5590;
assign w5592 = pi304 & ~w5591;
assign w5593 = pi314 & w5591;
assign v1537 = ~(w5592 | w5593);
assign w5594 = v1537;
assign v1538 = ~(pi247 | w5594);
assign w5595 = v1538;
assign w5596 = pi247 & pi280;
assign v1539 = ~(w5595 | w5596);
assign w5597 = v1539;
assign w5598 = ~w147 & w5542;
assign w5599 = w2730 & ~w5598;
assign w5600 = ~w5588 & w5599;
assign w5601 = pi282 & w1728;
assign w5602 = w3726 & ~w4960;
assign w5603 = w3728 & w4074;
assign w5604 = pi282 & w4076;
assign v1540 = ~(w5603 | w5604);
assign w5605 = v1540;
assign w5606 = ~w4961 & w5605;
assign w5607 = w1731 & ~w5602;
assign w5608 = ~w5606 & w5607;
assign v1541 = ~(w5601 | w5608);
assign w5609 = v1541;
assign w5610 = pi247 & ~pi283;
assign v1542 = ~(pi247 | w5259);
assign w5611 = v1542;
assign w5612 = ~w5590 & w5611;
assign v1543 = ~(w5610 | w5612);
assign w5613 = v1543;
assign v1544 = ~(pi247 | w5290);
assign w5614 = v1544;
assign w5615 = pi247 & ~pi284;
assign v1545 = ~(w5614 | w5615);
assign w5616 = v1545;
assign w5617 = w1260 & w5529;
assign v1546 = ~(w153 | w5529);
assign w5618 = v1546;
assign v1547 = ~(pi247 | w986);
assign w5619 = v1547;
assign w5620 = ~w5618 & w5619;
assign w5621 = ~w5617 & w5620;
assign w5622 = pi247 & ~pi285;
assign v1548 = ~(w5621 | w5622);
assign w5623 = v1548;
assign w5624 = pi247 & ~pi286;
assign w5625 = pi140 & w2897;
assign w5626 = pi303 & w2895;
assign w5627 = w5625 & w5626;
assign w5628 = w2896 & w5626;
assign w5629 = pi295 & w2038;
assign w5630 = pi289 & w5629;
assign w5631 = pi288 & w5630;
assign w5632 = pi290 & w5631;
assign w5633 = pi287 & w5632;
assign v1549 = ~(pi286 | w5633);
assign w5634 = v1549;
assign w5635 = pi286 & w5633;
assign v1550 = ~(w5628 | w5634);
assign w5636 = v1550;
assign w5637 = ~w5635 & w5636;
assign v1551 = ~(pi247 | w5627);
assign w5638 = v1551;
assign w5639 = ~w5637 & w5638;
assign w5640 = pi359 & ~w5624;
assign w5641 = ~w5639 & w5640;
assign w5642 = pi247 & ~pi287;
assign w5643 = pi139 & w2897;
assign w5644 = w5626 & w5643;
assign v1552 = ~(pi287 | w5632);
assign w5645 = v1552;
assign v1553 = ~(w5628 | w5633);
assign w5646 = v1553;
assign w5647 = ~w5645 & w5646;
assign v1554 = ~(pi247 | w5644);
assign w5648 = v1554;
assign w5649 = ~w5647 & w5648;
assign w5650 = pi359 & ~w5642;
assign w5651 = ~w5649 & w5650;
assign w5652 = pi247 & ~pi288;
assign w5653 = pi138 & w2897;
assign w5654 = w5626 & w5653;
assign v1555 = ~(pi288 | w5630);
assign w5655 = v1555;
assign v1556 = ~(w5628 | w5631);
assign w5656 = v1556;
assign w5657 = ~w5655 & w5656;
assign v1557 = ~(pi247 | w5654);
assign w5658 = v1557;
assign w5659 = ~w5657 & w5658;
assign w5660 = pi359 & ~w5652;
assign w5661 = ~w5659 & w5660;
assign w5662 = pi247 & ~pi289;
assign w5663 = pi141 & w2897;
assign w5664 = w5626 & w5663;
assign v1558 = ~(pi289 | w5629);
assign w5665 = v1558;
assign v1559 = ~(w5628 | w5630);
assign w5666 = v1559;
assign w5667 = ~w5665 & w5666;
assign v1560 = ~(pi247 | w5664);
assign w5668 = v1560;
assign w5669 = ~w5667 & w5668;
assign w5670 = pi359 & ~w5662;
assign w5671 = ~w5669 & w5670;
assign w5672 = pi247 & ~pi290;
assign w5673 = pi143 & w2897;
assign w5674 = w5626 & w5673;
assign v1561 = ~(pi290 | w5631);
assign w5675 = v1561;
assign v1562 = ~(w5628 | w5632);
assign w5676 = v1562;
assign w5677 = ~w5675 & w5676;
assign v1563 = ~(pi247 | w5674);
assign w5678 = v1563;
assign w5679 = ~w5677 & w5678;
assign w5680 = pi359 & ~w5672;
assign w5681 = ~w5679 & w5680;
assign w5682 = pi247 & ~pi291;
assign w5683 = pi367 & w982;
assign w5684 = ~pi196 & pi230;
assign w5685 = ~w1079 & w5684;
assign w5686 = w5683 & w5685;
assign w5687 = pi195 & ~pi331;
assign w5688 = pi333 & w5687;
assign w5689 = w982 & w5688;
assign v1564 = ~(pi247 | w5689);
assign w5690 = v1564;
assign w5691 = ~w5686 & w5690;
assign v1565 = ~(w4487 | w5691);
assign w5692 = v1565;
assign w5693 = w1109 & w1258;
assign w5694 = w982 & w5693;
assign v1566 = ~(pi291 | w5694);
assign w5695 = v1566;
assign w5696 = ~pi367 & w5694;
assign v1567 = ~(w983 | w5695);
assign w5697 = v1567;
assign w5698 = ~w5696 & w5697;
assign v1568 = ~(w5692 | w5698);
assign w5699 = v1568;
assign w5700 = pi359 & ~w5682;
assign w5701 = ~w5699 & w5700;
assign w5702 = pi247 & ~pi292;
assign w5703 = pi126 & w2897;
assign w5704 = w5626 & w5703;
assign v1569 = ~(pi292 | w983);
assign w5705 = v1569;
assign v1570 = ~(w2038 | w5705);
assign w5706 = v1570;
assign w5707 = ~w5628 & w5706;
assign v1571 = ~(pi247 | w5704);
assign w5708 = v1571;
assign w5709 = ~w5707 & w5708;
assign w5710 = pi359 & ~w5702;
assign w5711 = ~w5709 & w5710;
assign w5712 = ~w5542 & w5585;
assign w5713 = ~pi247 & w4089;
assign v1572 = ~(pi294 | w5713);
assign w5714 = v1572;
assign w5715 = ~pi247 & w983;
assign w5716 = ~w4089 & w5715;
assign v1573 = ~(pi294 | w983);
assign w5717 = v1573;
assign v1574 = ~(w5716 | w5717);
assign w5718 = v1574;
assign v1575 = ~(w986 | w5718);
assign w5719 = v1575;
assign w5720 = pi359 & ~w5714;
assign w5721 = ~w5719 & w5720;
assign w5722 = pi247 & ~pi295;
assign w5723 = pi142 & w2897;
assign w5724 = w5626 & w5723;
assign v1576 = ~(pi295 | w2038);
assign w5725 = v1576;
assign v1577 = ~(w5628 | w5629);
assign w5726 = v1577;
assign v1578 = ~(pi247 | w5726);
assign w5727 = v1578;
assign v1579 = ~(w5725 | w5727);
assign w5728 = v1579;
assign v1580 = ~(w5724 | w5728);
assign w5729 = v1580;
assign w5730 = pi359 & ~w5722;
assign w5731 = ~w5729 & w5730;
assign w5732 = pi247 & ~pi296;
assign w5733 = pi365 & w982;
assign w5734 = w5685 & w5733;
assign w5735 = w5690 & ~w5734;
assign v1581 = ~(w4487 | w5735);
assign w5736 = v1581;
assign v1582 = ~(pi296 | w5694);
assign w5737 = v1582;
assign w5738 = ~pi365 & w5694;
assign v1583 = ~(w983 | w5737);
assign w5739 = v1583;
assign w5740 = ~w5738 & w5739;
assign v1584 = ~(w5736 | w5740);
assign w5741 = v1584;
assign w5742 = pi359 & ~w5732;
assign w5743 = ~w5741 & w5742;
assign w5744 = pi247 & ~pi297;
assign w5745 = pi366 & w982;
assign w5746 = w5685 & w5745;
assign w5747 = w5690 & ~w5746;
assign v1585 = ~(w4487 | w5747);
assign w5748 = v1585;
assign v1586 = ~(pi297 | w5694);
assign w5749 = v1586;
assign w5750 = ~pi366 & w5694;
assign v1587 = ~(w983 | w5749);
assign w5751 = v1587;
assign w5752 = ~w5750 & w5751;
assign v1588 = ~(w5748 | w5752);
assign w5753 = v1588;
assign w5754 = pi359 & ~w5744;
assign w5755 = ~w5753 & w5754;
assign w5756 = pi247 & ~pi298;
assign w5757 = pi370 & w982;
assign w5758 = w5685 & w5757;
assign w5759 = w5690 & ~w5758;
assign v1589 = ~(w4487 | w5759);
assign w5760 = v1589;
assign v1590 = ~(pi298 | w5694);
assign w5761 = v1590;
assign w5762 = ~pi370 & w5694;
assign v1591 = ~(w983 | w5761);
assign w5763 = v1591;
assign w5764 = ~w5762 & w5763;
assign v1592 = ~(w5760 | w5764);
assign w5765 = v1592;
assign w5766 = pi359 & ~w5756;
assign w5767 = ~w5765 & w5766;
assign w5768 = pi247 & ~pi299;
assign w5769 = pi371 & w982;
assign w5770 = w5685 & w5769;
assign w5771 = w5690 & ~w5770;
assign v1593 = ~(w4487 | w5771);
assign w5772 = v1593;
assign v1594 = ~(pi299 | w5694);
assign w5773 = v1594;
assign w5774 = ~pi371 & w5694;
assign v1595 = ~(w983 | w5773);
assign w5775 = v1595;
assign w5776 = ~w5774 & w5775;
assign v1596 = ~(w5772 | w5776);
assign w5777 = v1596;
assign w5778 = pi359 & ~w5768;
assign w5779 = ~w5777 & w5778;
assign w5780 = pi247 & ~pi300;
assign w5781 = pi372 & w982;
assign w5782 = w5685 & w5781;
assign w5783 = w5690 & ~w5782;
assign v1597 = ~(w4487 | w5783);
assign w5784 = v1597;
assign v1598 = ~(pi300 | w5694);
assign w5785 = v1598;
assign w5786 = ~pi372 & w5694;
assign v1599 = ~(w983 | w5785);
assign w5787 = v1599;
assign w5788 = ~w5786 & w5787;
assign v1600 = ~(w5784 | w5788);
assign w5789 = v1600;
assign w5790 = pi359 & ~w5780;
assign w5791 = ~w5789 & w5790;
assign w5792 = pi302 & w4090;
assign w5793 = w5716 & ~w5792;
assign w5794 = w4091 & w5793;
assign w5795 = pi301 & ~w5715;
assign v1601 = ~(w5794 | w5795);
assign w5796 = v1601;
assign w5797 = pi359 & ~w5796;
assign w5798 = pi247 & ~pi302;
assign w5799 = pi369 & w982;
assign w5800 = w5685 & w5799;
assign w5801 = w5690 & ~w5800;
assign v1602 = ~(w4487 | w5801);
assign w5802 = v1602;
assign v1603 = ~(pi302 | w5694);
assign w5803 = v1603;
assign w5804 = ~pi369 & w5694;
assign v1604 = ~(w983 | w5803);
assign w5805 = v1604;
assign w5806 = ~w5804 & w5805;
assign v1605 = ~(w5802 | w5806);
assign w5807 = v1605;
assign w5808 = pi359 & ~w5798;
assign w5809 = ~w5807 & w5808;
assign w5810 = pi247 & ~pi303;
assign w5811 = pi368 & w982;
assign w5812 = w5685 & w5811;
assign w5813 = w5690 & ~w5812;
assign v1606 = ~(w4487 | w5813);
assign w5814 = v1606;
assign v1607 = ~(pi303 | w5694);
assign w5815 = v1607;
assign w5816 = ~pi368 & w5694;
assign v1608 = ~(w983 | w5815);
assign w5817 = v1608;
assign w5818 = ~w5816 & w5817;
assign v1609 = ~(w5814 | w5818);
assign w5819 = v1609;
assign w5820 = pi359 & ~w5810;
assign w5821 = ~w5819 & w5820;
assign w5822 = w16 & w47;
assign w5823 = w1051 & w5822;
assign w5824 = w4487 & w5823;
assign v1610 = ~(pi304 | w5824);
assign w5825 = v1610;
assign w5826 = pi304 & w5824;
assign w5827 = pi359 & ~w5825;
assign w5828 = ~w5826 & w5827;
assign w5829 = ~pi247 & w986;
assign v1611 = ~(pi305 | w5829);
assign w5830 = v1611;
assign w5831 = pi359 & ~w5830;
assign w5832 = ~w5793 & w5831;
assign w5833 = pi247 & ~pi307;
assign w5834 = w1109 & ~w5010;
assign w5835 = ~w11 & w1155;
assign w5836 = w4344 & ~w5835;
assign w5837 = pi132 & ~w5836;
assign w5838 = ~pi132 & w5836;
assign w5839 = w1134 & ~w5837;
assign w5840 = ~w5838 & w5839;
assign w5841 = ~pi296 & w108;
assign w5842 = w5836 & w5841;
assign w5843 = pi131 & ~w5842;
assign w5844 = ~pi131 & w5842;
assign w5845 = w1176 & ~w5843;
assign w5846 = ~w5844 & w5845;
assign v1612 = ~(w5840 | w5846);
assign w5847 = v1612;
assign w5848 = w101 & ~w5847;
assign w5849 = pi296 & ~w1000;
assign v1613 = ~(pi297 | w999);
assign w5850 = v1613;
assign v1614 = ~(w5849 | w5850);
assign w5851 = v1614;
assign v1615 = ~(w1134 | w1176);
assign w5852 = v1615;
assign v1616 = ~(pi291 | w614);
assign w5853 = v1616;
assign w5854 = ~w999 & w5853;
assign w5855 = ~pi302 & w83;
assign v1617 = ~(w1104 | w5855);
assign w5856 = v1617;
assign w5857 = ~w1139 & w5852;
assign w5858 = ~w5854 & w5857;
assign w5859 = w5856 & w5858;
assign w5860 = ~w5842 & w5851;
assign w5861 = w5859 & w5860;
assign w5862 = w0 & ~w5861;
assign w5863 = ~w5848 & w5862;
assign w5864 = pi301 & ~w85;
assign w5865 = ~w1233 & w5864;
assign w5866 = ~w1231 & w5865;
assign v1618 = ~(pi247 | w5834);
assign w5867 = v1618;
assign w5868 = ~w5866 & w5867;
assign w5869 = ~w5863 & w5868;
assign w5870 = pi359 & ~w5833;
assign w5871 = ~w5869 & w5870;
assign w5872 = pi308 & w1728;
assign w5873 = w9 & w32;
assign w5874 = w6 & ~w5873;
assign w5875 = ~w1037 & w5842;
assign w5876 = w5 & w749;
assign v1619 = ~(w69 | w1209);
assign w5877 = v1619;
assign w5878 = ~w5876 & w5877;
assign w5879 = ~w5842 & w5878;
assign w5880 = ~w121 & w5852;
assign w5881 = ~w5875 & w5880;
assign w5882 = ~w5879 & w5881;
assign v1620 = ~(w5874 | w5882);
assign w5883 = v1620;
assign w5884 = w0 & ~w5883;
assign v1621 = ~(w85 | w1230);
assign w5885 = v1621;
assign w5886 = ~w1243 & w5885;
assign w5887 = pi301 & ~w5886;
assign v1622 = ~(w5884 | w5887);
assign w5888 = v1622;
assign w5889 = w1731 & ~w5888;
assign v1623 = ~(w5872 | w5889);
assign w5890 = v1623;
assign v1624 = ~(pi247 | w4226);
assign w5891 = v1624;
assign w5892 = pi247 & pi309;
assign v1625 = ~(w5891 | w5892);
assign w5893 = v1625;
assign w5894 = pi247 & ~pi310;
assign w5895 = ~w98 & w5012;
assign w5896 = pi301 & ~w5895;
assign w5897 = w10 & w32;
assign w5898 = w122 & ~w1299;
assign v1626 = ~(w615 | w4088);
assign w5899 = v1626;
assign w5900 = w108 & ~w5899;
assign v1627 = ~(pi303 | w4143);
assign w5901 = v1627;
assign v1628 = ~(w48 | w5901);
assign w5902 = v1628;
assign w5903 = w47 & ~w5902;
assign w5904 = ~w1132 & w5849;
assign w5905 = pi297 & ~w83;
assign w5906 = ~w999 & w5905;
assign w5907 = ~w5854 & w5906;
assign w5908 = ~pi291 & w1000;
assign v1629 = ~(pi296 | w47);
assign w5909 = v1629;
assign w5910 = ~w1139 & w5909;
assign w5911 = ~w5907 & w5910;
assign w5912 = ~w5908 & w5911;
assign v1630 = ~(w5904 | w5912);
assign w5913 = v1630;
assign w5914 = pi297 & ~w5822;
assign v1631 = ~(w5850 | w5914);
assign w5915 = v1631;
assign v1632 = ~(w5900 | w5903);
assign w5916 = v1632;
assign w5917 = ~w5915 & w5916;
assign w5918 = ~w5913 & w5917;
assign v1633 = ~(w5842 | w5918);
assign w5919 = v1633;
assign w5920 = pi196 & w5842;
assign v1634 = ~(w1134 | w5920);
assign w5921 = v1634;
assign w5922 = ~w5919 & w5921;
assign v1635 = ~(w121 | w5922);
assign w5923 = v1635;
assign v1636 = ~(w1176 | w5897);
assign w5924 = v1636;
assign w5925 = ~w5898 & w5924;
assign w5926 = ~w5923 & w5925;
assign w5927 = w0 & ~w5926;
assign v1637 = ~(pi247 | w5545);
assign w5928 = v1637;
assign w5929 = ~w5896 & w5928;
assign w5930 = ~w5927 & w5929;
assign w5931 = pi359 & ~w5894;
assign w5932 = ~w5930 & w5931;
assign w5933 = w1284 & ~w4226;
assign w5934 = w4170 & w5933;
assign w5935 = pi304 & ~w5934;
assign w5936 = pi314 & w5934;
assign v1638 = ~(w5935 | w5936);
assign w5937 = v1638;
assign v1639 = ~(pi247 | w5937);
assign w5938 = v1639;
assign w5939 = pi247 & pi311;
assign v1640 = ~(w5938 | w5939);
assign w5940 = v1640;
assign w5941 = pi247 & ~pi312;
assign w5942 = ~pi247 & w4170;
assign w5943 = ~w5933 & w5942;
assign v1641 = ~(w5941 | w5943);
assign w5944 = v1641;
assign w5945 = pi313 & ~w5716;
assign w5946 = w4091 & w5715;
assign w5947 = w16 & w5946;
assign v1642 = ~(w5945 | w5947);
assign w5948 = v1642;
assign w5949 = pi359 & ~w5948;
assign w5950 = pi314 & ~w5716;
assign w5951 = w24 & w5946;
assign v1643 = ~(w5950 | w5951);
assign w5952 = v1643;
assign w5953 = pi359 & ~w5952;
assign w5954 = w2900 & w4487;
assign w5955 = ~pi181 & w5954;
assign w5956 = pi315 & ~w5954;
assign w5957 = pi359 & ~w5955;
assign w5958 = ~w5956 & w5957;
assign w5959 = pi138 & w5954;
assign w5960 = pi316 & ~w5954;
assign w5961 = pi359 & ~w5959;
assign w5962 = ~w5960 & w5961;
assign w5963 = pi139 & w5954;
assign w5964 = pi317 & ~w5954;
assign w5965 = pi359 & ~w5963;
assign w5966 = ~w5964 & w5965;
assign w5967 = pi178 & w5954;
assign w5968 = pi318 & ~w5954;
assign w5969 = pi359 & ~w5967;
assign w5970 = ~w5968 & w5969;
assign w5971 = pi142 & w5954;
assign w5972 = pi319 & ~w5954;
assign w5973 = pi359 & ~w5971;
assign w5974 = ~w5972 & w5973;
assign w5975 = pi129 & w5954;
assign w5976 = pi320 & ~w5954;
assign w5977 = pi359 & ~w5975;
assign w5978 = ~w5976 & w5977;
assign w5979 = ~pi180 & w5954;
assign w5980 = pi321 & ~w5954;
assign w5981 = pi359 & ~w5979;
assign w5982 = ~w5980 & w5981;
assign w5983 = pi132 & w5954;
assign w5984 = pi322 & ~w5954;
assign w5985 = pi359 & ~w5983;
assign w5986 = ~w5984 & w5985;
assign w5987 = pi102 & w5954;
assign w5988 = pi323 & ~w5954;
assign w5989 = pi359 & ~w5987;
assign w5990 = ~w5988 & w5989;
assign w5991 = pi184 & w5954;
assign w5992 = pi324 & ~w5954;
assign w5993 = pi359 & ~w5991;
assign w5994 = ~w5992 & w5993;
assign w5995 = pi131 & w5954;
assign w5996 = pi325 & ~w5954;
assign w5997 = pi359 & ~w5995;
assign w5998 = ~w5996 & w5997;
assign w5999 = pi126 & w5954;
assign w6000 = pi326 & ~w5954;
assign w6001 = pi359 & ~w5999;
assign w6002 = ~w6000 & w6001;
assign w6003 = pi141 & w5954;
assign w6004 = pi327 & ~w5954;
assign w6005 = pi359 & ~w6003;
assign w6006 = ~w6004 & w6005;
assign w6007 = pi143 & w5954;
assign w6008 = pi328 & ~w5954;
assign w6009 = pi359 & ~w6007;
assign w6010 = ~w6008 & w6009;
assign w6011 = pi140 & w5954;
assign w6012 = pi329 & ~w5954;
assign w6013 = pi359 & ~w6011;
assign w6014 = ~w6012 & w6013;
assign w6015 = pi133 & w5954;
assign w6016 = pi330 & ~w5954;
assign w6017 = pi359 & ~w6015;
assign w6018 = ~w6016 & w6017;
assign w6019 = ~pi247 & pi301;
assign w6020 = ~w5133 & w6019;
assign v1644 = ~(pi247 | w740);
assign w6021 = v1644;
assign w6022 = ~w1133 & w6021;
assign w6023 = w2893 & w6022;
assign w6024 = w5851 & w6023;
assign v1645 = ~(pi331 | w6024);
assign w6025 = v1645;
assign w6026 = pi359 & ~w6020;
assign w6027 = ~w6025 & w6026;
assign w6028 = ~pi247 & w5628;
assign v1646 = ~(pi332 | w6028);
assign w6029 = v1646;
assign w6030 = ~pi133 & w6028;
assign w6031 = pi359 & ~w6029;
assign w6032 = ~w6030 & w6031;
assign v1647 = ~(pi333 | w6020);
assign w6033 = v1647;
assign w6034 = pi359 & ~w6024;
assign w6035 = ~w6033 & w6034;
assign v1648 = ~(w148 | w983);
assign w6036 = v1648;
assign w6037 = pi359 & ~w6036;
assign w6038 = pi247 & ~pi335;
assign w6039 = w0 & ~w4157;
assign v1649 = ~(pi247 | w5130);
assign w6040 = v1649;
assign w6041 = ~w6039 & w6040;
assign w6042 = pi359 & ~w6038;
assign w6043 = ~w6041 & w6042;
assign w6044 = ~pi247 & w752;
assign w6045 = w2894 & w6044;
assign w6046 = w147 & w6045;
assign w6047 = pi336 & ~w6046;
assign w6048 = w5643 & w6045;
assign v1650 = ~(w6047 | w6048);
assign w6049 = v1650;
assign w6050 = pi359 & ~w6049;
assign w6051 = pi337 & ~w6046;
assign w6052 = w5663 & w6045;
assign v1651 = ~(w6051 | w6052);
assign w6053 = v1651;
assign w6054 = pi359 & ~w6053;
assign w6055 = pi338 & ~w6046;
assign w6056 = w5673 & w6045;
assign v1652 = ~(w6055 | w6056);
assign w6057 = v1652;
assign w6058 = pi359 & ~w6057;
assign v1653 = ~(pi339 | w6046);
assign w6059 = v1653;
assign w6060 = ~pi133 & w6046;
assign w6061 = pi359 & ~w6059;
assign w6062 = ~w6060 & w6061;
assign w6063 = pi340 & ~w6046;
assign w6064 = w5625 & w6045;
assign v1654 = ~(w6063 | w6064);
assign w6065 = v1654;
assign w6066 = pi359 & ~w6065;
assign w6067 = pi341 & ~w6046;
assign w6068 = w5703 & w6045;
assign v1655 = ~(w6067 | w6068);
assign w6069 = v1655;
assign w6070 = pi359 & ~w6069;
assign w6071 = pi342 & ~w6046;
assign w6072 = w5723 & w6045;
assign v1656 = ~(w6071 | w6072);
assign w6073 = v1656;
assign w6074 = pi359 & ~w6073;
assign w6075 = pi343 & ~w6046;
assign w6076 = w5653 & w6045;
assign v1657 = ~(w6075 | w6076);
assign w6077 = v1657;
assign w6078 = pi359 & ~w6077;
assign w6079 = pi344 & w1728;
assign w6080 = w1731 & w5578;
assign v1658 = ~(w6079 | w6080);
assign w6081 = v1658;
assign w6082 = pi131 & ~w120;
assign v1659 = ~(pi102 | pi297);
assign w6083 = v1659;
assign w6084 = pi302 & ~w6083;
assign w6085 = ~w6082 & w6084;
assign w6086 = pi359 & ~w6085;
assign w6087 = w131 & w6086;
assign w6088 = pi304 & w5620;
assign w6089 = ~pi247 & pi314;
assign w6090 = ~w5530 & w6089;
assign w6091 = pi247 & pi346;
assign v1660 = ~(w6090 | w6091);
assign w6092 = v1660;
assign w6093 = ~w6088 & w6092;
assign w6094 = pi347 & ~w982;
assign v1661 = ~(w5769 | w6094);
assign w6095 = v1661;
assign w6096 = pi359 & ~w6095;
assign w6097 = pi348 & ~w982;
assign v1662 = ~(w5811 | w6097);
assign w6098 = v1662;
assign w6099 = pi359 & ~w6098;
assign w6100 = pi349 & ~w982;
assign v1663 = ~(w5745 | w6100);
assign w6101 = v1663;
assign w6102 = pi359 & ~w6101;
assign w6103 = pi350 & ~w982;
assign v1664 = ~(w5781 | w6103);
assign w6104 = v1664;
assign w6105 = pi359 & ~w6104;
assign w6106 = pi351 & ~w982;
assign v1665 = ~(w5683 | w6106);
assign w6107 = v1665;
assign w6108 = pi359 & ~w6107;
assign w6109 = pi352 & ~w982;
assign v1666 = ~(w5799 | w6109);
assign w6110 = v1666;
assign w6111 = pi359 & ~w6110;
assign w6112 = pi353 & ~w982;
assign v1667 = ~(w5757 | w6112);
assign w6113 = v1667;
assign w6114 = pi359 & ~w6113;
assign w6115 = pi354 & ~w982;
assign v1668 = ~(w5733 | w6115);
assign w6116 = v1668;
assign w6117 = pi359 & ~w6116;
assign w6118 = pi357 & ~pi363;
assign v1669 = ~(pi355 | w6118);
assign w6119 = v1669;
assign w6120 = ~pi196 & pi359;
assign w6121 = ~w6119 & w6120;
assign w6122 = pi359 & ~pi364;
assign w6123 = pi359 & pi363;
assign w6124 = pi359 & ~pi362;
assign v1670 = ~(w10 | w7);
assign w6125 = v1670;
assign w6126 = w50 & w37;
assign w6127 = w73 & pi303;
assign w6128 = ~w34 & w0;
assign w6129 = (~pi301 & ~w98) | (~pi301 & w6136) | (~w98 & w6136);
assign v1671 = ~(w116 | w107);
assign w6130 = v1671;
assign w6131 = w85 & w120;
assign w6132 = w133 & ~w135;
assign v1672 = ~(w116 | w143);
assign w6133 = v1672;
assign w6134 = w4268 & w1082;
assign v1673 = ~(w4301 | w4298);
assign w6135 = v1673;
assign v1674 = ~(w99 | pi301);
assign w6136 = v1674;
assign w6137 = ~w0 & w6129;
assign v1675 = ~(w0 | w100);
assign w6138 = v1675;
assign w6139 = pi190 & pi301;
assign w6140 = w149 & ~w141;
assign v1676 = ~(w155 | w154);
assign w6141 = v1676;
assign w6142 = ~w152 & w7309;
assign w6143 = ~w152 & w7310;
assign w6144 = ~w152 & w7311;
assign v1677 = ~(w227 | w228);
assign w6145 = v1677;
assign w6146 = ~w152 & w7312;
assign w6147 = ~w152 & w7313;
assign w6148 = ~w152 & w7314;
assign w6149 = ~w152 & w7315;
assign v1678 = ~(w251 | w252);
assign w6150 = v1678;
assign w6151 = ~w152 & w7316;
assign w6152 = ~w152 & w7317;
assign v1679 = ~(w264 | w265);
assign w6153 = v1679;
assign w6154 = ~w152 & w7318;
assign w6155 = ~w152 & w7319;
assign w6156 = ~w152 & w7320;
assign w6157 = ~w152 & w7321;
assign w6158 = ~w152 & w7322;
assign v1680 = ~(w292 | w293);
assign w6159 = v1680;
assign w6160 = ~w152 & w7323;
assign w6161 = ~w152 & w7324;
assign w6162 = ~w152 & w7325;
assign v1681 = ~(w309 | w310);
assign w6163 = v1681;
assign w6164 = w317 & w97;
assign w6165 = w235 & w97;
assign w6166 = w276 & w97;
assign v1682 = ~(w351 | w352);
assign w6167 = v1682;
assign v1683 = ~(w367 | w368);
assign w6168 = v1683;
assign v1684 = ~(w96 | w147);
assign w6169 = v1684;
assign w6170 = w2999 & w3001;
assign v1685 = ~(w2999 | w3001);
assign w6171 = v1685;
assign v1686 = ~(w4295 | w4293);
assign w6172 = v1686;
assign w6173 = ~w177 & w7326;
assign w6174 = w178 & w6141;
assign w6175 = (~w154 & w183) | (~w154 & w7327) | (w183 & w7327);
assign w6176 = ~w184 & w6141;
assign w6177 = (~pi110 & w152) | (~pi110 & w7338) | (w152 & w7338);
assign w6178 = ~w152 & w7328;
assign v1687 = ~(w171 | pi101);
assign w6179 = v1687;
assign v1688 = ~(w171 | pi104);
assign w6180 = v1688;
assign w6181 = w176 & ~pi103;
assign v1689 = ~(w176 | pi105);
assign w6182 = v1689;
assign w6183 = w176 & ~pi148;
assign v1690 = ~(w176 | pi150);
assign w6184 = v1690;
assign w6185 = ~w152 & w7329;
assign w6186 = (~pi120 & w152) | (~pi120 & w7339) | (w152 & w7339);
assign w6187 = (~pi125 & w152) | (~pi125 & w7340) | (w152 & w7340);
assign w6188 = w176 & ~pi121;
assign v1691 = ~(w176 | pi122);
assign w6189 = v1691;
assign w6190 = (~pi156 & w152) | (~pi156 & w7341) | (w152 & w7341);
assign w6191 = ~w152 & w7330;
assign w6192 = w300 & w259;
assign w6193 = w176 & ~pi067;
assign v1692 = ~(w176 | pi072);
assign w6194 = v1692;
assign w6195 = w176 & ~pi084;
assign v1693 = ~(w176 | pi086);
assign w6196 = v1693;
assign w6197 = w509 & ~w503;
assign w6198 = ~w509 & w503;
assign w6199 = ~w300 & w380;
assign w6200 = w517 & w530;
assign w6201 = w496 & w6221;
assign w6202 = (w537 & ~w496) | (w537 & w6222) | (~w496 & w6222);
assign w6203 = ~w536 & w482;
assign w6204 = ~w547 & w548;
assign v1694 = ~(w866 | w864);
assign w6205 = v1694;
assign w6206 = ~w885 & w854;
assign w6207 = pi285 & pi160;
assign w6208 = ~pi285 & pi159;
assign w6209 = pi285 & pi155;
assign w6210 = ~pi285 & pi127;
assign w6211 = pi285 & pi157;
assign w6212 = ~pi285 & pi154;
assign w6213 = pi285 & pi158;
assign w6214 = ~pi285 & pi156;
assign w6215 = ~w1511 & w1573;
assign w6216 = ~w1511 & w2330;
assign w6217 = ~w1511 & w2407;
assign w6218 = ~w1511 & w2469;
assign v1695 = ~(w3007 | w3002);
assign w6219 = v1695;
assign v1696 = ~(w4290 | w4288);
assign w6220 = v1696;
assign v1697 = ~(w258 | w537);
assign w6221 = v1697;
assign w6222 = w258 & w537;
assign w6223 = w176 & ~pi111;
assign v1698 = ~(w176 | pi113);
assign w6224 = v1698;
assign w6225 = (~pi112 & w152) | (~pi112 & w7342) | (w152 & w7342);
assign v1699 = ~(w486 | w485);
assign w6226 = v1699;
assign w6227 = w499 & ~w217;
assign w6228 = ~w499 & w217;
assign w6229 = w6192 & ~w513;
assign w6230 = ~w6192 & w513;
assign w6231 = ~w526 & w524;
assign w6232 = w526 & ~w524;
assign v1700 = ~(w492 | w258);
assign w6233 = v1700;
assign w6234 = w491 & ~w482;
assign w6235 = w491 & ~w6203;
assign w6236 = ~w547 & w586;
assign w6237 = w547 & ~w586;
assign w6238 = w591 & ~w340;
assign w6239 = ~w1 & pi190;
assign w6240 = pi303 & pi301;
assign w6241 = w73 & pi298;
assign w6242 = w73 & pi302;
assign w6243 = (~pi301 & ~w75) | (~pi301 & w7331) | (~w75 & w7331);
assign w6244 = w133 & w144;
assign v1701 = ~(w147 | w141);
assign w6245 = v1701;
assign v1702 = ~(w149 | w145);
assign w6246 = v1702;
assign w6247 = (w134 & w7332) | (w134 & w7333) | (w7332 & w7333);
assign w6248 = (~w141 & w6140) | (~w141 & w145) | (w6140 & w145);
assign w6249 = w147 & w153;
assign w6250 = (w134 & w7343) | (w134 & w7344) | (w7343 & w7344);
assign w6251 = (~w154 & w6141) | (~w154 & w145) | (w6141 & w145);
assign w6252 = pi303 & pi296;
assign w6253 = w158 & w147;
assign w6254 = w158 & w164;
assign w6255 = pi314 & ~w151;
assign w6256 = (w6174 & w6173) | (w6174 & w143) | (w6173 & w143);
assign w6257 = (w6174 & w6173) | (w6174 & w145) | (w6173 & w145);
assign w6258 = w151 & w179;
assign w6259 = (w6176 & w6175) | (w6176 & w143) | (w6175 & w143);
assign w6260 = (w6176 & w6175) | (w6176 & w145) | (w6175 & w145);
assign w6261 = w151 & w185;
assign w6262 = w176 & ~pi155;
assign v1703 = ~(w176 | pi157);
assign w6263 = v1703;
assign w6264 = ~w6192 & w414;
assign v1704 = ~(w492 | w497);
assign w6265 = v1704;
assign w6266 = ~w517 & w520;
assign v1705 = ~(w492 | w493);
assign w6267 = v1705;
assign v1706 = ~(w343 | w363);
assign w6268 = v1706;
assign v1707 = ~(w492 | w299);
assign w6269 = v1707;
assign w6270 = w572 & w554;
assign w6271 = ~w552 & w6270;
assign v1708 = ~(w572 | w554);
assign w6272 = v1708;
assign w6273 = (~w572 & w552) | (~w572 & w6272) | (w552 & w6272);
assign v1709 = ~(w492 | w488);
assign w6274 = v1709;
assign w6275 = ~w577 & w576;
assign w6276 = w577 & ~w576;
assign w6277 = w582 & ~w548;
assign w6278 = w582 & ~w6204;
assign w6279 = ~w300 & w590;
assign w6280 = w300 & ~w590;
assign w6281 = w341 & ~w597;
assign w6282 = ~w341 & w597;
assign w6283 = ~w596 & w600;
assign w6284 = w606 & ~w502;
assign w6285 = ~w1 & w0;
assign w6286 = ~pi242 & pi000;
assign v1710 = ~(pi216 | pi198);
assign w6287 = v1710;
assign w6288 = w6287 & ~pi217;
assign w6289 = pi216 & pi198;
assign w6290 = pi202 & pi216;
assign w6291 = w629 & pi223;
assign v1711 = ~(w629 | pi223);
assign w6292 = v1711;
assign v1712 = ~(w641 | w633);
assign w6293 = v1712;
assign w6294 = pi132 & ~w628;
assign w6295 = ~w6287 & pi217;
assign w6296 = w646 & w628;
assign w6297 = w646 & ~w6294;
assign w6298 = pi132 & w648;
assign w6299 = pi132 & ~w638;
assign w6300 = w655 & w638;
assign w6301 = w655 & ~w6299;
assign w6302 = w658 & ~pi197;
assign v1713 = ~(pi202 | pi184);
assign w6303 = v1713;
assign v1714 = ~(pi202 | pi129);
assign w6304 = v1714;
assign w6305 = w669 & pi216;
assign v1715 = ~(w669 | pi216);
assign w6306 = v1715;
assign w6307 = pi132 & ~w648;
assign w6308 = ~w684 & pi129;
assign w6309 = w652 & ~w641;
assign w6310 = w622 & pi202;
assign w6311 = w690 & ~w697;
assign w6312 = ~pi241 & pi243;
assign w6313 = pi256 & pi243;
assign w6314 = pi241 & pi243;
assign w6315 = w734 & pi131;
assign w6316 = ~pi298 & pi274;
assign w6317 = pi303 & pi273;
assign w6318 = pi303 & pi275;
assign w6319 = ~pi298 & pi271;
assign w6320 = ~pi303 & pi264;
assign w6321 = pi298 & pi270;
assign w6322 = ~pi298 & pi197;
assign v1716 = ~(w773 | w774);
assign w6323 = v1716;
assign w6324 = ~pi303 & pi223;
assign v1717 = ~(pi256 | w809);
assign w6325 = v1717;
assign w6326 = pi256 & pi264;
assign v1718 = ~(w6326 | pi197);
assign w6327 = v1718;
assign w6328 = w826 & ~w815;
assign v1719 = ~(w860 | w858);
assign w6329 = v1719;
assign w6330 = w848 & w854;
assign w6331 = w848 & w6206;
assign v1720 = ~(w893 | w891);
assign w6332 = v1720;
assign w6333 = ~w898 & w899;
assign w6334 = ~w842 & w899;
assign w6335 = ~w842 & w6333;
assign w6336 = w842 & ~w899;
assign w6337 = w842 & ~w6333;
assign v1721 = ~(w827 | w6334);
assign w6338 = v1721;
assign v1722 = ~(w827 | w6335);
assign w6339 = v1722;
assign w6340 = w848 & ~w827;
assign w6341 = w924 & ~w923;
assign v1723 = ~(pi256 | w867);
assign w6342 = v1723;
assign w6343 = pi256 & pi271;
assign v1724 = ~(w6343 | pi225);
assign w6344 = v1724;
assign v1725 = ~(w818 | w877);
assign w6345 = v1725;
assign w6346 = w818 & w877;
assign w6347 = w935 & ~w933;
assign v1726 = ~(w898 | w827);
assign w6348 = v1726;
assign w6349 = ~w944 & w937;
assign v1727 = ~(w878 | w827);
assign w6350 = v1727;
assign v1728 = ~(pi256 | w849);
assign w6351 = v1728;
assign w6352 = pi256 & pi270;
assign v1729 = ~(w6352 | pi216);
assign w6353 = v1729;
assign w6354 = w885 & ~w854;
assign w6355 = ~w965 & w959;
assign w6356 = w970 & w948;
assign v1730 = ~(w903 | pi344);
assign w6357 = v1730;
assign w6358 = w972 & pi344;
assign w6359 = w972 & ~w6357;
assign w6360 = ~w698 & w976;
assign w6361 = ~w977 & w620;
assign v1731 = ~(w150 | w621);
assign w6362 = v1731;
assign w6363 = ~pi099 & pi361;
assign v1732 = ~(w982 | pi001);
assign w6364 = v1732;
assign w6365 = w986 & pi099;
assign v1733 = ~(w986 | pi099);
assign w6366 = v1733;
assign w6367 = pi302 & ~pi297;
assign w6368 = pi298 & ~pi300;
assign w6369 = w997 & ~w82;
assign w6370 = ~w1009 & w991;
assign v1734 = ~(w987 | pi098);
assign w6371 = v1734;
assign w6372 = w987 & pi098;
assign v1735 = ~(w38 | w8);
assign w6373 = v1735;
assign w6374 = w1028 & pi097;
assign v1736 = ~(w1028 | pi097);
assign w6375 = v1736;
assign w6376 = w982 & ~pi295;
assign w6377 = w1013 & w1035;
assign w6378 = w1037 & w71;
assign w6379 = ~w1046 & w9;
assign w6380 = w1039 & w0;
assign v1737 = ~(w1048 | w0);
assign w6381 = v1737;
assign v1738 = ~(w1048 | w6380);
assign w6382 = v1738;
assign v1739 = ~(w1013 | w1049);
assign w6383 = v1739;
assign w6384 = w0 & w71;
assign v1740 = ~(w1083 | w1080);
assign w6385 = v1740;
assign w6386 = w1096 & pi196;
assign w6387 = ~w1083 & w1101;
assign w6388 = w1106 & w986;
assign w6389 = w1111 & w1109;
assign w6390 = pi302 & pi297;
assign w6391 = w1128 & w1017;
assign w6392 = w1128 & ~pi297;
assign v1741 = ~(pi298 | pi300);
assign w6393 = v1741;
assign v1742 = ~(pi299 | w101);
assign w6394 = v1742;
assign w6395 = w1157 & ~w1152;
assign v1743 = ~(w77 | w1162);
assign w6396 = v1743;
assign w6397 = w1144 & w1164;
assign w6398 = w1171 & ~w1167;
assign w6399 = w73 & ~pi303;
assign v1744 = ~(w1191 | w1002);
assign w6400 = v1744;
assign v1745 = ~(w1 | w1185);
assign w6401 = v1745;
assign w6402 = w157 & pi291;
assign w6403 = ~w157 & w48;
assign w6404 = w1196 & w88;
assign v1746 = ~(pi301 | w1113);
assign w6405 = v1746;
assign v1747 = ~(w1255 | w986);
assign w6406 = v1747;
assign w6407 = w1108 & ~w1259;
assign v1748 = ~(w1248 | w1243);
assign w6408 = v1748;
assign w6409 = ~w1261 & pi301;
assign w6410 = w1208 & ~w1263;
assign w6411 = ~w0 & w1280;
assign w6412 = w986 & ~w1108;
assign w6413 = w1259 & w1284;
assign w6414 = pi190 & ~pi296;
assign w6415 = w1296 & w1261;
assign w6416 = w82 & w122;
assign w6417 = w1311 & w995;
assign w6418 = ~w1321 & w0;
assign w6419 = ~pi301 & w1326;
assign w6420 = ~w1328 & pi206;
assign w6421 = ~w1257 & pi130;
assign w6422 = ~w1283 & w1335;
assign w6423 = w1257 & pi349;
assign v1749 = ~(w1327 | w153);
assign w6424 = v1749;
assign v1750 = ~(w1340 | w1075);
assign w6425 = v1750;
assign w6426 = ~pi291 & pi301;
assign w6427 = w1343 & w2;
assign v1751 = ~(pi282 | pi276);
assign w6428 = v1751;
assign w6429 = w1283 & w1350;
assign w6430 = ~w1088 & w1103;
assign w6431 = w1052 & w1077;
assign w6432 = ~w1050 & w1359;
assign v1752 = ~(pi268 | w6382);
assign w6433 = v1752;
assign v1753 = ~(pi268 | w6381);
assign w6434 = v1753;
assign v1754 = ~(w1013 | w1364);
assign w6435 = v1754;
assign w6436 = ~pi285 & pi147;
assign w6437 = ~pi285 & pi149;
assign w6438 = ~pi285 & pi175;
assign w6439 = pi285 & pi148;
assign w6440 = ~pi285 & pi152;
assign w6441 = pi285 & pi150;
assign w6442 = pi285 & pi153;
assign w6443 = pi285 & pi151;
assign w6444 = ~w1257 & pi172;
assign v1755 = ~(w1764 | pi268);
assign w6445 = v1755;
assign w6446 = w1764 & pi268;
assign w6447 = w1283 & ~w1387;
assign v1756 = ~(w1340 | w1380);
assign w6448 = v1756;
assign w6449 = w1257 & pi351;
assign w6450 = ~w1328 & pi207;
assign v1757 = ~(w1392 | w1393);
assign w6451 = v1757;
assign w6452 = ~w1088 & w1384;
assign w6453 = w1052 & w1382;
assign v1758 = ~(w982 | pi002);
assign w6454 = v1758;
assign w6455 = w982 & ~pi289;
assign w6456 = w1013 & w1401;
assign w6457 = ~w1365 & w1403;
assign v1759 = ~(pi246 | w6382);
assign w6458 = v1759;
assign v1760 = ~(pi246 | w6381);
assign w6459 = v1760;
assign v1761 = ~(w1013 | w1408);
assign w6460 = v1761;
assign w6461 = ~pi285 & pi104;
assign w6462 = pi285 & pi109;
assign w6463 = pi285 & pi103;
assign w6464 = pi285 & pi107;
assign w6465 = ~pi285 & pi106;
assign w6466 = ~pi285 & pi108;
assign w6467 = ~pi285 & pi101;
assign w6468 = pi285 & pi105;
assign v1762 = ~(w1340 | w1424);
assign w6469 = v1762;
assign w6470 = w1764 & w1430;
assign w6471 = w6470 & pi259;
assign w6472 = w1283 & ~w1432;
assign w6473 = ~w1257 & pi144;
assign w6474 = w6471 & ~pi246;
assign w6475 = ~w1328 & pi210;
assign w6476 = w1257 & pi353;
assign v1763 = ~(w1439 | w1438);
assign w6477 = v1763;
assign w6478 = ~w1088 & w1428;
assign w6479 = w1052 & w1426;
assign v1764 = ~(w982 | pi003);
assign w6480 = v1764;
assign w6481 = w982 & ~pi287;
assign w6482 = w1013 & w1448;
assign w6483 = ~w1409 & w1450;
assign v1765 = ~(pi233 | w6382);
assign w6484 = v1765;
assign v1766 = ~(pi233 | w6381);
assign w6485 = v1766;
assign v1767 = ~(w1013 | w1455);
assign w6486 = v1767;
assign w6487 = ~pi285 & pi068;
assign w6488 = pi285 & pi071;
assign w6489 = ~pi285 & pi073;
assign w6490 = pi285 & pi069;
assign w6491 = ~pi285 & pi070;
assign w6492 = pi285 & pi072;
assign w6493 = pi285 & pi067;
assign w6494 = ~pi285 & pi066;
assign w6495 = ~w1257 & pi137;
assign w6496 = w6471 & pi246;
assign v1768 = ~(w6496 | pi233);
assign w6497 = v1768;
assign w6498 = w6496 & pi233;
assign w6499 = w1336 & ~w1477;
assign v1769 = ~(w1340 | w1471);
assign w6500 = v1769;
assign w6501 = w1257 & pi347;
assign w6502 = ~w1328 & pi211;
assign v1770 = ~(w1482 | w1483);
assign w6503 = v1770;
assign w6504 = ~w1088 & w1475;
assign w6505 = w1052 & w1473;
assign v1771 = ~(w982 | pi004);
assign w6506 = v1771;
assign w6507 = w982 & ~pi286;
assign w6508 = w1013 & w1491;
assign w6509 = ~w1456 & w1493;
assign v1772 = ~(pi099 | pi252);
assign w6510 = v1772;
assign w6511 = pi256 & ~pi243;
assign w6512 = pi239 & w1499;
assign v1773 = ~(w1510 | w145);
assign w6513 = v1773;
assign v1774 = ~(w147 | pi361);
assign w6514 = v1774;
assign w6515 = w166 & ~w1508;
assign v1775 = ~(w6515 | pi247);
assign w6516 = v1775;
assign w6517 = pi284 & pi283;
assign w6518 = w1526 & ~pi008;
assign w6519 = ~pi283 & pi284;
assign w6520 = w1529 & ~pi011;
assign v1776 = ~(pi283 | pi284);
assign w6521 = v1776;
assign w6522 = w1532 & ~pi005;
assign w6523 = w1532 & ~pi009;
assign w6524 = w1529 & ~pi007;
assign w6525 = w1526 & ~pi012;
assign w6526 = ~w998 & w0;
assign w6527 = w944 & ~pi243;
assign v1777 = ~(pi298 | pi269);
assign w6528 = v1777;
assign w6529 = pi298 & pi257;
assign w6530 = ~w658 & w701;
assign w6531 = w6313 & pi217;
assign v1778 = ~(w1559 | w1562);
assign w6532 = v1778;
assign v1779 = ~(w1568 | w1569);
assign w6533 = v1779;
assign v1780 = ~(w1551 | w1571);
assign w6534 = v1780;
assign w6535 = w1517 & ~w1573;
assign w6536 = w1517 & ~w6215;
assign v1781 = ~(w1516 | pi005);
assign w6537 = v1781;
assign w6538 = w1577 & ~w1573;
assign w6539 = w1577 & ~w6215;
assign v1782 = ~(w1516 | pi006);
assign w6540 = v1782;
assign w6541 = w1581 & ~w1573;
assign w6542 = w1581 & ~w6215;
assign v1783 = ~(w1516 | pi007);
assign w6543 = v1783;
assign w6544 = w1585 & ~w1573;
assign w6545 = w1585 & ~w6215;
assign v1784 = ~(w1516 | pi008);
assign w6546 = v1784;
assign w6547 = w1589 & ~w1573;
assign w6548 = w1589 & ~w6215;
assign v1785 = ~(w1516 | pi009);
assign w6549 = v1785;
assign w6550 = w1593 & ~w1573;
assign w6551 = w1593 & ~w6215;
assign v1786 = ~(w1516 | pi010);
assign w6552 = v1786;
assign w6553 = w1597 & ~w1573;
assign w6554 = w1597 & ~w6215;
assign v1787 = ~(w1516 | pi011);
assign w6555 = v1787;
assign w6556 = w1601 & ~w1573;
assign w6557 = w1601 & ~w6215;
assign w6558 = w965 & ~pi243;
assign v1788 = ~(pi298 | pi270);
assign w6559 = v1788;
assign w6560 = w6313 & pi216;
assign v1789 = ~(w1610 | w1613);
assign w6561 = v1789;
assign w6562 = w1617 & pi243;
assign w6563 = w1617 & ~w6558;
assign w6564 = w1618 & ~w6563;
assign w6565 = w1618 & ~w6562;
assign v1790 = ~(w1551 | w1621);
assign w6566 = v1790;
assign w6567 = w1529 & ~pi019;
assign w6568 = w1532 & ~pi017;
assign w6569 = w1532 & ~pi013;
assign w6570 = w1526 & ~pi016;
assign w6571 = w1526 & ~pi020;
assign w6572 = ~w1511 & w1639;
assign v1791 = ~(w1516 | pi013);
assign w6573 = v1791;
assign w6574 = w1577 & ~w1639;
assign w6575 = w1577 & ~w6572;
assign v1792 = ~(w1516 | pi014);
assign w6576 = v1792;
assign w6577 = w1581 & ~w1639;
assign w6578 = w1581 & ~w6572;
assign v1793 = ~(w1516 | pi015);
assign w6579 = v1793;
assign w6580 = w1585 & ~w1639;
assign w6581 = w1585 & ~w6572;
assign v1794 = ~(w1516 | pi016);
assign w6582 = v1794;
assign w6583 = w1589 & ~w1639;
assign w6584 = w1589 & ~w6572;
assign v1795 = ~(w1516 | pi017);
assign w6585 = v1795;
assign w6586 = w1593 & ~w1639;
assign w6587 = w1593 & ~w6572;
assign v1796 = ~(w1516 | pi018);
assign w6588 = v1796;
assign w6589 = w1597 & ~w1639;
assign w6590 = w1597 & ~w6572;
assign v1797 = ~(w1516 | pi019);
assign w6591 = v1797;
assign w6592 = w1601 & ~w1639;
assign w6593 = w1601 & ~w6572;
assign v1798 = ~(w1516 | pi020);
assign w6594 = v1798;
assign w6595 = w1529 & pi023;
assign w6596 = w1526 & pi028;
assign w6597 = w1529 & pi027;
assign w6598 = w1526 & pi024;
assign w6599 = w1532 & pi021;
assign w6600 = w1532 & pi025;
assign w6601 = pi298 & ~pi274;
assign w6602 = ~pi298 & pi257;
assign w6603 = w955 & ~pi243;
assign v1799 = ~(w1686 | w1689);
assign w6604 = v1799;
assign w6605 = w1693 & pi243;
assign w6606 = w1693 & ~w6603;
assign w6607 = w1694 & ~w6606;
assign w6608 = w1694 & ~w6605;
assign w6609 = ~w1551 & w1700;
assign v1800 = ~(w1511 | w1702);
assign w6610 = v1800;
assign w6611 = ~w1516 & pi021;
assign w6612 = w1577 & w1702;
assign w6613 = w1577 & ~w6610;
assign w6614 = ~w1516 & pi022;
assign w6615 = w1581 & w1702;
assign w6616 = w1581 & ~w6610;
assign w6617 = ~w1516 & pi023;
assign w6618 = w1585 & w1702;
assign w6619 = w1585 & ~w6610;
assign w6620 = ~w1516 & pi024;
assign w6621 = w1589 & w1702;
assign w6622 = w1589 & ~w6610;
assign w6623 = ~w1516 & pi025;
assign w6624 = w1593 & w1702;
assign w6625 = w1593 & ~w6610;
assign w6626 = ~w1516 & pi026;
assign w6627 = w1597 & w1702;
assign w6628 = w1597 & ~w6610;
assign w6629 = ~w1516 & pi027;
assign w6630 = w1601 & w1702;
assign w6631 = w1601 & ~w6610;
assign w6632 = ~w1516 & pi028;
assign w6633 = w982 & ~pi343;
assign v1801 = ~(pi099 | w982);
assign w6634 = v1801;
assign w6635 = pi348 & ~w6382;
assign w6636 = pi348 & ~w6381;
assign w6637 = ~w1013 & w1735;
assign w6638 = w1013 & pi029;
assign w6639 = ~w1013 & w7368;
assign v1802 = ~(pi285 | pi061);
assign w6640 = v1802;
assign w6641 = pi285 & ~pi060;
assign w6642 = pi285 & ~pi062;
assign w6643 = pi285 & ~pi058;
assign v1803 = ~(pi285 | pi057);
assign w6644 = v1803;
assign v1804 = ~(pi285 | pi059);
assign w6645 = v1804;
assign v1805 = ~(pi285 | pi063);
assign w6646 = v1805;
assign w6647 = pi285 & ~pi064;
assign v1806 = ~(w1340 | w1753);
assign w6648 = v1806;
assign w6649 = w1257 & pi138;
assign w6650 = ~w1328 & pi203;
assign w6651 = pi238 & pi232;
assign w6652 = w6651 & pi222;
assign w6653 = w6652 & pi229;
assign v1807 = ~(w6652 | pi229);
assign w6654 = v1807;
assign w6655 = w1283 & w1775;
assign w6656 = ~w1257 & pi186;
assign w6657 = w1083 & pi229;
assign w6658 = w1784 & pi343;
assign w6659 = ~w1756 & w1787;
assign w6660 = ~w1755 & w1790;
assign w6661 = w982 & ~pi338;
assign w6662 = pi352 & ~w6382;
assign w6663 = pi352 & ~w6381;
assign w6664 = ~w1013 & w1798;
assign w6665 = w1013 & pi030;
assign w6666 = pi285 & ~pi016;
assign w6667 = pi285 & ~pi018;
assign v1808 = ~(pi285 | pi017);
assign w6668 = v1808;
assign v1809 = ~(pi285 | pi019);
assign w6669 = v1809;
assign v1810 = ~(pi285 | pi013);
assign w6670 = v1810;
assign w6671 = pi285 & ~pi020;
assign w6672 = pi285 & ~pi014;
assign v1811 = ~(pi285 | pi015);
assign w6673 = v1811;
assign v1812 = ~(w1340 | w1815);
assign w6674 = v1812;
assign w6675 = ~w1257 & pi177;
assign w6676 = ~w1328 & pi204;
assign w6677 = w1283 & w1827;
assign w6678 = w1257 & pi143;
assign w6679 = w1083 & pi226;
assign w6680 = w1784 & pi338;
assign w6681 = ~w1756 & w1838;
assign w6682 = ~w1817 & w1841;
assign w6683 = w982 & ~pi336;
assign w6684 = pi353 & ~w6382;
assign w6685 = pi353 & ~w6381;
assign w6686 = ~w1013 & w1849;
assign w6687 = w1013 & pi031;
assign v1813 = ~(pi285 | pi056);
assign w6688 = v1813;
assign w6689 = pi285 & ~pi054;
assign v1814 = ~(pi285 | pi051);
assign w6690 = v1814;
assign v1815 = ~(pi285 | pi053);
assign w6691 = v1815;
assign w6692 = pi285 & ~pi055;
assign v1816 = ~(pi285 | pi049);
assign w6693 = v1816;
assign w6694 = pi285 & ~pi050;
assign w6695 = pi285 & ~pi052;
assign v1817 = ~(w1340 | w1866);
assign w6696 = v1817;
assign w6697 = ~w1257 & pi183;
assign w6698 = ~w1328 & pi205;
assign w6699 = pi226 & pi227;
assign v1818 = ~(pi226 | pi227);
assign w6700 = v1818;
assign w6701 = w1283 & w1878;
assign w6702 = w1257 & pi139;
assign w6703 = w1083 & pi227;
assign w6704 = w1784 & pi336;
assign w6705 = ~w1756 & w1889;
assign w6706 = ~w1868 & w1892;
assign w6707 = w982 & ~pi340;
assign w6708 = pi347 & ~w6382;
assign w6709 = pi347 & ~w6381;
assign w6710 = ~w1013 & w1900;
assign w6711 = w1013 & pi032;
assign v1819 = ~(pi285 | pi005);
assign w6712 = v1819;
assign v1820 = ~(pi285 | pi011);
assign w6713 = v1820;
assign v1821 = ~(pi285 | pi009);
assign w6714 = v1821;
assign v1822 = ~(pi285 | pi007);
assign w6715 = v1822;
assign w6716 = pi285 & ~pi006;
assign w6717 = pi285 & ~pi010;
assign w6718 = pi285 & ~pi012;
assign w6719 = pi285 & ~pi008;
assign v1823 = ~(w1340 | w1917);
assign w6720 = v1823;
assign w6721 = ~w1257 & pi117;
assign w6722 = ~w1328 & pi219;
assign v1824 = ~(w6699 | pi191);
assign w6723 = v1824;
assign w6724 = w6699 & pi191;
assign w6725 = w1283 & w1929;
assign w6726 = w1257 & pi140;
assign w6727 = w1083 & pi191;
assign w6728 = w1784 & pi340;
assign w6729 = ~w1756 & w1940;
assign w6730 = ~w1919 & w1943;
assign w6731 = w982 & ~pi337;
assign w6732 = w1013 & ~pi033;
assign w6733 = pi351 & ~w6382;
assign w6734 = pi351 & ~w6381;
assign v1825 = ~(w1013 | w1952);
assign w6735 = v1825;
assign w6736 = ~pi285 & pi021;
assign w6737 = ~pi285 & pi027;
assign w6738 = pi285 & pi028;
assign w6739 = pi285 & pi026;
assign w6740 = ~pi285 & pi025;
assign w6741 = pi285 & pi022;
assign w6742 = ~pi285 & pi023;
assign w6743 = pi285 & pi024;
assign v1826 = ~(w1340 | w1969);
assign w6744 = v1826;
assign w6745 = w1257 & pi141;
assign w6746 = ~w1328 & pi221;
assign v1827 = ~(w6651 | pi222);
assign w6747 = v1827;
assign w6748 = w1283 & w1980;
assign w6749 = ~w1257 & pi182;
assign w6750 = w1083 & pi222;
assign w6751 = w1784 & pi337;
assign w6752 = ~w1756 & w1991;
assign w6753 = ~w1971 & w1993;
assign w6754 = w982 & ~pi290;
assign w6755 = pi259 & ~w6382;
assign w6756 = pi259 & ~w6381;
assign w6757 = ~w1013 & w2001;
assign w6758 = w1013 & pi034;
assign w6759 = ~pi285 & pi110;
assign w6760 = pi285 & pi115;
assign w6761 = ~pi285 & pi100;
assign w6762 = pi285 & pi113;
assign w6763 = pi285 & pi116;
assign w6764 = ~pi285 & pi114;
assign w6765 = ~pi285 & pi112;
assign w6766 = pi285 & pi111;
assign v1828 = ~(pi259 | w1052);
assign w6767 = v1828;
assign v1829 = ~(w6470 | pi259);
assign w6768 = v1829;
assign v1830 = ~(w1340 | w2018);
assign w6769 = v1830;
assign w6770 = w1257 & pi352;
assign w6771 = ~w1328 & pi209;
assign v1831 = ~(pi146 | w2025);
assign w6772 = v1831;
assign v1832 = ~(w2026 | w2027);
assign w6773 = v1832;
assign w6774 = ~w1756 & w2022;
assign w6775 = ~w2020 & w2033;
assign w6776 = w982 & pi292;
assign w6777 = ~w982 & pi035;
assign w6778 = w1013 & ~w2040;
assign v1833 = ~(pi282 | w6382);
assign w6779 = v1833;
assign v1834 = ~(pi282 | w6381);
assign w6780 = v1834;
assign v1835 = ~(w1013 | w2042);
assign w6781 = v1835;
assign w6782 = pi285 & pi170;
assign w6783 = pi285 & pi171;
assign w6784 = ~pi285 & pi169;
assign w6785 = ~pi285 & pi167;
assign w6786 = ~pi285 & pi176;
assign w6787 = pi285 & pi168;
assign w6788 = pi285 & pi166;
assign w6789 = ~pi285 & pi165;
assign w6790 = ~w1257 & pi174;
assign v1836 = ~(w1340 | w2058);
assign w6791 = v1836;
assign w6792 = w1283 & w2065;
assign w6793 = ~w1328 & pi220;
assign w6794 = w1257 & pi354;
assign v1837 = ~(w1756 | w2061);
assign w6795 = v1837;
assign w6796 = w1052 & w2060;
assign w6797 = ~w2043 & w2077;
assign w6798 = w982 & ~pi288;
assign w6799 = pi265 & ~w6382;
assign w6800 = pi265 & ~w6381;
assign w6801 = ~w1013 & w2085;
assign w6802 = w1013 & pi036;
assign w6803 = pi285 & pi122;
assign w6804 = pi285 & pi118;
assign w6805 = pi285 & pi124;
assign w6806 = pi285 & pi121;
assign w6807 = ~pi285 & pi125;
assign w6808 = ~pi285 & pi123;
assign w6809 = ~pi285 & pi120;
assign w6810 = ~pi285 & pi119;
assign v1838 = ~(pi265 | w1052);
assign w6811 = v1838;
assign v1839 = ~(w6446 | pi265);
assign w6812 = v1839;
assign w6813 = w1283 & ~w1431;
assign v1840 = ~(w1340 | w2102);
assign w6814 = v1840;
assign w6815 = ~w1257 & pi173;
assign w6816 = ~w1328 & pi208;
assign v1841 = ~(pi348 | w2110);
assign w6817 = v1841;
assign v1842 = ~(w2111 | w2112);
assign w6818 = v1842;
assign w6819 = ~w1756 & w2105;
assign w6820 = ~w2104 & w2118;
assign w6821 = w982 & ~pi339;
assign w6822 = w1013 & ~pi037;
assign w6823 = pi350 & ~w6382;
assign w6824 = pi350 & ~w6381;
assign v1843 = ~(w1013 | w2127);
assign w6825 = v1843;
assign w6826 = pi285 & pi044;
assign w6827 = pi285 & pi046;
assign w6828 = pi285 & pi042;
assign w6829 = ~pi285 & pi043;
assign w6830 = ~pi285 & pi045;
assign w6831 = pi285 & pi048;
assign w6832 = ~pi285 & pi041;
assign w6833 = ~pi285 & pi047;
assign v1844 = ~(w1340 | w2144);
assign w6834 = v1844;
assign w6835 = ~w1257 & pi179;
assign w6836 = ~w1328 & pi218;
assign w6837 = ~w6724 & pi224;
assign w6838 = w6724 & ~pi224;
assign w6839 = w1283 & w2155;
assign w6840 = w1257 & pi133;
assign w6841 = w1083 & ~pi224;
assign w6842 = w1784 & pi339;
assign w6843 = ~w1756 & w2166;
assign w6844 = w2167 & ~w2166;
assign w6845 = w2167 & ~w6843;
assign w6846 = w2168 & ~w6845;
assign w6847 = w2168 & ~w6844;
assign w6848 = w982 & ~pi341;
assign w6849 = pi354 & ~w6382;
assign w6850 = pi354 & ~w6381;
assign w6851 = ~w1013 & w2176;
assign w6852 = w1013 & pi038;
assign w6853 = ~pi285 & pi090;
assign w6854 = pi285 & pi093;
assign w6855 = pi285 & pi091;
assign w6856 = pi285 & pi096;
assign w6857 = pi285 & pi094;
assign w6858 = ~pi285 & pi095;
assign w6859 = ~pi285 & pi081;
assign w6860 = ~pi285 & pi092;
assign v1845 = ~(w1340 | w2193);
assign w6861 = v1845;
assign w6862 = w1257 & pi126;
assign w6863 = ~w1328 & pi212;
assign w6864 = w1283 & w2204;
assign w6865 = ~w1257 & pi187;
assign w6866 = w1083 & pi238;
assign w6867 = w1784 & pi341;
assign w6868 = ~w1756 & w2215;
assign w6869 = ~w2195 & w2218;
assign w6870 = w982 & ~pi332;
assign w6871 = ~pi285 & pi083;
assign w6872 = ~pi285 & pi089;
assign w6873 = ~pi285 & pi087;
assign w6874 = pi285 & pi088;
assign w6875 = ~pi285 & pi085;
assign w6876 = pi285 & pi082;
assign w6877 = pi285 & pi086;
assign w6878 = pi285 & pi084;
assign v1846 = ~(pi244 | w1052);
assign w6879 = v1846;
assign v1847 = ~(w1340 | w2240);
assign w6880 = v1847;
assign w6881 = w1336 & pi244;
assign w6882 = ~w1328 & pi200;
assign w6883 = w1257 & pi350;
assign w6884 = w2250 & ~w2249;
assign w6885 = w2246 & w1756;
assign w6886 = ~w2243 & w2242;
assign w6887 = pi244 & ~w6382;
assign w6888 = pi244 & ~w6381;
assign w6889 = ~w1013 & w2254;
assign v1848 = ~(pi039 | w1732);
assign w6890 = v1848;
assign w6891 = w2257 & ~w2242;
assign w6892 = w2257 & ~w6886;
assign w6893 = w2259 & ~w6892;
assign w6894 = w2259 & ~w6891;
assign w6895 = w982 & ~pi342;
assign w6896 = pi349 & ~w6382;
assign w6897 = pi349 & ~w6381;
assign w6898 = ~w1013 & w2265;
assign w6899 = w1013 & pi040;
assign w6900 = ~pi285 & pi076;
assign w6901 = ~pi285 & pi079;
assign w6902 = pi285 & pi075;
assign w6903 = pi285 & pi080;
assign v1849 = ~(w1340 | w2282);
assign w6904 = v1849;
assign w6905 = ~w1328 & pi199;
assign v1850 = ~(pi238 | pi232);
assign w6906 = v1850;
assign w6907 = w1283 & w2292;
assign w6908 = w1257 & pi142;
assign v1851 = ~(pi185 | w2285);
assign w6909 = v1851;
assign w6910 = w1083 & pi232;
assign w6911 = w1784 & pi342;
assign w6912 = ~w1756 & w2303;
assign w6913 = ~w2284 & w2306;
assign w6914 = w6313 & pi223;
assign w6915 = ~w690 & w701;
assign w6916 = w837 & ~pi243;
assign w6917 = pi303 & pi257;
assign w6918 = w2318 & pi242;
assign v1852 = ~(w2325 | w2326);
assign w6919 = v1852;
assign v1853 = ~(w1551 | w2328);
assign w6920 = v1853;
assign v1854 = ~(w162 | w2328);
assign w6921 = v1854;
assign w6922 = ~w162 & w6920;
assign w6923 = w1529 & pi043;
assign w6924 = w1526 & pi048;
assign w6925 = w1526 & pi044;
assign w6926 = w1532 & pi045;
assign w6927 = w1529 & pi047;
assign w6928 = w1532 & pi041;
assign w6929 = ~w1511 & w2371;
assign w6930 = w1529 & ~pi056;
assign w6931 = w1532 & ~pi049;
assign w6932 = w1526 & ~pi054;
assign w6933 = w1529 & ~pi051;
assign w6934 = w1526 & ~pi052;
assign w6935 = w1532 & ~pi053;
assign w6936 = w6313 & pi198;
assign w6937 = ~w701 & w2393;
assign w6938 = w844 & w735;
assign w6939 = ~w2398 & pi242;
assign w6940 = pi243 & w2400;
assign w6941 = w2403 & w1551;
assign v1855 = ~(w2405 | w1551);
assign w6942 = v1855;
assign v1856 = ~(w2405 | w6941);
assign w6943 = v1856;
assign v1857 = ~(w162 | w6942);
assign w6944 = v1857;
assign v1858 = ~(w162 | w6943);
assign w6945 = v1858;
assign w6946 = w1517 & ~w2407;
assign w6947 = w1517 & ~w6217;
assign v1859 = ~(w1516 | pi049);
assign w6948 = v1859;
assign w6949 = w1577 & ~w2407;
assign w6950 = w1577 & ~w6217;
assign v1860 = ~(w1516 | pi050);
assign w6951 = v1860;
assign w6952 = w1581 & ~w2407;
assign w6953 = w1581 & ~w6217;
assign v1861 = ~(w1516 | pi051);
assign w6954 = v1861;
assign w6955 = w1585 & ~w2407;
assign w6956 = w1585 & ~w6217;
assign v1862 = ~(w1516 | pi052);
assign w6957 = v1862;
assign w6958 = w1589 & ~w2407;
assign w6959 = w1589 & ~w6217;
assign v1863 = ~(w1516 | pi053);
assign w6960 = v1863;
assign w6961 = w1601 & ~w2407;
assign w6962 = w1601 & ~w6217;
assign v1864 = ~(w1516 | pi054);
assign w6963 = v1864;
assign w6964 = w1593 & ~w2407;
assign w6965 = w1593 & ~w6217;
assign v1865 = ~(w1516 | pi055);
assign w6966 = v1865;
assign w6967 = w1597 & ~w2407;
assign w6968 = w1597 & ~w6217;
assign w6969 = w1529 & ~pi059;
assign w6970 = w1529 & ~pi063;
assign w6971 = w1532 & ~pi061;
assign w6972 = w1532 & ~pi057;
assign w6973 = w1526 & ~pi060;
assign w6974 = w1526 & ~pi064;
assign w6975 = w2445 & w162;
assign v1866 = ~(pi303 | pi272);
assign w6976 = v1866;
assign w6977 = w2458 & w2462;
assign w6978 = pi243 & w2463;
assign w6979 = pi242 & w2463;
assign w6980 = pi242 & w6978;
assign w6981 = w1552 & ~w2466;
assign v1867 = ~(w1551 | w162);
assign w6982 = v1867;
assign v1868 = ~(w2447 | w2469);
assign w6983 = v1868;
assign v1869 = ~(w2447 | w6218);
assign w6984 = v1869;
assign w6985 = ~w1516 & pi057;
assign w6986 = ~w1516 & pi058;
assign w6987 = ~w1516 & pi059;
assign w6988 = ~w1516 & pi060;
assign w6989 = ~w1516 & pi061;
assign w6990 = ~w1516 & pi062;
assign w6991 = ~w1516 & pi063;
assign w6992 = ~w1516 & pi064;
assign w6993 = w1529 & pi076;
assign w6994 = w1529 & pi079;
assign w6995 = w1532 & pi078;
assign w6996 = w1526 & pi080;
assign w6997 = w1532 & pi074;
assign w6998 = w1526 & pi077;
assign w6999 = pi298 & ~pi271;
assign w7000 = pi243 & w2522;
assign v1870 = ~(pi242 | w2524);
assign w7001 = v1870;
assign w7002 = w1552 & ~w2526;
assign w7003 = ~w1551 & w2529;
assign v1871 = ~(w1511 | w2531);
assign w7004 = v1871;
assign w7005 = ~w1516 & pi065;
assign w7006 = ~pi239 & w1499;
assign w7007 = w166 & ~w2536;
assign w7008 = w1526 & pi072;
assign w7009 = w1526 & pi071;
assign w7010 = w1532 & pi066;
assign w7011 = w1532 & pi073;
assign w7012 = w1529 & pi068;
assign w7013 = w1529 & pi070;
assign w7014 = w2552 & w162;
assign w7015 = ~w1551 & w2558;
assign v1872 = ~(w2559 | w2555);
assign w7016 = v1872;
assign v1873 = ~(w2538 | pi066);
assign w7017 = v1873;
assign v1874 = ~(w2538 | pi067);
assign w7018 = v1874;
assign v1875 = ~(w2538 | pi068);
assign w7019 = v1875;
assign v1876 = ~(w2538 | pi069);
assign w7020 = v1876;
assign v1877 = ~(w2538 | pi070);
assign w7021 = v1877;
assign v1878 = ~(w2538 | pi071);
assign w7022 = v1878;
assign v1879 = ~(w2538 | pi072);
assign w7023 = v1879;
assign v1880 = ~(w2538 | pi073);
assign w7024 = v1880;
assign w7025 = w1517 & w2531;
assign w7026 = w1517 & ~w7004;
assign w7027 = ~w1516 & pi074;
assign w7028 = w1577 & w2531;
assign w7029 = w1577 & ~w7004;
assign w7030 = ~w1516 & pi075;
assign w7031 = w1581 & w2531;
assign w7032 = w1581 & ~w7004;
assign w7033 = ~w1516 & pi076;
assign w7034 = w1585 & w2531;
assign w7035 = w1585 & ~w7004;
assign w7036 = ~w1516 & pi077;
assign w7037 = w1589 & w2531;
assign w7038 = w1589 & ~w7004;
assign w7039 = ~w1516 & pi078;
assign w7040 = w1597 & w2531;
assign w7041 = w1597 & ~w7004;
assign w7042 = ~w1516 & pi079;
assign w7043 = w1601 & w2531;
assign w7044 = w1601 & ~w7004;
assign w7045 = ~w1516 & pi080;
assign w7046 = w1526 & pi096;
assign w7047 = w1529 & pi095;
assign w7048 = w1529 & pi092;
assign w7049 = w1532 & pi081;
assign w7050 = w1526 & pi093;
assign w7051 = w1532 & pi090;
assign w7052 = w779 & w736;
assign w7053 = pi303 & ~pi264;
assign w7054 = ~pi303 & pi257;
assign w7055 = ~w2644 & w2645;
assign v1881 = ~(w162 | w2629);
assign w7056 = v1881;
assign w7057 = ~w1511 & w2651;
assign w7058 = w2628 & w1589;
assign v1882 = ~(w1516 | pi081);
assign w7059 = v1882;
assign v1883 = ~(w1551 | w2657);
assign w7060 = v1883;
assign w7061 = w1529 & pi085;
assign w7062 = w1532 & pi087;
assign w7063 = w1526 & pi082;
assign w7064 = w1532 & pi083;
assign w7065 = w1529 & pi089;
assign w7066 = w1526 & pi086;
assign w7067 = ~w2671 & w162;
assign w7068 = w162 & ~w2674;
assign w7069 = ~w2675 & w2580;
assign w7070 = ~w2538 & pi082;
assign w7071 = ~w2675 & w2539;
assign w7072 = ~w2538 & pi083;
assign w7073 = ~w2675 & w2564;
assign w7074 = ~w2538 & pi084;
assign w7075 = ~w2675 & w2568;
assign w7076 = ~w2538 & pi085;
assign w7077 = ~w2675 & w2584;
assign w7078 = ~w2538 & pi086;
assign w7079 = ~w2675 & w2588;
assign w7080 = ~w2538 & pi087;
assign w7081 = ~w2675 & w2572;
assign w7082 = ~w2538 & pi088;
assign w7083 = ~w2675 & w2576;
assign w7084 = ~w1516 & pi090;
assign w7085 = ~w2628 & w1517;
assign w7086 = w2628 & w1577;
assign v1884 = ~(w1516 | pi091);
assign w7087 = v1884;
assign w7088 = w2628 & w1581;
assign v1885 = ~(w1516 | pi092);
assign w7089 = v1885;
assign w7090 = w2628 & w1585;
assign v1886 = ~(w1516 | pi093);
assign w7091 = v1886;
assign w7092 = w2628 & w1593;
assign v1887 = ~(w1516 | pi094);
assign w7093 = v1887;
assign w7094 = w2628 & w1597;
assign v1888 = ~(w1516 | pi095);
assign w7095 = v1888;
assign w7096 = w2628 & w1601;
assign v1889 = ~(w1013 | pi356);
assign w7097 = v1889;
assign v1890 = ~(w38 | pi237);
assign w7098 = v1890;
assign w7099 = ~pi190 & pi301;
assign w7100 = w1233 & w2726;
assign w7101 = pi252 & ~w2723;
assign w7102 = pi361 & ~w2733;
assign w7103 = w1013 & w2734;
assign w7104 = w2731 & pi097;
assign v1891 = ~(w2731 | pi097);
assign w7105 = v1891;
assign w7106 = w146 & ~w2723;
assign w7107 = w146 & w7101;
assign v1892 = ~(w7104 | pi098);
assign w7108 = v1892;
assign v1893 = ~(w2741 | pi099);
assign w7109 = v1893;
assign w7110 = pi356 & ~w2741;
assign v1894 = ~(pi356 | w2733);
assign w7111 = v1894;
assign w7112 = pi359 & pi099;
assign w7113 = pi359 & ~w7109;
assign w7114 = w1529 & pi114;
assign w7115 = w1532 & pi100;
assign w7116 = w1526 & pi113;
assign w7117 = w1526 & pi115;
assign w7118 = w1529 & pi112;
assign w7119 = w1532 & pi110;
assign w7120 = w2767 & w162;
assign w7121 = ~w1551 & w2772;
assign v1895 = ~(w2773 | w2769);
assign w7122 = v1895;
assign v1896 = ~(w2538 | pi100);
assign w7123 = v1896;
assign w7124 = w1529 & pi108;
assign w7125 = w1526 & pi105;
assign w7126 = w1526 & pi109;
assign w7127 = w1532 & pi106;
assign w7128 = w1529 & pi104;
assign w7129 = w1532 & pi101;
assign v1897 = ~(w2797 | w2793);
assign w7130 = v1897;
assign v1898 = ~(w2538 | pi101);
assign w7131 = v1898;
assign v1899 = ~(pi251 | pi240);
assign w7132 = v1899;
assign w7133 = ~pi239 & w2804;
assign w7134 = ~w1696 & w2805;
assign w7135 = w130 & pi000;
assign v1900 = ~(pi242 | w745);
assign w7136 = v1900;
assign v1901 = ~(w841 | w899);
assign w7137 = v1901;
assign v1902 = ~(w841 | w6333);
assign w7138 = v1902;
assign w7139 = w911 & ~w926;
assign w7140 = w944 & ~w937;
assign w7141 = w965 & ~w959;
assign w7142 = w2813 & ~pi344;
assign w7143 = ~w2834 & w2835;
assign w7144 = w734 & pi102;
assign w7145 = ~w690 & w697;
assign w7146 = ~w658 & pi197;
assign w7147 = w643 & ~pi129;
assign w7148 = w643 & ~w6308;
assign w7149 = w2875 & w2873;
assign v1903 = ~(w2875 | w2873);
assign w7150 = v1903;
assign w7151 = w2869 & w701;
assign v1904 = ~(w762 | w2849);
assign w7152 = v1904;
assign w7153 = w2863 & w2886;
assign w7154 = ~w1013 & w2891;
assign w7155 = pi301 & pi296;
assign w7156 = w7155 & w751;
assign w7157 = ~w2895 & pi193;
assign w7158 = w2903 & w2905;
assign w7159 = w2810 & w2907;
assign v1905 = ~(w2929 | w2807);
assign w7160 = v1905;
assign w7161 = ~w2930 & w2931;
assign v1906 = ~(w2538 | pi103);
assign w7162 = v1906;
assign v1907 = ~(w2538 | pi104);
assign w7163 = v1907;
assign v1908 = ~(w2538 | pi105);
assign w7164 = v1908;
assign v1909 = ~(w2538 | pi106);
assign w7165 = v1909;
assign v1910 = ~(w2538 | pi107);
assign w7166 = v1910;
assign v1911 = ~(w2538 | pi108);
assign w7167 = v1911;
assign v1912 = ~(w2538 | pi109);
assign w7168 = v1912;
assign v1913 = ~(w2538 | pi110);
assign w7169 = v1913;
assign v1914 = ~(w2538 | pi111);
assign w7170 = v1914;
assign v1915 = ~(w2538 | pi112);
assign w7171 = v1915;
assign v1916 = ~(w2538 | pi113);
assign w7172 = v1916;
assign v1917 = ~(w2538 | pi114);
assign w7173 = v1917;
assign v1918 = ~(w2538 | pi115);
assign w7174 = v1918;
assign v1919 = ~(w2538 | pi116);
assign w7175 = v1919;
assign v1920 = ~(pi099 | pi350);
assign w7176 = v1920;
assign w7177 = pi099 & pi117;
assign v1921 = ~(w147 | w2983);
assign w7178 = v1921;
assign v1922 = ~(w2980 | w2984);
assign w7179 = v1922;
assign w7180 = pi099 & pi185;
assign v1923 = ~(w147 | w2988);
assign w7181 = v1923;
assign w7182 = pi099 & pi187;
assign v1924 = ~(w147 | w2991);
assign w7183 = v1924;
assign v1925 = ~(pi099 | pi353);
assign w7184 = v1925;
assign w7185 = pi099 & pi144;
assign v1926 = ~(w147 | w2996);
assign w7186 = v1926;
assign v1927 = ~(pi099 | pi349);
assign w7187 = v1927;
assign w7188 = pi099 & pi130;
assign v1928 = ~(w147 | w3000);
assign w7189 = v1928;
assign w7190 = pi099 & pi174;
assign w7191 = ~pi099 & pi354;
assign v1929 = ~(w3006 | w3005);
assign w7192 = v1929;
assign v1930 = ~(pi099 | pi351);
assign w7193 = v1930;
assign w7194 = pi099 & pi172;
assign v1931 = ~(w147 | w3012);
assign w7195 = v1931;
assign v1932 = ~(pi099 | pi348);
assign w7196 = v1932;
assign w7197 = pi099 & pi173;
assign v1933 = ~(w147 | w3017);
assign w7198 = v1933;
assign v1934 = ~(w3010 | w3013);
assign w7199 = v1934;
assign w7200 = w3016 & w3018;
assign v1935 = ~(pi099 | pi352);
assign w7201 = v1935;
assign w7202 = pi099 & pi146;
assign v1936 = ~(w147 | w3025);
assign w7203 = v1936;
assign w7204 = ~w3021 & w3028;
assign v1937 = ~(w3024 | w3026);
assign w7205 = v1937;
assign w7206 = w2994 & w2997;
assign w7207 = w3030 & w3033;
assign w7208 = pi099 & pi135;
assign v1938 = ~(w147 | w3036);
assign w7209 = v1938;
assign v1939 = ~(pi099 | pi347);
assign w7210 = v1939;
assign w7211 = pi099 & pi137;
assign v1940 = ~(w147 | w3041);
assign w7212 = v1940;
assign v1941 = ~(w2980 | w3037);
assign w7213 = v1941;
assign v1942 = ~(w3039 | w3042);
assign w7214 = v1942;
assign v1943 = ~(w3047 | w3046);
assign w7215 = v1943;
assign w7216 = ~w3048 & w3050;
assign v1944 = ~(w2980 | w2989);
assign w7217 = v1944;
assign v1945 = ~(w2980 | w2992);
assign w7218 = v1945;
assign w7219 = w3053 & ~w3050;
assign w7220 = w3053 & ~w7216;
assign w7221 = pi099 & pi183;
assign v1946 = ~(w147 | w3055);
assign w7222 = v1946;
assign w7223 = pi099 & pi186;
assign v1947 = ~(w147 | w3058);
assign w7224 = v1947;
assign w7225 = pi099 & pi177;
assign v1948 = ~(w147 | w3061);
assign w7226 = v1948;
assign w7227 = pi099 & pi182;
assign v1949 = ~(w147 | w3066);
assign w7228 = v1949;
assign v1950 = ~(w3057 | w3068);
assign w7229 = v1950;
assign w7230 = w3069 & ~w7219;
assign w7231 = w3069 & ~w7220;
assign v1951 = ~(w2980 | w3067);
assign w7232 = v1951;
assign v1952 = ~(w2980 | w3056);
assign w7233 = v1952;
assign v1953 = ~(w2980 | w3059);
assign w7234 = v1953;
assign v1954 = ~(w2980 | w3062);
assign w7235 = v1954;
assign v1955 = ~(w3071 | w3070);
assign w7236 = v1955;
assign v1956 = ~(w164 | w982);
assign w7237 = v1956;
assign w7238 = w3081 & ~w3084;
assign v1957 = ~(w3084 | w1732);
assign w7239 = v1957;
assign w7240 = ~w3086 & w3091;
assign w7241 = ~pi239 & w3092;
assign w7242 = ~w3093 & w1731;
assign w7243 = w1526 & pi124;
assign w7244 = w1526 & pi122;
assign w7245 = w1529 & pi125;
assign w7246 = w1529 & pi119;
assign w7247 = w1532 & pi120;
assign w7248 = w1532 & pi123;
assign w7249 = w517 & ~w520;
assign w7250 = w3117 & w3119;
assign w7251 = w3115 & w2572;
assign v1958 = ~(w2538 | pi118);
assign w7252 = v1958;
assign w7253 = w3115 & w2576;
assign v1959 = ~(w2538 | pi119);
assign w7254 = v1959;
assign w7255 = w3115 & w2539;
assign v1960 = ~(w2538 | pi120);
assign w7256 = v1960;
assign w7257 = w3115 & w2564;
assign v1961 = ~(w2538 | pi121);
assign w7258 = v1961;
assign w7259 = w3115 & w2584;
assign v1962 = ~(w2538 | pi122);
assign w7260 = v1962;
assign w7261 = w3115 & w2588;
assign v1963 = ~(w2538 | pi123);
assign w7262 = v1963;
assign w7263 = w3115 & w2580;
assign v1964 = ~(w2538 | pi124);
assign w7264 = v1964;
assign w7265 = w3115 & w2568;
assign w7266 = w3146 & ~pi239;
assign w7267 = ~w2647 & w3147;
assign w7268 = ~w2895 & pi341;
assign w7269 = w2450 & pi292;
assign w7270 = w3152 & w2897;
assign w7271 = ~w1013 & w3156;
assign w7272 = ~w2901 & pi126;
assign w7273 = pi126 & ~w3154;
assign w7274 = w2898 & w3162;
assign w7275 = w1529 & pi159;
assign w7276 = w1529 & pi156;
assign w7277 = w1532 & pi154;
assign w7278 = w1526 & pi160;
assign w7279 = w1532 & pi127;
assign w7280 = w1526 & pi157;
assign w7281 = w3179 & w162;
assign w7282 = ~w1551 & w3189;
assign w7283 = w3188 & ~w3182;
assign v1965 = ~(w2538 | pi127);
assign w7284 = v1965;
assign w7285 = w3146 & pi239;
assign w7286 = ~w7285 & w1502;
assign w7287 = pi189 & pi301;
assign v1966 = ~(w3198 | pi273);
assign w7288 = v1966;
assign w7289 = w3198 & ~w3202;
assign v1967 = ~(w3196 | w3205);
assign w7290 = v1967;
assign v1968 = ~(w7285 | w1502);
assign w7291 = v1968;
assign v1969 = ~(w2901 | pi129);
assign w7292 = v1969;
assign v1970 = ~(w1013 | w3222);
assign w7293 = v1970;
assign w7294 = w130 & w1501;
assign w7295 = w3217 & w3229;
assign w7296 = pi239 & w3092;
assign w7297 = ~pi099 & pi130;
assign w7298 = ~w3087 & w3241;
assign v1971 = ~(w3235 | pi247);
assign w7299 = v1971;
assign w7300 = w2805 & ~w1569;
assign w7301 = w2805 & w6533;
assign v1972 = ~(w977 | w2810);
assign w7302 = v1972;
assign w7303 = w3254 & w2810;
assign w7304 = w3254 & ~w7302;
assign v1973 = ~(w3258 | w7303);
assign w7305 = v1973;
assign v1974 = ~(w3258 | w7304);
assign w7306 = v1974;
assign w7307 = ~w2647 & w2805;
assign w7308 = pi132 & w701;
assign w7309 = w156 & w7345;
assign w7310 = w156 & w7346;
assign w7311 = w156 & w7347;
assign w7312 = w170 & pi109;
assign w7313 = w170 & pi107;
assign w7314 = w170 & ~pi106;
assign w7315 = w170 & ~pi108;
assign w7316 = w156 & w7348;
assign w7317 = w156 & w7349;
assign w7318 = w156 & w7350;
assign w7319 = w156 & w7351;
assign w7320 = w156 & w7352;
assign w7321 = w156 & w7353;
assign w7322 = w156 & w7354;
assign w7323 = w156 & w7355;
assign w7324 = w156 & w7356;
assign w7325 = w156 & w7357;
assign v1975 = ~(w162 | w154);
assign w7326 = v1975;
assign w7327 = w162 & ~w154;
assign w7328 = w156 & w7358;
assign w7329 = w156 & w7359;
assign w7330 = w156 & w7360;
assign v1976 = ~(w73 | pi301);
assign w7331 = v1976;
assign w7332 = w6140 & ~w141;
assign w7333 = (~w141 & w6140) | (~w141 & ~w142) | (w6140 & ~w142);
assign w7334 = w610 & w608;
assign v1977 = ~(w3016 | w3018);
assign w7335 = v1977;
assign w7336 = w3024 & w3026;
assign v1978 = ~(w4316 | w4285);
assign w7337 = v1978;
assign v1979 = ~(w170 | pi110);
assign w7338 = v1979;
assign v1980 = ~(w170 | pi120);
assign w7339 = v1980;
assign v1981 = ~(w170 | pi125);
assign w7340 = v1981;
assign v1982 = ~(w170 | pi156);
assign w7341 = v1982;
assign v1983 = ~(w170 | pi112);
assign w7342 = v1983;
assign w7343 = w6141 & ~w154;
assign w7344 = (~w154 & w6141) | (~w154 & ~w142) | (w6141 & ~w142);
assign w7345 = w169 & pi116;
assign w7346 = w169 & pi115;
assign w7347 = w169 & ~pi100;
assign w7348 = w169 & pi151;
assign w7349 = w169 & pi153;
assign w7350 = w169 & ~pi152;
assign w7351 = w169 & pi124;
assign w7352 = w169 & pi118;
assign w7353 = w169 & ~pi123;
assign w7354 = w169 & ~pi119;
assign w7355 = w169 & pi158;
assign w7356 = w169 & pi160;
assign w7357 = w169 & ~pi159;
assign w7358 = w169 & ~pi114;
assign w7359 = w169 & ~pi175;
assign w7360 = w169 & ~pi127;
assign v1984 = ~(w581 | w546);
assign w7361 = v1984;
assign w7362 = ~w581 & w6277;
assign w7363 = (~w116 & ~w149) | (~w116 & w6246) | (~w149 & w6246);
assign w7364 = (w546 & ~w6277) | (w546 & ~w6278) | (~w6277 & ~w6278);
assign w7365 = (~w854 & ~w6206) | (~w854 & ~w884) | (~w6206 & ~w884);
assign w7366 = (~w620 & ~w6361) | (~w620 & ~w973) | (~w6361 & ~w973);
assign w7367 = (~w0 & ~w6380) | (~w0 & ~w1047) | (~w6380 & ~w1047);
assign w7368 = ~w1048 & w7367;
assign w7369 = (~w116 & ~w1510) | (~w116 & w6513) | (~w1510 & w6513);
assign w7370 = (pi243 & ~w6527) | (pi243 & ~w947) | (~w6527 & ~w947);
assign w7371 = (w1571 & ~w6534) | (w1571 & ~w1570) | (~w6534 & ~w1570);
assign w7372 = (~w6565 & ~w6564) | (~w6565 & ~w968) | (~w6564 & ~w968);
assign w7373 = (w1621 & ~w6566) | (w1621 & ~w1620) | (~w6566 & ~w1620);
assign w7374 = (~w1790 & ~w6660) | (~w1790 & ~w1788) | (~w6660 & ~w1788);
assign w7375 = (~w1841 & ~w6682) | (~w1841 & ~w1839) | (~w6682 & ~w1839);
assign w7376 = (~w1892 & ~w6706) | (~w1892 & ~w1890) | (~w6706 & ~w1890);
assign w7377 = (~w1943 & ~w6730) | (~w1943 & ~w1941) | (~w6730 & ~w1941);
assign w7378 = (~w1993 & ~w6753) | (~w1993 & ~w1992) | (~w6753 & ~w1992);
assign w7379 = (~w2033 & ~w6775) | (~w2033 & ~w2031) | (~w6775 & ~w2031);
assign w7380 = (~w2118 & ~w6820) | (~w2118 & ~w2116) | (~w6820 & ~w2116);
assign w7381 = (~w6847 & ~w6846) | (~w6847 & ~w2162) | (~w6846 & ~w2162);
assign w7382 = (~w2218 & ~w6869) | (~w2218 & ~w2216) | (~w6869 & ~w2216);
assign w7383 = (~w2306 & ~w6913) | (~w2306 & ~w2304) | (~w6913 & ~w2304);
assign w7384 = (pi243 & ~w6916) | (pi243 & ~w902) | (~w6916 & ~w902);
assign w7385 = (~w2330 & ~w6216) | (~w2330 & ~w575) | (~w6216 & ~w575);
assign w7386 = (~w2400 & ~w6940) | (~w2400 & ~w916) | (~w6940 & ~w916);
assign w7387 = (~w6979 & ~w6980) | (~w6979 & ~w926) | (~w6980 & ~w926);
assign w7388 = (~w1551 & ~w6941) | (~w1551 & ~w2402) | (~w6941 & ~w2402);
assign w7389 = (w899 & w6333) | (w899 & ~w887) | (w6333 & ~w887);
assign w7390 = (~w2835 & ~w7143) | (~w2835 & ~w2833) | (~w7143 & ~w2833);
assign w7391 = (~w2931 & ~w7161) | (~w2931 & ~w2908) | (~w7161 & ~w2908);
assign w7392 = (~w3050 & ~w7216) | (~w3050 & ~w3045) | (~w7216 & ~w3045);
assign w7393 = (~w7230 & ~w7231) | (~w7230 & ~w3045) | (~w7231 & ~w3045);
assign w7394 = (~w3091 & ~w7240) | (~w3091 & ~w3080) | (~w7240 & ~w3080);
assign w7395 = (~w3162 & ~w7274) | (~w3162 & ~w3161) | (~w7274 & ~w3161);
assign w7396 = (~w7300 & ~w7301) | (~w7300 & ~w1567) | (~w7301 & ~w1567);
assign one = 1;
assign po000 = pi194;// level 0
assign po001 = pi281;// level 0
assign po002 = pi279;// level 0
assign po003 = pi293;// level 0
assign po004 = pi306;// level 0
assign po005 = pi334;// level 0
assign po006 = pi230;// level 0
assign po007 = ~pi247;// level 0
assign po008 = pi035;// level 0
assign po009 = pi001;// level 0
assign po010 = pi002;// level 0
assign po011 = pi036;// level 0
assign po012 = pi034;// level 0
assign po013 = pi003;// level 0
assign po014 = pi004;// level 0
assign po015 = pi039;// level 0
assign po016 = pi038;// level 0
assign po017 = pi040;// level 0
assign po018 = pi033;// level 0
assign po019 = pi029;// level 0
assign po020 = pi030;// level 0
assign po021 = pi031;// level 0
assign po022 = pi032;// level 0
assign po023 = pi037;// level 0
assign po024 = pi161;// level 0
assign po025 = pi162;// level 0
assign po026 = pi163;// level 0
assign po027 = pi164;// level 0
assign po028 = pi145;// level 0
assign po029 = pi128;// level 0
assign po030 = pi136;// level 0
assign po031 = pi134;// level 0
assign po032 = one;// level 0
assign po033 = pi360;// level 0
assign po034 = w980;// level 30
assign po035 = pi247;// level 0
assign po036 = pi000;// level 0
assign po037 = w1362;// level 22
assign po038 = w1406;// level 22
assign po039 = w1453;// level 22
assign po040 = w1496;// level 22
assign po041 = ~w1576;// level 28
assign po042 = ~w1580;// level 28
assign po043 = ~w1584;// level 28
assign po044 = ~w1588;// level 28
assign po045 = ~w1592;// level 28
assign po046 = ~w1596;// level 28
assign po047 = ~w1600;// level 28
assign po048 = ~w1604;// level 28
assign po049 = ~w1643;// level 28
assign po050 = ~w1646;// level 27
assign po051 = ~w1649;// level 27
assign po052 = ~w1652;// level 27
assign po053 = ~w1655;// level 27
assign po054 = ~w1658;// level 27
assign po055 = ~w1661;// level 27
assign po056 = ~w1664;// level 27
assign po057 = ~w1706;// level 28
assign po058 = ~w1709;// level 27
assign po059 = ~w1712;// level 27
assign po060 = ~w1715;// level 27
assign po061 = ~w1718;// level 27
assign po062 = ~w1721;// level 27
assign po063 = ~w1724;// level 27
assign po064 = ~w1727;// level 27
assign po065 = ~w1794;// level 22
assign po066 = ~w1845;// level 22
assign po067 = ~w1896;// level 22
assign po068 = ~w1947;// level 22
assign po069 = ~w1997;// level 22
assign po070 = ~w2037;// level 22
assign po071 = w2081;// level 22
assign po072 = ~w2122;// level 22
assign po073 = ~w2172;// level 21
assign po074 = ~w2222;// level 22
assign po075 = ~w2261;// level 21
assign po076 = ~w2310;// level 22
assign po077 = pi041;// level 0
assign po078 = w1516;// level 13
assign po079 = ~w2333;// level 28
assign po080 = pi042;// level 0
assign po081 = ~w2336;// level 28
assign po082 = pi043;// level 0
assign po083 = ~w2356;// level 28
assign po084 = pi044;// level 0
assign po085 = ~w2359;// level 28
assign po086 = pi045;// level 0
assign po087 = ~w2362;// level 28
assign po088 = pi046;// level 0
assign po089 = ~w2365;// level 28
assign po090 = pi047;// level 0
assign po091 = ~w2369;// level 28
assign po092 = pi048;// level 0
assign po093 = w2373;// level 27
assign po094 = ~w2410;// level 28
assign po095 = ~w2413;// level 28
assign po096 = ~w2416;// level 28
assign po097 = ~w2419;// level 28
assign po098 = ~w2422;// level 28
assign po099 = ~w2425;// level 28
assign po100 = ~w2428;// level 28
assign po101 = ~w2431;// level 28
assign po102 = w2473;// level 29
assign po103 = w2476;// level 29
assign po104 = w2479;// level 29
assign po105 = w2482;// level 29
assign po106 = w2485;// level 29
assign po107 = w2488;// level 29
assign po108 = w2491;// level 29
assign po109 = w2494;// level 29
assign po110 = ~w2535;// level 28
assign po111 = w2563;// level 27
assign po112 = w2567;// level 27
assign po113 = w2571;// level 27
assign po114 = w2575;// level 27
assign po115 = w2579;// level 27
assign po116 = w2583;// level 27
assign po117 = w2587;// level 27
assign po118 = w2591;// level 27
assign po119 = ~w2594;// level 27
assign po120 = ~w2597;// level 27
assign po121 = ~w2600;// level 27
assign po122 = ~w2603;// level 27
assign po123 = ~w2606;// level 27
assign po124 = ~w2609;// level 27
assign po125 = ~w2612;// level 27
assign po126 = w2655;// level 27
assign po127 = ~w2678;// level 27
assign po128 = ~w2681;// level 27
assign po129 = ~w2684;// level 27
assign po130 = ~w2687;// level 27
assign po131 = ~w2690;// level 27
assign po132 = ~w2693;// level 27
assign po133 = ~w2696;// level 27
assign po134 = ~w2699;// level 27
assign po135 = ~w2702;// level 27
assign po136 = w2705;// level 27
assign po137 = w2708;// level 27
assign po138 = w2711;// level 27
assign po139 = w2714;// level 27
assign po140 = w2717;// level 27
assign po141 = w2720;// level 27
assign po142 = w2740;// level 15
assign po143 = w2746;// level 14
assign po144 = w2753;// level 15
assign po145 = w2777;// level 27
assign po146 = w2801;// level 27
assign po147 = ~w2936;// level 27
assign po148 = w2939;// level 27
assign po149 = w2942;// level 27
assign po150 = w2945;// level 27
assign po151 = w2948;// level 27
assign po152 = w2951;// level 27
assign po153 = w2954;// level 27
assign po154 = w2957;// level 27
assign po155 = w2960;// level 27
assign po156 = w2963;// level 27
assign po157 = w2966;// level 27
assign po158 = w2969;// level 27
assign po159 = w2972;// level 27
assign po160 = w2975;// level 27
assign po161 = w2978;// level 27
assign po162 = w3099;// level 25
assign po163 = w3123;// level 25
assign po164 = w3126;// level 25
assign po165 = w3129;// level 25
assign po166 = w3132;// level 25
assign po167 = w3135;// level 25
assign po168 = w3138;// level 25
assign po169 = w3141;// level 25
assign po170 = w3144;// level 25
assign po171 = ~w3166;// level 16
assign po172 = w3195;// level 24
assign po173 = ~w3211;// level 20
assign po174 = w3233;// level 16
assign po175 = ~w3248;// level 18
assign po176 = ~w3264;// level 21
assign po177 = ~w3302;// level 20
assign po178 = ~w3320;// level 19
assign po179 = ~w3330;// level 19
assign po180 = ~w3353;// level 25
assign po181 = ~w3364;// level 19
assign po182 = ~w3381;// level 24
assign po183 = ~w3399;// level 18
assign po184 = ~w3417;// level 20
assign po185 = ~w3435;// level 19
assign po186 = ~w3453;// level 18
assign po187 = ~w3471;// level 18
assign po188 = ~w3489;// level 18
assign po189 = ~w3504;// level 23
assign po190 = ~w3515;// level 18
assign po191 = ~w3533;// level 23
assign po192 = w3560;// level 27
assign po193 = w3563;// level 27
assign po194 = w3566;// level 27
assign po195 = w3569;// level 27
assign po196 = w3572;// level 27
assign po197 = w3575;// level 27
assign po198 = w3578;// level 27
assign po199 = w3581;// level 24
assign po200 = w3584;// level 24
assign po201 = w3587;// level 24
assign po202 = w3590;// level 24
assign po203 = w3593;// level 24
assign po204 = w3596;// level 24
assign po205 = w3599;// level 24
assign po206 = ~w3610;// level 14
assign po207 = ~w3621;// level 15
assign po208 = ~w3631;// level 15
assign po209 = ~w3642;// level 18
assign po210 = w3665;// level 23
assign po211 = w3668;// level 23
assign po212 = w3671;// level 23
assign po213 = w3674;// level 23
assign po214 = w3677;// level 23
assign po215 = w3680;// level 23
assign po216 = w3683;// level 23
assign po217 = ~w3702;// level 19
assign po218 = ~w3722;// level 21
assign po219 = ~w3738;// level 18
assign po220 = w3741;// level 27
assign po221 = w3744;// level 23
assign po222 = w3766;// level 28
assign po223 = ~w3792;// level 20
assign po224 = ~w3832;// level 30
assign po225 = ~w3866;// level 21
assign po226 = ~w3898;// level 24
assign po227 = ~w3915;// level 28
assign po228 = ~w3940;// level 30
assign po229 = w3967;// level 20
assign po230 = ~w3986;// level 27
assign po231 = ~w4003;// level 28
assign po232 = ~w4020;// level 26
assign po233 = ~w4050;// level 22
assign po234 = ~w4063;// level 22
assign po235 = w4072;// level 20
assign po236 = ~w4087;// level 25
assign po237 = w4112;// level 21
assign po238 = w4117;// level 21
assign po239 = ~w4122;// level 21
assign po240 = w4125;// level 22
assign po241 = w4129;// level 22
assign po242 = ~w4251;// level 24
assign po243 = ~w4266;// level 23
assign po244 = w4372;// level 26
assign po245 = w4395;// level 23
assign po246 = w4400;// level 21
assign po247 = ~w4415;// level 23
assign po248 = w4449;// level 26
assign po249 = w4485;// level 27
assign po250 = w4518;// level 29
assign po251 = w4540;// level 17
assign po252 = w4562;// level 17
assign po253 = ~w4582;// level 19
assign po254 = w4605;// level 19
assign po255 = w4630;// level 21
assign po256 = w4652;// level 21
assign po257 = w4675;// level 23
assign po258 = w4679;// level 21
assign po259 = w4683;// level 21
assign po260 = ~w4698;// level 23
assign po261 = ~w4713;// level 23
assign po262 = ~w4728;// level 24
assign po263 = w4760;// level 26
assign po264 = w4786;// level 30
assign po265 = w4808;// level 17
assign po266 = ~w4823;// level 23
assign po267 = ~w4832;// level 25
assign po268 = ~w4847;// level 24
assign po269 = ~w4856;// level 27
assign po270 = ~w4871;// level 23
assign po271 = ~w4880;// level 27
assign po272 = ~w4889;// level 27
assign po273 = w4895;// level 15
assign po274 = ~w4904;// level 25
assign po275 = w4909;// level 14
assign po276 = ~w4941;// level 14
assign po277 = ~w4950;// level 25
assign po278 = ~w4969;// level 22
assign po279 = ~w4973;// level 15
assign po280 = ~w4976;// level 20
assign po281 = ~w4979;// level 20
assign po282 = w4980;// level 1
assign po283 = ~w4989;// level 24
assign po284 = ~w4993;// level 15
assign po285 = ~w4997;// level 14
assign po286 = ~w5060;// level 18
assign po287 = ~w5068;// level 14
assign po288 = ~w5075;// level 14
assign po289 = ~w5084;// level 23
assign po290 = ~w5087;// level 20
assign po291 = ~w5102;// level 22
assign po292 = w5103;// level 13
assign po293 = ~w5106;// level 20
assign po294 = ~w5109;// level 20
assign po295 = ~w5112;// level 20
assign po296 = ~w5116;// level 14
assign po297 = w5119;// level 12
assign po298 = ~w5122;// level 20
assign po299 = ~w5125;// level 20
assign po300 = ~w5128;// level 20
assign po301 = ~w5155;// level 18
assign po302 = ~w5180;// level 15
assign po303 = ~w5183;// level 20
assign po304 = ~w5198;// level 22
assign po305 = ~w5201;// level 19
assign po306 = ~w5204;// level 19
assign po307 = ~w5207;// level 19
assign po308 = ~w5210;// level 20
assign po309 = ~w5334;// level 23
assign po310 = ~w5349;// level 21
assign po311 = ~w5352;// level 19
assign po312 = ~w5355;// level 19
assign po313 = ~w5364;// level 18
assign po314 = w5392;// level 22
assign po315 = w5413;// level 22
assign po316 = w5434;// level 22
assign po317 = w5455;// level 22
assign po318 = w5476;// level 22
assign po319 = w5497;// level 22
assign po320 = w5518;// level 22
assign po321 = ~w5527;// level 17
assign po322 = w5533;// level 14
assign po323 = ~w5539;// level 18
assign po324 = ~w5589;// level 17
assign po325 = ~w5597;// level 20
assign po326 = ~w5600;// level 17
assign po327 = ~w5609;// level 15
assign po328 = w5613;// level 17
assign po329 = w5616;// level 16
assign po330 = w5623;// level 16
assign po331 = w5641;// level 14
assign po332 = w5651;// level 13
assign po333 = w5661;// level 11
assign po334 = w5671;// level 10
assign po335 = w5681;// level 12
assign po336 = w5701;// level 9
assign po337 = w5711;// level 9
assign po338 = ~w5712;// level 16
assign po339 = w5721;// level 9
assign po340 = w5731;// level 10
assign po341 = w5743;// level 9
assign po342 = w5755;// level 9
assign po343 = w5767;// level 9
assign po344 = w5779;// level 9
assign po345 = w5791;// level 9
assign po346 = w5797;// level 10
assign po347 = w5809;// level 9
assign po348 = w5821;// level 9
assign po349 = w5828;// level 9
assign po350 = w5832;// level 8
assign po351 = ~w5587;// level 13
assign po352 = w5871;// level 13
assign po353 = ~w5890;// level 13
assign po354 = ~w5893;// level 14
assign po355 = w5932;// level 15
assign po356 = ~w5940;// level 18
assign po357 = w5944;// level 15
assign po358 = w5949;// level 9
assign po359 = w5953;// level 9
assign po360 = ~w5958;// level 9
assign po361 = ~w5962;// level 9
assign po362 = ~w5966;// level 9
assign po363 = ~w5970;// level 9
assign po364 = ~w5974;// level 9
assign po365 = ~w5978;// level 9
assign po366 = ~w5982;// level 9
assign po367 = ~w5986;// level 9
assign po368 = ~w5990;// level 9
assign po369 = ~w5994;// level 9
assign po370 = ~w5998;// level 9
assign po371 = ~w6002;// level 9
assign po372 = ~w6006;// level 9
assign po373 = ~w6010;// level 9
assign po374 = ~w6014;// level 9
assign po375 = ~w6018;// level 9
assign po376 = w6027;// level 8
assign po377 = w6032;// level 9
assign po378 = w6035;// level 8
assign po379 = ~w6037;// level 6
assign po380 = w6043;// level 8
assign po381 = w6050;// level 8
assign po382 = w6054;// level 8
assign po383 = w6058;// level 8
assign po384 = w6062;// level 8
assign po385 = w6066;// level 8
assign po386 = w6070;// level 8
assign po387 = w6074;// level 8
assign po388 = w6078;// level 8
assign po389 = ~w6081;// level 6
assign po390 = w6087;// level 5
assign po391 = ~w6093;// level 9
assign po392 = w6096;// level 5
assign po393 = w6099;// level 5
assign po394 = w6102;// level 5
assign po395 = w6105;// level 5
assign po396 = w6108;// level 5
assign po397 = w6111;// level 5
assign po398 = w6114;// level 5
assign po399 = w6117;// level 5
assign po400 = w6121;// level 3
assign po401 = w6122;// level 1
assign po402 = w6123;// level 1
assign po403 = w6124;// level 1
endmodule
