// Benchmark "hamming" written by ABC on Wed Apr 29 17:31:55 2015

module hamming ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    po0, po1, po2, po3, po4, po5, po6  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199;
  output po0, po1, po2, po3, po4, po5, po6;
  wire n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
    n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
    n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
    n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
    n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
    n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
    n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
    n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
    n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
    n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
    n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
    n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
    n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
    n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
    n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
    n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
    n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
    n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
    n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
    n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
    n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
    n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
    n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
    n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
    n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
    n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
    n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
    n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
    n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
    n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
    n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
    n3563, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818;
  assign n208 = pi096 & ~pi196;
  assign n209 = ~pi096 & pi196;
  assign n210 = ~n208 & ~n209;
  assign n211 = pi063 & ~pi163;
  assign n212 = ~pi063 & pi163;
  assign n213 = ~n211 & ~n212;
  assign n214 = pi064 & ~pi164;
  assign n215 = ~pi064 & pi164;
  assign n216 = ~n214 & ~n215;
  assign n217 = ~n213 & n216;
  assign n218 = n213 & ~n216;
  assign n219 = ~n217 & ~n218;
  assign n220 = pi065 & ~pi165;
  assign n221 = ~pi065 & pi165;
  assign n222 = ~n220 & ~n221;
  assign n223 = pi066 & ~pi166;
  assign n224 = ~pi066 & pi166;
  assign n225 = ~n223 & ~n224;
  assign n226 = n222 & n225;
  assign n227 = ~n222 & ~n225;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~n219 & n228;
  assign n230 = n219 & ~n228;
  assign n231 = ~n229 & ~n230;
  assign n232 = pi062 & ~pi162;
  assign n233 = ~pi062 & pi162;
  assign n234 = ~n232 & ~n233;
  assign n235 = pi002 & ~pi102;
  assign n236 = ~pi002 & pi102;
  assign n237 = ~n235 & ~n236;
  assign n238 = pi003 & ~pi103;
  assign n239 = ~pi003 & pi103;
  assign n240 = ~n238 & ~n239;
  assign n241 = n237 & n240;
  assign n242 = ~n237 & ~n240;
  assign n243 = ~n241 & ~n242;
  assign n244 = pi000 & ~pi100;
  assign n245 = ~pi000 & pi100;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi001 & ~pi101;
  assign n248 = ~pi001 & pi101;
  assign n249 = ~n247 & ~n248;
  assign n250 = n246 & n249;
  assign n251 = ~n246 & ~n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = ~n243 & n252;
  assign n254 = n243 & ~n252;
  assign n255 = ~n253 & ~n254;
  assign n256 = pi005 & ~pi105;
  assign n257 = ~pi005 & pi105;
  assign n258 = ~n256 & ~n257;
  assign n259 = pi006 & ~pi106;
  assign n260 = ~pi006 & pi106;
  assign n261 = ~n259 & ~n260;
  assign n262 = n258 & n261;
  assign n263 = ~n258 & ~n261;
  assign n264 = pi007 & ~pi107;
  assign n265 = ~pi007 & pi107;
  assign n266 = ~n264 & ~n265;
  assign n267 = pi004 & ~pi104;
  assign n268 = ~pi004 & pi104;
  assign n269 = ~n267 & ~n268;
  assign n270 = n266 & n269;
  assign n271 = ~n263 & n270;
  assign n272 = ~n262 & n271;
  assign n273 = ~n255 & n272;
  assign n274 = ~n262 & ~n263;
  assign n275 = n266 & ~n269;
  assign n276 = ~n274 & n275;
  assign n277 = ~n255 & n276;
  assign n278 = ~n273 & ~n277;
  assign n279 = n270 & ~n274;
  assign n280 = ~n253 & n279;
  assign n281 = ~n254 & n280;
  assign n282 = ~n263 & n275;
  assign n283 = ~n262 & n282;
  assign n284 = ~n253 & n283;
  assign n285 = ~n254 & n284;
  assign n286 = ~n281 & ~n285;
  assign n287 = n278 & n286;
  assign n288 = ~n266 & n269;
  assign n289 = ~n274 & n288;
  assign n290 = ~n255 & n289;
  assign n291 = ~n266 & ~n269;
  assign n292 = ~n263 & n291;
  assign n293 = ~n262 & n292;
  assign n294 = ~n255 & n293;
  assign n295 = ~n290 & ~n294;
  assign n296 = ~n263 & n288;
  assign n297 = ~n262 & n296;
  assign n298 = ~n253 & n297;
  assign n299 = ~n254 & n298;
  assign n300 = ~n274 & n291;
  assign n301 = ~n253 & n300;
  assign n302 = ~n254 & n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = n295 & n303;
  assign n305 = pi014 & ~pi114;
  assign n306 = ~pi014 & pi114;
  assign n307 = ~n305 & ~n306;
  assign n308 = pi013 & ~pi113;
  assign n309 = ~pi013 & pi113;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~n307 & ~n310;
  assign n312 = n307 & n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = pi011 & ~pi111;
  assign n315 = ~pi011 & pi111;
  assign n316 = ~n314 & ~n315;
  assign n317 = pi012 & ~pi112;
  assign n318 = ~pi012 & pi112;
  assign n319 = ~n317 & ~n318;
  assign n320 = n316 & n319;
  assign n321 = ~n316 & ~n319;
  assign n322 = ~n320 & ~n321;
  assign n323 = n313 & ~n322;
  assign n324 = pi010 & ~pi110;
  assign n325 = ~pi010 & pi110;
  assign n326 = ~n324 & ~n325;
  assign n327 = pi009 & ~pi109;
  assign n328 = ~pi009 & pi109;
  assign n329 = ~n327 & ~n328;
  assign n330 = pi008 & ~pi108;
  assign n331 = ~pi008 & pi108;
  assign n332 = ~n330 & ~n331;
  assign n333 = ~n329 & n332;
  assign n334 = n329 & ~n332;
  assign n335 = ~n333 & ~n334;
  assign n336 = ~n326 & ~n335;
  assign n337 = ~n313 & n322;
  assign n338 = ~n336 & ~n337;
  assign n339 = ~n323 & n338;
  assign n340 = pi015 & ~pi115;
  assign n341 = ~pi015 & pi115;
  assign n342 = ~n340 & ~n341;
  assign n343 = n326 & ~n333;
  assign n344 = ~n334 & n343;
  assign n345 = n342 & ~n344;
  assign n346 = n339 & n345;
  assign n347 = n304 & n346;
  assign n348 = n287 & n347;
  assign n349 = n287 & n304;
  assign n350 = ~n323 & ~n337;
  assign n351 = ~n336 & n345;
  assign n352 = ~n350 & n351;
  assign n353 = ~n349 & n352;
  assign n354 = ~n336 & ~n344;
  assign n355 = ~n337 & n342;
  assign n356 = ~n323 & n355;
  assign n357 = ~n354 & n356;
  assign n358 = ~n349 & n357;
  assign n359 = ~n353 & ~n358;
  assign n360 = ~n348 & n359;
  assign n361 = ~n342 & ~n354;
  assign n362 = ~n350 & n361;
  assign n363 = ~n349 & n362;
  assign n364 = pi031 & ~pi131;
  assign n365 = ~pi031 & pi131;
  assign n366 = ~n364 & ~n365;
  assign n367 = pi032 & ~pi132;
  assign n368 = ~pi032 & pi132;
  assign n369 = ~n367 & ~n368;
  assign n370 = ~n366 & ~n369;
  assign n371 = n366 & n369;
  assign n372 = pi033 & ~pi133;
  assign n373 = ~pi033 & pi133;
  assign n374 = ~n372 & ~n373;
  assign n375 = ~n371 & n374;
  assign n376 = ~n370 & n375;
  assign n377 = ~n370 & ~n371;
  assign n378 = ~n374 & ~n377;
  assign n379 = ~n376 & ~n378;
  assign n380 = pi035 & ~pi135;
  assign n381 = ~pi035 & pi135;
  assign n382 = ~n380 & ~n381;
  assign n383 = pi036 & ~pi136;
  assign n384 = ~pi036 & pi136;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n382 & ~n385;
  assign n387 = n382 & n385;
  assign n388 = pi034 & ~pi134;
  assign n389 = ~pi034 & pi134;
  assign n390 = ~n388 & ~n389;
  assign n391 = ~n387 & n390;
  assign n392 = ~n386 & n391;
  assign n393 = ~n386 & ~n387;
  assign n394 = ~n390 & ~n393;
  assign n395 = ~n392 & ~n394;
  assign n396 = n379 & n395;
  assign n397 = ~n379 & ~n395;
  assign n398 = ~n396 & ~n397;
  assign n399 = pi041 & ~pi141;
  assign n400 = ~pi041 & pi141;
  assign n401 = ~n399 & ~n400;
  assign n402 = pi016 & ~pi116;
  assign n403 = ~pi016 & pi116;
  assign n404 = ~n402 & ~n403;
  assign n405 = ~n401 & n404;
  assign n406 = n401 & ~n404;
  assign n407 = ~n405 & ~n406;
  assign n408 = ~n398 & ~n407;
  assign n409 = ~n396 & n407;
  assign n410 = ~n397 & n409;
  assign n411 = ~n408 & ~n410;
  assign n412 = ~n363 & ~n411;
  assign n413 = ~n342 & ~n344;
  assign n414 = ~n336 & n413;
  assign n415 = ~n350 & n414;
  assign n416 = n304 & n415;
  assign n417 = n287 & n416;
  assign n418 = ~n337 & ~n342;
  assign n419 = ~n323 & n418;
  assign n420 = ~n354 & n419;
  assign n421 = n304 & n420;
  assign n422 = n287 & n421;
  assign n423 = ~n417 & ~n422;
  assign n424 = n339 & n413;
  assign n425 = ~n349 & n424;
  assign n426 = n342 & ~n354;
  assign n427 = ~n350 & n426;
  assign n428 = n304 & n427;
  assign n429 = n287 & n428;
  assign n430 = ~n425 & ~n429;
  assign n431 = n423 & n430;
  assign n432 = n412 & n431;
  assign n433 = n360 & n432;
  assign n434 = ~n353 & ~n429;
  assign n435 = ~n348 & ~n358;
  assign n436 = n434 & n435;
  assign n437 = ~n363 & ~n417;
  assign n438 = ~n422 & ~n425;
  assign n439 = n437 & n438;
  assign n440 = n436 & n439;
  assign n441 = n411 & ~n440;
  assign n442 = ~n433 & ~n441;
  assign n443 = pi021 & ~pi121;
  assign n444 = ~pi021 & pi121;
  assign n445 = ~n443 & ~n444;
  assign n446 = pi019 & ~pi119;
  assign n447 = ~pi019 & pi119;
  assign n448 = ~n446 & ~n447;
  assign n449 = pi020 & ~pi120;
  assign n450 = ~pi020 & pi120;
  assign n451 = ~n449 & ~n450;
  assign n452 = ~n448 & ~n451;
  assign n453 = n448 & n451;
  assign n454 = ~n452 & ~n453;
  assign n455 = pi017 & ~pi117;
  assign n456 = ~pi017 & pi117;
  assign n457 = ~n455 & ~n456;
  assign n458 = pi018 & ~pi118;
  assign n459 = ~pi018 & pi118;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n457 & ~n460;
  assign n462 = n457 & n460;
  assign n463 = ~n461 & ~n462;
  assign n464 = ~n454 & n463;
  assign n465 = n454 & ~n463;
  assign n466 = ~n464 & ~n465;
  assign n467 = ~n445 & ~n466;
  assign n468 = n445 & ~n464;
  assign n469 = ~n465 & n468;
  assign n470 = ~n467 & ~n469;
  assign n471 = pi023 & ~pi123;
  assign n472 = ~pi023 & pi123;
  assign n473 = ~n471 & ~n472;
  assign n474 = pi024 & ~pi124;
  assign n475 = ~pi024 & pi124;
  assign n476 = ~n474 & ~n475;
  assign n477 = ~n473 & ~n476;
  assign n478 = n473 & n476;
  assign n479 = pi022 & ~pi122;
  assign n480 = ~pi022 & pi122;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n478 & n481;
  assign n483 = ~n477 & n482;
  assign n484 = ~n477 & ~n478;
  assign n485 = ~n481 & ~n484;
  assign n486 = ~n483 & ~n485;
  assign n487 = pi025 & ~pi125;
  assign n488 = ~pi025 & pi125;
  assign n489 = ~n487 & ~n488;
  assign n490 = pi026 & ~pi126;
  assign n491 = ~pi026 & pi126;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n489 & ~n492;
  assign n494 = n489 & n492;
  assign n495 = pi027 & ~pi127;
  assign n496 = ~pi027 & pi127;
  assign n497 = ~n495 & ~n496;
  assign n498 = ~n494 & n497;
  assign n499 = ~n493 & n498;
  assign n500 = ~n493 & ~n494;
  assign n501 = ~n497 & ~n500;
  assign n502 = ~n499 & ~n501;
  assign n503 = ~n486 & ~n502;
  assign n504 = n486 & n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = n470 & n505;
  assign n507 = ~n470 & ~n505;
  assign n508 = pi028 & ~pi128;
  assign n509 = ~pi028 & pi128;
  assign n510 = ~n508 & ~n509;
  assign n511 = pi030 & ~pi130;
  assign n512 = ~pi030 & pi130;
  assign n513 = ~n511 & ~n512;
  assign n514 = pi029 & ~pi129;
  assign n515 = ~pi029 & pi129;
  assign n516 = ~n514 & ~n515;
  assign n517 = ~n513 & n516;
  assign n518 = n513 & ~n516;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~n510 & ~n519;
  assign n521 = n510 & ~n517;
  assign n522 = ~n518 & n521;
  assign n523 = ~n520 & ~n522;
  assign n524 = ~n507 & ~n523;
  assign n525 = ~n506 & n524;
  assign n526 = ~n506 & ~n507;
  assign n527 = n523 & ~n526;
  assign n528 = ~n525 & ~n527;
  assign n529 = pi039 & ~pi139;
  assign n530 = ~pi039 & pi139;
  assign n531 = ~n529 & ~n530;
  assign n532 = pi040 & ~pi140;
  assign n533 = ~pi040 & pi140;
  assign n534 = ~n532 & ~n533;
  assign n535 = ~n531 & ~n534;
  assign n536 = n531 & n534;
  assign n537 = ~n535 & ~n536;
  assign n538 = pi037 & ~pi137;
  assign n539 = ~pi037 & pi137;
  assign n540 = ~n538 & ~n539;
  assign n541 = pi038 & ~pi138;
  assign n542 = ~pi038 & pi138;
  assign n543 = ~n541 & ~n542;
  assign n544 = n540 & n543;
  assign n545 = ~n540 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n537 & n546;
  assign n548 = ~n528 & n547;
  assign n549 = pi058 & ~pi158;
  assign n550 = ~pi058 & pi158;
  assign n551 = ~n549 & ~n550;
  assign n552 = pi049 & ~pi149;
  assign n553 = ~pi049 & pi149;
  assign n554 = ~n552 & ~n553;
  assign n555 = pi050 & ~pi150;
  assign n556 = ~pi050 & pi150;
  assign n557 = ~n555 & ~n556;
  assign n558 = n554 & n557;
  assign n559 = ~n554 & ~n557;
  assign n560 = pi051 & ~pi151;
  assign n561 = ~pi051 & pi151;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~n559 & n562;
  assign n564 = ~n558 & n563;
  assign n565 = ~n558 & ~n559;
  assign n566 = ~n562 & ~n565;
  assign n567 = ~n564 & ~n566;
  assign n568 = pi042 & ~pi142;
  assign n569 = ~pi042 & pi142;
  assign n570 = ~n568 & ~n569;
  assign n571 = pi045 & ~pi145;
  assign n572 = ~pi045 & pi145;
  assign n573 = ~n571 & ~n572;
  assign n574 = ~n570 & n573;
  assign n575 = n570 & ~n573;
  assign n576 = ~n574 & ~n575;
  assign n577 = pi043 & ~pi143;
  assign n578 = ~pi043 & pi143;
  assign n579 = ~n577 & ~n578;
  assign n580 = pi044 & ~pi144;
  assign n581 = ~pi044 & pi144;
  assign n582 = ~n580 & ~n581;
  assign n583 = n579 & n582;
  assign n584 = ~n579 & ~n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~n576 & n585;
  assign n587 = n576 & ~n585;
  assign n588 = ~n586 & ~n587;
  assign n589 = pi047 & ~pi147;
  assign n590 = ~pi047 & pi147;
  assign n591 = ~n589 & ~n590;
  assign n592 = pi048 & ~pi148;
  assign n593 = ~pi048 & pi148;
  assign n594 = ~n592 & ~n593;
  assign n595 = n591 & n594;
  assign n596 = ~n591 & ~n594;
  assign n597 = pi046 & ~pi146;
  assign n598 = ~pi046 & pi146;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~n596 & n599;
  assign n601 = ~n595 & n600;
  assign n602 = ~n595 & ~n596;
  assign n603 = ~n599 & ~n602;
  assign n604 = ~n601 & ~n603;
  assign n605 = ~n588 & n604;
  assign n606 = n588 & ~n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n567 & ~n607;
  assign n609 = n567 & ~n605;
  assign n610 = ~n606 & n609;
  assign n611 = ~n608 & ~n610;
  assign n612 = pi052 & ~pi152;
  assign n613 = ~pi052 & pi152;
  assign n614 = ~n612 & ~n613;
  assign n615 = pi055 & ~pi155;
  assign n616 = ~pi055 & pi155;
  assign n617 = ~n615 & ~n616;
  assign n618 = pi056 & ~pi156;
  assign n619 = ~pi056 & pi156;
  assign n620 = ~n618 & ~n619;
  assign n621 = ~n617 & ~n620;
  assign n622 = n617 & n620;
  assign n623 = pi057 & ~pi157;
  assign n624 = ~pi057 & pi157;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~n622 & n625;
  assign n627 = ~n621 & n626;
  assign n628 = ~n621 & ~n622;
  assign n629 = ~n625 & ~n628;
  assign n630 = ~n627 & ~n629;
  assign n631 = pi053 & ~pi153;
  assign n632 = ~pi053 & pi153;
  assign n633 = ~n631 & ~n632;
  assign n634 = pi054 & ~pi154;
  assign n635 = ~pi054 & pi154;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n633 & ~n636;
  assign n638 = n633 & n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = ~n630 & n639;
  assign n641 = ~n627 & ~n639;
  assign n642 = ~n629 & n641;
  assign n643 = ~n640 & ~n642;
  assign n644 = ~n614 & ~n643;
  assign n645 = n614 & ~n640;
  assign n646 = ~n642 & n645;
  assign n647 = ~n644 & ~n646;
  assign n648 = ~n611 & n647;
  assign n649 = n611 & ~n647;
  assign n650 = ~n648 & ~n649;
  assign n651 = n551 & ~n650;
  assign n652 = ~n548 & n651;
  assign n653 = n537 & ~n546;
  assign n654 = ~n528 & n653;
  assign n655 = ~n537 & ~n546;
  assign n656 = ~n525 & n655;
  assign n657 = ~n527 & n656;
  assign n658 = n537 & n546;
  assign n659 = ~n525 & n658;
  assign n660 = ~n527 & n659;
  assign n661 = ~n657 & ~n660;
  assign n662 = ~n654 & n661;
  assign n663 = n652 & n662;
  assign n664 = n442 & n663;
  assign n665 = ~n551 & ~n648;
  assign n666 = ~n649 & n665;
  assign n667 = ~n548 & n666;
  assign n668 = n662 & n667;
  assign n669 = n442 & n668;
  assign n670 = ~n664 & ~n669;
  assign n671 = ~n551 & ~n650;
  assign n672 = ~n548 & n671;
  assign n673 = n662 & n672;
  assign n674 = ~n442 & n673;
  assign n675 = n551 & ~n648;
  assign n676 = ~n649 & n675;
  assign n677 = ~n548 & n676;
  assign n678 = n662 & n677;
  assign n679 = ~n442 & n678;
  assign n680 = ~n674 & ~n679;
  assign n681 = n670 & n680;
  assign n682 = ~n433 & n671;
  assign n683 = ~n548 & ~n657;
  assign n684 = ~n654 & ~n660;
  assign n685 = n683 & n684;
  assign n686 = ~n441 & ~n685;
  assign n687 = n682 & n686;
  assign n688 = ~n433 & n676;
  assign n689 = n686 & n688;
  assign n690 = ~n687 & ~n689;
  assign n691 = n651 & ~n685;
  assign n692 = ~n442 & n691;
  assign n693 = n666 & ~n685;
  assign n694 = ~n442 & n693;
  assign n695 = ~n692 & ~n694;
  assign n696 = n690 & n695;
  assign n697 = n681 & n696;
  assign n698 = pi059 & ~pi159;
  assign n699 = ~pi059 & pi159;
  assign n700 = ~n698 & ~n699;
  assign n701 = pi060 & ~pi160;
  assign n702 = ~pi060 & pi160;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~n700 & ~n703;
  assign n705 = n700 & n703;
  assign n706 = pi061 & ~pi161;
  assign n707 = ~pi061 & pi161;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n705 & n708;
  assign n710 = ~n704 & n709;
  assign n711 = ~n704 & ~n705;
  assign n712 = ~n708 & ~n711;
  assign n713 = ~n710 & ~n712;
  assign n714 = ~n697 & ~n713;
  assign n715 = ~n669 & ~n674;
  assign n716 = ~n679 & n715;
  assign n717 = ~n687 & n713;
  assign n718 = ~n689 & ~n692;
  assign n719 = ~n664 & ~n694;
  assign n720 = n718 & n719;
  assign n721 = n717 & n720;
  assign n722 = n716 & n721;
  assign n723 = ~n714 & ~n722;
  assign n724 = ~n234 & ~n723;
  assign n725 = n234 & ~n714;
  assign n726 = ~n722 & n725;
  assign n727 = ~n724 & ~n726;
  assign n728 = n231 & ~n727;
  assign n729 = ~n231 & ~n724;
  assign n730 = ~n726 & n729;
  assign n731 = pi067 & ~pi167;
  assign n732 = ~pi067 & pi167;
  assign n733 = ~n731 & ~n732;
  assign n734 = pi068 & ~pi168;
  assign n735 = ~pi068 & pi168;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~n733 & ~n736;
  assign n738 = n733 & n736;
  assign n739 = pi070 & ~pi170;
  assign n740 = ~pi070 & pi170;
  assign n741 = ~n739 & ~n740;
  assign n742 = pi069 & ~pi169;
  assign n743 = ~pi069 & pi169;
  assign n744 = ~n742 & ~n743;
  assign n745 = n741 & n744;
  assign n746 = ~n738 & n745;
  assign n747 = ~n737 & n746;
  assign n748 = ~n730 & n747;
  assign n749 = ~n728 & n748;
  assign n750 = ~n728 & ~n730;
  assign n751 = n741 & ~n744;
  assign n752 = ~n738 & n751;
  assign n753 = ~n737 & n752;
  assign n754 = ~n750 & n753;
  assign n755 = ~n737 & ~n738;
  assign n756 = n751 & ~n755;
  assign n757 = ~n730 & n756;
  assign n758 = ~n728 & n757;
  assign n759 = ~n754 & ~n758;
  assign n760 = ~n749 & n759;
  assign n761 = ~n741 & n744;
  assign n762 = ~n738 & n761;
  assign n763 = ~n737 & n762;
  assign n764 = ~n750 & n763;
  assign n765 = ~n755 & n761;
  assign n766 = ~n730 & n765;
  assign n767 = ~n728 & n766;
  assign n768 = ~n764 & ~n767;
  assign n769 = ~n741 & ~n744;
  assign n770 = ~n738 & n769;
  assign n771 = ~n737 & n770;
  assign n772 = ~n730 & n771;
  assign n773 = ~n728 & n772;
  assign n774 = n745 & ~n755;
  assign n775 = ~n750 & n774;
  assign n776 = ~n773 & ~n775;
  assign n777 = n768 & n776;
  assign n778 = ~n755 & n769;
  assign n779 = ~n750 & n778;
  assign n780 = pi071 & ~pi171;
  assign n781 = ~pi071 & pi171;
  assign n782 = ~n780 & ~n781;
  assign n783 = pi072 & ~pi172;
  assign n784 = ~pi072 & pi172;
  assign n785 = ~n783 & ~n784;
  assign n786 = n782 & n785;
  assign n787 = ~n782 & ~n785;
  assign n788 = pi073 & ~pi173;
  assign n789 = ~pi073 & pi173;
  assign n790 = ~n788 & ~n789;
  assign n791 = pi074 & ~pi174;
  assign n792 = ~pi074 & pi174;
  assign n793 = ~n791 & ~n792;
  assign n794 = ~n790 & ~n793;
  assign n795 = ~n787 & n794;
  assign n796 = ~n786 & n795;
  assign n797 = ~n779 & n796;
  assign n798 = n777 & n797;
  assign n799 = n760 & n798;
  assign n800 = n790 & n793;
  assign n801 = ~n787 & n800;
  assign n802 = ~n786 & n801;
  assign n803 = ~n779 & n802;
  assign n804 = n777 & n803;
  assign n805 = n760 & n804;
  assign n806 = ~n754 & ~n775;
  assign n807 = ~n749 & ~n758;
  assign n808 = n806 & n807;
  assign n809 = ~n764 & ~n779;
  assign n810 = ~n767 & ~n773;
  assign n811 = n809 & n810;
  assign n812 = n808 & n811;
  assign n813 = ~n786 & ~n787;
  assign n814 = n794 & ~n813;
  assign n815 = ~n812 & n814;
  assign n816 = ~n805 & ~n815;
  assign n817 = ~n799 & n816;
  assign n818 = ~n794 & ~n800;
  assign n819 = n813 & n818;
  assign n820 = ~n812 & n819;
  assign n821 = n800 & ~n813;
  assign n822 = ~n812 & n821;
  assign n823 = ~n820 & ~n822;
  assign n824 = ~n813 & n818;
  assign n825 = ~n779 & n824;
  assign n826 = n777 & n825;
  assign n827 = n760 & n826;
  assign n828 = pi075 & ~pi175;
  assign n829 = ~pi075 & pi175;
  assign n830 = ~n828 & ~n829;
  assign n831 = pi076 & ~pi176;
  assign n832 = ~pi076 & pi176;
  assign n833 = ~n831 & ~n832;
  assign n834 = n830 & ~n833;
  assign n835 = ~n827 & n834;
  assign n836 = n823 & n835;
  assign n837 = n817 & n836;
  assign n838 = ~n830 & n833;
  assign n839 = ~n827 & n838;
  assign n840 = n823 & n839;
  assign n841 = n817 & n840;
  assign n842 = pi077 & ~pi177;
  assign n843 = ~pi077 & pi177;
  assign n844 = ~n842 & ~n843;
  assign n845 = pi078 & ~pi178;
  assign n846 = ~pi078 & pi178;
  assign n847 = ~n845 & ~n846;
  assign n848 = n844 & n847;
  assign n849 = ~n844 & ~n847;
  assign n850 = ~n848 & ~n849;
  assign n851 = pi079 & ~pi179;
  assign n852 = ~pi079 & pi179;
  assign n853 = ~n851 & ~n852;
  assign n854 = pi080 & ~pi180;
  assign n855 = ~pi080 & pi180;
  assign n856 = ~n854 & ~n855;
  assign n857 = ~n853 & ~n856;
  assign n858 = n853 & n856;
  assign n859 = ~n857 & ~n858;
  assign n860 = n850 & ~n859;
  assign n861 = ~n850 & n859;
  assign n862 = pi081 & ~pi181;
  assign n863 = ~pi081 & pi181;
  assign n864 = ~n862 & ~n863;
  assign n865 = pi082 & ~pi182;
  assign n866 = ~pi082 & pi182;
  assign n867 = ~n865 & ~n866;
  assign n868 = ~n864 & n867;
  assign n869 = n864 & ~n867;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n861 & n870;
  assign n872 = ~n860 & n871;
  assign n873 = ~n860 & ~n861;
  assign n874 = ~n870 & ~n873;
  assign n875 = ~n872 & ~n874;
  assign n876 = ~n841 & ~n875;
  assign n877 = ~n837 & n876;
  assign n878 = ~n820 & ~n827;
  assign n879 = ~n805 & ~n822;
  assign n880 = ~n799 & ~n815;
  assign n881 = n879 & n880;
  assign n882 = n878 & n881;
  assign n883 = n830 & n833;
  assign n884 = ~n882 & n883;
  assign n885 = ~n830 & ~n833;
  assign n886 = ~n882 & n885;
  assign n887 = ~n884 & ~n886;
  assign n888 = n877 & n887;
  assign n889 = ~n837 & ~n841;
  assign n890 = ~n884 & n889;
  assign n891 = ~n886 & n890;
  assign n892 = n875 & ~n891;
  assign n893 = ~n888 & ~n892;
  assign n894 = pi086 & ~pi186;
  assign n895 = ~pi086 & pi186;
  assign n896 = ~n894 & ~n895;
  assign n897 = pi085 & ~pi185;
  assign n898 = ~pi085 & pi185;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~n896 & ~n899;
  assign n901 = n896 & n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = pi083 & ~pi183;
  assign n904 = ~pi083 & pi183;
  assign n905 = ~n903 & ~n904;
  assign n906 = pi084 & ~pi184;
  assign n907 = ~pi084 & pi184;
  assign n908 = ~n906 & ~n907;
  assign n909 = ~n905 & ~n908;
  assign n910 = ~n902 & n909;
  assign n911 = ~n893 & n910;
  assign n912 = ~n905 & n908;
  assign n913 = ~n900 & n912;
  assign n914 = ~n901 & n913;
  assign n915 = ~n893 & n914;
  assign n916 = n905 & ~n908;
  assign n917 = ~n900 & n916;
  assign n918 = ~n901 & n917;
  assign n919 = ~n893 & n918;
  assign n920 = ~n915 & ~n919;
  assign n921 = ~n911 & n920;
  assign n922 = ~n900 & n909;
  assign n923 = ~n901 & n922;
  assign n924 = ~n888 & n923;
  assign n925 = ~n892 & n924;
  assign n926 = ~n902 & n912;
  assign n927 = ~n888 & n926;
  assign n928 = ~n892 & n927;
  assign n929 = ~n902 & n916;
  assign n930 = ~n888 & n929;
  assign n931 = ~n892 & n930;
  assign n932 = ~n928 & ~n931;
  assign n933 = ~n925 & n932;
  assign n934 = n905 & n908;
  assign n935 = ~n902 & n934;
  assign n936 = ~n893 & n935;
  assign n937 = ~n900 & n934;
  assign n938 = ~n901 & n937;
  assign n939 = ~n888 & n938;
  assign n940 = ~n892 & n939;
  assign n941 = pi087 & ~pi187;
  assign n942 = ~pi087 & pi187;
  assign n943 = ~n941 & ~n942;
  assign n944 = pi088 & ~pi188;
  assign n945 = ~pi088 & pi188;
  assign n946 = ~n944 & ~n945;
  assign n947 = n943 & n946;
  assign n948 = ~n943 & ~n946;
  assign n949 = ~n947 & ~n948;
  assign n950 = pi089 & ~pi189;
  assign n951 = ~pi089 & pi189;
  assign n952 = ~n950 & ~n951;
  assign n953 = pi090 & ~pi190;
  assign n954 = ~pi090 & pi190;
  assign n955 = ~n953 & ~n954;
  assign n956 = ~n952 & n955;
  assign n957 = ~n949 & n956;
  assign n958 = ~n940 & n957;
  assign n959 = ~n936 & n958;
  assign n960 = n933 & n959;
  assign n961 = n921 & n960;
  assign n962 = n952 & n955;
  assign n963 = ~n947 & n962;
  assign n964 = ~n948 & n963;
  assign n965 = ~n940 & n964;
  assign n966 = ~n936 & n965;
  assign n967 = n933 & n966;
  assign n968 = n921 & n967;
  assign n969 = ~n961 & ~n968;
  assign n970 = n952 & ~n955;
  assign n971 = ~n949 & n970;
  assign n972 = ~n940 & n971;
  assign n973 = ~n936 & n972;
  assign n974 = n933 & n973;
  assign n975 = n921 & n974;
  assign n976 = ~n952 & ~n955;
  assign n977 = ~n947 & n976;
  assign n978 = ~n948 & n977;
  assign n979 = ~n940 & n978;
  assign n980 = ~n936 & n979;
  assign n981 = n933 & n980;
  assign n982 = n921 & n981;
  assign n983 = ~n975 & ~n982;
  assign n984 = n969 & n983;
  assign n985 = ~n928 & ~n940;
  assign n986 = ~n925 & ~n931;
  assign n987 = n985 & n986;
  assign n988 = ~n915 & ~n936;
  assign n989 = ~n911 & ~n919;
  assign n990 = n988 & n989;
  assign n991 = n987 & n990;
  assign n992 = ~n949 & n962;
  assign n993 = ~n991 & n992;
  assign n994 = ~n947 & n956;
  assign n995 = ~n948 & n994;
  assign n996 = ~n991 & n995;
  assign n997 = ~n993 & ~n996;
  assign n998 = ~n949 & n976;
  assign n999 = ~n991 & n998;
  assign n1000 = ~n947 & n970;
  assign n1001 = ~n948 & n1000;
  assign n1002 = ~n991 & n1001;
  assign n1003 = ~n999 & ~n1002;
  assign n1004 = n997 & n1003;
  assign n1005 = n984 & n1004;
  assign n1006 = pi092 & ~pi192;
  assign n1007 = ~pi092 & pi192;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = pi093 & ~pi193;
  assign n1010 = ~pi093 & pi193;
  assign n1011 = ~n1009 & ~n1010;
  assign n1012 = pi091 & ~pi191;
  assign n1013 = ~pi091 & pi191;
  assign n1014 = ~n1012 & ~n1013;
  assign n1015 = n1011 & n1014;
  assign n1016 = ~n1008 & n1015;
  assign n1017 = ~n1005 & n1016;
  assign n1018 = ~n1011 & ~n1014;
  assign n1019 = ~n1008 & n1018;
  assign n1020 = ~n1005 & n1019;
  assign n1021 = n1008 & n1011;
  assign n1022 = ~n1014 & n1021;
  assign n1023 = ~n1005 & n1022;
  assign n1024 = ~n1020 & ~n1023;
  assign n1025 = ~n1017 & n1024;
  assign n1026 = ~n996 & ~n999;
  assign n1027 = ~n1002 & n1026;
  assign n1028 = ~n968 & ~n975;
  assign n1029 = ~n982 & n1028;
  assign n1030 = n1011 & ~n1014;
  assign n1031 = ~n1008 & n1030;
  assign n1032 = ~n961 & n1031;
  assign n1033 = ~n993 & n1032;
  assign n1034 = n1029 & n1033;
  assign n1035 = n1027 & n1034;
  assign n1036 = ~n1011 & n1014;
  assign n1037 = ~n1008 & n1036;
  assign n1038 = ~n961 & n1037;
  assign n1039 = ~n993 & n1038;
  assign n1040 = n1029 & n1039;
  assign n1041 = n1027 & n1040;
  assign n1042 = n1008 & n1014;
  assign n1043 = n1011 & n1042;
  assign n1044 = ~n961 & n1043;
  assign n1045 = ~n993 & n1044;
  assign n1046 = n1029 & n1045;
  assign n1047 = n1027 & n1046;
  assign n1048 = ~n1041 & ~n1047;
  assign n1049 = ~n1035 & n1048;
  assign n1050 = n1008 & ~n1011;
  assign n1051 = n1014 & n1050;
  assign n1052 = ~n1005 & n1051;
  assign n1053 = pi094 & ~pi194;
  assign n1054 = ~pi094 & pi194;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = ~n1014 & n1050;
  assign n1057 = ~n961 & n1056;
  assign n1058 = ~n993 & n1057;
  assign n1059 = n1029 & n1058;
  assign n1060 = n1027 & n1059;
  assign n1061 = ~n1055 & ~n1060;
  assign n1062 = ~n1052 & n1061;
  assign n1063 = n1049 & n1062;
  assign n1064 = n1025 & n1063;
  assign n1065 = ~n1041 & ~n1060;
  assign n1066 = ~n1035 & ~n1047;
  assign n1067 = n1065 & n1066;
  assign n1068 = ~n1020 & ~n1052;
  assign n1069 = ~n1017 & ~n1023;
  assign n1070 = n1068 & n1069;
  assign n1071 = n1067 & n1070;
  assign n1072 = n1055 & ~n1071;
  assign n1073 = ~n1064 & ~n1072;
  assign n1074 = pi095 & ~pi195;
  assign n1075 = ~pi095 & pi195;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = ~n1073 & n1076;
  assign n1078 = ~n1064 & ~n1076;
  assign n1079 = ~n1072 & n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = n210 & ~n1080;
  assign n1082 = ~n210 & ~n1079;
  assign n1083 = ~n1077 & n1082;
  assign n1084 = pi097 & ~pi197;
  assign n1085 = ~pi097 & pi197;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1083 & ~n1086;
  assign n1088 = ~n1081 & n1087;
  assign n1089 = ~n1081 & ~n1083;
  assign n1090 = n1086 & ~n1089;
  assign n1091 = ~n1088 & ~n1090;
  assign n1092 = pi098 & ~pi198;
  assign n1093 = ~pi098 & pi198;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = ~n1091 & n1094;
  assign n1096 = ~n1088 & ~n1094;
  assign n1097 = ~n1090 & n1096;
  assign n1098 = pi099 & ~pi199;
  assign n1099 = ~pi099 & pi199;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n1097 & ~n1100;
  assign n1102 = ~n1095 & n1101;
  assign n1103 = ~n1095 & ~n1097;
  assign n1104 = n1100 & ~n1103;
  assign po0 = ~n1102 & ~n1104;
  assign n1106 = ~n1090 & ~n1094;
  assign n1107 = ~n1088 & ~n1106;
  assign n1108 = ~n1005 & ~n1014;
  assign n1109 = ~n961 & n1014;
  assign n1110 = ~n993 & n1109;
  assign n1111 = n1029 & n1110;
  assign n1112 = n1027 & n1111;
  assign n1113 = ~n1008 & ~n1112;
  assign n1114 = ~n1108 & ~n1113;
  assign n1115 = ~n433 & n685;
  assign n1116 = ~n441 & n1115;
  assign n1117 = ~n442 & ~n685;
  assign n1118 = ~n611 & ~n1117;
  assign n1119 = ~n1116 & n1118;
  assign n1120 = ~n1116 & ~n1117;
  assign n1121 = n611 & ~n1120;
  assign n1122 = ~n1119 & ~n1121;
  assign n1123 = n614 & ~n1122;
  assign n1124 = ~n614 & ~n1119;
  assign n1125 = ~n1121 & n1124;
  assign n1126 = n639 & ~n1125;
  assign n1127 = ~n1123 & n1126;
  assign n1128 = ~n1123 & ~n1125;
  assign n1129 = ~n639 & ~n1128;
  assign n1130 = ~n1127 & ~n1129;
  assign n1131 = ~n621 & ~n1130;
  assign n1132 = ~n622 & ~n1131;
  assign n1133 = ~n637 & ~n1127;
  assign n1134 = ~n562 & ~n1122;
  assign n1135 = ~n1125 & ~n1134;
  assign n1136 = ~n1133 & ~n1135;
  assign n1137 = ~n637 & ~n1125;
  assign n1138 = ~n1134 & n1137;
  assign n1139 = ~n1127 & n1138;
  assign n1140 = ~n1136 & ~n1139;
  assign n1141 = ~n1132 & n1140;
  assign n1142 = n1132 & ~n1140;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n396 & n404;
  assign n1145 = ~n397 & n1144;
  assign n1146 = ~n525 & n1145;
  assign n1147 = ~n527 & n1146;
  assign n1148 = ~n440 & n1147;
  assign n1149 = ~n348 & ~n525;
  assign n1150 = ~n527 & n1149;
  assign n1151 = n359 & n430;
  assign n1152 = ~n398 & n404;
  assign n1153 = ~n363 & n1152;
  assign n1154 = n423 & n1153;
  assign n1155 = n1151 & n1154;
  assign n1156 = n1150 & n1155;
  assign n1157 = ~n1148 & ~n1156;
  assign n1158 = ~n396 & ~n404;
  assign n1159 = ~n397 & n1158;
  assign n1160 = ~n363 & n1159;
  assign n1161 = n423 & n1160;
  assign n1162 = n1151 & n1161;
  assign n1163 = n1150 & n1162;
  assign n1164 = ~n398 & ~n404;
  assign n1165 = ~n525 & n1164;
  assign n1166 = ~n527 & n1165;
  assign n1167 = ~n440 & n1166;
  assign n1168 = ~n1163 & ~n1167;
  assign n1169 = n1157 & n1168;
  assign n1170 = ~n363 & n1145;
  assign n1171 = ~n528 & n1170;
  assign n1172 = n431 & n1171;
  assign n1173 = n360 & n1172;
  assign n1174 = ~n528 & n1152;
  assign n1175 = ~n440 & n1174;
  assign n1176 = ~n1173 & ~n1175;
  assign n1177 = ~n528 & n1159;
  assign n1178 = ~n440 & n1177;
  assign n1179 = ~n363 & n1164;
  assign n1180 = ~n528 & n1179;
  assign n1181 = n431 & n1180;
  assign n1182 = n360 & n1181;
  assign n1183 = ~n1178 & ~n1182;
  assign n1184 = n1176 & n1183;
  assign n1185 = n1169 & n1184;
  assign n1186 = ~n386 & ~n1185;
  assign n1187 = ~n387 & ~n1186;
  assign n1188 = ~n1156 & ~n1163;
  assign n1189 = ~n1167 & n1188;
  assign n1190 = ~n1175 & ~n1178;
  assign n1191 = ~n1148 & ~n1182;
  assign n1192 = n1190 & n1191;
  assign n1193 = ~n545 & ~n1173;
  assign n1194 = n1192 & n1193;
  assign n1195 = n1189 & n1194;
  assign n1196 = ~n544 & ~n1195;
  assign n1197 = ~n1187 & n1196;
  assign n1198 = n1187 & ~n1196;
  assign n1199 = ~n1197 & ~n1198;
  assign n1200 = ~n433 & ~n570;
  assign n1201 = n686 & n1200;
  assign n1202 = n570 & ~n685;
  assign n1203 = ~n442 & n1202;
  assign n1204 = ~n1201 & ~n1203;
  assign n1205 = ~n548 & ~n570;
  assign n1206 = n662 & n1205;
  assign n1207 = ~n442 & n1206;
  assign n1208 = ~n548 & n570;
  assign n1209 = n662 & n1208;
  assign n1210 = n442 & n1209;
  assign n1211 = ~n1207 & ~n1210;
  assign n1212 = n1204 & n1211;
  assign n1213 = ~n584 & ~n1212;
  assign n1214 = ~n401 & ~n1120;
  assign n1215 = ~n570 & ~n1117;
  assign n1216 = ~n1116 & n1215;
  assign n1217 = ~n583 & ~n1216;
  assign n1218 = ~n1214 & n1217;
  assign n1219 = ~n1213 & n1218;
  assign n1220 = ~n1199 & n1219;
  assign n1221 = ~n583 & ~n1213;
  assign n1222 = ~n1214 & ~n1216;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1199 & n1223;
  assign n1225 = ~n1220 & ~n1224;
  assign n1226 = n1221 & ~n1222;
  assign n1227 = n1199 & n1226;
  assign n1228 = ~n1197 & n1222;
  assign n1229 = ~n1198 & ~n1221;
  assign n1230 = n1228 & n1229;
  assign n1231 = ~n1227 & ~n1230;
  assign n1232 = n1225 & n1231;
  assign n1233 = ~n573 & ~n585;
  assign n1234 = ~n1201 & n1233;
  assign n1235 = ~n1203 & ~n1207;
  assign n1236 = ~n1210 & n1235;
  assign n1237 = n1234 & n1236;
  assign n1238 = ~n588 & n599;
  assign n1239 = ~n586 & ~n599;
  assign n1240 = ~n587 & n1239;
  assign n1241 = ~n1238 & ~n1240;
  assign n1242 = ~n685 & ~n1241;
  assign n1243 = ~n442 & n1242;
  assign n1244 = ~n548 & ~n1241;
  assign n1245 = n662 & n1244;
  assign n1246 = n442 & n1245;
  assign n1247 = ~n1243 & ~n1246;
  assign n1248 = ~n433 & n1241;
  assign n1249 = n686 & n1248;
  assign n1250 = ~n548 & n1241;
  assign n1251 = n662 & n1250;
  assign n1252 = ~n442 & n1251;
  assign n1253 = ~n1249 & ~n1252;
  assign n1254 = n1247 & n1253;
  assign n1255 = ~n599 & ~n1254;
  assign n1256 = ~n573 & ~n583;
  assign n1257 = ~n584 & n1256;
  assign n1258 = ~n1212 & n1257;
  assign n1259 = ~n1255 & ~n1258;
  assign n1260 = ~n1237 & n1259;
  assign n1261 = ~n596 & ~n1241;
  assign n1262 = ~n685 & n1261;
  assign n1263 = ~n442 & n1262;
  assign n1264 = ~n595 & ~n1263;
  assign n1265 = ~n596 & ~n1238;
  assign n1266 = ~n1240 & n1265;
  assign n1267 = ~n548 & n1266;
  assign n1268 = n662 & n1267;
  assign n1269 = ~n442 & n1268;
  assign n1270 = ~n548 & n1261;
  assign n1271 = n662 & n1270;
  assign n1272 = n442 & n1271;
  assign n1273 = ~n433 & n1266;
  assign n1274 = n686 & n1273;
  assign n1275 = ~n1272 & ~n1274;
  assign n1276 = ~n1269 & n1275;
  assign n1277 = n1264 & n1276;
  assign n1278 = ~n1260 & ~n1277;
  assign n1279 = ~n558 & ~n596;
  assign n1280 = ~n595 & n1279;
  assign n1281 = ~n1254 & n1280;
  assign n1282 = ~n558 & ~n602;
  assign n1283 = ~n1243 & n1282;
  assign n1284 = ~n1246 & ~n1249;
  assign n1285 = ~n1252 & n1284;
  assign n1286 = n1283 & n1285;
  assign n1287 = ~n559 & ~n1286;
  assign n1288 = ~n1281 & n1287;
  assign n1289 = ~n1237 & ~n1258;
  assign n1290 = ~n1255 & n1277;
  assign n1291 = n1289 & n1290;
  assign n1292 = ~n1288 & ~n1291;
  assign n1293 = ~n1278 & n1292;
  assign n1294 = ~n1277 & ~n1281;
  assign n1295 = n1287 & n1294;
  assign n1296 = ~n1260 & n1295;
  assign n1297 = ~n559 & ~n595;
  assign n1298 = ~n1263 & n1297;
  assign n1299 = n1276 & n1298;
  assign n1300 = ~n1255 & n1299;
  assign n1301 = ~n1281 & ~n1286;
  assign n1302 = n1289 & n1301;
  assign n1303 = n1300 & n1302;
  assign n1304 = ~n1296 & ~n1303;
  assign n1305 = ~n1293 & n1304;
  assign n1306 = ~n1232 & ~n1305;
  assign n1307 = n1232 & n1305;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = ~n1143 & n1308;
  assign n1310 = n1143 & ~n1308;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = n404 & ~n467;
  assign n1313 = ~n469 & n1312;
  assign n1314 = ~n363 & n1313;
  assign n1315 = n431 & n1314;
  assign n1316 = n360 & n1315;
  assign n1317 = ~n404 & ~n467;
  assign n1318 = ~n469 & n1317;
  assign n1319 = ~n440 & n1318;
  assign n1320 = ~n1316 & ~n1319;
  assign n1321 = n404 & ~n470;
  assign n1322 = ~n440 & n1321;
  assign n1323 = ~n404 & ~n470;
  assign n1324 = ~n363 & n1323;
  assign n1325 = n431 & n1324;
  assign n1326 = n360 & n1325;
  assign n1327 = ~n1322 & ~n1326;
  assign n1328 = n1320 & n1327;
  assign n1329 = n481 & ~n1328;
  assign n1330 = n404 & ~n481;
  assign n1331 = ~n467 & n1330;
  assign n1332 = ~n469 & n1331;
  assign n1333 = ~n440 & n1332;
  assign n1334 = ~n404 & ~n481;
  assign n1335 = ~n467 & n1334;
  assign n1336 = ~n469 & n1335;
  assign n1337 = ~n363 & n1336;
  assign n1338 = n431 & n1337;
  assign n1339 = n360 & n1338;
  assign n1340 = ~n1333 & ~n1339;
  assign n1341 = ~n470 & n1330;
  assign n1342 = ~n363 & n1341;
  assign n1343 = n431 & n1342;
  assign n1344 = n360 & n1343;
  assign n1345 = ~n470 & n1334;
  assign n1346 = ~n440 & n1345;
  assign n1347 = ~n1344 & ~n1346;
  assign n1348 = n1340 & n1347;
  assign n1349 = ~n1329 & n1348;
  assign n1350 = ~n477 & ~n1349;
  assign n1351 = ~n478 & ~n1350;
  assign n1352 = ~n329 & ~n332;
  assign n1353 = ~n349 & n1352;
  assign n1354 = ~n277 & ~n281;
  assign n1355 = ~n285 & n1354;
  assign n1356 = ~n294 & ~n299;
  assign n1357 = ~n273 & ~n302;
  assign n1358 = n1356 & n1357;
  assign n1359 = ~n290 & n333;
  assign n1360 = n1358 & n1359;
  assign n1361 = n1355 & n1360;
  assign n1362 = ~n1353 & ~n1361;
  assign n1363 = n329 & n332;
  assign n1364 = ~n326 & ~n1363;
  assign n1365 = ~n349 & n1364;
  assign n1366 = ~n326 & ~n334;
  assign n1367 = ~n290 & n1366;
  assign n1368 = n1358 & n1367;
  assign n1369 = n1355 & n1368;
  assign n1370 = ~n1365 & ~n1369;
  assign n1371 = n1362 & n1370;
  assign n1372 = ~n273 & ~n332;
  assign n1373 = n1355 & n1372;
  assign n1374 = n304 & ~n1373;
  assign n1375 = ~n262 & ~n269;
  assign n1376 = ~n253 & n1375;
  assign n1377 = ~n254 & n1376;
  assign n1378 = ~n262 & n269;
  assign n1379 = ~n255 & n1378;
  assign n1380 = ~n263 & ~n1379;
  assign n1381 = ~n1377 & n1380;
  assign n1382 = n237 & ~n251;
  assign n1383 = ~n250 & ~n1382;
  assign n1384 = n269 & ~n1383;
  assign n1385 = ~n255 & n1384;
  assign n1386 = ~n250 & ~n269;
  assign n1387 = ~n1382 & n1386;
  assign n1388 = ~n255 & n1387;
  assign n1389 = n242 & n251;
  assign n1390 = n241 & n250;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1388 & n1391;
  assign n1393 = ~n1385 & n1392;
  assign n1394 = ~n1381 & n1393;
  assign n1395 = n1381 & ~n1393;
  assign n1396 = ~n1394 & ~n1395;
  assign n1397 = ~n1374 & n1396;
  assign n1398 = n1374 & ~n1396;
  assign n1399 = ~n1397 & ~n1398;
  assign n1400 = ~n1371 & n1399;
  assign n1401 = n1371 & ~n1399;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = ~n321 & ~n344;
  assign n1404 = ~n336 & n1403;
  assign n1405 = ~n290 & n1404;
  assign n1406 = n1358 & n1405;
  assign n1407 = n1355 & n1406;
  assign n1408 = ~n321 & ~n354;
  assign n1409 = ~n349 & n1408;
  assign n1410 = ~n320 & ~n1409;
  assign n1411 = ~n1407 & n1410;
  assign n1412 = ~n312 & ~n322;
  assign n1413 = ~n344 & n1412;
  assign n1414 = ~n336 & n1413;
  assign n1415 = ~n349 & n1414;
  assign n1416 = ~n354 & n1412;
  assign n1417 = ~n290 & n1416;
  assign n1418 = n1358 & n1417;
  assign n1419 = n1355 & n1418;
  assign n1420 = ~n312 & ~n320;
  assign n1421 = ~n311 & ~n1420;
  assign n1422 = ~n1419 & n1421;
  assign n1423 = ~n1415 & n1422;
  assign n1424 = ~n1411 & n1423;
  assign n1425 = ~n311 & ~n1419;
  assign n1426 = ~n1415 & n1425;
  assign n1427 = n1411 & ~n1426;
  assign n1428 = ~n1424 & ~n1427;
  assign n1429 = n1402 & ~n1428;
  assign n1430 = ~n1402 & n1428;
  assign n1431 = ~n404 & ~n429;
  assign n1432 = n360 & n1431;
  assign n1433 = n439 & ~n1432;
  assign n1434 = ~n1430 & ~n1433;
  assign n1435 = ~n1429 & n1434;
  assign n1436 = ~n1429 & ~n1430;
  assign n1437 = n1433 & ~n1436;
  assign n1438 = ~n1435 & ~n1437;
  assign n1439 = ~n404 & ~n461;
  assign n1440 = ~n363 & n1439;
  assign n1441 = n431 & n1440;
  assign n1442 = n360 & n1441;
  assign n1443 = n404 & ~n461;
  assign n1444 = ~n440 & n1443;
  assign n1445 = ~n462 & ~n1444;
  assign n1446 = ~n1442 & n1445;
  assign n1447 = n404 & ~n452;
  assign n1448 = ~n463 & n1447;
  assign n1449 = ~n440 & n1448;
  assign n1450 = ~n453 & ~n1449;
  assign n1451 = ~n404 & ~n452;
  assign n1452 = n463 & n1451;
  assign n1453 = ~n440 & n1452;
  assign n1454 = ~n463 & n1451;
  assign n1455 = ~n363 & n1454;
  assign n1456 = n431 & n1455;
  assign n1457 = n360 & n1456;
  assign n1458 = n463 & n1447;
  assign n1459 = ~n363 & n1458;
  assign n1460 = n431 & n1459;
  assign n1461 = n360 & n1460;
  assign n1462 = ~n1457 & ~n1461;
  assign n1463 = ~n1453 & n1462;
  assign n1464 = n1450 & n1463;
  assign n1465 = ~n1446 & n1464;
  assign n1466 = ~n1438 & n1465;
  assign n1467 = n1446 & ~n1464;
  assign n1468 = ~n1438 & n1467;
  assign n1469 = ~n1466 & ~n1468;
  assign n1470 = ~n1444 & ~n1453;
  assign n1471 = ~n1442 & n1470;
  assign n1472 = ~n453 & ~n462;
  assign n1473 = ~n1449 & n1472;
  assign n1474 = n1462 & n1473;
  assign n1475 = n1471 & n1474;
  assign n1476 = ~n1435 & n1475;
  assign n1477 = ~n1437 & n1476;
  assign n1478 = ~n1435 & ~n1446;
  assign n1479 = ~n1437 & ~n1464;
  assign n1480 = n1478 & n1479;
  assign n1481 = ~n1477 & ~n1480;
  assign n1482 = n1469 & n1481;
  assign n1483 = n1351 & n1482;
  assign n1484 = ~n483 & ~n494;
  assign n1485 = ~n485 & n1484;
  assign n1486 = ~n1316 & n1485;
  assign n1487 = ~n1319 & ~n1322;
  assign n1488 = ~n1326 & n1487;
  assign n1489 = n1486 & n1488;
  assign n1490 = ~n486 & ~n494;
  assign n1491 = ~n1328 & n1490;
  assign n1492 = ~n493 & ~n1491;
  assign n1493 = ~n1489 & n1492;
  assign n1494 = ~n445 & ~n1328;
  assign n1495 = n1348 & ~n1494;
  assign n1496 = ~n1493 & n1495;
  assign n1497 = n1493 & ~n1495;
  assign n1498 = ~n1496 & ~n1497;
  assign n1499 = ~n1483 & n1498;
  assign n1500 = ~n1351 & ~n1482;
  assign n1501 = ~n404 & ~n440;
  assign n1502 = ~n363 & n404;
  assign n1503 = n431 & n1502;
  assign n1504 = n360 & n1503;
  assign n1505 = n528 & ~n1504;
  assign n1506 = ~n1501 & n1505;
  assign n1507 = ~n1501 & ~n1504;
  assign n1508 = ~n528 & ~n1507;
  assign n1509 = ~n1506 & ~n1508;
  assign n1510 = ~n513 & ~n1509;
  assign n1511 = n404 & ~n526;
  assign n1512 = ~n363 & n1511;
  assign n1513 = n431 & n1512;
  assign n1514 = n360 & n1513;
  assign n1515 = ~n510 & ~n516;
  assign n1516 = ~n1514 & n1515;
  assign n1517 = ~n404 & ~n507;
  assign n1518 = ~n506 & n1517;
  assign n1519 = ~n363 & n1518;
  assign n1520 = n431 & n1519;
  assign n1521 = n360 & n1520;
  assign n1522 = ~n404 & ~n526;
  assign n1523 = ~n440 & n1522;
  assign n1524 = n404 & ~n507;
  assign n1525 = ~n506 & n1524;
  assign n1526 = ~n440 & n1525;
  assign n1527 = ~n1523 & ~n1526;
  assign n1528 = ~n1521 & n1527;
  assign n1529 = n1516 & n1528;
  assign n1530 = ~n1514 & ~n1523;
  assign n1531 = ~n1521 & ~n1526;
  assign n1532 = n1530 & n1531;
  assign n1533 = n510 & ~n516;
  assign n1534 = ~n1532 & n1533;
  assign n1535 = ~n1529 & ~n1534;
  assign n1536 = ~n1510 & n1535;
  assign n1537 = ~n510 & ~n1532;
  assign n1538 = ~n497 & ~n1514;
  assign n1539 = n1528 & n1538;
  assign n1540 = ~n1537 & ~n1539;
  assign n1541 = ~n370 & ~n528;
  assign n1542 = ~n1507 & n1541;
  assign n1543 = ~n370 & ~n525;
  assign n1544 = ~n527 & n1543;
  assign n1545 = ~n1504 & n1544;
  assign n1546 = ~n1501 & n1545;
  assign n1547 = ~n371 & ~n1546;
  assign n1548 = ~n1542 & n1547;
  assign n1549 = ~n1540 & n1548;
  assign n1550 = ~n1536 & n1549;
  assign n1551 = ~n1540 & ~n1548;
  assign n1552 = n1536 & n1551;
  assign n1553 = ~n1550 & ~n1552;
  assign n1554 = n1535 & n1540;
  assign n1555 = ~n1510 & n1548;
  assign n1556 = n1554 & n1555;
  assign n1557 = n1540 & ~n1548;
  assign n1558 = ~n1536 & n1557;
  assign n1559 = ~n1556 & ~n1558;
  assign n1560 = n1553 & n1559;
  assign n1561 = ~n1500 & ~n1560;
  assign n1562 = n1499 & n1561;
  assign n1563 = ~n1483 & ~n1500;
  assign n1564 = ~n1498 & ~n1560;
  assign n1565 = ~n1563 & n1564;
  assign n1566 = ~n1562 & ~n1565;
  assign n1567 = n1498 & n1560;
  assign n1568 = ~n1563 & n1567;
  assign n1569 = ~n1498 & n1560;
  assign n1570 = n1563 & n1569;
  assign n1571 = ~n1568 & ~n1570;
  assign n1572 = n1566 & n1571;
  assign n1573 = n546 & ~n1185;
  assign n1574 = ~n546 & ~n1173;
  assign n1575 = n1192 & n1574;
  assign n1576 = n1189 & n1575;
  assign n1577 = ~n1573 & ~n1576;
  assign n1578 = ~n535 & ~n1577;
  assign n1579 = ~n536 & ~n1578;
  assign n1580 = ~n374 & ~n390;
  assign n1581 = n378 & ~n1506;
  assign n1582 = ~n1508 & n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584 = ~n371 & ~n390;
  assign n1585 = ~n370 & n1584;
  assign n1586 = ~n1509 & n1585;
  assign n1587 = ~n377 & ~n390;
  assign n1588 = ~n1506 & n1587;
  assign n1589 = ~n1508 & n1588;
  assign n1590 = ~n371 & ~n374;
  assign n1591 = ~n370 & n1590;
  assign n1592 = ~n1509 & n1591;
  assign n1593 = ~n1589 & ~n1592;
  assign n1594 = ~n1586 & n1593;
  assign n1595 = n1583 & n1594;
  assign n1596 = ~n1579 & n1595;
  assign n1597 = n1579 & ~n1595;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n1572 & ~n1598;
  assign n1600 = ~n1562 & n1598;
  assign n1601 = ~n1565 & ~n1568;
  assign n1602 = ~n1570 & n1601;
  assign n1603 = n1600 & n1602;
  assign n1604 = ~n1599 & ~n1603;
  assign n1605 = ~n1311 & n1604;
  assign n1606 = n1311 & ~n1604;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = ~n687 & ~n704;
  assign n1609 = n720 & n1608;
  assign n1610 = n716 & n1609;
  assign n1611 = ~n705 & ~n1610;
  assign n1612 = n650 & ~n1117;
  assign n1613 = ~n1116 & n1612;
  assign n1614 = ~n650 & ~n1120;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n551 & ~n1615;
  assign n1617 = ~n625 & ~n1613;
  assign n1618 = ~n1614 & n1617;
  assign n1619 = ~n1616 & ~n1618;
  assign n1620 = ~n1611 & n1619;
  assign n1621 = n1611 & ~n1619;
  assign n1622 = ~n1620 & ~n1621;
  assign n1623 = ~n234 & ~n714;
  assign n1624 = ~n722 & n1623;
  assign n1625 = ~n697 & n712;
  assign n1626 = ~n705 & ~n708;
  assign n1627 = ~n704 & n1626;
  assign n1628 = ~n687 & n1627;
  assign n1629 = n720 & n1628;
  assign n1630 = n716 & n1629;
  assign n1631 = ~n1625 & ~n1630;
  assign n1632 = ~n1624 & n1631;
  assign n1633 = ~n1622 & n1632;
  assign n1634 = n1622 & ~n1632;
  assign n1635 = ~n1633 & ~n1634;
  assign n1636 = ~n1607 & n1635;
  assign n1637 = ~n1605 & ~n1635;
  assign n1638 = ~n1606 & n1637;
  assign n1639 = ~n1636 & ~n1638;
  assign n1640 = n213 & ~n724;
  assign n1641 = ~n726 & n1640;
  assign n1642 = ~n213 & ~n727;
  assign n1643 = ~n216 & ~n227;
  assign n1644 = ~n1642 & n1643;
  assign n1645 = ~n1641 & n1644;
  assign n1646 = ~n1639 & n1645;
  assign n1647 = ~n1607 & ~n1622;
  assign n1648 = ~n1605 & n1622;
  assign n1649 = ~n1606 & n1648;
  assign n1650 = ~n1647 & ~n1649;
  assign n1651 = n1632 & ~n1642;
  assign n1652 = ~n213 & ~n1631;
  assign n1653 = ~n727 & n1652;
  assign n1654 = ~n1651 & ~n1653;
  assign n1655 = ~n1650 & n1654;
  assign n1656 = ~n1647 & ~n1654;
  assign n1657 = ~n1649 & n1656;
  assign n1658 = ~n1655 & ~n1657;
  assign n1659 = ~n1646 & ~n1658;
  assign n1660 = ~n216 & ~n1642;
  assign n1661 = ~n1641 & n1660;
  assign n1662 = ~n1636 & n1661;
  assign n1663 = ~n1638 & n1662;
  assign n1664 = ~n1641 & ~n1642;
  assign n1665 = n216 & ~n1664;
  assign n1666 = ~n226 & ~n1661;
  assign n1667 = ~n1665 & n1666;
  assign n1668 = ~n227 & ~n1667;
  assign n1669 = ~n1663 & n1668;
  assign n1670 = ~n1659 & n1669;
  assign n1671 = n1646 & ~n1655;
  assign n1672 = ~n1657 & n1671;
  assign n1673 = ~n216 & n227;
  assign n1674 = ~n1642 & n1673;
  assign n1675 = ~n1641 & n1674;
  assign n1676 = ~n1639 & n1675;
  assign n1677 = ~n1672 & n1676;
  assign n1678 = ~n1670 & n1677;
  assign n1679 = ~n1670 & ~n1672;
  assign n1680 = ~n1636 & n1675;
  assign n1681 = ~n1638 & n1680;
  assign n1682 = n1654 & ~n1668;
  assign n1683 = ~n1650 & n1682;
  assign n1684 = ~n1654 & ~n1668;
  assign n1685 = ~n1647 & n1684;
  assign n1686 = ~n1649 & n1685;
  assign n1687 = ~n1683 & ~n1686;
  assign n1688 = ~n1681 & n1687;
  assign n1689 = ~n1679 & n1688;
  assign n1690 = ~n1678 & ~n1689;
  assign n1691 = ~n779 & ~n782;
  assign n1692 = n777 & n1691;
  assign n1693 = n760 & n1692;
  assign n1694 = n782 & ~n812;
  assign n1695 = ~n785 & ~n1694;
  assign n1696 = ~n1693 & ~n1695;
  assign n1697 = ~n737 & ~n750;
  assign n1698 = ~n738 & ~n1697;
  assign n1699 = ~n811 & ~n1698;
  assign n1700 = ~n750 & n755;
  assign n1701 = ~n730 & ~n755;
  assign n1702 = ~n728 & n1701;
  assign n1703 = ~n1700 & ~n1702;
  assign n1704 = ~n744 & ~n1698;
  assign n1705 = ~n1703 & n1704;
  assign n1706 = ~n744 & ~n1703;
  assign n1707 = n1698 & ~n1706;
  assign n1708 = ~n1705 & ~n1707;
  assign n1709 = n811 & ~n1708;
  assign n1710 = ~n1699 & ~n1709;
  assign n1711 = ~n1696 & ~n1710;
  assign n1712 = ~n1693 & ~n1699;
  assign n1713 = ~n1695 & n1712;
  assign n1714 = ~n1709 & n1713;
  assign n1715 = ~n1675 & ~n1714;
  assign n1716 = ~n1711 & n1715;
  assign n1717 = n1687 & n1716;
  assign n1718 = ~n1675 & ~n1683;
  assign n1719 = ~n1686 & n1718;
  assign n1720 = ~n1711 & ~n1714;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1717 & ~n1721;
  assign n1723 = ~n849 & ~n891;
  assign n1724 = ~n848 & ~n1723;
  assign n1725 = ~n1722 & n1724;
  assign n1726 = ~n1690 & n1725;
  assign n1727 = ~n1678 & ~n1722;
  assign n1728 = ~n1724 & n1727;
  assign n1729 = ~n1689 & n1728;
  assign n1730 = ~n1726 & ~n1729;
  assign n1731 = ~n848 & ~n1717;
  assign n1732 = ~n1723 & n1731;
  assign n1733 = ~n1721 & n1732;
  assign n1734 = n1690 & n1733;
  assign n1735 = n1722 & ~n1724;
  assign n1736 = ~n1690 & n1735;
  assign n1737 = ~n1734 & ~n1736;
  assign n1738 = n1730 & n1737;
  assign n1739 = n850 & ~n891;
  assign n1740 = n834 & ~n850;
  assign n1741 = ~n882 & n1740;
  assign n1742 = n838 & ~n850;
  assign n1743 = ~n882 & n1742;
  assign n1744 = ~n850 & n883;
  assign n1745 = ~n827 & n1744;
  assign n1746 = n823 & n1745;
  assign n1747 = n817 & n1746;
  assign n1748 = ~n850 & n885;
  assign n1749 = ~n827 & n1748;
  assign n1750 = n823 & n1749;
  assign n1751 = n817 & n1750;
  assign n1752 = ~n1747 & ~n1751;
  assign n1753 = ~n1743 & n1752;
  assign n1754 = ~n1741 & n1753;
  assign n1755 = ~n1739 & n1754;
  assign n1756 = n859 & ~n1755;
  assign n1757 = ~n859 & ~n1747;
  assign n1758 = ~n1751 & n1757;
  assign n1759 = ~n1741 & ~n1743;
  assign n1760 = n1758 & n1759;
  assign n1761 = ~n1739 & n1760;
  assign n1762 = ~n864 & ~n1761;
  assign n1763 = ~n1756 & n1762;
  assign n1764 = ~n864 & ~n867;
  assign n1765 = ~n867 & ~n1761;
  assign n1766 = ~n1756 & n1765;
  assign n1767 = ~n1764 & ~n1766;
  assign n1768 = ~n1763 & n1767;
  assign n1769 = ~n858 & ~n1755;
  assign n1770 = ~n857 & ~n1769;
  assign n1771 = ~n812 & n813;
  assign n1772 = ~n779 & ~n813;
  assign n1773 = n777 & n1772;
  assign n1774 = n760 & n1773;
  assign n1775 = ~n794 & ~n1774;
  assign n1776 = ~n1771 & n1775;
  assign n1777 = ~n800 & ~n1776;
  assign n1778 = n830 & ~n882;
  assign n1779 = ~n833 & ~n1778;
  assign n1780 = ~n827 & ~n830;
  assign n1781 = n823 & n1780;
  assign n1782 = n817 & n1781;
  assign n1783 = ~n1779 & ~n1782;
  assign n1784 = ~n1777 & ~n1783;
  assign n1785 = ~n1771 & ~n1774;
  assign n1786 = n794 & ~n830;
  assign n1787 = ~n1785 & n1786;
  assign n1788 = n1777 & ~n1787;
  assign n1789 = ~n1779 & n1788;
  assign n1790 = ~n1784 & ~n1789;
  assign n1791 = ~n1770 & n1790;
  assign n1792 = ~n857 & ~n1790;
  assign n1793 = ~n1769 & n1792;
  assign n1794 = ~n1791 & ~n1793;
  assign n1795 = ~n1768 & n1794;
  assign n1796 = ~n1738 & n1795;
  assign n1797 = ~n893 & ~n905;
  assign n1798 = ~n888 & n905;
  assign n1799 = ~n892 & n1798;
  assign n1800 = ~n908 & ~n1799;
  assign n1801 = ~n1797 & ~n1800;
  assign n1802 = ~n1796 & ~n1801;
  assign n1803 = ~n1768 & ~n1794;
  assign n1804 = n1738 & n1803;
  assign n1805 = n1768 & ~n1794;
  assign n1806 = ~n1738 & n1805;
  assign n1807 = n1737 & ~n1791;
  assign n1808 = ~n1763 & ~n1793;
  assign n1809 = n1767 & n1808;
  assign n1810 = n1730 & n1809;
  assign n1811 = n1807 & n1810;
  assign n1812 = ~n1806 & ~n1811;
  assign n1813 = ~n1804 & n1812;
  assign n1814 = n1802 & n1813;
  assign n1815 = ~n1796 & ~n1806;
  assign n1816 = ~n1804 & ~n1811;
  assign n1817 = n1815 & n1816;
  assign n1818 = n1801 & ~n1817;
  assign n1819 = ~n949 & ~n991;
  assign n1820 = ~n940 & n949;
  assign n1821 = ~n936 & n1820;
  assign n1822 = n933 & n1821;
  assign n1823 = n921 & n1822;
  assign n1824 = n952 & ~n1823;
  assign n1825 = ~n1819 & n1824;
  assign n1826 = ~n955 & ~n1825;
  assign n1827 = ~n1819 & ~n1823;
  assign n1828 = ~n952 & ~n1827;
  assign n1829 = ~n947 & ~n991;
  assign n1830 = ~n948 & ~n1829;
  assign n1831 = ~n1797 & ~n1799;
  assign n1832 = n908 & ~n1831;
  assign n1833 = ~n1797 & n1800;
  assign n1834 = ~n901 & ~n1833;
  assign n1835 = ~n1832 & n1834;
  assign n1836 = ~n900 & ~n1835;
  assign n1837 = ~n1830 & ~n1836;
  assign n1838 = ~n1828 & n1837;
  assign n1839 = ~n1826 & n1838;
  assign n1840 = ~n1818 & n1839;
  assign n1841 = ~n1814 & n1840;
  assign n1842 = ~n1814 & ~n1818;
  assign n1843 = ~n1830 & n1836;
  assign n1844 = ~n1828 & n1843;
  assign n1845 = ~n1826 & n1844;
  assign n1846 = ~n1842 & n1845;
  assign n1847 = ~n1841 & ~n1846;
  assign n1848 = ~n900 & ~n948;
  assign n1849 = ~n1835 & n1848;
  assign n1850 = ~n1829 & n1849;
  assign n1851 = ~n1828 & n1850;
  assign n1852 = ~n1826 & n1851;
  assign n1853 = ~n1818 & n1852;
  assign n1854 = ~n1814 & n1853;
  assign n1855 = n1830 & ~n1836;
  assign n1856 = ~n1828 & n1855;
  assign n1857 = ~n1826 & n1856;
  assign n1858 = ~n1842 & n1857;
  assign n1859 = ~n1854 & ~n1858;
  assign n1860 = n1847 & n1859;
  assign n1861 = ~n1826 & ~n1828;
  assign n1862 = n1843 & ~n1861;
  assign n1863 = ~n1818 & n1862;
  assign n1864 = ~n1814 & n1863;
  assign n1865 = n1837 & ~n1861;
  assign n1866 = ~n1842 & n1865;
  assign n1867 = ~n1864 & ~n1866;
  assign n1868 = n1855 & ~n1861;
  assign n1869 = ~n1818 & n1868;
  assign n1870 = ~n1814 & n1869;
  assign n1871 = n1850 & ~n1861;
  assign n1872 = ~n1842 & n1871;
  assign n1873 = ~n1870 & ~n1872;
  assign n1874 = n1867 & n1873;
  assign n1875 = n1860 & n1874;
  assign n1876 = n1114 & ~n1875;
  assign n1877 = n1055 & ~n1060;
  assign n1878 = ~n1041 & n1877;
  assign n1879 = n1068 & n1878;
  assign n1880 = ~n1023 & n1066;
  assign n1881 = ~n1017 & n1880;
  assign n1882 = ~n1879 & n1881;
  assign n1883 = ~n1846 & ~n1854;
  assign n1884 = ~n1858 & n1883;
  assign n1885 = ~n1114 & ~n1864;
  assign n1886 = ~n1866 & ~n1870;
  assign n1887 = ~n1841 & ~n1872;
  assign n1888 = n1886 & n1887;
  assign n1889 = n1885 & n1888;
  assign n1890 = n1884 & n1889;
  assign n1891 = n1882 & ~n1890;
  assign n1892 = ~n1876 & n1891;
  assign n1893 = ~n1882 & n1885;
  assign n1894 = n1888 & n1893;
  assign n1895 = n1884 & n1894;
  assign n1896 = n1114 & ~n1882;
  assign n1897 = ~n1875 & n1896;
  assign n1898 = ~n1895 & ~n1897;
  assign n1899 = n1083 & n1898;
  assign n1900 = ~n1892 & n1899;
  assign n1901 = ~n1892 & n1898;
  assign n1902 = n1079 & ~n1901;
  assign n1903 = ~n1079 & ~n1895;
  assign n1904 = ~n1897 & n1903;
  assign n1905 = ~n1892 & n1904;
  assign n1906 = ~n1083 & ~n1905;
  assign n1907 = ~n1902 & n1906;
  assign n1908 = ~n1900 & ~n1907;
  assign n1909 = ~n1107 & n1908;
  assign n1910 = n1107 & ~n1908;
  assign n1911 = ~n1909 & ~n1910;
  assign n1912 = ~n1102 & ~n1911;
  assign n1913 = n1102 & ~n1909;
  assign n1914 = ~n1910 & n1913;
  assign n1915 = n1096 & ~n1900;
  assign n1916 = ~n1090 & n1915;
  assign n1917 = ~n1907 & n1916;
  assign n1918 = ~n1914 & ~n1917;
  assign po1 = ~n1912 & n1918;
  assign n1920 = n1024 & n1062;
  assign n1921 = n1049 & n1920;
  assign n1922 = ~n1017 & ~n1108;
  assign n1923 = ~n1113 & n1922;
  assign n1924 = ~n1864 & n1923;
  assign n1925 = n1921 & n1924;
  assign n1926 = n1888 & n1925;
  assign n1927 = n1884 & n1926;
  assign n1928 = n1063 & ~n1114;
  assign n1929 = n1025 & n1928;
  assign n1930 = ~n1875 & n1929;
  assign n1931 = ~n1079 & ~n1930;
  assign n1932 = ~n1927 & n1931;
  assign n1933 = ~n1052 & n1065;
  assign n1934 = ~n1020 & n1933;
  assign n1935 = ~n1114 & ~n1934;
  assign n1936 = ~n1875 & n1935;
  assign n1937 = ~n1858 & ~n1934;
  assign n1938 = n1883 & n1937;
  assign n1939 = n1114 & ~n1864;
  assign n1940 = n1888 & n1939;
  assign n1941 = n1938 & n1940;
  assign n1942 = ~n1936 & ~n1941;
  assign n1943 = n1898 & n1942;
  assign n1944 = ~n1932 & n1943;
  assign n1945 = ~n1818 & n1836;
  assign n1946 = ~n1814 & n1945;
  assign n1947 = ~n1836 & ~n1842;
  assign n1948 = ~n943 & ~n991;
  assign n1949 = ~n1830 & ~n1948;
  assign n1950 = ~n1947 & n1949;
  assign n1951 = ~n1946 & n1950;
  assign n1952 = ~n1946 & ~n1947;
  assign n1953 = n1830 & ~n1952;
  assign n1954 = ~n1830 & ~n1947;
  assign n1955 = ~n1946 & n1954;
  assign n1956 = ~n1861 & ~n1955;
  assign n1957 = ~n1953 & n1956;
  assign n1958 = ~n1951 & ~n1957;
  assign n1959 = n1676 & ~n1683;
  assign n1960 = ~n1686 & n1959;
  assign n1961 = ~n1679 & ~n1960;
  assign n1962 = ~n1676 & ~n1719;
  assign n1963 = n1698 & ~n1962;
  assign n1964 = ~n1961 & n1963;
  assign n1965 = ~n1658 & n1698;
  assign n1966 = ~n1659 & ~n1698;
  assign n1967 = ~n1965 & n1966;
  assign n1968 = ~n1639 & n1668;
  assign n1969 = ~n226 & ~n1665;
  assign n1970 = ~n227 & ~n1661;
  assign n1971 = ~n1969 & n1970;
  assign n1972 = n1706 & ~n1971;
  assign n1973 = ~n1968 & n1972;
  assign n1974 = ~n1672 & n1973;
  assign n1975 = ~n1676 & ~n1698;
  assign n1976 = n1688 & ~n1975;
  assign n1977 = ~n1974 & ~n1976;
  assign n1978 = n1967 & n1977;
  assign n1979 = n1706 & ~n1975;
  assign n1980 = ~n1688 & ~n1979;
  assign n1981 = ~n1706 & ~n1974;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n1978 & n1982;
  assign n1984 = ~n1964 & ~n1983;
  assign n1985 = ~n1466 & n1495;
  assign n1986 = ~n1468 & ~n1477;
  assign n1987 = ~n1480 & n1986;
  assign n1988 = n1985 & n1987;
  assign n1989 = ~n1482 & ~n1495;
  assign n1990 = ~n1351 & ~n1989;
  assign n1991 = ~n1988 & n1990;
  assign n1992 = ~n478 & ~n1333;
  assign n1993 = ~n1339 & ~n1344;
  assign n1994 = ~n1346 & n1993;
  assign n1995 = n1992 & n1994;
  assign n1996 = ~n1494 & n1995;
  assign n1997 = ~n1350 & n1996;
  assign n1998 = n1482 & n1997;
  assign n1999 = ~n478 & ~n1495;
  assign n2000 = ~n1350 & n1999;
  assign n2001 = ~n1482 & n2000;
  assign n2002 = n1493 & ~n2001;
  assign n2003 = ~n1998 & n2002;
  assign n2004 = ~n1991 & ~n2003;
  assign n2005 = ~n1433 & ~n1442;
  assign n2006 = n1445 & n2005;
  assign n2007 = n1436 & n2006;
  assign n2008 = ~n363 & ~n462;
  assign n2009 = n423 & ~n425;
  assign n2010 = n2008 & n2009;
  assign n2011 = ~n1432 & n2010;
  assign n2012 = ~n1444 & n2011;
  assign n2013 = ~n1442 & n2012;
  assign n2014 = ~n1436 & n2013;
  assign n2015 = ~n2007 & ~n2014;
  assign n2016 = ~n457 & ~n1507;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = ~n1464 & ~n1494;
  assign n2019 = ~n2017 & n2018;
  assign n2020 = ~n1437 & n1478;
  assign n2021 = n2015 & ~n2020;
  assign n2022 = ~n445 & ~n453;
  assign n2023 = ~n1449 & n2022;
  assign n2024 = n1463 & n2023;
  assign n2025 = ~n1328 & n2024;
  assign n2026 = ~n2017 & ~n2025;
  assign n2027 = ~n2021 & n2026;
  assign n2028 = ~n2019 & ~n2027;
  assign n2029 = ~n1348 & ~n1446;
  assign n2030 = ~n1464 & n2029;
  assign n2031 = ~n1438 & n2030;
  assign n2032 = ~n1348 & n1475;
  assign n2033 = ~n1438 & n2032;
  assign n2034 = ~n2031 & ~n2033;
  assign n2035 = n1464 & n2029;
  assign n2036 = n1438 & n2035;
  assign n2037 = ~n1348 & n1446;
  assign n2038 = ~n1435 & n2037;
  assign n2039 = n1479 & n2038;
  assign n2040 = ~n2036 & ~n2039;
  assign n2041 = n2034 & n2040;
  assign n2042 = ~n1436 & n2016;
  assign n2043 = n1433 & ~n2042;
  assign n2044 = ~n1388 & ~n1389;
  assign n2045 = ~n1394 & n2044;
  assign n2046 = n1362 & ~n1398;
  assign n2047 = ~n1370 & n2046;
  assign n2048 = n304 & ~n1396;
  assign n2049 = ~n290 & ~n1363;
  assign n2050 = n1358 & n2049;
  assign n2051 = n1355 & n2050;
  assign n2052 = ~n1353 & ~n2051;
  assign n2053 = ~n1397 & n2052;
  assign n2054 = ~n2048 & ~n2053;
  assign n2055 = ~n2047 & ~n2054;
  assign n2056 = ~n2045 & ~n2055;
  assign n2057 = n2045 & ~n2047;
  assign n2058 = ~n2054 & n2057;
  assign n2059 = ~n2056 & ~n2058;
  assign n2060 = ~n1424 & ~n1430;
  assign n2061 = ~n2059 & n2060;
  assign n2062 = n2059 & ~n2060;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = n1436 & ~n2016;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n2043 & n2065;
  assign n2067 = ~n2043 & ~n2064;
  assign n2068 = n2063 & ~n2067;
  assign n2069 = ~n2066 & ~n2068;
  assign n2070 = ~n2041 & ~n2069;
  assign n2071 = n2028 & n2070;
  assign n2072 = n2041 & ~n2069;
  assign n2073 = ~n2028 & n2072;
  assign n2074 = ~n2071 & ~n2073;
  assign n2075 = ~n2041 & n2069;
  assign n2076 = ~n2028 & n2075;
  assign n2077 = ~n2019 & ~n2066;
  assign n2078 = ~n2068 & n2077;
  assign n2079 = ~n2027 & n2041;
  assign n2080 = n2078 & n2079;
  assign n2081 = ~n2076 & ~n2080;
  assign n2082 = n2074 & n2081;
  assign n2083 = ~n2004 & n2082;
  assign n2084 = n2004 & ~n2082;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = ~n1536 & ~n1540;
  assign n2087 = n1499 & ~n1500;
  assign n2088 = ~n1498 & ~n1563;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = ~n1510 & n1554;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2086 & ~n2091;
  assign n2093 = ~n2085 & ~n2092;
  assign n2094 = ~n370 & n374;
  assign n2095 = ~n1509 & n2094;
  assign n2096 = ~n374 & ~n1506;
  assign n2097 = ~n1508 & n2096;
  assign n2098 = n371 & ~n2097;
  assign n2099 = ~n2095 & ~n2098;
  assign n2100 = ~n2093 & n2099;
  assign n2101 = n2085 & n2092;
  assign n2102 = ~n2086 & ~n2090;
  assign n2103 = ~n2089 & ~n2102;
  assign n2104 = n370 & ~n374;
  assign n2105 = ~n1506 & n2104;
  assign n2106 = ~n1508 & n2105;
  assign n2107 = ~n2087 & n2102;
  assign n2108 = ~n2088 & n2107;
  assign n2109 = ~n2106 & ~n2108;
  assign n2110 = ~n2103 & n2109;
  assign n2111 = ~n2101 & ~n2110;
  assign n2112 = n2100 & n2111;
  assign n2113 = ~n2093 & ~n2101;
  assign n2114 = n2099 & ~n2110;
  assign n2115 = ~n2113 & ~n2114;
  assign n2116 = ~n2112 & ~n2115;
  assign n2117 = n377 & ~n1506;
  assign n2118 = ~n1508 & n2117;
  assign n2119 = ~n377 & ~n1509;
  assign n2120 = ~n2118 & ~n2119;
  assign n2121 = ~n374 & ~n2120;
  assign n2122 = n374 & ~n2118;
  assign n2123 = ~n2119 & n2122;
  assign n2124 = ~n2121 & ~n2123;
  assign n2125 = ~n390 & ~n2124;
  assign n2126 = ~n1562 & n2125;
  assign n2127 = n1602 & n2126;
  assign n2128 = n1498 & ~n1595;
  assign n2129 = ~n1483 & n2128;
  assign n2130 = n1561 & n2129;
  assign n2131 = ~n1498 & ~n1595;
  assign n2132 = ~n1560 & n2131;
  assign n2133 = ~n1563 & n2132;
  assign n2134 = ~n2130 & ~n2133;
  assign n2135 = n1560 & n2128;
  assign n2136 = ~n1563 & n2135;
  assign n2137 = n1560 & n2131;
  assign n2138 = n1563 & n2137;
  assign n2139 = ~n2136 & ~n2138;
  assign n2140 = n2134 & n2139;
  assign n2141 = n1498 & n1595;
  assign n2142 = ~n1560 & n2141;
  assign n2143 = ~n1563 & n2142;
  assign n2144 = ~n1498 & n1595;
  assign n2145 = ~n1483 & n2144;
  assign n2146 = n1561 & n2145;
  assign n2147 = ~n2143 & ~n2146;
  assign n2148 = n1560 & n2141;
  assign n2149 = n1563 & n2148;
  assign n2150 = n1560 & n2144;
  assign n2151 = ~n1563 & n2150;
  assign n2152 = ~n2149 & ~n2151;
  assign n2153 = n2147 & n2152;
  assign n2154 = n2140 & n2153;
  assign n2155 = n1187 & ~n2154;
  assign n2156 = ~n2127 & ~n2155;
  assign n2157 = n531 & ~n1196;
  assign n2158 = n544 & ~n1173;
  assign n2159 = n1192 & n2158;
  assign n2160 = n1189 & n2159;
  assign n2161 = ~n1187 & ~n2160;
  assign n2162 = ~n2157 & n2161;
  assign n2163 = ~n2154 & n2162;
  assign n2164 = ~n2133 & ~n2136;
  assign n2165 = ~n2138 & n2164;
  assign n2166 = n1187 & ~n2160;
  assign n2167 = ~n2157 & n2166;
  assign n2168 = ~n2143 & n2167;
  assign n2169 = ~n2146 & ~n2149;
  assign n2170 = ~n2130 & ~n2151;
  assign n2171 = n2169 & n2170;
  assign n2172 = n2168 & n2171;
  assign n2173 = n2165 & n2172;
  assign n2174 = ~n531 & n545;
  assign n2175 = ~n1185 & n2174;
  assign n2176 = ~n2173 & ~n2175;
  assign n2177 = ~n2163 & n2176;
  assign n2178 = ~n2156 & n2177;
  assign n2179 = ~n2116 & n2178;
  assign n2180 = ~n1199 & ~n1222;
  assign n2181 = ~n1198 & n1228;
  assign n2182 = ~n2180 & ~n2181;
  assign n2183 = ~n1599 & n2182;
  assign n2184 = ~n1603 & n2183;
  assign n2185 = ~n1604 & ~n2182;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n573 & n584;
  assign n2188 = ~n1201 & n2187;
  assign n2189 = n1236 & n2188;
  assign n2190 = ~n2186 & ~n2189;
  assign n2191 = ~n1212 & ~n1256;
  assign n2192 = n573 & n582;
  assign n2193 = n579 & n2192;
  assign n2194 = ~n2191 & ~n2193;
  assign n2195 = ~n584 & ~n2194;
  assign n2196 = ~n2190 & ~n2195;
  assign n2197 = ~n2179 & n2196;
  assign n2198 = n2156 & ~n2177;
  assign n2199 = ~n2116 & n2198;
  assign n2200 = ~n2127 & ~n2175;
  assign n2201 = ~n2173 & n2200;
  assign n2202 = ~n2155 & ~n2163;
  assign n2203 = n2201 & n2202;
  assign n2204 = ~n2112 & n2203;
  assign n2205 = ~n2115 & n2204;
  assign n2206 = ~n2199 & ~n2205;
  assign n2207 = ~n2112 & ~n2156;
  assign n2208 = ~n2115 & ~n2177;
  assign n2209 = n2207 & n2208;
  assign n2210 = n1199 & ~n2143;
  assign n2211 = n2171 & n2210;
  assign n2212 = n2165 & n2211;
  assign n2213 = ~n1199 & ~n2154;
  assign n2214 = ~n531 & ~n1573;
  assign n2215 = ~n1576 & n2214;
  assign n2216 = n1579 & ~n2215;
  assign n2217 = ~n2213 & n2216;
  assign n2218 = ~n2212 & n2217;
  assign n2219 = n1199 & ~n1604;
  assign n2220 = ~n1199 & ~n1599;
  assign n2221 = ~n1603 & n2220;
  assign n2222 = ~n1222 & ~n2221;
  assign n2223 = ~n2219 & n2222;
  assign n2224 = ~n2218 & ~n2223;
  assign n2225 = ~n2209 & ~n2224;
  assign n2226 = n2206 & n2225;
  assign n2227 = n2197 & n2226;
  assign n2228 = ~n1278 & ~n1291;
  assign n2229 = ~n1598 & ~n2228;
  assign n2230 = n1232 & n2229;
  assign n2231 = ~n1572 & n2230;
  assign n2232 = n1598 & ~n2228;
  assign n2233 = n1232 & n2232;
  assign n2234 = n1572 & n2233;
  assign n2235 = ~n2231 & ~n2234;
  assign n2236 = ~n1232 & ~n1570;
  assign n2237 = n1601 & n2236;
  assign n2238 = ~n1562 & n2229;
  assign n2239 = n2237 & n2238;
  assign n2240 = ~n1232 & n2232;
  assign n2241 = ~n1572 & n2240;
  assign n2242 = ~n2239 & ~n2241;
  assign n2243 = n2235 & n2242;
  assign n2244 = ~n1224 & ~n1227;
  assign n2245 = ~n1230 & ~n1278;
  assign n2246 = n2244 & n2245;
  assign n2247 = ~n1220 & ~n1291;
  assign n2248 = ~n1598 & n2247;
  assign n2249 = n2246 & n2248;
  assign n2250 = n1572 & n2249;
  assign n2251 = n1598 & n2247;
  assign n2252 = n2246 & n2251;
  assign n2253 = ~n1572 & n2252;
  assign n2254 = ~n2250 & ~n2253;
  assign n2255 = ~n1598 & n2228;
  assign n2256 = ~n1232 & n2255;
  assign n2257 = ~n1572 & n2256;
  assign n2258 = n1598 & n2228;
  assign n2259 = ~n1562 & n2258;
  assign n2260 = n2237 & n2259;
  assign n2261 = ~n2257 & ~n2260;
  assign n2262 = n2254 & n2261;
  assign n2263 = n2243 & n2262;
  assign n2264 = n1288 & ~n2263;
  assign n2265 = ~n2234 & ~n2239;
  assign n2266 = ~n2241 & n2265;
  assign n2267 = ~n1288 & ~n2250;
  assign n2268 = ~n2253 & ~n2257;
  assign n2269 = ~n2231 & ~n2260;
  assign n2270 = n2268 & n2269;
  assign n2271 = n2267 & n2270;
  assign n2272 = n2266 & n2271;
  assign n2273 = ~n1134 & ~n2272;
  assign n2274 = ~n2264 & ~n2273;
  assign n2275 = ~n602 & ~n1254;
  assign n2276 = n602 & ~n1243;
  assign n2277 = n1285 & n2276;
  assign n2278 = ~n554 & ~n2277;
  assign n2279 = ~n2275 & n2278;
  assign n2280 = ~n2250 & n2279;
  assign n2281 = n2270 & n2280;
  assign n2282 = n2266 & n2281;
  assign n2283 = n1232 & ~n1598;
  assign n2284 = ~n1572 & n2283;
  assign n2285 = n1232 & ~n1565;
  assign n2286 = n1571 & n2285;
  assign n2287 = n1600 & n2286;
  assign n2288 = ~n2284 & ~n2287;
  assign n2289 = ~n1562 & ~n1598;
  assign n2290 = n2237 & n2289;
  assign n2291 = ~n1232 & n1598;
  assign n2292 = ~n1572 & n2291;
  assign n2293 = ~n2290 & ~n2292;
  assign n2294 = n2288 & n2293;
  assign n2295 = n1255 & ~n2294;
  assign n2296 = n1291 & ~n2294;
  assign n2297 = ~n1260 & n1277;
  assign n2298 = ~n2284 & n2297;
  assign n2299 = ~n2287 & ~n2290;
  assign n2300 = ~n2292 & n2299;
  assign n2301 = n2298 & n2300;
  assign n2302 = ~n2296 & ~n2301;
  assign n2303 = ~n2295 & n2302;
  assign n2304 = n2282 & n2303;
  assign n2305 = ~n2274 & n2304;
  assign n2306 = ~n2227 & ~n2305;
  assign n2307 = ~n2179 & n2224;
  assign n2308 = ~n2196 & ~n2209;
  assign n2309 = n2206 & n2308;
  assign n2310 = n2307 & n2309;
  assign n2311 = ~n2179 & ~n2199;
  assign n2312 = ~n2205 & ~n2209;
  assign n2313 = n2311 & n2312;
  assign n2314 = ~n2196 & ~n2224;
  assign n2315 = ~n2313 & n2314;
  assign n2316 = ~n2195 & ~n2218;
  assign n2317 = ~n2190 & n2316;
  assign n2318 = ~n2223 & n2317;
  assign n2319 = ~n2313 & n2318;
  assign n2320 = ~n2315 & ~n2319;
  assign n2321 = ~n2310 & n2320;
  assign n2322 = n2306 & n2321;
  assign n2323 = ~n1135 & ~n1288;
  assign n2324 = ~n1133 & n2323;
  assign n2325 = ~n2250 & n2324;
  assign n2326 = n2270 & n2325;
  assign n2327 = n2266 & n2326;
  assign n2328 = ~n1127 & n1137;
  assign n2329 = ~n1134 & n1288;
  assign n2330 = ~n2328 & n2329;
  assign n2331 = ~n2250 & n2330;
  assign n2332 = n2270 & n2331;
  assign n2333 = n2266 & n2332;
  assign n2334 = ~n1135 & n1288;
  assign n2335 = ~n1133 & n2334;
  assign n2336 = ~n2263 & n2335;
  assign n2337 = ~n2333 & ~n2336;
  assign n2338 = ~n2327 & n2337;
  assign n2339 = n1135 & ~n1306;
  assign n2340 = ~n1307 & n2339;
  assign n2341 = ~n1135 & ~n1308;
  assign n2342 = ~n2340 & ~n2341;
  assign n2343 = ~n1604 & ~n2342;
  assign n2344 = n1604 & n2342;
  assign n2345 = n621 & ~n625;
  assign n2346 = ~n639 & n2345;
  assign n2347 = ~n1125 & n2346;
  assign n2348 = ~n1123 & n2347;
  assign n2349 = ~n1133 & ~n2348;
  assign n2350 = ~n2344 & n2349;
  assign n2351 = ~n2343 & n2350;
  assign n2352 = ~n1132 & ~n1618;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~n2343 & ~n2344;
  assign n2355 = ~n1129 & n2345;
  assign n2356 = n1133 & ~n2355;
  assign n2357 = ~n2354 & n2356;
  assign n2358 = ~n1134 & ~n1288;
  assign n2359 = ~n2328 & n2358;
  assign n2360 = ~n2263 & n2359;
  assign n2361 = ~n2357 & ~n2360;
  assign n2362 = n2353 & n2361;
  assign n2363 = n2338 & n2362;
  assign n2364 = n2353 & ~n2357;
  assign n2365 = ~n2333 & ~n2360;
  assign n2366 = ~n2327 & ~n2336;
  assign n2367 = n2365 & n2366;
  assign n2368 = ~n2364 & ~n2367;
  assign n2369 = ~n2363 & ~n2368;
  assign n2370 = ~n2274 & n2303;
  assign n2371 = ~n2264 & ~n2282;
  assign n2372 = ~n2273 & n2371;
  assign n2373 = ~n2303 & n2372;
  assign n2374 = ~n2370 & ~n2373;
  assign n2375 = ~n2369 & n2374;
  assign n2376 = n2369 & ~n2374;
  assign n2377 = ~n2375 & ~n2376;
  assign n2378 = ~n1647 & ~n1651;
  assign n2379 = ~n1649 & n2378;
  assign n2380 = ~n1618 & ~n1620;
  assign n2381 = ~n1605 & n2380;
  assign n2382 = ~n1606 & n2381;
  assign n2383 = ~n1607 & n1621;
  assign n2384 = ~n1653 & ~n2383;
  assign n2385 = ~n2382 & n2384;
  assign n2386 = ~n2379 & n2385;
  assign n2387 = ~n2377 & n2386;
  assign n2388 = ~n2322 & n2387;
  assign n2389 = ~n2382 & ~n2383;
  assign n2390 = ~n1653 & ~n2389;
  assign n2391 = ~n2379 & n2390;
  assign n2392 = ~n2315 & n2391;
  assign n2393 = ~n2310 & ~n2319;
  assign n2394 = n2392 & n2393;
  assign n2395 = n2306 & n2394;
  assign n2396 = ~n2377 & n2395;
  assign n2397 = ~n2227 & ~n2315;
  assign n2398 = n2393 & n2397;
  assign n2399 = ~n2305 & n2385;
  assign n2400 = ~n2379 & n2399;
  assign n2401 = ~n2375 & n2400;
  assign n2402 = ~n2376 & n2401;
  assign n2403 = n2398 & n2402;
  assign n2404 = ~n2396 & ~n2403;
  assign n2405 = ~n2388 & n2404;
  assign n2406 = ~n1653 & ~n2379;
  assign n2407 = ~n2310 & ~n2406;
  assign n2408 = n2320 & n2407;
  assign n2409 = ~n2305 & ~n2389;
  assign n2410 = ~n2227 & n2409;
  assign n2411 = ~n2375 & n2410;
  assign n2412 = ~n2376 & n2411;
  assign n2413 = n2408 & n2412;
  assign n2414 = ~n1639 & n1661;
  assign n2415 = ~n1686 & ~n2414;
  assign n2416 = n1718 & n2415;
  assign n2417 = ~n2413 & n2416;
  assign n2418 = ~n2389 & ~n2406;
  assign n2419 = ~n2377 & n2418;
  assign n2420 = ~n2322 & n2419;
  assign n2421 = n2389 & ~n2406;
  assign n2422 = ~n2375 & n2421;
  assign n2423 = ~n2376 & n2422;
  assign n2424 = ~n2322 & n2423;
  assign n2425 = ~n2420 & ~n2424;
  assign n2426 = ~n2305 & n2389;
  assign n2427 = ~n2227 & n2426;
  assign n2428 = n2408 & n2427;
  assign n2429 = ~n2377 & n2428;
  assign n2430 = ~n2375 & n2391;
  assign n2431 = ~n2376 & n2430;
  assign n2432 = ~n2322 & n2431;
  assign n2433 = ~n2429 & ~n2432;
  assign n2434 = n2425 & n2433;
  assign n2435 = n2417 & n2434;
  assign n2436 = n2405 & n2435;
  assign n2437 = ~n2396 & ~n2432;
  assign n2438 = ~n2388 & ~n2403;
  assign n2439 = n2437 & n2438;
  assign n2440 = ~n2413 & ~n2420;
  assign n2441 = ~n2424 & ~n2429;
  assign n2442 = n2440 & n2441;
  assign n2443 = n2439 & n2442;
  assign n2444 = ~n2416 & ~n2443;
  assign n2445 = ~n2436 & ~n2444;
  assign n2446 = ~n1984 & ~n2445;
  assign n2447 = n1984 & ~n2436;
  assign n2448 = ~n2444 & n2447;
  assign n2449 = ~n2446 & ~n2448;
  assign n2450 = ~n1968 & ~n1971;
  assign n2451 = ~n1672 & n2450;
  assign n2452 = n1966 & ~n2451;
  assign n2453 = ~n1719 & n1975;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = ~n1976 & ~n2454;
  assign n2456 = ~n811 & ~n1964;
  assign n2457 = ~n2455 & n2456;
  assign n2458 = ~n1693 & ~n2457;
  assign n2459 = n787 & ~n811;
  assign n2460 = ~n1672 & n1708;
  assign n2461 = ~n1670 & n2460;
  assign n2462 = ~n1962 & n2461;
  assign n2463 = ~n1708 & ~n1960;
  assign n2464 = ~n1679 & n2463;
  assign n2465 = ~n1676 & ~n1708;
  assign n2466 = ~n1719 & n2465;
  assign n2467 = n1675 & ~n1705;
  assign n2468 = ~n1707 & n2467;
  assign n2469 = ~n1639 & n2468;
  assign n2470 = ~n1683 & n2469;
  assign n2471 = ~n1686 & n2470;
  assign n2472 = ~n1962 & n2471;
  assign n2473 = ~n2466 & ~n2472;
  assign n2474 = ~n2464 & n2473;
  assign n2475 = ~n2462 & n2474;
  assign n2476 = n1695 & ~n2475;
  assign n2477 = ~n2459 & ~n2476;
  assign n2478 = n2458 & ~n2477;
  assign n2479 = ~n1690 & n1722;
  assign n2480 = ~n1689 & n1727;
  assign n2481 = n1777 & ~n2480;
  assign n2482 = ~n2479 & n2481;
  assign n2483 = ~n1777 & n1782;
  assign n2484 = ~n1722 & n2483;
  assign n2485 = ~n1690 & n2484;
  assign n2486 = ~n1717 & n2483;
  assign n2487 = ~n1721 & n2486;
  assign n2488 = ~n1678 & n2487;
  assign n2489 = ~n1689 & n2488;
  assign n2490 = ~n2485 & ~n2489;
  assign n2491 = ~n1678 & n1787;
  assign n2492 = ~n1722 & n2491;
  assign n2493 = ~n1689 & n2492;
  assign n2494 = ~n1717 & n1787;
  assign n2495 = ~n1721 & n2494;
  assign n2496 = ~n1690 & n2495;
  assign n2497 = ~n2493 & ~n2496;
  assign n2498 = n2490 & n2497;
  assign n2499 = ~n2482 & n2498;
  assign n2500 = ~n2478 & n2499;
  assign n2501 = n811 & ~n2466;
  assign n2502 = ~n2472 & n2501;
  assign n2503 = ~n2464 & n2502;
  assign n2504 = ~n2462 & n2503;
  assign n2505 = ~n2458 & ~n2504;
  assign n2506 = ~n2500 & n2505;
  assign n2507 = ~n2449 & n2506;
  assign n2508 = ~n2446 & ~n2505;
  assign n2509 = ~n2448 & ~n2500;
  assign n2510 = n2508 & n2509;
  assign n2511 = ~n2507 & ~n2510;
  assign n2512 = ~n2493 & ~n2504;
  assign n2513 = ~n2496 & n2512;
  assign n2514 = ~n2482 & n2490;
  assign n2515 = n2513 & n2514;
  assign n2516 = ~n2458 & n2515;
  assign n2517 = ~n2478 & n2516;
  assign n2518 = n2449 & n2517;
  assign n2519 = n2500 & ~n2505;
  assign n2520 = ~n2449 & n2519;
  assign n2521 = ~n2518 & ~n2520;
  assign n2522 = n2511 & n2521;
  assign n2523 = ~n2479 & ~n2480;
  assign n2524 = ~n1777 & ~n2523;
  assign n2525 = ~n833 & ~n1782;
  assign n2526 = ~n1778 & n2525;
  assign n2527 = ~n2482 & n2526;
  assign n2528 = ~n2524 & n2527;
  assign n2529 = ~n2482 & ~n2524;
  assign n2530 = n1783 & ~n2529;
  assign n2531 = ~n1783 & ~n2482;
  assign n2532 = ~n2524 & n2531;
  assign n2533 = n1724 & ~n2532;
  assign n2534 = ~n2530 & n2533;
  assign n2535 = ~n2528 & ~n2534;
  assign n2536 = ~n2522 & n2535;
  assign n2537 = n1797 & ~n1817;
  assign n2538 = ~n1738 & n1790;
  assign n2539 = ~n1726 & ~n1790;
  assign n2540 = ~n1729 & ~n1734;
  assign n2541 = ~n1736 & n2540;
  assign n2542 = n2539 & n2541;
  assign n2543 = ~n2538 & ~n2542;
  assign n2544 = n1770 & ~n2543;
  assign n2545 = ~n1770 & ~n2538;
  assign n2546 = ~n2542 & n2545;
  assign n2547 = ~n1756 & ~n1761;
  assign n2548 = n864 & ~n2547;
  assign n2549 = ~n867 & ~n1763;
  assign n2550 = ~n2548 & n2549;
  assign n2551 = ~n2546 & n2550;
  assign n2552 = ~n2544 & n2551;
  assign n2553 = ~n2537 & ~n2552;
  assign n2554 = n858 & ~n1747;
  assign n2555 = ~n1751 & n2554;
  assign n2556 = n1759 & n2555;
  assign n2557 = ~n1739 & n2556;
  assign n2558 = ~n864 & ~n2557;
  assign n2559 = n1770 & ~n2558;
  assign n2560 = ~n2538 & ~n2559;
  assign n2561 = ~n2542 & n2560;
  assign n2562 = ~n853 & ~n864;
  assign n2563 = ~n856 & n2562;
  assign n2564 = ~n1755 & n2563;
  assign n2565 = ~n2561 & ~n2564;
  assign n2566 = ~n2553 & ~n2565;
  assign n2567 = ~n2536 & n2566;
  assign n2568 = n2521 & ~n2535;
  assign n2569 = n2511 & n2568;
  assign n2570 = n901 & ~n1833;
  assign n2571 = ~n1801 & ~n2570;
  assign n2572 = ~n1836 & n2571;
  assign n2573 = n1816 & ~n2572;
  assign n2574 = n1815 & n2573;
  assign n2575 = ~n900 & n908;
  assign n2576 = ~n1831 & n2575;
  assign n2577 = ~n1801 & ~n1836;
  assign n2578 = n2570 & ~n2577;
  assign n2579 = ~n2576 & ~n2578;
  assign n2580 = ~n2537 & n2579;
  assign n2581 = ~n2574 & n2580;
  assign n2582 = ~n943 & ~n1801;
  assign n2583 = ~n991 & n2582;
  assign n2584 = ~n1796 & n2583;
  assign n2585 = n1813 & n2584;
  assign n2586 = n900 & ~n943;
  assign n2587 = ~n1833 & n2586;
  assign n2588 = ~n1832 & n2587;
  assign n2589 = ~n943 & ~n1797;
  assign n2590 = ~n1800 & n2589;
  assign n2591 = ~n991 & n2590;
  assign n2592 = ~n1817 & n2591;
  assign n2593 = ~n2588 & ~n2592;
  assign n2594 = ~n2585 & n2593;
  assign n2595 = ~n2581 & n2594;
  assign n2596 = ~n2569 & ~n2595;
  assign n2597 = n2567 & n2596;
  assign n2598 = ~n2536 & ~n2569;
  assign n2599 = ~n2537 & ~n2565;
  assign n2600 = ~n2552 & n2599;
  assign n2601 = n2594 & n2600;
  assign n2602 = ~n2581 & n2601;
  assign n2603 = n2598 & n2602;
  assign n2604 = ~n2597 & ~n2603;
  assign n2605 = ~n2564 & ~n2588;
  assign n2606 = ~n2561 & n2605;
  assign n2607 = ~n2592 & n2606;
  assign n2608 = ~n2585 & n2607;
  assign n2609 = ~n2581 & n2608;
  assign n2610 = ~n2553 & n2609;
  assign n2611 = n2598 & n2610;
  assign n2612 = ~n2537 & n2565;
  assign n2613 = ~n2552 & n2612;
  assign n2614 = ~n2536 & n2613;
  assign n2615 = n2596 & n2614;
  assign n2616 = ~n2611 & ~n2615;
  assign n2617 = n2604 & n2616;
  assign n2618 = ~n2565 & ~n2585;
  assign n2619 = n2593 & n2618;
  assign n2620 = ~n2581 & n2619;
  assign n2621 = ~n2553 & n2620;
  assign n2622 = ~n2598 & n2621;
  assign n2623 = ~n2595 & n2600;
  assign n2624 = ~n2598 & n2623;
  assign n2625 = ~n2622 & ~n2624;
  assign n2626 = ~n2553 & n2565;
  assign n2627 = ~n2595 & n2626;
  assign n2628 = ~n2598 & n2627;
  assign n2629 = ~n2537 & n2606;
  assign n2630 = ~n2585 & ~n2592;
  assign n2631 = n2629 & n2630;
  assign n2632 = ~n2552 & n2631;
  assign n2633 = ~n2581 & n2632;
  assign n2634 = ~n2598 & n2633;
  assign n2635 = ~n2628 & ~n2634;
  assign n2636 = n2625 & n2635;
  assign n2637 = n2617 & n2636;
  assign n2638 = n1958 & ~n2637;
  assign n2639 = ~n1958 & n2637;
  assign n2640 = ~n1876 & ~n1934;
  assign n2641 = ~n1890 & ~n2640;
  assign n2642 = ~n2639 & ~n2641;
  assign n2643 = ~n2638 & n2642;
  assign n2644 = ~n2638 & ~n2639;
  assign n2645 = n2641 & ~n2644;
  assign n2646 = ~n2643 & ~n2645;
  assign n2647 = ~n1944 & ~n2646;
  assign n2648 = n1944 & ~n2641;
  assign n2649 = ~n2644 & n2648;
  assign n2650 = ~n1890 & ~n1936;
  assign n2651 = ~n1941 & n2650;
  assign n2652 = n1898 & ~n2640;
  assign n2653 = n2651 & n2652;
  assign n2654 = ~n1932 & n2653;
  assign n2655 = n2644 & n2654;
  assign n2656 = ~n2649 & ~n2655;
  assign n2657 = ~n2647 & n2656;
  assign n2658 = ~n1902 & ~n1905;
  assign n2659 = ~n1088 & ~n1900;
  assign n2660 = ~n2658 & ~n2659;
  assign n2661 = ~n2657 & ~n2660;
  assign n2662 = n2656 & n2660;
  assign n2663 = ~n2647 & n2662;
  assign n2664 = ~n2661 & ~n2663;
  assign n2665 = ~n1918 & n2664;
  assign n2666 = n1918 & ~n2664;
  assign po2 = ~n2665 & ~n2666;
  assign n2668 = n2656 & ~n2663;
  assign n2669 = ~n2665 & n2668;
  assign n2670 = ~n841 & ~n844;
  assign n2671 = ~n837 & n2670;
  assign n2672 = n887 & n2671;
  assign n2673 = ~n2532 & n2672;
  assign n2674 = ~n2530 & n2673;
  assign n2675 = ~n2507 & n2674;
  assign n2676 = ~n2510 & ~n2518;
  assign n2677 = ~n2520 & n2676;
  assign n2678 = n2675 & n2677;
  assign n2679 = ~n2507 & n2528;
  assign n2680 = n2677 & n2679;
  assign n2681 = ~n2678 & ~n2680;
  assign n2682 = ~n2115 & n2207;
  assign n2683 = ~n2116 & n2156;
  assign n2684 = ~n2177 & ~n2683;
  assign n2685 = ~n2682 & n2684;
  assign n2686 = ~n385 & ~n1173;
  assign n2687 = n1192 & n2686;
  assign n2688 = n1189 & n2687;
  assign n2689 = ~n2154 & n2688;
  assign n2690 = ~n2112 & n2689;
  assign n2691 = ~n2115 & n2690;
  assign n2692 = ~n2685 & ~n2691;
  assign n2693 = n2206 & ~n2209;
  assign n2694 = ~n536 & ~n579;
  assign n2695 = ~n1201 & n2694;
  assign n2696 = n1236 & n2695;
  assign n2697 = ~n1222 & n2696;
  assign n2698 = ~n1578 & n2697;
  assign n2699 = ~n2215 & n2698;
  assign n2700 = ~n2213 & n2699;
  assign n2701 = ~n2212 & n2700;
  assign n2702 = ~n2179 & ~n2701;
  assign n2703 = n2693 & n2702;
  assign n2704 = ~n579 & ~n1201;
  assign n2705 = n1236 & n2704;
  assign n2706 = ~n2184 & n2705;
  assign n2707 = ~n2185 & n2706;
  assign n2708 = n2224 & ~n2707;
  assign n2709 = ~n2703 & ~n2708;
  assign n2710 = n2692 & ~n2709;
  assign n2711 = ~n2692 & n2709;
  assign n2712 = ~n1540 & ~n2089;
  assign n2713 = n1540 & ~n2087;
  assign n2714 = ~n2088 & n2713;
  assign n2715 = n1510 & n1535;
  assign n2716 = ~n2714 & n2715;
  assign n2717 = ~n2712 & n2716;
  assign n2718 = ~n2085 & n2717;
  assign n2719 = ~n2712 & ~n2714;
  assign n2720 = n1535 & ~n2719;
  assign n2721 = ~n1535 & ~n2714;
  assign n2722 = ~n2712 & n2721;
  assign n2723 = ~n366 & ~n1506;
  assign n2724 = ~n1508 & n2723;
  assign n2725 = ~n2722 & n2724;
  assign n2726 = ~n2720 & n2725;
  assign n2727 = ~n2085 & n2092;
  assign n2728 = ~n2083 & n2712;
  assign n2729 = ~n2084 & n2728;
  assign n2730 = ~n2727 & ~n2729;
  assign n2731 = n2726 & ~n2730;
  assign n2732 = ~n2718 & ~n2731;
  assign n2733 = n2112 & ~n2726;
  assign n2734 = n390 & ~n2121;
  assign n2735 = ~n2123 & n2734;
  assign n2736 = ~n382 & ~n2125;
  assign n2737 = ~n2735 & n2736;
  assign n2738 = ~n2154 & n2737;
  assign n2739 = ~n2127 & ~n2738;
  assign n2740 = ~n2112 & ~n2739;
  assign n2741 = ~n2115 & n2740;
  assign n2742 = ~n2733 & ~n2741;
  assign n2743 = ~n2732 & n2742;
  assign n2744 = n2732 & ~n2742;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~n2073 & ~n2076;
  assign n2747 = ~n2080 & n2746;
  assign n2748 = ~n486 & ~n1328;
  assign n2749 = n486 & ~n1316;
  assign n2750 = n1488 & n2749;
  assign n2751 = ~n2748 & ~n2750;
  assign n2752 = ~n489 & ~n2751;
  assign n2753 = ~n2071 & ~n2752;
  assign n2754 = ~n1991 & n2753;
  assign n2755 = ~n1988 & ~n1989;
  assign n2756 = n1351 & ~n2755;
  assign n2757 = ~n2003 & ~n2756;
  assign n2758 = n2754 & n2757;
  assign n2759 = n2747 & n2758;
  assign n2760 = n1539 & ~n2089;
  assign n2761 = ~n2085 & n2760;
  assign n2762 = ~n2759 & ~n2761;
  assign n2763 = n2056 & ~n2064;
  assign n2764 = ~n2063 & n2763;
  assign n2765 = ~n2043 & n2764;
  assign n2766 = ~n2068 & ~n2765;
  assign n2767 = n2077 & n2766;
  assign n2768 = ~n2058 & n2060;
  assign n2769 = ~n2056 & ~n2768;
  assign n2770 = ~n2066 & n2769;
  assign n2771 = ~n2027 & ~n2770;
  assign n2772 = n2767 & n2771;
  assign n2773 = ~n2027 & n2078;
  assign n2774 = ~n2765 & ~n2770;
  assign n2775 = ~n2773 & ~n2774;
  assign n2776 = ~n2772 & ~n2775;
  assign n2777 = ~n473 & ~n1333;
  assign n2778 = n1994 & n2777;
  assign n2779 = ~n1329 & n2778;
  assign n2780 = ~n2755 & n2779;
  assign n2781 = n2041 & ~n2780;
  assign n2782 = ~n2028 & ~n2069;
  assign n2783 = ~n2773 & ~n2782;
  assign n2784 = ~n2781 & n2783;
  assign n2785 = n2776 & ~n2784;
  assign n2786 = ~n2776 & n2784;
  assign n2787 = ~n2752 & ~n2756;
  assign n2788 = ~n1991 & ~n2780;
  assign n2789 = n2082 & n2788;
  assign n2790 = ~n2787 & n2789;
  assign n2791 = ~n2786 & n2790;
  assign n2792 = ~n2785 & n2791;
  assign n2793 = ~n2785 & ~n2786;
  assign n2794 = ~n2790 & ~n2793;
  assign n2795 = ~n2792 & ~n2794;
  assign n2796 = ~n2762 & n2795;
  assign n2797 = n2762 & ~n2795;
  assign n2798 = ~n2796 & ~n2797;
  assign n2799 = n1537 & ~n2089;
  assign n2800 = ~n2722 & ~n2799;
  assign n2801 = ~n2085 & ~n2800;
  assign n2802 = ~n2798 & n2801;
  assign n2803 = ~n2796 & ~n2801;
  assign n2804 = ~n2797 & n2803;
  assign n2805 = ~n2802 & ~n2804;
  assign n2806 = ~n2745 & n2805;
  assign n2807 = n2745 & ~n2805;
  assign n2808 = ~n2806 & ~n2807;
  assign n2809 = ~n2711 & n2808;
  assign n2810 = ~n2710 & n2809;
  assign n2811 = ~n2710 & ~n2711;
  assign n2812 = ~n2808 & ~n2811;
  assign n2813 = ~n2810 & ~n2812;
  assign n2814 = ~n1289 & ~n2284;
  assign n2815 = n2300 & n2814;
  assign n2816 = n1289 & ~n2294;
  assign n2817 = ~n2815 & ~n2816;
  assign n2818 = ~n591 & ~n1243;
  assign n2819 = n1285 & n2818;
  assign n2820 = ~n2817 & n2819;
  assign n2821 = ~n2227 & n2820;
  assign n2822 = n2321 & n2821;
  assign n2823 = n2307 & n2693;
  assign n2824 = ~n2224 & ~n2313;
  assign n2825 = n2196 & ~n2707;
  assign n2826 = ~n2824 & n2825;
  assign n2827 = ~n2823 & n2826;
  assign n2828 = ~n2227 & n2295;
  assign n2829 = n2321 & n2828;
  assign n2830 = ~n2827 & ~n2829;
  assign n2831 = ~n2822 & n2830;
  assign n2832 = ~n2813 & n2831;
  assign n2833 = n2813 & ~n2831;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = ~n2302 & ~n2819;
  assign n2836 = ~n2282 & ~n2835;
  assign n2837 = ~n2227 & ~n2836;
  assign n2838 = n2321 & n2837;
  assign n2839 = n2303 & n2372;
  assign n2840 = ~n2227 & n2839;
  assign n2841 = n2321 & n2840;
  assign n2842 = n2373 & ~n2398;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = ~n2838 & n2843;
  assign n2845 = n2374 & ~n2398;
  assign n2846 = ~n2227 & ~n2282;
  assign n2847 = ~n2310 & ~n2374;
  assign n2848 = n2320 & n2847;
  assign n2849 = n2846 & n2848;
  assign n2850 = ~n2845 & ~n2849;
  assign n2851 = ~n637 & ~n2354;
  assign n2852 = ~n1133 & ~n2344;
  assign n2853 = ~n2343 & n2852;
  assign n2854 = ~n617 & ~n1127;
  assign n2855 = ~n1129 & n2854;
  assign n2856 = ~n2853 & n2855;
  assign n2857 = ~n2851 & n2856;
  assign n2858 = n1125 & ~n2264;
  assign n2859 = ~n2272 & n2858;
  assign n2860 = ~n633 & ~n1125;
  assign n2861 = ~n1123 & n2860;
  assign n2862 = ~n2344 & n2861;
  assign n2863 = ~n2343 & n2862;
  assign n2864 = ~n2853 & ~n2863;
  assign n2865 = ~n2859 & n2864;
  assign n2866 = ~n2857 & n2865;
  assign n2867 = ~n2859 & ~n2863;
  assign n2868 = ~n1133 & ~n2861;
  assign n2869 = ~n2344 & n2868;
  assign n2870 = ~n2343 & n2869;
  assign n2871 = n2857 & ~n2859;
  assign n2872 = ~n2870 & ~n2871;
  assign n2873 = ~n2867 & ~n2872;
  assign n2874 = ~n2866 & ~n2873;
  assign n2875 = ~n2850 & n2874;
  assign n2876 = ~n2844 & n2875;
  assign n2877 = ~n2834 & n2876;
  assign n2878 = n2844 & ~n2875;
  assign n2879 = ~n2834 & n2878;
  assign n2880 = ~n2877 & ~n2879;
  assign n2881 = ~n2841 & n2874;
  assign n2882 = ~n2838 & ~n2842;
  assign n2883 = n2881 & n2882;
  assign n2884 = ~n2850 & n2883;
  assign n2885 = ~n2832 & n2884;
  assign n2886 = ~n2833 & n2885;
  assign n2887 = ~n2844 & ~n2875;
  assign n2888 = ~n2832 & n2887;
  assign n2889 = ~n2833 & n2888;
  assign n2890 = ~n2886 & ~n2889;
  assign n2891 = n2880 & n2890;
  assign n2892 = ~n222 & ~n1661;
  assign n2893 = ~n1665 & n2892;
  assign n2894 = ~n1658 & n2893;
  assign n2895 = ~n2414 & ~n2894;
  assign n2896 = ~n2413 & ~n2895;
  assign n2897 = n2434 & n2896;
  assign n2898 = n2405 & n2897;
  assign n2899 = ~n2322 & ~n2377;
  assign n2900 = n2306 & ~n2375;
  assign n2901 = ~n2376 & n2900;
  assign n2902 = n2321 & n2901;
  assign n2903 = ~n2389 & ~n2902;
  assign n2904 = ~n2899 & n2903;
  assign n2905 = ~n2899 & ~n2902;
  assign n2906 = n2389 & ~n2905;
  assign n2907 = ~n1639 & n1642;
  assign n2908 = ~n2906 & n2907;
  assign n2909 = ~n2904 & n2908;
  assign n2910 = ~n2898 & ~n2909;
  assign n2911 = ~n2282 & ~n2374;
  assign n2912 = ~n2227 & n2367;
  assign n2913 = ~n2911 & n2912;
  assign n2914 = n2321 & n2913;
  assign n2915 = n2364 & ~n2857;
  assign n2916 = ~n2914 & n2915;
  assign n2917 = n2367 & ~n2374;
  assign n2918 = ~n2398 & n2917;
  assign n2919 = ~n2282 & ~n2367;
  assign n2920 = ~n2227 & n2919;
  assign n2921 = n2848 & n2920;
  assign n2922 = ~n2367 & ~n2370;
  assign n2923 = ~n2373 & n2922;
  assign n2924 = ~n2398 & n2923;
  assign n2925 = ~n2921 & ~n2924;
  assign n2926 = ~n2918 & n2925;
  assign n2927 = n2916 & n2926;
  assign n2928 = ~n1605 & n1616;
  assign n2929 = ~n1606 & n2928;
  assign n2930 = ~n1143 & ~n1619;
  assign n2931 = ~n1141 & n1619;
  assign n2932 = ~n1142 & n2931;
  assign n2933 = ~n2930 & ~n2932;
  assign n2934 = ~n2264 & ~n2933;
  assign n2935 = ~n2272 & n2934;
  assign n2936 = ~n2264 & ~n2272;
  assign n2937 = n2933 & ~n2936;
  assign n2938 = ~n2935 & ~n2937;
  assign n2939 = ~n697 & ~n700;
  assign n2940 = ~n2938 & n2939;
  assign n2941 = ~n2929 & ~n2940;
  assign n2942 = ~n2227 & n2369;
  assign n2943 = ~n2911 & n2942;
  assign n2944 = n2321 & n2943;
  assign n2945 = ~n2941 & ~n2944;
  assign n2946 = n2376 & ~n2398;
  assign n2947 = ~n2369 & n2847;
  assign n2948 = n2320 & n2846;
  assign n2949 = n2947 & n2948;
  assign n2950 = n2375 & ~n2398;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~n2946 & n2951;
  assign n2953 = n2945 & n2952;
  assign n2954 = ~n2927 & ~n2953;
  assign n2955 = ~n2389 & ~n2929;
  assign n2956 = ~n2940 & n2955;
  assign n2957 = ~n2902 & n2956;
  assign n2958 = ~n2899 & n2957;
  assign n2959 = ~n2944 & ~n2949;
  assign n2960 = ~n2946 & ~n2950;
  assign n2961 = n2959 & n2960;
  assign n2962 = ~n1631 & ~n1647;
  assign n2963 = ~n1649 & n2962;
  assign n2964 = ~n2389 & n2963;
  assign n2965 = ~n2961 & n2964;
  assign n2966 = ~n1649 & ~n2383;
  assign n2967 = ~n2382 & n2966;
  assign n2968 = n2962 & n2967;
  assign n2969 = ~n2944 & n2968;
  assign n2970 = n2952 & n2969;
  assign n2971 = ~n2965 & ~n2970;
  assign n2972 = ~n2958 & n2971;
  assign n2973 = ~n2954 & n2972;
  assign n2974 = ~n2910 & n2973;
  assign n2975 = ~n2891 & n2974;
  assign n2976 = n2954 & ~n2972;
  assign n2977 = ~n2910 & n2976;
  assign n2978 = ~n2891 & n2977;
  assign n2979 = ~n2975 & ~n2978;
  assign n2980 = ~n2879 & ~n2886;
  assign n2981 = ~n2889 & ~n2972;
  assign n2982 = n2980 & n2981;
  assign n2983 = ~n2877 & ~n2954;
  assign n2984 = ~n2910 & n2983;
  assign n2985 = n2982 & n2984;
  assign n2986 = n2954 & n2972;
  assign n2987 = ~n2910 & n2986;
  assign n2988 = n2891 & n2987;
  assign n2989 = ~n2985 & ~n2988;
  assign n2990 = n2979 & n2989;
  assign n2991 = ~n1639 & n1971;
  assign n2992 = ~n1659 & n2991;
  assign n2993 = ~n1960 & n2992;
  assign n2994 = ~n730 & ~n733;
  assign n2995 = ~n728 & n2994;
  assign n2996 = ~n1962 & n2995;
  assign n2997 = ~n2993 & n2996;
  assign n2998 = ~n1961 & n2997;
  assign n2999 = ~n1984 & ~n2998;
  assign n3000 = ~n2445 & n2999;
  assign n3001 = ~n2443 & n2895;
  assign n3002 = ~n2898 & n2998;
  assign n3003 = ~n3001 & n3002;
  assign n3004 = ~n1719 & n2895;
  assign n3005 = ~n2413 & n3004;
  assign n3006 = n2434 & n3005;
  assign n3007 = n2405 & n3006;
  assign n3008 = n2898 & ~n3007;
  assign n3009 = ~n3003 & n3008;
  assign n3010 = ~n3000 & n3009;
  assign n3011 = n2990 & n3010;
  assign n3012 = ~n3003 & ~n3007;
  assign n3013 = ~n3000 & n3012;
  assign n3014 = ~n2990 & ~n3013;
  assign n3015 = ~n3011 & ~n3014;
  assign n3016 = ~n2446 & n2505;
  assign n3017 = ~n2448 & n3016;
  assign n3018 = ~n2449 & ~n2505;
  assign n3019 = ~n790 & ~n1785;
  assign n3020 = ~n2480 & n3019;
  assign n3021 = ~n2479 & n3020;
  assign n3022 = ~n2478 & ~n3021;
  assign n3023 = ~n3018 & ~n3022;
  assign n3024 = ~n3017 & ~n3023;
  assign n3025 = n3015 & ~n3024;
  assign n3026 = n2890 & n2972;
  assign n3027 = n1624 & ~n1647;
  assign n3028 = ~n1649 & n3027;
  assign n3029 = ~n2907 & ~n3028;
  assign n3030 = ~n2906 & ~n3029;
  assign n3031 = ~n2904 & n3030;
  assign n3032 = ~n2954 & ~n3031;
  assign n3033 = n2880 & n3032;
  assign n3034 = n3026 & n3033;
  assign n3035 = n2890 & ~n2972;
  assign n3036 = ~n2954 & n3031;
  assign n3037 = n2880 & n3036;
  assign n3038 = n3035 & n3037;
  assign n3039 = ~n3034 & ~n3038;
  assign n3040 = ~n2904 & ~n2965;
  assign n3041 = ~n2958 & ~n2970;
  assign n3042 = n3040 & n3041;
  assign n3043 = n2954 & n3030;
  assign n3044 = n3042 & n3043;
  assign n3045 = n2891 & n3044;
  assign n3046 = ~n2889 & ~n3031;
  assign n3047 = ~n2972 & n3046;
  assign n3048 = ~n2877 & n2954;
  assign n3049 = n2980 & n3048;
  assign n3050 = n3047 & n3049;
  assign n3051 = ~n3045 & ~n3050;
  assign n3052 = n3039 & n3051;
  assign n3053 = ~n2972 & n3032;
  assign n3054 = ~n2891 & n3053;
  assign n3055 = ~n2954 & n3030;
  assign n3056 = n3042 & n3055;
  assign n3057 = ~n2891 & n3056;
  assign n3058 = ~n3054 & ~n3057;
  assign n3059 = n2954 & n3031;
  assign n3060 = ~n2972 & n3059;
  assign n3061 = ~n2891 & n3060;
  assign n3062 = n2986 & ~n3031;
  assign n3063 = ~n2891 & n3062;
  assign n3064 = ~n3061 & ~n3063;
  assign n3065 = n3058 & n3064;
  assign n3066 = n3052 & n3065;
  assign n3067 = ~n2898 & ~n3013;
  assign n3068 = ~n3066 & n3067;
  assign n3069 = n3013 & n3065;
  assign n3070 = n2990 & n3052;
  assign n3071 = n3069 & n3070;
  assign n3072 = ~n3068 & ~n3071;
  assign n3073 = n3025 & n3072;
  assign n3074 = ~n2681 & n3073;
  assign n3075 = ~n2478 & n2505;
  assign n3076 = ~n2446 & n3075;
  assign n3077 = ~n2448 & n3076;
  assign n3078 = ~n2478 & ~n2505;
  assign n3079 = ~n2449 & n3078;
  assign n3080 = ~n2498 & ~n3079;
  assign n3081 = ~n3077 & n3080;
  assign n3082 = n1777 & ~n3019;
  assign n3083 = ~n2480 & n3082;
  assign n3084 = ~n2479 & n3083;
  assign n3085 = ~n3018 & n3084;
  assign n3086 = ~n3017 & n3085;
  assign n3087 = ~n3081 & ~n3086;
  assign n3088 = n2681 & ~n3087;
  assign n3089 = n3073 & n3088;
  assign n3090 = n3015 & ~n3068;
  assign n3091 = ~n3071 & n3090;
  assign n3092 = ~n2681 & n3024;
  assign n3093 = ~n3091 & n3092;
  assign n3094 = ~n3089 & ~n3093;
  assign n3095 = ~n3074 & n3094;
  assign n3096 = ~n3024 & n3087;
  assign n3097 = n2681 & n3096;
  assign n3098 = ~n3091 & n3097;
  assign n3099 = ~n847 & ~n1747;
  assign n3100 = ~n1751 & n3099;
  assign n3101 = n1759 & n3100;
  assign n3102 = ~n1739 & n3101;
  assign n3103 = ~n2532 & n3102;
  assign n3104 = ~n2530 & n3103;
  assign n3105 = ~n2507 & n3104;
  assign n3106 = n2677 & n3105;
  assign n3107 = ~n853 & ~n1755;
  assign n3108 = ~n2538 & n3107;
  assign n3109 = ~n2542 & n3108;
  assign n3110 = ~n2536 & n3109;
  assign n3111 = ~n2569 & n3110;
  assign n3112 = ~n3106 & ~n3111;
  assign n3113 = ~n3098 & n3112;
  assign n3114 = ~n2678 & n3024;
  assign n3115 = ~n2680 & ~n3087;
  assign n3116 = n3114 & n3115;
  assign n3117 = ~n3091 & n3116;
  assign n3118 = ~n2678 & ~n3071;
  assign n3119 = ~n2680 & n3118;
  assign n3120 = ~n3014 & ~n3081;
  assign n3121 = ~n3086 & n3120;
  assign n3122 = ~n3011 & n3024;
  assign n3123 = ~n3068 & n3122;
  assign n3124 = n3121 & n3123;
  assign n3125 = n3119 & n3124;
  assign n3126 = ~n3117 & ~n3125;
  assign n3127 = n3113 & n3126;
  assign n3128 = n3095 & n3127;
  assign n3129 = ~n3098 & ~n3117;
  assign n3130 = ~n3089 & ~n3125;
  assign n3131 = n3129 & n3130;
  assign n3132 = ~n833 & ~n853;
  assign n3133 = ~n848 & n3132;
  assign n3134 = ~n849 & n3133;
  assign n3135 = ~n1782 & n3134;
  assign n3136 = ~n1778 & n3135;
  assign n3137 = ~n1779 & n3136;
  assign n3138 = ~n2482 & n3137;
  assign n3139 = ~n2524 & n3138;
  assign n3140 = ~n844 & ~n853;
  assign n3141 = ~n1754 & n3140;
  assign n3142 = ~n1778 & ~n1782;
  assign n3143 = n833 & ~n3142;
  assign n3144 = n3140 & ~n3143;
  assign n3145 = ~n1782 & n3132;
  assign n3146 = ~n1778 & n3145;
  assign n3147 = ~n3144 & ~n3146;
  assign n3148 = ~n1755 & ~n3147;
  assign n3149 = ~n2482 & n3148;
  assign n3150 = ~n2524 & n3149;
  assign n3151 = ~n3141 & ~n3150;
  assign n3152 = ~n3139 & n3151;
  assign n3153 = ~n2507 & ~n3152;
  assign n3154 = ~n2530 & ~n2532;
  assign n3155 = ~n2482 & n3136;
  assign n3156 = ~n2524 & n3155;
  assign n3157 = ~n3154 & ~n3156;
  assign n3158 = ~n2520 & ~n3157;
  assign n3159 = n2676 & n3158;
  assign n3160 = n3153 & n3159;
  assign n3161 = ~n3106 & ~n3160;
  assign n3162 = ~n3111 & n3161;
  assign n3163 = ~n3074 & ~n3093;
  assign n3164 = ~n3162 & n3163;
  assign n3165 = ~n3131 & n3164;
  assign n3166 = ~n3128 & ~n3165;
  assign n3167 = ~n2598 & n2600;
  assign n3168 = ~n2598 & n2626;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n2569 & n2614;
  assign n3171 = n2567 & ~n2569;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = n3169 & n3172;
  assign n3174 = ~n2581 & ~n2594;
  assign n3175 = ~n3173 & n3174;
  assign n3176 = ~n899 & ~n1833;
  assign n3177 = ~n1832 & n3176;
  assign n3178 = ~n1836 & ~n3177;
  assign n3179 = ~n1842 & n3178;
  assign n3180 = ~n3173 & n3179;
  assign n3181 = ~n3175 & ~n3180;
  assign n3182 = n2565 & ~n2598;
  assign n3183 = ~n2536 & ~n2565;
  assign n3184 = ~n2569 & n3183;
  assign n3185 = ~n3182 & ~n3184;
  assign n3186 = n2553 & ~n3185;
  assign n3187 = ~n2546 & ~n2565;
  assign n3188 = ~n2536 & n3187;
  assign n3189 = ~n2569 & n3188;
  assign n3190 = ~n856 & ~n2547;
  assign n3191 = ~n2538 & n3190;
  assign n3192 = ~n2542 & n3191;
  assign n3193 = ~n2536 & n3192;
  assign n3194 = ~n2569 & n3193;
  assign n3195 = ~n3189 & ~n3194;
  assign n3196 = ~n2536 & n2626;
  assign n3197 = ~n2569 & n3196;
  assign n3198 = n2566 & ~n2598;
  assign n3199 = ~n1817 & n1833;
  assign n3200 = ~n3177 & ~n3199;
  assign n3201 = ~n909 & ~n1796;
  assign n3202 = n1813 & n3201;
  assign n3203 = ~n2537 & ~n3202;
  assign n3204 = ~n3200 & n3203;
  assign n3205 = ~n3198 & ~n3204;
  assign n3206 = ~n3197 & n3205;
  assign n3207 = ~n3195 & ~n3206;
  assign n3208 = ~n3186 & n3207;
  assign n3209 = n3181 & n3208;
  assign n3210 = ~n3166 & n3209;
  assign n3211 = ~n3165 & ~n3181;
  assign n3212 = ~n3128 & n3208;
  assign n3213 = n3211 & n3212;
  assign n3214 = ~n3210 & ~n3213;
  assign n3215 = n3195 & ~n3206;
  assign n3216 = ~n3186 & n3215;
  assign n3217 = n3181 & n3216;
  assign n3218 = n3166 & n3217;
  assign n3219 = ~n3181 & n3216;
  assign n3220 = ~n3166 & n3219;
  assign n3221 = ~n3218 & ~n3220;
  assign n3222 = n3214 & n3221;
  assign n3223 = ~n3175 & ~n3195;
  assign n3224 = ~n3186 & ~n3206;
  assign n3225 = ~n3180 & ~n3224;
  assign n3226 = n3223 & n3225;
  assign n3227 = n3166 & n3226;
  assign n3228 = ~n3195 & ~n3224;
  assign n3229 = ~n3181 & n3228;
  assign n3230 = ~n3166 & n3229;
  assign n3231 = ~n3227 & ~n3230;
  assign n3232 = ~n3175 & n3195;
  assign n3233 = n3225 & n3232;
  assign n3234 = ~n3166 & n3233;
  assign n3235 = n3195 & ~n3224;
  assign n3236 = ~n3128 & n3235;
  assign n3237 = n3211 & n3236;
  assign n3238 = ~n3234 & ~n3237;
  assign n3239 = n3231 & n3238;
  assign n3240 = n3222 & n3239;
  assign n3241 = n1108 & ~n1864;
  assign n3242 = n1888 & n3241;
  assign n3243 = n1884 & n3242;
  assign n3244 = ~n2638 & n3243;
  assign n3245 = ~n2603 & ~n2611;
  assign n3246 = ~n2615 & n3245;
  assign n3247 = n1951 & ~n2622;
  assign n3248 = ~n2624 & ~n2628;
  assign n3249 = ~n2597 & ~n2634;
  assign n3250 = n3248 & n3249;
  assign n3251 = n3247 & n3250;
  assign n3252 = n3246 & n3251;
  assign n3253 = n3244 & ~n3252;
  assign n3254 = ~n3240 & n3253;
  assign n3255 = n2639 & ~n3240;
  assign n3256 = ~n3213 & ~n3218;
  assign n3257 = ~n3220 & n3256;
  assign n3258 = ~n2639 & ~n3244;
  assign n3259 = ~n3227 & n3258;
  assign n3260 = ~n3230 & ~n3234;
  assign n3261 = ~n3210 & ~n3237;
  assign n3262 = n3260 & n3261;
  assign n3263 = n3259 & n3262;
  assign n3264 = n3257 & n3263;
  assign n3265 = ~n3255 & ~n3264;
  assign n3266 = ~n3254 & n3265;
  assign n3267 = ~n1942 & ~n2639;
  assign n3268 = ~n2638 & n3267;
  assign n3269 = ~n1108 & n1113;
  assign n3270 = ~n1864 & n3269;
  assign n3271 = n1888 & n3270;
  assign n3272 = n1884 & n3271;
  assign n3273 = ~n2639 & n3272;
  assign n3274 = ~n2638 & n3273;
  assign n3275 = ~n3268 & ~n3274;
  assign n3276 = ~n3266 & n3275;
  assign n3277 = ~n3255 & ~n3275;
  assign n3278 = ~n3254 & ~n3264;
  assign n3279 = n3277 & n3278;
  assign n3280 = ~n3276 & ~n3279;
  assign n3281 = ~n2669 & n3280;
  assign n3282 = n2669 & ~n3280;
  assign po3 = ~n3281 & ~n3282;
  assign n3284 = ~n3038 & ~n3045;
  assign n3285 = ~n3050 & n3284;
  assign n3286 = n3007 & ~n3054;
  assign n3287 = ~n3057 & ~n3061;
  assign n3288 = ~n3034 & ~n3063;
  assign n3289 = n3287 & n3288;
  assign n3290 = n3286 & n3289;
  assign n3291 = n3285 & n3290;
  assign n3292 = n2982 & n3048;
  assign n3293 = ~n2906 & n3028;
  assign n3294 = ~n2904 & n3293;
  assign n3295 = ~n2954 & ~n2972;
  assign n3296 = ~n2891 & n3295;
  assign n3297 = ~n3294 & ~n3296;
  assign n3298 = ~n3292 & n3297;
  assign n3299 = ~n2891 & n2954;
  assign n3300 = ~n2889 & n2980;
  assign n3301 = n2983 & n3300;
  assign n3302 = ~n3299 & ~n3301;
  assign n3303 = n2972 & ~n3302;
  assign n3304 = ~n3298 & ~n3303;
  assign n3305 = n2990 & ~n3304;
  assign n3306 = ~n3291 & n3305;
  assign n3307 = ~n2850 & ~n2866;
  assign n3308 = ~n2844 & ~n3307;
  assign n3309 = ~n2832 & n3308;
  assign n3310 = ~n2833 & n3309;
  assign n3311 = n2844 & ~n3307;
  assign n3312 = ~n2834 & n3311;
  assign n3313 = n2929 & ~n2944;
  assign n3314 = n2952 & n3313;
  assign n3315 = ~n3312 & n3314;
  assign n3316 = ~n3310 & n3315;
  assign n3317 = n2367 & ~n2867;
  assign n3318 = n2364 & ~n3317;
  assign n3319 = ~n2914 & n3318;
  assign n3320 = n2926 & n3319;
  assign n3321 = ~n2844 & n3320;
  assign n3322 = ~n2834 & n3321;
  assign n3323 = ~n2841 & ~n2921;
  assign n3324 = ~n2918 & ~n2924;
  assign n3325 = n3323 & n3324;
  assign n3326 = n2882 & n3319;
  assign n3327 = n3325 & n3326;
  assign n3328 = ~n2832 & n3327;
  assign n3329 = ~n2833 & n3328;
  assign n3330 = ~n3322 & ~n3329;
  assign n3331 = n2363 & ~n2867;
  assign n3332 = ~n2841 & n3331;
  assign n3333 = n2882 & n3332;
  assign n3334 = ~n2850 & n3333;
  assign n3335 = ~n2834 & n3334;
  assign n3336 = ~n2850 & n3331;
  assign n3337 = ~n2844 & n3336;
  assign n3338 = ~n2832 & n3337;
  assign n3339 = ~n2833 & n3338;
  assign n3340 = ~n3335 & ~n3339;
  assign n3341 = n3330 & n3340;
  assign n3342 = ~n3316 & n3341;
  assign n3343 = n2940 & ~n2944;
  assign n3344 = n2952 & n3343;
  assign n3345 = ~n2877 & n3344;
  assign n3346 = n3300 & n3345;
  assign n3347 = ~n3342 & n3346;
  assign n3348 = n3342 & ~n3346;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = ~n2832 & ~n2844;
  assign n3351 = ~n2833 & n3350;
  assign n3352 = ~n2850 & ~n2867;
  assign n3353 = ~n2850 & n2853;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = ~n2834 & n2844;
  assign n3356 = ~n3354 & ~n3355;
  assign n3357 = ~n3351 & n3356;
  assign n3358 = ~n2832 & ~n2843;
  assign n3359 = ~n2833 & n3358;
  assign n3360 = ~n3357 & ~n3359;
  assign n3361 = ~n2822 & ~n2838;
  assign n3362 = n2295 & ~n3361;
  assign n3363 = n2813 & ~n3362;
  assign n3364 = ~n2730 & n2739;
  assign n3365 = ~n2112 & ~n3364;
  assign n3366 = n2726 & ~n3365;
  assign n3367 = ~n2744 & ~n3366;
  assign n3368 = n2805 & ~n3367;
  assign n3369 = ~n2732 & ~n2742;
  assign n3370 = ~n2805 & n3369;
  assign n3371 = ~n3368 & ~n3370;
  assign n3372 = n2718 & ~n2802;
  assign n3373 = ~n2804 & n3372;
  assign n3374 = n2712 & ~n2795;
  assign n3375 = n2722 & ~n2798;
  assign n3376 = ~n3374 & ~n3375;
  assign n3377 = ~n2085 & ~n3376;
  assign n3378 = ~n2759 & ~n2790;
  assign n3379 = ~n2793 & n3378;
  assign n3380 = ~n2041 & ~n2773;
  assign n3381 = ~n2782 & n3380;
  assign n3382 = n2776 & ~n3381;
  assign n3383 = ~n3379 & n3382;
  assign n3384 = n2017 & ~n2063;
  assign n3385 = ~n2765 & ~n3384;
  assign n3386 = ~n2770 & n3385;
  assign n3387 = ~n3382 & n3386;
  assign n3388 = n2056 & ~n3386;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3383 & n3389;
  assign n3391 = ~n3377 & n3390;
  assign n3392 = ~n3373 & n3391;
  assign n3393 = ~n3371 & n3392;
  assign n3394 = n3371 & ~n3392;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = ~n2710 & n2808;
  assign n3397 = ~n2711 & ~n3396;
  assign n3398 = n3395 & n3397;
  assign n3399 = n2830 & n3361;
  assign n3400 = ~n3395 & ~n3397;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~n3398 & n3401;
  assign n3403 = n3363 & n3402;
  assign n3404 = n3363 & ~n3399;
  assign n3405 = ~n3398 & ~n3400;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = ~n3403 & ~n3406;
  assign n3408 = ~n3360 & ~n3407;
  assign n3409 = ~n3359 & ~n3403;
  assign n3410 = ~n3406 & n3409;
  assign n3411 = ~n3357 & n3410;
  assign n3412 = ~n3408 & ~n3411;
  assign n3413 = ~n3349 & n3412;
  assign n3414 = n3349 & ~n3412;
  assign n3415 = ~n3413 & ~n3414;
  assign n3416 = n3306 & ~n3415;
  assign n3417 = ~n3306 & n3415;
  assign n3418 = n1964 & ~n2445;
  assign n3419 = ~n3054 & n3418;
  assign n3420 = n3289 & n3419;
  assign n3421 = n3285 & n3420;
  assign n3422 = ~n3417 & ~n3421;
  assign n3423 = ~n3416 & n3422;
  assign n3424 = ~n3416 & ~n3417;
  assign n3425 = n3421 & ~n3424;
  assign n3426 = ~n2446 & n2457;
  assign n3427 = ~n2448 & n3426;
  assign n3428 = ~n3091 & n3427;
  assign n3429 = ~n3425 & ~n3428;
  assign n3430 = ~n3423 & n3429;
  assign n3431 = ~n3423 & ~n3425;
  assign n3432 = n3428 & ~n3431;
  assign n3433 = n1693 & ~n2475;
  assign n3434 = ~n2446 & n3433;
  assign n3435 = ~n2448 & n3434;
  assign n3436 = ~n3091 & n3435;
  assign n3437 = ~n2898 & ~n3066;
  assign n3438 = ~n1964 & n1983;
  assign n3439 = ~n2445 & n3438;
  assign n3440 = ~n2975 & n3439;
  assign n3441 = ~n2978 & ~n2985;
  assign n3442 = ~n2988 & n3441;
  assign n3443 = n3440 & n3442;
  assign n3444 = ~n3437 & n3443;
  assign n3445 = ~n2446 & n2478;
  assign n3446 = ~n2448 & n3445;
  assign n3447 = ~n3091 & n3446;
  assign n3448 = ~n3444 & ~n3447;
  assign n3449 = ~n3436 & n3448;
  assign n3450 = n2482 & ~n3018;
  assign n3451 = ~n3017 & n3450;
  assign n3452 = ~n3091 & n3451;
  assign n3453 = ~n3449 & ~n3452;
  assign n3454 = ~n3432 & n3453;
  assign n3455 = ~n3430 & n3454;
  assign n3456 = ~n3112 & n3130;
  assign n3457 = n3129 & n3456;
  assign n3458 = ~n3098 & n3194;
  assign n3459 = n3126 & n3458;
  assign n3460 = n3095 & n3459;
  assign n3461 = n3024 & ~n3091;
  assign n3462 = ~n3073 & ~n3461;
  assign n3463 = n3081 & ~n3462;
  assign n3464 = ~n3162 & n3194;
  assign n3465 = n3163 & ~n3464;
  assign n3466 = ~n3463 & n3465;
  assign n3467 = ~n3460 & n3466;
  assign n3468 = ~n3457 & n3467;
  assign n3469 = ~n3455 & n3468;
  assign n3470 = ~n3444 & n3451;
  assign n3471 = ~n3091 & n3470;
  assign n3472 = ~n3447 & n3471;
  assign n3473 = ~n3436 & n3472;
  assign n3474 = ~n3432 & n3473;
  assign n3475 = ~n3430 & n3474;
  assign n3476 = ~n3430 & ~n3432;
  assign n3477 = ~n3436 & ~n3452;
  assign n3478 = n3448 & n3477;
  assign n3479 = ~n3476 & n3478;
  assign n3480 = ~n3449 & n3452;
  assign n3481 = ~n3476 & n3480;
  assign n3482 = ~n3479 & ~n3481;
  assign n3483 = ~n3475 & n3482;
  assign n3484 = n3469 & n3483;
  assign n3485 = ~n3455 & ~n3479;
  assign n3486 = ~n3475 & ~n3481;
  assign n3487 = n3485 & n3486;
  assign n3488 = ~n3468 & ~n3487;
  assign n3489 = ~n3484 & ~n3488;
  assign n3490 = ~n3189 & ~n3198;
  assign n3491 = ~n3197 & n3490;
  assign n3492 = ~n3166 & ~n3491;
  assign n3493 = ~n3166 & n3194;
  assign n3494 = ~n856 & ~n2564;
  assign n3495 = ~n2547 & n3494;
  assign n3496 = ~n2538 & n3495;
  assign n3497 = ~n2542 & n3496;
  assign n3498 = ~n2561 & n3497;
  assign n3499 = ~n2536 & n3498;
  assign n3500 = ~n2569 & n3499;
  assign n3501 = ~n3128 & ~n3500;
  assign n3502 = ~n3165 & n3501;
  assign n3503 = ~n3182 & n3199;
  assign n3504 = ~n3184 & n3503;
  assign n3505 = ~n3502 & n3504;
  assign n3506 = ~n3493 & n3505;
  assign n3507 = ~n3492 & ~n3506;
  assign n3508 = ~n3489 & n3507;
  assign n3509 = n3489 & ~n3507;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = n1947 & ~n3173;
  assign n3512 = ~n3166 & n3511;
  assign n3513 = ~n3128 & n3195;
  assign n3514 = ~n3165 & n3513;
  assign n3515 = ~n3166 & ~n3195;
  assign n3516 = ~n3224 & ~n3515;
  assign n3517 = ~n3514 & n3516;
  assign n3518 = ~n3514 & ~n3515;
  assign n3519 = n3224 & ~n3518;
  assign n3520 = ~n3517 & ~n3519;
  assign n3521 = n3175 & ~n3520;
  assign n3522 = ~n3512 & ~n3521;
  assign n3523 = n1828 & ~n1955;
  assign n3524 = ~n1953 & n3523;
  assign n3525 = n2636 & n3524;
  assign n3526 = n2617 & n3525;
  assign n3527 = ~n3240 & n3526;
  assign n3528 = ~n3240 & n3252;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530 = n3522 & n3529;
  assign n3531 = n3510 & ~n3530;
  assign n3532 = ~n3510 & n3530;
  assign n3533 = ~n1951 & ~n2622;
  assign n3534 = ~n3524 & n3533;
  assign n3535 = n3250 & n3534;
  assign n3536 = ~n1958 & n3246;
  assign n3537 = n3535 & n3536;
  assign n3538 = ~n3240 & n3537;
  assign n3539 = n2656 & ~n3268;
  assign n3540 = n3274 & ~n3539;
  assign n3541 = n2656 & n3275;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = ~n3254 & ~n3542;
  assign n3544 = n3265 & ~n3543;
  assign n3545 = ~n3538 & ~n3544;
  assign n3546 = ~n3532 & n3545;
  assign n3547 = ~n3531 & n3546;
  assign n3548 = ~n3531 & ~n3532;
  assign n3549 = n3537 & ~n3539;
  assign n3550 = ~n3240 & n3549;
  assign n3551 = ~n3255 & n3550;
  assign n3552 = n3278 & n3551;
  assign n3553 = ~n3545 & ~n3552;
  assign n3554 = ~n3548 & n3553;
  assign n3555 = ~n3547 & ~n3554;
  assign n3556 = ~n1917 & ~n2660;
  assign n3557 = ~n1914 & n3556;
  assign n3558 = n2657 & ~n3557;
  assign n3559 = ~n3279 & n3558;
  assign n3560 = ~n3276 & n3559;
  assign n3561 = ~n3555 & n3560;
  assign n3562 = ~n3547 & ~n3560;
  assign n3563 = ~n3554 & n3562;
  assign po4 = n3561 | n3563;
  assign n3565 = ~n3254 & ~n3274;
  assign n3566 = n3265 & ~n3565;
  assign n3567 = ~n3548 & n3566;
  assign n3568 = n1900 & ~n2649;
  assign n3569 = ~n2655 & n3568;
  assign n3570 = ~n2647 & n3569;
  assign n3571 = ~n3279 & n3570;
  assign n3572 = ~n3276 & n3571;
  assign n3573 = ~n3255 & ~n3539;
  assign n3574 = n3278 & n3573;
  assign n3575 = ~n3572 & ~n3574;
  assign n3576 = ~n3567 & n3575;
  assign n3577 = n3538 & ~n3548;
  assign n3578 = ~n3538 & ~n3566;
  assign n3579 = ~n3532 & n3578;
  assign n3580 = ~n3531 & n3579;
  assign n3581 = ~n3577 & ~n3580;
  assign n3582 = ~n3576 & n3581;
  assign n3583 = n1911 & ~n2647;
  assign n3584 = n1101 & n2656;
  assign n3585 = ~n1095 & n3584;
  assign n3586 = ~n3556 & n3585;
  assign n3587 = n3583 & n3586;
  assign n3588 = ~n3279 & n3587;
  assign n3589 = ~n3276 & n3588;
  assign n3590 = ~n3555 & ~n3589;
  assign n3591 = ~n1102 & ~n1909;
  assign n3592 = ~n1910 & n2657;
  assign n3593 = ~n3591 & n3592;
  assign n3594 = ~n3279 & n3593;
  assign n3595 = ~n3276 & n3594;
  assign n3596 = ~n3547 & ~n3595;
  assign n3597 = ~n3554 & n3596;
  assign n3598 = ~n3590 & ~n3597;
  assign n3599 = ~n3582 & n3598;
  assign n3600 = ~n3087 & ~n3462;
  assign n3601 = ~n3073 & n3087;
  assign n3602 = ~n3461 & n3601;
  assign n3603 = n2680 & ~n3602;
  assign n3604 = ~n3600 & n3603;
  assign n3605 = ~n3455 & n3604;
  assign n3606 = n3483 & n3605;
  assign n3607 = n3449 & ~n3476;
  assign n3608 = ~n3432 & ~n3449;
  assign n3609 = ~n3430 & n3608;
  assign n3610 = n3600 & ~n3609;
  assign n3611 = ~n3607 & n3610;
  assign n3612 = ~n3606 & ~n3611;
  assign n3613 = n3129 & n3163;
  assign n3614 = n3456 & n3613;
  assign n3615 = n2678 & ~n3462;
  assign n3616 = ~n3464 & ~n3615;
  assign n3617 = ~n3460 & n3616;
  assign n3618 = ~n3614 & n3617;
  assign n3619 = n3486 & ~n3618;
  assign n3620 = n3485 & n3619;
  assign n3621 = ~n3612 & ~n3620;
  assign n3622 = n3612 & n3620;
  assign n3623 = ~n3621 & ~n3622;
  assign n3624 = ~n3348 & ~n3412;
  assign n3625 = n2813 & ~n2830;
  assign n3626 = ~n3405 & n3625;
  assign n3627 = ~n2810 & n2827;
  assign n3628 = ~n2812 & n3627;
  assign n3629 = ~n3406 & ~n3628;
  assign n3630 = ~n3626 & ~n3629;
  assign n3631 = ~n3411 & ~n3630;
  assign n3632 = ~n3395 & n3397;
  assign n3633 = ~n3628 & n3632;
  assign n3634 = ~n3370 & ~n3373;
  assign n3635 = n3391 & n3634;
  assign n3636 = ~n3368 & n3635;
  assign n3637 = ~n3633 & ~n3636;
  assign n3638 = ~n3347 & ~n3637;
  assign n3639 = ~n3631 & n3638;
  assign n3640 = ~n3624 & n3639;
  assign n3641 = ~n3417 & n3640;
  assign n3642 = ~n3421 & ~n3444;
  assign n3643 = ~n3416 & ~n3642;
  assign n3644 = n3641 & n3643;
  assign n3645 = n3424 & ~n3642;
  assign n3646 = n3415 & ~n3640;
  assign n3647 = ~n3306 & n3646;
  assign n3648 = ~n3641 & ~n3647;
  assign n3649 = ~n3645 & n3648;
  assign n3650 = ~n3644 & ~n3649;
  assign n3651 = ~n3432 & ~n3436;
  assign n3652 = ~n3430 & ~n3651;
  assign n3653 = ~n3650 & ~n3652;
  assign n3654 = ~n3430 & n3650;
  assign n3655 = ~n3651 & n3654;
  assign n3656 = ~n3653 & ~n3655;
  assign n3657 = ~n3432 & n3447;
  assign n3658 = ~n3430 & n3657;
  assign n3659 = ~n3018 & n3021;
  assign n3660 = ~n3017 & n3659;
  assign n3661 = ~n3091 & n3660;
  assign n3662 = ~n3609 & n3661;
  assign n3663 = ~n3607 & n3662;
  assign n3664 = ~n3658 & ~n3663;
  assign n3665 = ~n3656 & n3664;
  assign n3666 = n3656 & ~n3664;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = ~n3182 & ~n3194;
  assign n3669 = ~n3184 & n3668;
  assign n3670 = ~n3166 & ~n3669;
  assign n3671 = n2552 & ~n3670;
  assign n3672 = ~n3166 & n3189;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = ~n3502 & ~n3673;
  assign n3675 = ~n3489 & n3674;
  assign n3676 = ~n3667 & n3675;
  assign n3677 = ~n3623 & n3676;
  assign n3678 = ~n3667 & ~n3675;
  assign n3679 = n3623 & n3678;
  assign n3680 = ~n3677 & ~n3679;
  assign n3681 = n3667 & n3675;
  assign n3682 = n3623 & n3681;
  assign n3683 = n3667 & ~n3675;
  assign n3684 = ~n3623 & n3683;
  assign n3685 = ~n3682 & ~n3684;
  assign n3686 = n3680 & n3685;
  assign n3687 = n1833 & ~n1836;
  assign n3688 = ~n1817 & n3687;
  assign n3689 = ~n2537 & n3688;
  assign n3690 = ~n1842 & n3689;
  assign n3691 = ~n2552 & n3690;
  assign n3692 = ~n3194 & n3691;
  assign n3693 = n3185 & n3692;
  assign n3694 = ~n3166 & n3693;
  assign n3695 = ~n3506 & ~n3694;
  assign n3696 = ~n3484 & n3492;
  assign n3697 = ~n3488 & n3696;
  assign n3698 = ~n3489 & ~n3492;
  assign n3699 = n1955 & ~n3504;
  assign n3700 = ~n902 & ~n948;
  assign n3701 = ~n908 & ~n947;
  assign n3702 = ~n3700 & n3701;
  assign n3703 = ~n1799 & n3702;
  assign n3704 = ~n1797 & n3703;
  assign n3705 = ~n1836 & n3704;
  assign n3706 = ~n1817 & n3705;
  assign n3707 = ~n2553 & n3706;
  assign n3708 = ~n3185 & n3707;
  assign n3709 = ~n3699 & ~n3708;
  assign n3710 = ~n3185 & n3706;
  assign n3711 = n3173 & ~n3710;
  assign n3712 = ~n3709 & ~n3711;
  assign n3713 = ~n3520 & n3712;
  assign n3714 = ~n3694 & ~n3713;
  assign n3715 = ~n3698 & n3714;
  assign n3716 = ~n3697 & n3715;
  assign n3717 = ~n3695 & ~n3716;
  assign n3718 = ~n3512 & ~n3713;
  assign n3719 = ~n3697 & ~n3698;
  assign n3720 = ~n3718 & ~n3719;
  assign n3721 = n2537 & ~n3182;
  assign n3722 = ~n3184 & n3721;
  assign n3723 = ~n3502 & n3722;
  assign n3724 = ~n3493 & n3723;
  assign n3725 = ~n3698 & n3724;
  assign n3726 = ~n3697 & n3725;
  assign n3727 = ~n3720 & ~n3726;
  assign n3728 = ~n3717 & n3727;
  assign n3729 = ~n3686 & n3728;
  assign n3730 = n3686 & ~n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~n3508 & n3718;
  assign n3733 = ~n3509 & n3732;
  assign n3734 = n3527 & ~n3733;
  assign n3735 = ~n3577 & ~n3734;
  assign n3736 = ~n3731 & n3735;
  assign n3737 = n3731 & ~n3735;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = n3599 & n3738;
  assign n3740 = n3582 & ~n3736;
  assign n3741 = ~n3598 & ~n3737;
  assign n3742 = n3740 & n3741;
  assign n3743 = ~n3739 & ~n3742;
  assign n3744 = n3582 & ~n3590;
  assign n3745 = ~n3597 & n3744;
  assign n3746 = ~n3738 & n3745;
  assign n3747 = ~n3582 & ~n3598;
  assign n3748 = ~n3738 & n3747;
  assign n3749 = ~n3746 & ~n3748;
  assign po5 = ~n3743 | ~n3749;
  assign n3751 = ~n1918 & n2657;
  assign n3752 = ~n3279 & n3751;
  assign n3753 = ~n3276 & n3752;
  assign n3754 = ~n3577 & n3753;
  assign n3755 = ~n3580 & n3754;
  assign n3756 = ~n3576 & n3755;
  assign n3757 = ~n3590 & n3756;
  assign n3758 = n3738 & n3757;
  assign n3759 = n3254 & ~n3548;
  assign n3760 = n3735 & ~n3759;
  assign n3761 = ~n3731 & ~n3760;
  assign n3762 = ~n3717 & ~n3720;
  assign n3763 = ~n3686 & ~n3762;
  assign n3764 = ~n3614 & ~n3615;
  assign n3765 = ~n3455 & ~n3764;
  assign n3766 = n3483 & n3765;
  assign n3767 = n3612 & ~n3766;
  assign n3768 = n3667 & n3767;
  assign n3769 = n3189 & ~n3489;
  assign n3770 = ~n3189 & ~n3484;
  assign n3771 = ~n3488 & n3770;
  assign n3772 = ~n3769 & ~n3771;
  assign n3773 = n3515 & ~n3772;
  assign n3774 = ~n3768 & n3773;
  assign n3775 = ~n3197 & ~n3198;
  assign n3776 = ~n3166 & ~n3775;
  assign n3777 = ~n3489 & n3776;
  assign n3778 = n3667 & n3777;
  assign n3779 = ~n3623 & n3778;
  assign n3780 = ~n3656 & n3663;
  assign n3781 = ~n3652 & ~n3658;
  assign n3782 = ~n3645 & ~n3648;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = ~n3417 & ~n3640;
  assign n3785 = n3643 & n3784;
  assign n3786 = ~n3304 & ~n3415;
  assign n3787 = n2990 & ~n3291;
  assign n3788 = ~n3640 & ~n3787;
  assign n3789 = ~n3786 & n3788;
  assign n3790 = ~n3785 & ~n3789;
  assign n3791 = ~n3783 & n3790;
  assign n3792 = ~n3780 & n3791;
  assign n3793 = ~n3779 & n3792;
  assign n3794 = n3612 & ~n3665;
  assign n3795 = ~n3666 & n3794;
  assign n3796 = n3766 & ~n3795;
  assign n3797 = n3612 & ~n3777;
  assign n3798 = ~n3622 & ~n3667;
  assign n3799 = ~n3797 & n3798;
  assign n3800 = ~n3796 & ~n3799;
  assign n3801 = n3793 & n3800;
  assign n3802 = ~n3774 & n3801;
  assign n3803 = ~n3763 & n3802;
  assign n3804 = ~n3761 & n3803;
  assign n3805 = ~n3758 & n3804;
  assign n3806 = ~n3590 & n3753;
  assign n3807 = ~n3582 & n3806;
  assign n3808 = ~n3738 & n3807;
  assign n3809 = ~n3279 & n3566;
  assign n3810 = ~n3548 & n3809;
  assign n3811 = n2663 & ~n3279;
  assign n3812 = ~n3276 & n3811;
  assign n3813 = ~n3574 & ~n3812;
  assign n3814 = n3581 & ~n3813;
  assign n3815 = ~n3567 & ~n3814;
  assign n3816 = ~n3810 & ~n3815;
  assign n3817 = ~n3738 & n3816;
  assign n3818 = ~n3808 & ~n3817;
  assign po6 = ~n3805 | ~n3818;
endmodule


