// Benchmark "i2c" written by ABC on Wed Apr 29 13:48:26 2015

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n473,
    n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n486,
    n487, n488, n489, n490, n491, n492, n494, n495, n496, n497, n498, n499,
    n501, n502, n503, n504, n505, n506, n507, n509, n510, n511, n512, n513,
    n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
    n528, n529, n530, n531, n532, n533, n534, n536, n537, n538, n539, n540,
    n541, n542, n543, n545, n546, n547, n548, n549, n550, n551, n552, n553,
    n554, n556, n557, n558, n559, n560, n561, n563, n564, n565, n566, n567,
    n568, n569, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n601, n602, n603, n604, n605, n606,
    n608, n609, n610, n611, n612, n613, n615, n616, n617, n618, n619, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n638, n639, n640, n642, n643, n644, n645, n646, n647,
    n649, n650, n652, n653, n654, n655, n656, n657, n658, n659, n660, n662,
    n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
    n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705, n706, n707, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n764, n765, n766, n767, n768, n769, n771, n772, n773, n774, n775, n776,
    n778, n779, n780, n781, n782, n783, n785, n786, n787, n788, n789, n790,
    n792, n793, n794, n795, n796, n797, n799, n800, n801, n802, n803, n804,
    n806, n807, n808, n809, n810, n811, n813, n814, n815, n816, n817, n818,
    n820, n821, n822, n823, n824, n825, n826, n827, n829, n830, n831, n832,
    n833, n834, n835, n836, n838, n839, n840, n841, n842, n843, n844, n845,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n857, n858, n859,
    n860, n861, n862, n863, n864, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n876, n877, n878, n879, n880, n881, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n903, n904, n905, n906, n907, n908, n909, n910, n911, n913,
    n914, n915, n916, n917, n918, n919, n920, n921, n923, n924, n925, n926,
    n927, n928, n929, n930, n931, n932, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n944, n945, n946, n947, n949, n950, n951, n952, n953,
    n954, n956, n957, n958, n959, n960, n961, n963, n965, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n992, n993, n994, n995, n996,
    n997, n998, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
    n1008, n1010, n1011, n1012, n1014, n1015, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1031,
    n1032, n1033, n1034, n1035, n1036, n1038, n1039, n1040, n1041, n1042,
    n1043, n1045, n1046, n1047, n1048, n1049, n1050, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1060, n1061, n1062, n1063, n1064, n1065,
    n1067, n1068, n1069, n1070, n1071, n1072, n1074, n1075, n1076, n1077,
    n1078, n1079, n1081, n1082, n1083, n1084, n1085, n1086, n1088, n1089,
    n1090, n1091, n1092, n1093, n1095, n1096, n1097, n1098, n1099, n1100,
    n1102, n1103, n1104, n1105, n1106, n1107, n1109, n1110, n1111, n1112,
    n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1123, n1124,
    n1125, n1126, n1127, n1128, n1130, n1131, n1132, n1133, n1134, n1135,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1146, n1147,
    n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158,
    n1160, n1161, n1162, n1163, n1164, n1165, n1167, n1168, n1169, n1170,
    n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
    n1193, n1194, n1195, n1196, n1197, n1198, n1200, n1201, n1202, n1203,
    n1204, n1205, n1207, n1208, n1209, n1210, n1211, n1212, n1214, n1215,
    n1216, n1217, n1218, n1219, n1221, n1222, n1223, n1224, n1225, n1226,
    n1228, n1229, n1230, n1231, n1232, n1233, n1235, n1236, n1237, n1238,
    n1239, n1240, n1242, n1243, n1244, n1245, n1246, n1247, n1249, n1250,
    n1251, n1252, n1253, n1254, n1256, n1257, n1258, n1259, n1260, n1261,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1272, n1273,
    n1274, n1275, n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284,
    n1285, n1286, n1288, n1289, n1290, n1291, n1292, n1293, n1295, n1296,
    n1297, n1298, n1299, n1300, n1302, n1303, n1304, n1305, n1306, n1307,
    n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1375, n1376, n1377, n1378, n1379, n1380, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
    n1408, n1409, n1410, n1412, n1413, n1414, n1415, n1417, n1418, n1419,
    n1420, n1422, n1423, n1424, n1426, n1427, n1429, n1430, n1431, n1433,
    n1434, n1435, n1438, n1439, n1440, n1442, n1444, n1445, n1447, n1452,
    n1453, n1455;
  assign n291 = ~pi000 & ~pi054;
  assign n292 = ~pi005 & ~pi022;
  assign n293 = pi056 & ~n292;
  assign n294 = ~pi009 & ~pi011;
  assign n295 = ~pi005 & ~pi012;
  assign n296 = ~pi011 & n295;
  assign n297 = ~pi017 & ~pi018;
  assign n298 = ~pi016 & n297;
  assign n299 = ~pi013 & ~pi014;
  assign n300 = ~pi007 & n299;
  assign n301 = ~pi008 & n300;
  assign n302 = ~pi004 & ~pi006;
  assign n303 = ~pi010 & n302;
  assign n304 = ~pi019 & ~pi021;
  assign n305 = n303 & n304;
  assign n306 = n301 & n305;
  assign n307 = n298 & n306;
  assign n308 = n296 & n307;
  assign n309 = n294 & ~n308;
  assign n310 = n293 & n309;
  assign n311 = n294 & n308;
  assign n312 = pi000 & n292;
  assign n313 = ~n293 & ~n312;
  assign n314 = n311 & ~n313;
  assign n315 = ~n310 & ~n314;
  assign n316 = n292 & ~n294;
  assign n317 = pi056 & n316;
  assign n318 = n308 & n317;
  assign n319 = ~n308 & n317;
  assign n320 = pi054 & ~n319;
  assign n321 = ~n318 & n320;
  assign n322 = n315 & n321;
  assign n323 = ~pi017 & ~pi019;
  assign n324 = ~pi009 & ~pi022;
  assign n325 = ~pi011 & n324;
  assign n326 = ~pi010 & ~pi014;
  assign n327 = ~pi016 & ~pi018;
  assign n328 = n295 & n327;
  assign n329 = n326 & n328;
  assign n330 = n325 & n329;
  assign n331 = n302 & n330;
  assign n332 = ~pi007 & ~pi013;
  assign n333 = ~pi021 & n332;
  assign n334 = n331 & n333;
  assign n335 = ~pi008 & ~pi021;
  assign n336 = ~pi013 & n335;
  assign n337 = n331 & n336;
  assign n338 = ~n334 & ~n337;
  assign n339 = n325 & n328;
  assign n340 = n302 & n339;
  assign n341 = ~pi007 & n340;
  assign n342 = pi013 & pi014;
  assign n343 = ~pi010 & ~n342;
  assign n344 = ~n299 & ~n343;
  assign n345 = n341 & ~n344;
  assign n346 = n335 & n345;
  assign n347 = n338 & ~n346;
  assign n348 = n323 & ~n347;
  assign n349 = ~n292 & ~n294;
  assign n350 = n292 & n294;
  assign n351 = ~n349 & ~n350;
  assign n352 = ~n311 & ~n351;
  assign n353 = ~pi008 & ~pi019;
  assign n354 = n331 & n332;
  assign n355 = n353 & n354;
  assign n356 = ~pi017 & n355;
  assign n357 = n352 & ~n356;
  assign n358 = ~n348 & n357;
  assign n359 = n322 & ~n358;
  assign n360 = ~n291 & ~n359;
  assign n361 = ~pi003 & ~pi129;
  assign po015 = n360 | ~n361;
  assign n363 = pi001 & pi054;
  assign n364 = pi017 & n363;
  assign n365 = ~pi014 & n303;
  assign n366 = ~pi012 & ~pi018;
  assign n367 = ~pi016 & n304;
  assign n368 = ~pi013 & n367;
  assign n369 = ~pi011 & ~pi022;
  assign n370 = ~pi009 & n369;
  assign n371 = ~pi005 & n370;
  assign n372 = ~pi008 & ~pi017;
  assign n373 = ~pi007 & n372;
  assign n374 = n371 & n373;
  assign n375 = n368 & n374;
  assign n376 = n366 & n375;
  assign n377 = n365 & n376;
  assign n378 = n364 & ~n377;
  assign n379 = pi017 & n377;
  assign n380 = ~pi017 & ~n377;
  assign n381 = ~n379 & ~n380;
  assign n382 = pi054 & ~n381;
  assign n383 = ~n378 & ~n382;
  assign n384 = ~pi004 & ~pi010;
  assign n385 = n299 & n384;
  assign n386 = ~pi005 & ~pi011;
  assign n387 = ~pi022 & n386;
  assign n388 = ~n325 & ~n387;
  assign n389 = ~pi012 & ~n388;
  assign n390 = ~n371 & ~n389;
  assign n391 = ~pi006 & n327;
  assign n392 = ~n390 & n391;
  assign n393 = n385 & n392;
  assign n394 = ~pi005 & n369;
  assign n395 = ~pi009 & ~pi016;
  assign n396 = n366 & n395;
  assign n397 = n394 & n396;
  assign n398 = ~pi013 & n365;
  assign n399 = ~n365 & ~n385;
  assign n400 = ~n398 & n399;
  assign n401 = n397 & ~n400;
  assign n402 = ~n393 & ~n401;
  assign n403 = n397 & n398;
  assign n404 = pi007 & ~n403;
  assign n405 = ~n402 & ~n404;
  assign n406 = n323 & n335;
  assign n407 = ~n378 & n406;
  assign n408 = n405 & n407;
  assign n409 = ~n383 & ~n408;
  assign n410 = ~pi017 & n377;
  assign n411 = n363 & n410;
  assign n412 = pi001 & ~pi054;
  assign n413 = ~n411 & ~n412;
  assign n414 = ~n409 & n413;
  assign po016 = ~n361 | ~n414;
  assign n416 = ~pi046 & ~pi050;
  assign n417 = ~pi041 & ~pi043;
  assign n418 = n416 & n417;
  assign n419 = ~pi042 & ~pi044;
  assign n420 = ~pi038 & ~pi040;
  assign n421 = n419 & n420;
  assign n422 = n418 & n421;
  assign n423 = ~pi015 & ~pi049;
  assign n424 = ~pi002 & ~pi020;
  assign n425 = n423 & n424;
  assign n426 = ~pi024 & ~pi045;
  assign n427 = ~pi047 & ~pi048;
  assign n428 = n426 & n427;
  assign n429 = n425 & n428;
  assign n430 = n422 & n429;
  assign n431 = pi082 & ~n430;
  assign n432 = pi122 & pi127;
  assign n433 = ~pi002 & n432;
  assign n434 = pi065 & ~n432;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~n431 & n435;
  assign n437 = ~pi015 & ~pi024;
  assign n438 = ~pi045 & ~pi047;
  assign n439 = ~pi043 & ~pi048;
  assign n440 = ~pi040 & n419;
  assign n441 = ~pi041 & n416;
  assign n442 = ~pi038 & n441;
  assign n443 = n440 & n442;
  assign n444 = n439 & n443;
  assign n445 = n438 & n444;
  assign n446 = ~pi020 & ~pi049;
  assign n447 = n445 & n446;
  assign n448 = n437 & n447;
  assign n449 = ~pi002 & n448;
  assign n450 = pi002 & ~n448;
  assign n451 = ~n449 & ~n450;
  assign n452 = n431 & ~n451;
  assign n453 = ~n436 & ~n452;
  assign po017 = ~pi129 & ~n453;
  assign n455 = ~pi113 & ~pi123;
  assign n456 = pi000 & n455;
  assign n457 = ~pi017 & n371;
  assign n458 = ~pi006 & ~pi012;
  assign n459 = ~pi014 & n384;
  assign n460 = n327 & n459;
  assign n461 = ~pi013 & n460;
  assign n462 = n458 & n461;
  assign n463 = n457 & n462;
  assign n464 = ~pi061 & ~pi118;
  assign n465 = ~n463 & n464;
  assign n466 = ~pi007 & ~pi008;
  assign n467 = ~pi021 & n466;
  assign n468 = ~pi019 & n467;
  assign n469 = n464 & ~n468;
  assign n470 = ~n465 & ~n469;
  assign n471 = ~n456 & n470;
  assign po018 = ~pi129 & ~n471;
  assign n473 = ~pi014 & n332;
  assign n474 = n303 & n397;
  assign n475 = n406 & n474;
  assign n476 = n473 & n475;
  assign n477 = pi054 & n304;
  assign n478 = n301 & n477;
  assign n479 = n302 & n397;
  assign n480 = n478 & n479;
  assign n481 = ~n476 & n480;
  assign n482 = ~pi017 & n481;
  assign n483 = pi004 & ~pi054;
  assign n484 = ~n482 & ~n483;
  assign po019 = n361 & ~n484;
  assign n486 = ~pi025 & pi028;
  assign n487 = pi054 & ~pi059;
  assign n488 = n486 & n487;
  assign n489 = n476 & n488;
  assign n490 = ~pi029 & n489;
  assign n491 = pi005 & ~pi054;
  assign n492 = ~n490 & ~n491;
  assign po020 = n361 & ~n492;
  assign n494 = pi025 & ~pi028;
  assign n495 = ~pi029 & n476;
  assign n496 = n487 & n495;
  assign n497 = n494 & n496;
  assign n498 = pi006 & ~pi054;
  assign n499 = ~n497 & ~n498;
  assign po021 = n361 & ~n499;
  assign n501 = ~pi017 & pi054;
  assign n502 = n473 & n474;
  assign n503 = ~n476 & n502;
  assign n504 = n304 & n503;
  assign n505 = n501 & n504;
  assign n506 = pi007 & ~pi054;
  assign n507 = ~n505 & ~n506;
  assign po022 = n361 & ~n507;
  assign n509 = ~pi008 & pi054;
  assign n510 = n503 & n509;
  assign n511 = n323 & n510;
  assign n512 = pi008 & ~pi054;
  assign n513 = ~n511 & ~n512;
  assign po023 = n361 & ~n513;
  assign n515 = ~pi054 & n361;
  assign n516 = pi009 & n515;
  assign n517 = ~pi017 & n304;
  assign n518 = pi054 & n361;
  assign n519 = ~n476 & n518;
  assign n520 = n324 & n519;
  assign n521 = n301 & n520;
  assign n522 = n517 & n521;
  assign n523 = ~pi016 & n303;
  assign n524 = n295 & n523;
  assign n525 = ~pi018 & n524;
  assign n526 = n522 & n525;
  assign po024 = n516 | n526;
  assign n528 = pi054 & n332;
  assign n529 = n323 & n474;
  assign n530 = ~n476 & n529;
  assign n531 = n335 & n530;
  assign n532 = n528 & n531;
  assign n533 = pi010 & ~pi054;
  assign n534 = ~n532 & ~n533;
  assign po025 = n361 & ~n534;
  assign n536 = pi011 & n515;
  assign n537 = n365 & n467;
  assign n538 = ~pi013 & n537;
  assign n539 = n323 & n538;
  assign n540 = n294 & n328;
  assign n541 = n518 & n540;
  assign n542 = ~n476 & n541;
  assign n543 = n539 & n542;
  assign po026 = n536 | n543;
  assign n545 = pi012 & n515;
  assign n546 = ~pi010 & n299;
  assign n547 = ~pi016 & n302;
  assign n548 = n518 & n547;
  assign n549 = n371 & n467;
  assign n550 = ~pi012 & n549;
  assign n551 = n323 & n550;
  assign n552 = n548 & n551;
  assign n553 = n546 & n552;
  assign n554 = ~n476 & n553;
  assign po027 = n545 | n554;
  assign n556 = ~pi025 & ~pi028;
  assign n557 = pi029 & n556;
  assign n558 = n476 & n557;
  assign n559 = n487 & n558;
  assign n560 = pi013 & ~pi054;
  assign n561 = ~n559 & ~n560;
  assign po028 = n361 & ~n561;
  assign n563 = ~pi014 & pi054;
  assign n564 = n474 & n517;
  assign n565 = ~n476 & n564;
  assign n566 = n466 & n565;
  assign n567 = n563 & n566;
  assign n568 = pi014 & ~pi054;
  assign n569 = ~n567 & ~n568;
  assign po029 = n361 & ~n569;
  assign n571 = ~pi049 & n426;
  assign n572 = ~pi048 & n571;
  assign n573 = ~pi044 & ~pi050;
  assign n574 = ~pi042 & n573;
  assign n575 = ~pi038 & n574;
  assign n576 = ~pi040 & n575;
  assign n577 = ~pi046 & ~pi047;
  assign n578 = n576 & n577;
  assign n579 = n417 & n578;
  assign n580 = n572 & n579;
  assign n581 = pi015 & n580;
  assign n582 = ~pi015 & ~n580;
  assign n583 = ~n581 & ~n582;
  assign n584 = n431 & n583;
  assign n585 = ~pi070 & ~n432;
  assign n586 = pi015 & n432;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n431 & ~n587;
  assign n589 = ~n584 & ~n588;
  assign po030 = ~pi129 & ~n589;
  assign n591 = pi016 & n515;
  assign n592 = n366 & n371;
  assign n593 = ~pi017 & n592;
  assign n594 = ~pi013 & ~pi016;
  assign n595 = n466 & n594;
  assign n596 = n459 & n595;
  assign n597 = n304 & n596;
  assign n598 = n593 & n597;
  assign n599 = n519 & n598;
  assign po031 = n591 | n599;
  assign n601 = n476 & n556;
  assign n602 = pi054 & n601;
  assign n603 = ~pi029 & n602;
  assign n604 = pi059 & n603;
  assign n605 = pi017 & ~pi054;
  assign n606 = ~n604 & ~n605;
  assign po032 = n361 & ~n606;
  assign n608 = pi018 & n515;
  assign n609 = ~pi008 & n303;
  assign n610 = n473 & n593;
  assign n611 = n304 & n610;
  assign n612 = n609 & n611;
  assign n613 = n519 & n612;
  assign po033 = n608 | n613;
  assign n615 = n335 & ~n476;
  assign n616 = n502 & n615;
  assign n617 = ~pi019 & n518;
  assign n618 = n616 & n617;
  assign n619 = pi019 & n515;
  assign po034 = n618 | n619;
  assign n621 = pi020 & n432;
  assign n622 = ~pi071 & ~n432;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~n431 & ~n623;
  assign n625 = n423 & n426;
  assign n626 = n416 & n421;
  assign n627 = ~pi041 & ~pi047;
  assign n628 = n626 & n627;
  assign n629 = n439 & n628;
  assign n630 = n625 & n629;
  assign n631 = pi020 & ~n630;
  assign n632 = ~pi020 & n625;
  assign n633 = n629 & n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = n431 & ~n634;
  assign n636 = ~n624 & ~n635;
  assign po035 = ~pi129 & ~n636;
  assign n638 = ~pi017 & n518;
  assign n639 = n616 & n638;
  assign n640 = pi021 & n515;
  assign po036 = n639 | n640;
  assign n642 = pi022 & n515;
  assign n643 = n325 & n467;
  assign n644 = n462 & n643;
  assign n645 = ~n476 & n644;
  assign n646 = n323 & n645;
  assign n647 = n518 & n646;
  assign po037 = n642 | n647;
  assign n649 = pi061 & ~pi129;
  assign n650 = ~pi023 & pi055;
  assign po038 = n649 & ~n650;
  assign n652 = ~pi024 & n445;
  assign n653 = pi024 & ~n445;
  assign n654 = ~n652 & ~n653;
  assign n655 = n431 & ~n654;
  assign n656 = pi024 & n432;
  assign n657 = ~pi063 & ~n432;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n431 & ~n658;
  assign n660 = ~n655 & ~n659;
  assign po039 = ~pi129 & ~n660;
  assign n662 = ~pi026 & pi027;
  assign n663 = ~pi053 & ~pi058;
  assign n664 = n662 & n663;
  assign n665 = ~pi085 & n664;
  assign n666 = ~pi039 & ~pi052;
  assign n667 = ~pi051 & n666;
  assign n668 = pi116 & n667;
  assign n669 = n665 & n668;
  assign n670 = pi026 & ~pi027;
  assign n671 = n663 & n670;
  assign n672 = ~pi085 & n671;
  assign n673 = pi116 & ~n667;
  assign n674 = n672 & n673;
  assign n675 = ~n669 & ~n674;
  assign n676 = ~pi026 & ~pi027;
  assign n677 = ~pi058 & n676;
  assign n678 = ~pi053 & n677;
  assign n679 = pi085 & n678;
  assign n680 = ~n665 & ~n679;
  assign n681 = pi025 & ~pi116;
  assign n682 = ~n680 & n681;
  assign n683 = pi116 & n679;
  assign n684 = pi100 & n683;
  assign n685 = ~n682 & ~n684;
  assign n686 = ~pi097 & ~pi100;
  assign n687 = ~pi095 & n686;
  assign n688 = ~pi110 & ~n687;
  assign n689 = ~pi085 & n678;
  assign n690 = n688 & n689;
  assign n691 = ~pi096 & n690;
  assign n692 = pi100 & n691;
  assign n693 = ~n688 & n689;
  assign n694 = pi025 & n693;
  assign n695 = ~n692 & ~n694;
  assign n696 = ~pi026 & ~pi085;
  assign n697 = ~pi027 & n696;
  assign n698 = ~pi058 & n697;
  assign n699 = pi053 & n698;
  assign n700 = ~pi053 & pi058;
  assign n701 = n697 & n700;
  assign n702 = ~n699 & ~n701;
  assign n703 = ~n672 & n702;
  assign n704 = n681 & ~n703;
  assign n705 = n695 & ~n704;
  assign n706 = n685 & n705;
  assign n707 = n675 & n706;
  assign po040 = n361 & ~n707;
  assign n709 = ~n672 & ~n679;
  assign n710 = pi026 & ~n709;
  assign n711 = ~pi116 & n710;
  assign n712 = ~n674 & ~n711;
  assign n713 = ~n684 & n712;
  assign n714 = pi026 & n689;
  assign n715 = ~n688 & n714;
  assign n716 = n713 & ~n715;
  assign n717 = ~n692 & n716;
  assign po041 = n361 & ~n717;
  assign n719 = ~pi100 & pi116;
  assign n720 = n679 & n719;
  assign n721 = n665 & n673;
  assign n722 = pi027 & ~n680;
  assign n723 = ~pi116 & n722;
  assign n724 = ~n721 & ~n723;
  assign n725 = ~n720 & n724;
  assign n726 = pi027 & n689;
  assign n727 = ~n688 & n726;
  assign n728 = n725 & ~n727;
  assign n729 = ~pi096 & ~pi100;
  assign n730 = n690 & n729;
  assign n731 = pi095 & n730;
  assign n732 = n728 & ~n731;
  assign po042 = n361 & ~n732;
  assign n734 = pi028 & ~n688;
  assign n735 = n689 & n734;
  assign n736 = pi028 & ~pi116;
  assign n737 = ~n720 & ~n736;
  assign n738 = ~n709 & ~n737;
  assign n739 = n668 & n672;
  assign n740 = ~n738 & ~n739;
  assign n741 = ~n665 & n702;
  assign n742 = n736 & ~n741;
  assign n743 = ~n721 & ~n742;
  assign n744 = n740 & n743;
  assign n745 = ~n731 & n744;
  assign n746 = ~n735 & n745;
  assign po043 = n361 & ~n746;
  assign n748 = pi029 & ~n688;
  assign n749 = n689 & n748;
  assign n750 = ~pi095 & n730;
  assign n751 = pi116 & n701;
  assign n752 = pi097 & n751;
  assign n753 = ~n679 & ~n701;
  assign n754 = pi029 & ~pi116;
  assign n755 = ~n753 & n754;
  assign n756 = ~n752 & ~n755;
  assign n757 = ~n750 & n756;
  assign n758 = ~n749 & n757;
  assign n759 = ~n672 & ~n699;
  assign n760 = ~n665 & n759;
  assign n761 = n754 & ~n760;
  assign n762 = n758 & ~n761;
  assign po044 = n361 & ~n762;
  assign n764 = pi088 & pi106;
  assign n765 = pi060 & pi109;
  assign n766 = pi030 & ~pi109;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~pi106 & ~n767;
  assign n769 = ~n764 & ~n768;
  assign po045 = ~pi129 & ~n769;
  assign n771 = pi089 & pi106;
  assign n772 = pi031 & ~pi109;
  assign n773 = pi030 & pi109;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~pi106 & ~n774;
  assign n776 = ~n771 & ~n775;
  assign po046 = ~pi129 & ~n776;
  assign n778 = pi099 & pi106;
  assign n779 = pi032 & ~pi109;
  assign n780 = pi031 & pi109;
  assign n781 = ~n779 & ~n780;
  assign n782 = ~pi106 & ~n781;
  assign n783 = ~n778 & ~n782;
  assign po047 = ~pi129 & ~n783;
  assign n785 = pi090 & pi106;
  assign n786 = pi033 & ~pi109;
  assign n787 = pi032 & pi109;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~pi106 & ~n788;
  assign n790 = ~n785 & ~n789;
  assign po048 = ~pi129 & ~n790;
  assign n792 = pi091 & pi106;
  assign n793 = pi034 & ~pi109;
  assign n794 = pi033 & pi109;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~pi106 & ~n795;
  assign n797 = ~n792 & ~n796;
  assign po049 = ~pi129 & ~n797;
  assign n799 = pi092 & pi106;
  assign n800 = pi035 & ~pi109;
  assign n801 = pi034 & pi109;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~pi106 & ~n802;
  assign n804 = ~n799 & ~n803;
  assign po050 = ~pi129 & ~n804;
  assign n806 = pi098 & pi106;
  assign n807 = pi036 & ~pi109;
  assign n808 = pi035 & pi109;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~pi106 & ~n809;
  assign n811 = ~n806 & ~n810;
  assign po051 = ~pi129 & ~n811;
  assign n813 = pi093 & pi106;
  assign n814 = pi037 & ~pi109;
  assign n815 = pi036 & pi109;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~pi106 & ~n816;
  assign n818 = ~n813 & ~n817;
  assign po052 = ~pi129 & ~n818;
  assign n820 = pi038 & ~n440;
  assign n821 = ~n421 & ~n820;
  assign n822 = n431 & ~n821;
  assign n823 = ~pi074 & ~n432;
  assign n824 = pi038 & n432;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n431 & ~n825;
  assign n827 = ~n822 & ~n826;
  assign po053 = ~pi129 & ~n827;
  assign n829 = pi106 & ~pi129;
  assign n830 = ~pi039 & ~pi109;
  assign n831 = ~pi051 & ~pi052;
  assign n832 = pi039 & ~n831;
  assign n833 = ~n667 & ~n832;
  assign n834 = pi109 & n833;
  assign n835 = ~n830 & ~n834;
  assign n836 = ~pi129 & n835;
  assign po054 = n829 | n836;
  assign n838 = pi040 & n432;
  assign n839 = ~pi073 & ~n432;
  assign n840 = ~n838 & ~n839;
  assign n841 = ~n431 & ~n840;
  assign n842 = pi040 & ~n419;
  assign n843 = ~n440 & ~n842;
  assign n844 = n431 & ~n843;
  assign n845 = ~n841 & ~n844;
  assign po055 = ~pi129 & ~n845;
  assign n847 = ~pi076 & ~n432;
  assign n848 = pi041 & n432;
  assign n849 = ~n847 & ~n848;
  assign n850 = ~n431 & ~n849;
  assign n851 = ~pi041 & ~n626;
  assign n852 = pi041 & n626;
  assign n853 = ~n851 & ~n852;
  assign n854 = n431 & n853;
  assign n855 = ~n850 & ~n854;
  assign po056 = ~pi129 & ~n855;
  assign n857 = pi042 & n432;
  assign n858 = ~pi072 & ~n432;
  assign n859 = ~n857 & ~n858;
  assign n860 = ~n431 & ~n859;
  assign n861 = pi042 & pi044;
  assign n862 = ~n419 & ~n861;
  assign n863 = n431 & ~n862;
  assign n864 = ~n860 & ~n863;
  assign po057 = ~pi129 & ~n864;
  assign n866 = pi043 & n432;
  assign n867 = ~pi077 & ~n432;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n431 & ~n868;
  assign n870 = ~pi043 & ~n443;
  assign n871 = pi043 & n443;
  assign n872 = ~n870 & ~n871;
  assign n873 = n431 & n872;
  assign n874 = ~n869 & ~n873;
  assign po058 = ~pi129 & ~n874;
  assign n876 = pi044 & n432;
  assign n877 = ~pi067 & ~n432;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~n431 & ~n878;
  assign n880 = ~pi044 & n431;
  assign n881 = ~n879 & ~n880;
  assign po059 = ~pi129 & ~n881;
  assign n883 = pi045 & n432;
  assign n884 = ~pi068 & ~n432;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n431 & ~n885;
  assign n887 = pi045 & ~n629;
  assign n888 = ~pi045 & n629;
  assign n889 = ~n887 & ~n888;
  assign n890 = n431 & ~n889;
  assign n891 = ~n886 & ~n890;
  assign po060 = ~pi129 & ~n891;
  assign n893 = pi046 & n576;
  assign n894 = ~pi046 & ~n576;
  assign n895 = ~n893 & ~n894;
  assign n896 = n431 & n895;
  assign n897 = pi046 & n432;
  assign n898 = ~pi075 & ~n432;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~n431 & ~n899;
  assign n901 = ~n896 & ~n900;
  assign po061 = ~pi129 & ~n901;
  assign n903 = pi047 & n432;
  assign n904 = ~pi064 & ~n432;
  assign n905 = ~n903 & ~n904;
  assign n906 = ~n431 & ~n905;
  assign n907 = pi047 & n422;
  assign n908 = ~pi047 & ~n422;
  assign n909 = ~n907 & ~n908;
  assign n910 = n431 & n909;
  assign n911 = ~n906 & ~n910;
  assign po062 = ~pi129 & ~n911;
  assign n913 = pi048 & n432;
  assign n914 = ~pi062 & ~n432;
  assign n915 = ~n913 & ~n914;
  assign n916 = ~n431 & ~n915;
  assign n917 = ~pi048 & n579;
  assign n918 = pi048 & ~n579;
  assign n919 = ~n917 & ~n918;
  assign n920 = n431 & ~n919;
  assign n921 = ~n916 & ~n920;
  assign po063 = ~pi129 & ~n921;
  assign n923 = pi049 & n432;
  assign n924 = ~pi069 & ~n432;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n431 & ~n925;
  assign n927 = n422 & n428;
  assign n928 = pi049 & ~n927;
  assign n929 = ~pi049 & n927;
  assign n930 = ~n928 & ~n929;
  assign n931 = n431 & ~n930;
  assign n932 = ~n926 & ~n931;
  assign po064 = ~pi129 & ~n932;
  assign n934 = pi050 & n421;
  assign n935 = ~pi050 & ~n421;
  assign n936 = ~n934 & ~n935;
  assign n937 = n431 & n936;
  assign n938 = pi050 & n432;
  assign n939 = ~pi066 & ~n432;
  assign n940 = ~n938 & ~n939;
  assign n941 = ~n431 & ~n940;
  assign n942 = ~n937 & ~n941;
  assign po065 = ~pi129 & ~n942;
  assign n944 = pi051 & pi109;
  assign n945 = ~pi051 & ~pi109;
  assign n946 = ~n944 & ~n945;
  assign n947 = ~pi129 & n946;
  assign po066 = n829 | n947;
  assign n949 = ~pi052 & ~pi109;
  assign n950 = pi051 & pi052;
  assign n951 = ~n831 & ~n950;
  assign n952 = pi109 & n951;
  assign n953 = ~n949 & ~n952;
  assign n954 = ~pi129 & n953;
  assign po067 = n829 | n954;
  assign n956 = pi053 & n693;
  assign n957 = pi053 & ~n702;
  assign n958 = ~pi116 & n957;
  assign n959 = ~n956 & ~n958;
  assign n960 = ~n750 & n959;
  assign n961 = ~n752 & n960;
  assign po068 = n361 & ~n961;
  assign n963 = ~n431 & ~n432;
  assign po069 = pi129 | n963;
  assign n965 = pi114 & ~pi122;
  assign po129 = pi123 | pi129;
  assign po070 = n965 & ~po129;
  assign n968 = pi094 & pi116;
  assign n969 = pi037 & ~pi116;
  assign n970 = ~n968 & ~n969;
  assign n971 = n672 & ~n970;
  assign n972 = pi037 & n689;
  assign n973 = ~n971 & ~n972;
  assign n974 = ~pi094 & ~pi116;
  assign n975 = n701 & ~n974;
  assign n976 = n973 & ~n975;
  assign n977 = ~n665 & ~n699;
  assign n978 = ~n679 & n977;
  assign n979 = pi037 & ~n978;
  assign n980 = n976 & ~n979;
  assign po071 = n361 & ~n980;
  assign n982 = pi057 & ~n760;
  assign n983 = pi057 & ~pi116;
  assign n984 = pi060 & pi116;
  assign n985 = ~n983 & ~n984;
  assign n986 = n701 & ~n985;
  assign n987 = ~n679 & ~n689;
  assign n988 = pi057 & ~n987;
  assign n989 = ~n986 & ~n988;
  assign n990 = ~n982 & n989;
  assign po072 = n361 & ~n990;
  assign n992 = pi058 & ~pi116;
  assign n993 = ~n665 & ~n701;
  assign n994 = n992 & ~n993;
  assign n995 = ~n669 & ~n994;
  assign n996 = n672 & n992;
  assign n997 = n995 & ~n996;
  assign n998 = ~n739 & n997;
  assign po073 = n361 & ~n998;
  assign n1000 = pi059 & ~pi116;
  assign n1001 = ~n703 & n1000;
  assign n1002 = pi059 & ~n688;
  assign n1003 = pi096 & n688;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = n689 & ~n1004;
  assign n1006 = ~n680 & n1000;
  assign n1007 = ~n1005 & ~n1006;
  assign n1008 = ~n1001 & n1007;
  assign po074 = n361 & ~n1008;
  assign n1010 = ~pi117 & ~pi122;
  assign n1011 = pi060 & ~n1010;
  assign n1012 = pi123 & n1010;
  assign po075 = n1011 | n1012;
  assign n1014 = ~pi114 & ~pi122;
  assign n1015 = pi123 & ~pi129;
  assign po076 = n1014 & n1015;
  assign n1017 = pi131 & pi133;
  assign n1018 = pi132 & n1017;
  assign n1019 = ~pi137 & ~pi138;
  assign n1020 = ~pi136 & n1019;
  assign n1021 = pi136 & n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = ~n1020 & ~n1022;
  assign n1024 = ~pi062 & ~n1023;
  assign n1025 = pi140 & n1021;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = n1018 & ~n1026;
  assign n1028 = ~pi062 & ~n1018;
  assign n1029 = ~n1027 & ~n1028;
  assign po077 = pi129 | ~n1029;
  assign n1031 = ~pi063 & ~n1023;
  assign n1032 = pi142 & n1021;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = n1018 & ~n1033;
  assign n1035 = ~pi063 & ~n1018;
  assign n1036 = ~n1034 & ~n1035;
  assign po078 = pi129 | ~n1036;
  assign n1038 = ~pi064 & ~n1023;
  assign n1039 = pi139 & n1021;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = n1018 & ~n1040;
  assign n1042 = ~pi064 & ~n1018;
  assign n1043 = ~n1041 & ~n1042;
  assign po079 = pi129 | ~n1043;
  assign n1045 = ~pi065 & ~n1023;
  assign n1046 = pi146 & n1021;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = n1018 & ~n1047;
  assign n1049 = ~pi065 & ~n1018;
  assign n1050 = ~n1048 & ~n1049;
  assign po080 = pi129 | ~n1050;
  assign n1052 = ~n1021 & ~n1022;
  assign n1053 = ~pi066 & ~n1052;
  assign n1054 = pi143 & n1020;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1018 & ~n1055;
  assign n1057 = ~pi066 & ~n1018;
  assign n1058 = ~n1056 & ~n1057;
  assign po081 = pi129 | ~n1058;
  assign n1060 = ~pi067 & ~n1052;
  assign n1061 = pi139 & n1020;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = n1018 & ~n1062;
  assign n1064 = ~pi067 & ~n1018;
  assign n1065 = ~n1063 & ~n1064;
  assign po082 = pi129 | ~n1065;
  assign n1067 = ~pi068 & ~n1023;
  assign n1068 = pi141 & n1021;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = n1018 & ~n1069;
  assign n1071 = ~pi068 & ~n1018;
  assign n1072 = ~n1070 & ~n1071;
  assign po083 = pi129 | ~n1072;
  assign n1074 = ~pi069 & ~n1023;
  assign n1075 = pi143 & n1021;
  assign n1076 = ~n1074 & ~n1075;
  assign n1077 = n1018 & ~n1076;
  assign n1078 = ~pi069 & ~n1018;
  assign n1079 = ~n1077 & ~n1078;
  assign po084 = pi129 | ~n1079;
  assign n1081 = ~pi070 & ~n1023;
  assign n1082 = pi144 & n1021;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = n1018 & ~n1083;
  assign n1085 = ~pi070 & ~n1018;
  assign n1086 = ~n1084 & ~n1085;
  assign po085 = pi129 | ~n1086;
  assign n1088 = ~pi071 & ~n1023;
  assign n1089 = pi145 & n1021;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = n1018 & ~n1090;
  assign n1092 = ~pi071 & ~n1018;
  assign n1093 = ~n1091 & ~n1092;
  assign po086 = pi129 | ~n1093;
  assign n1095 = ~pi072 & ~n1052;
  assign n1096 = pi140 & n1020;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = n1018 & ~n1097;
  assign n1099 = ~pi072 & ~n1018;
  assign n1100 = ~n1098 & ~n1099;
  assign po087 = pi129 | ~n1100;
  assign n1102 = ~pi073 & ~n1052;
  assign n1103 = pi141 & n1020;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = n1018 & ~n1104;
  assign n1106 = ~pi073 & ~n1018;
  assign n1107 = ~n1105 & ~n1106;
  assign po088 = pi129 | ~n1107;
  assign n1109 = ~pi074 & ~n1052;
  assign n1110 = pi142 & n1020;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n1018 & ~n1111;
  assign n1113 = ~pi074 & ~n1018;
  assign n1114 = ~n1112 & ~n1113;
  assign po089 = pi129 | ~n1114;
  assign n1116 = ~pi075 & ~n1052;
  assign n1117 = pi144 & n1020;
  assign n1118 = ~n1116 & ~n1117;
  assign n1119 = n1018 & ~n1118;
  assign n1120 = ~pi075 & ~n1018;
  assign n1121 = ~n1119 & ~n1120;
  assign po090 = pi129 | ~n1121;
  assign n1123 = ~pi076 & ~n1052;
  assign n1124 = pi145 & n1020;
  assign n1125 = ~n1123 & ~n1124;
  assign n1126 = n1018 & ~n1125;
  assign n1127 = ~pi076 & ~n1018;
  assign n1128 = ~n1126 & ~n1127;
  assign po091 = pi129 | ~n1128;
  assign n1130 = ~pi077 & ~n1052;
  assign n1131 = pi146 & n1020;
  assign n1132 = ~n1130 & ~n1131;
  assign n1133 = n1018 & ~n1132;
  assign n1134 = ~pi077 & ~n1018;
  assign n1135 = ~n1133 & ~n1134;
  assign po092 = pi129 | ~n1135;
  assign n1137 = pi137 & ~pi138;
  assign n1138 = ~pi136 & n1137;
  assign n1139 = pi078 & ~n1138;
  assign n1140 = pi142 & n1138;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = n1018 & ~n1141;
  assign n1143 = pi078 & ~n1018;
  assign n1144 = ~n1142 & ~n1143;
  assign po093 = ~pi129 & ~n1144;
  assign n1146 = pi079 & ~n1138;
  assign n1147 = pi143 & n1138;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = n1018 & ~n1148;
  assign n1150 = pi079 & ~n1018;
  assign n1151 = ~n1149 & ~n1150;
  assign po094 = ~pi129 & ~n1151;
  assign n1153 = pi080 & ~n1138;
  assign n1154 = pi144 & n1138;
  assign n1155 = ~n1153 & ~n1154;
  assign n1156 = n1018 & ~n1155;
  assign n1157 = pi080 & ~n1018;
  assign n1158 = ~n1156 & ~n1157;
  assign po095 = ~pi129 & ~n1158;
  assign n1160 = pi081 & ~n1138;
  assign n1161 = pi145 & n1138;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = n1018 & ~n1162;
  assign n1164 = pi081 & ~n1018;
  assign n1165 = ~n1163 & ~n1164;
  assign po096 = ~pi129 & ~n1165;
  assign n1167 = pi082 & ~n1138;
  assign n1168 = pi146 & n1138;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = n1018 & ~n1169;
  assign n1171 = pi082 & ~n1018;
  assign n1172 = ~n1170 & ~n1171;
  assign po097 = ~pi129 & ~n1172;
  assign n1174 = pi087 & n1138;
  assign n1175 = ~pi062 & n1021;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~pi072 & n1020;
  assign n1178 = pi137 & pi138;
  assign n1179 = ~pi136 & n1178;
  assign n1180 = ~pi115 & n1179;
  assign n1181 = ~pi137 & pi138;
  assign n1182 = pi136 & n1181;
  assign n1183 = pi089 & n1182;
  assign n1184 = ~n1180 & ~n1183;
  assign n1185 = ~pi136 & n1181;
  assign n1186 = pi119 & n1185;
  assign n1187 = pi136 & n1137;
  assign n1188 = pi031 & n1187;
  assign n1189 = ~n1186 & ~n1188;
  assign n1190 = n1184 & n1189;
  assign n1191 = ~n1177 & n1190;
  assign po098 = ~n1176 | ~n1191;
  assign n1193 = pi084 & ~n1138;
  assign n1194 = pi141 & n1138;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = n1018 & ~n1195;
  assign n1197 = pi084 & ~n1018;
  assign n1198 = ~n1196 & ~n1197;
  assign po099 = ~pi129 & ~n1198;
  assign n1200 = pi085 & n679;
  assign n1201 = ~pi116 & n1200;
  assign n1202 = pi085 & ~n688;
  assign n1203 = ~n1003 & ~n1202;
  assign n1204 = n689 & ~n1203;
  assign n1205 = ~n1201 & ~n1204;
  assign po100 = n361 & ~n1205;
  assign n1207 = pi086 & ~n1138;
  assign n1208 = pi139 & n1138;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n1018 & ~n1209;
  assign n1211 = pi086 & ~n1018;
  assign n1212 = ~n1210 & ~n1211;
  assign po101 = ~pi129 & ~n1212;
  assign n1214 = pi087 & ~n1138;
  assign n1215 = pi140 & n1138;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = n1018 & ~n1216;
  assign n1218 = pi087 & ~n1018;
  assign n1219 = ~n1217 & ~n1218;
  assign po102 = ~pi129 & ~n1219;
  assign n1221 = pi088 & ~n1187;
  assign n1222 = pi139 & n1187;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = n1018 & ~n1223;
  assign n1225 = pi088 & ~n1018;
  assign n1226 = ~n1224 & ~n1225;
  assign po103 = ~pi129 & ~n1226;
  assign n1228 = pi089 & ~n1187;
  assign n1229 = pi140 & n1187;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = n1018 & ~n1230;
  assign n1232 = pi089 & ~n1018;
  assign n1233 = ~n1231 & ~n1232;
  assign po104 = ~pi129 & ~n1233;
  assign n1235 = pi090 & ~n1187;
  assign n1236 = pi142 & n1187;
  assign n1237 = ~n1235 & ~n1236;
  assign n1238 = n1018 & ~n1237;
  assign n1239 = pi090 & ~n1018;
  assign n1240 = ~n1238 & ~n1239;
  assign po105 = ~pi129 & ~n1240;
  assign n1242 = pi091 & ~n1187;
  assign n1243 = pi143 & n1187;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = n1018 & ~n1244;
  assign n1246 = pi091 & ~n1018;
  assign n1247 = ~n1245 & ~n1246;
  assign po106 = ~pi129 & ~n1247;
  assign n1249 = pi092 & ~n1187;
  assign n1250 = pi144 & n1187;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = n1018 & ~n1251;
  assign n1253 = pi092 & ~n1018;
  assign n1254 = ~n1252 & ~n1253;
  assign po107 = ~pi129 & ~n1254;
  assign n1256 = pi093 & ~n1187;
  assign n1257 = pi146 & n1187;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = n1018 & ~n1258;
  assign n1260 = pi093 & ~n1018;
  assign n1261 = ~n1259 & ~n1260;
  assign po108 = ~pi129 & ~n1261;
  assign n1263 = pi082 & n1181;
  assign n1264 = ~pi136 & n1263;
  assign n1265 = pi142 & n1264;
  assign n1266 = pi094 & ~n1264;
  assign n1267 = ~n1265 & ~n1266;
  assign n1268 = n1018 & ~n1267;
  assign n1269 = pi094 & ~n1018;
  assign n1270 = ~n1268 & ~n1269;
  assign po109 = ~pi129 & ~n1270;
  assign n1272 = ~pi003 & ~pi110;
  assign n1273 = ~n1018 & n1272;
  assign n1274 = pi095 & n1273;
  assign n1275 = ~pi143 & n1264;
  assign n1276 = ~pi095 & ~n1264;
  assign n1277 = ~n1275 & ~n1276;
  assign n1278 = n1018 & n1277;
  assign n1279 = ~n1274 & ~n1278;
  assign po110 = ~pi129 & ~n1279;
  assign n1281 = pi096 & n1273;
  assign n1282 = ~pi146 & n1264;
  assign n1283 = ~pi096 & ~n1264;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = n1018 & n1284;
  assign n1286 = ~n1281 & ~n1285;
  assign po111 = ~pi129 & ~n1286;
  assign n1288 = pi097 & n1273;
  assign n1289 = pi145 & n1264;
  assign n1290 = pi097 & ~n1264;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = n1018 & ~n1291;
  assign n1293 = ~n1288 & ~n1292;
  assign po112 = ~pi129 & ~n1293;
  assign n1295 = pi098 & ~n1187;
  assign n1296 = pi145 & n1187;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n1018 & ~n1297;
  assign n1299 = pi098 & ~n1018;
  assign n1300 = ~n1298 & ~n1299;
  assign po113 = ~pi129 & ~n1300;
  assign n1302 = pi099 & ~n1187;
  assign n1303 = pi141 & n1187;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n1018 & ~n1304;
  assign n1306 = pi099 & ~n1018;
  assign n1307 = ~n1305 & ~n1306;
  assign po114 = ~pi129 & ~n1307;
  assign n1309 = pi100 & n1273;
  assign n1310 = ~pi144 & n1264;
  assign n1311 = ~pi100 & ~n1264;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = n1018 & n1312;
  assign n1314 = ~n1309 & ~n1313;
  assign po115 = ~pi129 & ~n1314;
  assign n1316 = pi082 & n1138;
  assign n1317 = ~pi065 & n1021;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = ~pi077 & n1020;
  assign n1320 = pi096 & n1179;
  assign n1321 = pi093 & n1182;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = pi124 & n1185;
  assign n1324 = pi037 & n1187;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = n1322 & n1325;
  assign n1327 = ~n1319 & n1326;
  assign po116 = ~n1318 | ~n1327;
  assign n1329 = pi079 & n1138;
  assign n1330 = ~pi069 & n1021;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = ~pi066 & n1020;
  assign n1333 = pi095 & n1179;
  assign n1334 = pi091 & n1182;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = pi034 & n1187;
  assign n1337 = n1335 & ~n1336;
  assign n1338 = ~n1332 & n1337;
  assign po117 = ~n1331 | ~n1338;
  assign n1340 = pi078 & n1138;
  assign n1341 = ~pi063 & n1021;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = ~pi074 & n1020;
  assign n1344 = pi094 & n1179;
  assign n1345 = pi090 & n1182;
  assign n1346 = ~n1344 & ~n1345;
  assign n1347 = pi033 & n1187;
  assign n1348 = n1346 & ~n1347;
  assign n1349 = ~n1343 & n1348;
  assign po118 = ~n1342 | ~n1349;
  assign n1351 = pi084 & n1138;
  assign n1352 = ~pi068 & n1021;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~pi073 & n1020;
  assign n1355 = ~pi112 & n1179;
  assign n1356 = pi099 & n1182;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = pi032 & n1187;
  assign n1359 = n1357 & ~n1358;
  assign n1360 = ~n1354 & n1359;
  assign po119 = ~n1353 | ~n1360;
  assign n1362 = pi080 & n1138;
  assign n1363 = ~pi070 & n1021;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = ~pi075 & n1020;
  assign n1366 = pi100 & n1179;
  assign n1367 = pi092 & n1182;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = pi125 & n1185;
  assign n1370 = pi035 & n1187;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = n1368 & n1371;
  assign n1373 = ~n1365 & n1372;
  assign po120 = ~n1364 | ~n1373;
  assign n1375 = n663 & n697;
  assign n1376 = pi085 & ~n1375;
  assign n1377 = pi116 & n1376;
  assign n1378 = ~pi085 & n1375;
  assign n1379 = n688 & n1378;
  assign n1380 = ~n1377 & ~n1379;
  assign po121 = n361 & ~n1380;
  assign n1382 = ~pi071 & n1021;
  assign n1383 = ~pi076 & n1020;
  assign n1384 = ~n1382 & ~n1383;
  assign n1385 = pi081 & n1138;
  assign n1386 = pi097 & n1179;
  assign n1387 = pi098 & n1182;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = pi023 & n1185;
  assign n1390 = pi036 & n1187;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = n1388 & n1391;
  assign n1393 = ~n1385 & n1392;
  assign po122 = ~n1384 | ~n1393;
  assign n1395 = pi111 & n1179;
  assign n1396 = pi088 & n1182;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = pi030 & n1187;
  assign n1399 = pi120 & n1185;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = pi086 & n1138;
  assign n1402 = ~pi064 & n1021;
  assign n1403 = ~n1401 & ~n1402;
  assign n1404 = ~pi067 & n1020;
  assign n1405 = n1403 & ~n1404;
  assign n1406 = n1400 & n1405;
  assign po123 = ~n1397 | ~n1406;
  assign n1408 = n662 & n673;
  assign n1409 = pi116 & n670;
  assign n1410 = ~n1408 & ~n1409;
  assign po124 = n361 & ~n1410;
  assign n1412 = pi116 & n361;
  assign n1413 = ~pi097 & n700;
  assign n1414 = pi053 & ~pi058;
  assign n1415 = ~n1413 & ~n1414;
  assign po125 = n1412 & ~n1415;
  assign n1417 = pi139 & n1264;
  assign n1418 = pi111 & ~n1264;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = ~pi129 & n1018;
  assign po126 = ~n1419 & n1420;
  assign n1422 = pi141 & n1264;
  assign n1423 = ~pi112 & ~n1264;
  assign n1424 = ~n1422 & ~n1423;
  assign po127 = n1420 & ~n1424;
  assign n1426 = ~pi113 & n515;
  assign n1427 = ~n369 & n518;
  assign po128 = n1426 | n1427;
  assign n1429 = pi140 & n1264;
  assign n1430 = ~pi115 & ~n1264;
  assign n1431 = ~n1429 & ~n1430;
  assign po130 = n1420 & ~n1431;
  assign n1433 = ~pi007 & ~pi009;
  assign n1434 = ~pi004 & ~pi012;
  assign n1435 = n1433 & n1434;
  assign po131 = n518 & ~n1435;
  assign po132 = ~pi122 | pi129;
  assign n1438 = n487 & n557;
  assign n1439 = ~pi054 & pi118;
  assign n1440 = ~n1438 & ~n1439;
  assign po133 = ~pi129 & ~n1440;
  assign n1442 = ~pi095 & ~pi100;
  assign po134 = ~pi129 & ~n1442;
  assign n1444 = ~pi111 & ~pi129;
  assign n1445 = ~pi120 & n1272;
  assign po135 = n1444 & ~n1445;
  assign n1447 = pi081 & pi120;
  assign po136 = ~pi129 & n1447;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi057 & ~pi129;
  assign n1452 = ~pi096 & pi125;
  assign n1453 = ~pi003 & ~n1452;
  assign po140 = ~pi129 & ~n1453;
  assign n1455 = pi132 & pi133;
  assign po141 = ~pi126 & n1455;
  assign po012 = 1'b1;
  assign po000 = pi108;
  assign po001 = pi083;
  assign po002 = pi104;
  assign po003 = pi103;
  assign po004 = pi102;
  assign po005 = pi105;
  assign po006 = pi107;
  assign po007 = pi101;
  assign po008 = pi126;
  assign po009 = pi121;
  assign po010 = pi001;
  assign po011 = pi000;
  assign po013 = pi130;
  assign po014 = pi128;
endmodule


